magic
tech gf180mcuD
magscale 1 5
timestamp 1764970766
<< metal1 >>
rect 336 6677 31864 6694
rect 336 6651 2233 6677
rect 2259 6651 2285 6677
rect 2311 6651 2337 6677
rect 2363 6651 12233 6677
rect 12259 6651 12285 6677
rect 12311 6651 12337 6677
rect 12363 6651 22233 6677
rect 22259 6651 22285 6677
rect 22311 6651 22337 6677
rect 22363 6651 31864 6677
rect 336 6634 31864 6651
rect 1863 6593 1889 6599
rect 1863 6561 1889 6567
rect 2983 6593 3009 6599
rect 2983 6561 3009 6567
rect 3767 6593 3793 6599
rect 3767 6561 3793 6567
rect 4887 6593 4913 6599
rect 4887 6561 4913 6567
rect 5671 6593 5697 6599
rect 5671 6561 5697 6567
rect 8695 6593 8721 6599
rect 8695 6561 8721 6567
rect 9479 6593 9505 6599
rect 9479 6561 9505 6567
rect 10599 6593 10625 6599
rect 10599 6561 10625 6567
rect 11383 6593 11409 6599
rect 11383 6561 11409 6567
rect 12503 6593 12529 6599
rect 12503 6561 12529 6567
rect 13287 6593 13313 6599
rect 26055 6593 26081 6599
rect 25433 6567 25439 6593
rect 25465 6567 25471 6593
rect 13287 6561 13313 6567
rect 26055 6561 26081 6567
rect 27455 6593 27481 6599
rect 27455 6561 27481 6567
rect 28239 6593 28265 6599
rect 28239 6561 28265 6567
rect 31263 6593 31289 6599
rect 31263 6561 31289 6567
rect 7457 6511 7463 6537
rect 7489 6511 7495 6537
rect 30249 6511 30255 6537
rect 30281 6511 30287 6537
rect 25607 6481 25633 6487
rect 849 6455 855 6481
rect 881 6455 887 6481
rect 2137 6455 2143 6481
rect 2169 6455 2175 6481
rect 3201 6455 3207 6481
rect 3233 6455 3239 6481
rect 3985 6455 3991 6481
rect 4017 6455 4023 6481
rect 5161 6455 5167 6481
rect 5193 6455 5199 6481
rect 5945 6455 5951 6481
rect 5977 6455 5983 6481
rect 6449 6455 6455 6481
rect 6481 6455 6487 6481
rect 7849 6455 7855 6481
rect 7881 6455 7887 6481
rect 8969 6455 8975 6481
rect 9001 6455 9007 6481
rect 9753 6455 9759 6481
rect 9785 6455 9791 6481
rect 10873 6455 10879 6481
rect 10905 6455 10911 6481
rect 11657 6455 11663 6481
rect 11689 6455 11695 6481
rect 12721 6455 12727 6481
rect 12753 6455 12759 6481
rect 13561 6455 13567 6481
rect 13593 6455 13599 6481
rect 14457 6455 14463 6481
rect 14489 6455 14495 6481
rect 25769 6455 25775 6481
rect 25801 6455 25807 6481
rect 27169 6455 27175 6481
rect 27201 6455 27207 6481
rect 27953 6455 27959 6481
rect 27985 6455 27991 6481
rect 29073 6455 29079 6481
rect 29105 6455 29111 6481
rect 29857 6455 29863 6481
rect 29889 6455 29895 6481
rect 30977 6455 30983 6481
rect 31009 6455 31015 6481
rect 25607 6449 25633 6455
rect 1247 6425 1273 6431
rect 1247 6393 1273 6399
rect 6959 6425 6985 6431
rect 6959 6393 6985 6399
rect 13959 6425 13985 6431
rect 29409 6399 29415 6425
rect 29441 6399 29447 6425
rect 13959 6393 13985 6399
rect 336 6285 31864 6302
rect 336 6259 1903 6285
rect 1929 6259 1955 6285
rect 1981 6259 2007 6285
rect 2033 6259 11903 6285
rect 11929 6259 11955 6285
rect 11981 6259 12007 6285
rect 12033 6259 21903 6285
rect 21929 6259 21955 6285
rect 21981 6259 22007 6285
rect 22033 6259 31864 6285
rect 336 6242 31864 6259
rect 3487 6201 3513 6207
rect 3487 6169 3513 6175
rect 4271 6201 4297 6207
rect 4271 6169 4297 6175
rect 5055 6201 5081 6207
rect 5055 6169 5081 6175
rect 5839 6201 5865 6207
rect 5839 6169 5865 6175
rect 8191 6201 8217 6207
rect 8191 6169 8217 6175
rect 8975 6201 9001 6207
rect 8975 6169 9001 6175
rect 9927 6201 9953 6207
rect 9927 6169 9953 6175
rect 11215 6201 11241 6207
rect 11215 6169 11241 6175
rect 11999 6201 12025 6207
rect 11999 6169 12025 6175
rect 12559 6201 12585 6207
rect 12559 6169 12585 6175
rect 26279 6201 26305 6207
rect 26279 6169 26305 6175
rect 27063 6201 27089 6207
rect 27063 6169 27089 6175
rect 27847 6201 27873 6207
rect 27847 6169 27873 6175
rect 28631 6201 28657 6207
rect 28631 6169 28657 6175
rect 14911 6145 14937 6151
rect 1801 6119 1807 6145
rect 1833 6119 1839 6145
rect 7513 6119 7519 6145
rect 7545 6119 7551 6145
rect 13449 6119 13455 6145
rect 13481 6119 13487 6145
rect 14911 6113 14937 6119
rect 15191 6145 15217 6151
rect 15191 6113 15217 6119
rect 15583 6145 15609 6151
rect 15583 6113 15609 6119
rect 17487 6145 17513 6151
rect 30305 6119 30311 6145
rect 30337 6119 30343 6145
rect 31089 6119 31095 6145
rect 31121 6119 31127 6145
rect 17487 6113 17513 6119
rect 15471 6089 15497 6095
rect 6057 6063 6063 6089
rect 6089 6063 6095 6089
rect 9193 6063 9199 6089
rect 9225 6063 9231 6089
rect 9417 6063 9423 6089
rect 9449 6063 9455 6089
rect 13729 6063 13735 6089
rect 13761 6063 13767 6089
rect 15471 6057 15497 6063
rect 17599 6089 17625 6095
rect 17599 6057 17625 6063
rect 20679 6089 20705 6095
rect 26049 6063 26055 6089
rect 26081 6063 26087 6089
rect 26777 6063 26783 6089
rect 26809 6063 26815 6089
rect 20679 6057 20705 6063
rect 17879 6033 17905 6039
rect 2193 6007 2199 6033
rect 2225 6007 2231 6033
rect 3761 6007 3767 6033
rect 3793 6007 3799 6033
rect 4545 6007 4551 6033
rect 4577 6007 4583 6033
rect 5329 6007 5335 6033
rect 5361 6007 5367 6033
rect 7065 6007 7071 6033
rect 7097 6007 7103 6033
rect 8465 6007 8471 6033
rect 8497 6007 8503 6033
rect 11489 6007 11495 6033
rect 11521 6007 11527 6033
rect 12273 6007 12279 6033
rect 12305 6007 12311 6033
rect 13057 6007 13063 6033
rect 13089 6007 13095 6033
rect 17879 6001 17905 6007
rect 20287 6033 20313 6039
rect 20287 6001 20313 6007
rect 20399 6033 20425 6039
rect 20399 6001 20425 6007
rect 21799 6033 21825 6039
rect 29583 6033 29609 6039
rect 27561 6007 27567 6033
rect 27593 6007 27599 6033
rect 28345 6007 28351 6033
rect 28377 6007 28383 6033
rect 29913 6007 29919 6033
rect 29945 6007 29951 6033
rect 30697 6007 30703 6033
rect 30729 6007 30735 6033
rect 21799 6001 21825 6007
rect 29583 6001 29609 6007
rect 14519 5977 14545 5983
rect 14519 5945 14545 5951
rect 14631 5977 14657 5983
rect 14631 5945 14657 5951
rect 21407 5977 21433 5983
rect 21407 5945 21433 5951
rect 21519 5977 21545 5983
rect 21519 5945 21545 5951
rect 29135 5977 29161 5983
rect 29135 5945 29161 5951
rect 29303 5977 29329 5983
rect 29303 5945 29329 5951
rect 336 5893 31864 5910
rect 336 5867 2233 5893
rect 2259 5867 2285 5893
rect 2311 5867 2337 5893
rect 2363 5867 12233 5893
rect 12259 5867 12285 5893
rect 12311 5867 12337 5893
rect 12363 5867 22233 5893
rect 22259 5867 22285 5893
rect 22311 5867 22337 5893
rect 22363 5867 31864 5893
rect 336 5850 31864 5867
rect 2311 5809 2337 5815
rect 2311 5777 2337 5783
rect 3879 5809 3905 5815
rect 3879 5777 3905 5783
rect 5447 5809 5473 5815
rect 5447 5777 5473 5783
rect 9311 5809 9337 5815
rect 9311 5777 9337 5783
rect 10151 5809 10177 5815
rect 10151 5777 10177 5783
rect 26503 5809 26529 5815
rect 26503 5777 26529 5783
rect 27287 5809 27313 5815
rect 27287 5777 27313 5783
rect 28239 5809 28265 5815
rect 28239 5777 28265 5783
rect 29023 5809 29049 5815
rect 29023 5777 29049 5783
rect 29807 5809 29833 5815
rect 29807 5777 29833 5783
rect 30591 5809 30617 5815
rect 30591 5777 30617 5783
rect 23087 5753 23113 5759
rect 10425 5727 10431 5753
rect 10457 5727 10463 5753
rect 23087 5721 23113 5727
rect 1191 5697 1217 5703
rect 14015 5697 14041 5703
rect 2585 5671 2591 5697
rect 2617 5671 2623 5697
rect 3257 5671 3263 5697
rect 3289 5671 3295 5697
rect 4153 5671 4159 5697
rect 4185 5671 4191 5697
rect 5721 5671 5727 5697
rect 5753 5671 5759 5697
rect 6505 5671 6511 5697
rect 6537 5671 6543 5697
rect 6729 5671 6735 5697
rect 6761 5671 6767 5697
rect 7457 5671 7463 5697
rect 7489 5671 7495 5697
rect 9025 5671 9031 5697
rect 9057 5671 9063 5697
rect 11153 5671 11159 5697
rect 11185 5671 11191 5697
rect 11993 5671 11999 5697
rect 12025 5671 12031 5697
rect 13617 5671 13623 5697
rect 13649 5671 13655 5697
rect 1191 5665 1217 5671
rect 14015 5665 14041 5671
rect 23367 5697 23393 5703
rect 26217 5671 26223 5697
rect 26249 5671 26255 5697
rect 27001 5671 27007 5697
rect 27033 5671 27039 5697
rect 28009 5671 28015 5697
rect 28041 5671 28047 5697
rect 28737 5671 28743 5697
rect 28769 5671 28775 5697
rect 29521 5671 29527 5697
rect 29553 5671 29559 5697
rect 30361 5671 30367 5697
rect 30393 5671 30399 5697
rect 31313 5671 31319 5697
rect 31345 5671 31351 5697
rect 23367 5665 23393 5671
rect 1359 5641 1385 5647
rect 7183 5641 7209 5647
rect 961 5615 967 5641
rect 993 5615 999 5641
rect 3033 5615 3039 5641
rect 3065 5615 3071 5641
rect 6169 5615 6175 5641
rect 6201 5615 6207 5641
rect 1359 5609 1385 5615
rect 7183 5609 7209 5615
rect 7967 5641 7993 5647
rect 7967 5609 7993 5615
rect 10711 5641 10737 5647
rect 13119 5641 13145 5647
rect 11545 5615 11551 5641
rect 11577 5615 11583 5641
rect 10711 5609 10737 5615
rect 13119 5609 13145 5615
rect 13847 5641 13873 5647
rect 23479 5641 23505 5647
rect 14233 5615 14239 5641
rect 14265 5615 14271 5641
rect 13847 5609 13873 5615
rect 23479 5609 23505 5615
rect 31095 5641 31121 5647
rect 31095 5609 31121 5615
rect 31487 5641 31513 5647
rect 31487 5609 31513 5615
rect 336 5501 31864 5518
rect 336 5475 1903 5501
rect 1929 5475 1955 5501
rect 1981 5475 2007 5501
rect 2033 5475 11903 5501
rect 11929 5475 11955 5501
rect 11981 5475 12007 5501
rect 12033 5475 21903 5501
rect 21929 5475 21955 5501
rect 21981 5475 22007 5501
rect 22033 5475 31864 5501
rect 336 5458 31864 5475
rect 4047 5417 4073 5423
rect 4047 5385 4073 5391
rect 4831 5417 4857 5423
rect 4831 5385 4857 5391
rect 5615 5417 5641 5423
rect 5615 5385 5641 5391
rect 7183 5417 7209 5423
rect 7183 5385 7209 5391
rect 8135 5417 8161 5423
rect 8135 5385 8161 5391
rect 8919 5417 8945 5423
rect 8919 5385 8945 5391
rect 9535 5417 9561 5423
rect 9535 5385 9561 5391
rect 11103 5417 11129 5423
rect 11103 5385 11129 5391
rect 11999 5417 12025 5423
rect 11999 5385 12025 5391
rect 10767 5361 10793 5367
rect 30759 5361 30785 5367
rect 3425 5335 3431 5361
rect 3457 5335 3463 5361
rect 27673 5335 27679 5361
rect 27705 5335 27711 5361
rect 28569 5335 28575 5361
rect 28601 5335 28607 5361
rect 29409 5335 29415 5361
rect 29441 5335 29447 5361
rect 10767 5329 10793 5335
rect 30759 5329 30785 5335
rect 3649 5279 3655 5305
rect 3681 5279 3687 5305
rect 4545 5279 4551 5305
rect 4577 5279 4583 5305
rect 5329 5279 5335 5305
rect 5361 5279 5367 5305
rect 8633 5279 8639 5305
rect 8665 5279 8671 5305
rect 9977 5279 9983 5305
rect 10009 5279 10015 5305
rect 11601 5279 11607 5305
rect 11633 5279 11639 5305
rect 21569 5279 21575 5305
rect 21601 5279 21607 5305
rect 29017 5279 29023 5305
rect 29049 5279 29055 5305
rect 30305 5279 30311 5305
rect 30337 5279 30343 5305
rect 31145 5279 31151 5305
rect 31177 5279 31183 5305
rect 6399 5249 6425 5255
rect 6113 5223 6119 5249
rect 6145 5223 6151 5249
rect 6399 5217 6425 5223
rect 6791 5249 6817 5255
rect 21799 5249 21825 5255
rect 7681 5223 7687 5249
rect 7713 5223 7719 5249
rect 7849 5223 7855 5249
rect 7881 5223 7887 5249
rect 12497 5223 12503 5249
rect 12529 5223 12535 5249
rect 28065 5223 28071 5249
rect 28097 5223 28103 5249
rect 28233 5223 28239 5249
rect 28265 5223 28271 5249
rect 31425 5223 31431 5249
rect 31457 5223 31463 5249
rect 6791 5217 6817 5223
rect 21799 5217 21825 5223
rect 6511 5193 6537 5199
rect 6511 5161 6537 5167
rect 10375 5193 10401 5199
rect 10375 5161 10401 5167
rect 10487 5193 10513 5199
rect 10487 5161 10513 5167
rect 21407 5193 21433 5199
rect 21407 5161 21433 5167
rect 336 5109 31864 5126
rect 336 5083 2233 5109
rect 2259 5083 2285 5109
rect 2311 5083 2337 5109
rect 2363 5083 12233 5109
rect 12259 5083 12285 5109
rect 12311 5083 12337 5109
rect 12363 5083 22233 5109
rect 22259 5083 22285 5109
rect 22311 5083 22337 5109
rect 22363 5083 31864 5109
rect 336 5066 31864 5083
rect 3767 5025 3793 5031
rect 3767 4993 3793 4999
rect 3879 5025 3905 5031
rect 3879 4993 3905 4999
rect 4159 4969 4185 4975
rect 30137 4943 30143 4969
rect 30169 4943 30175 4969
rect 30529 4943 30535 4969
rect 30561 4943 30567 4969
rect 4159 4937 4185 4943
rect 27959 4913 27985 4919
rect 5777 4887 5783 4913
rect 5809 4887 5815 4913
rect 7513 4887 7519 4913
rect 7545 4887 7551 4913
rect 28681 4887 28687 4913
rect 28713 4887 28719 4913
rect 29409 4887 29415 4913
rect 29441 4887 29447 4913
rect 30977 4887 30983 4913
rect 31009 4887 31015 4913
rect 27959 4881 27985 4887
rect 5279 4857 5305 4863
rect 5279 4825 5305 4831
rect 7071 4857 7097 4863
rect 7071 4825 7097 4831
rect 27735 4857 27761 4863
rect 27735 4825 27761 4831
rect 28239 4857 28265 4863
rect 28239 4825 28265 4831
rect 28407 4857 28433 4863
rect 29863 4857 29889 4863
rect 28961 4831 28967 4857
rect 28993 4831 28999 4857
rect 31369 4831 31375 4857
rect 31401 4831 31407 4857
rect 28407 4825 28433 4831
rect 29863 4825 29889 4831
rect 336 4717 31864 4734
rect 336 4691 1903 4717
rect 1929 4691 1955 4717
rect 1981 4691 2007 4717
rect 2033 4691 11903 4717
rect 11929 4691 11955 4717
rect 11981 4691 12007 4717
rect 12033 4691 21903 4717
rect 21929 4691 21955 4717
rect 21981 4691 22007 4717
rect 22033 4691 31864 4717
rect 336 4674 31864 4691
rect 29359 4633 29385 4639
rect 29359 4601 29385 4607
rect 30759 4633 30785 4639
rect 30759 4601 30785 4607
rect 2199 4577 2225 4583
rect 1409 4551 1415 4577
rect 1441 4551 1447 4577
rect 2199 4545 2225 4551
rect 8919 4577 8945 4583
rect 8919 4545 8945 4551
rect 10711 4577 10737 4583
rect 10711 4545 10737 4551
rect 11103 4577 11129 4583
rect 11103 4545 11129 4551
rect 14911 4577 14937 4583
rect 14911 4545 14937 4551
rect 20231 4577 20257 4583
rect 20231 4545 20257 4551
rect 20623 4577 20649 4583
rect 20623 4545 20649 4551
rect 23703 4577 23729 4583
rect 23703 4545 23729 4551
rect 24095 4577 24121 4583
rect 28345 4551 28351 4577
rect 28377 4551 28383 4577
rect 28793 4551 28799 4577
rect 28825 4551 28831 4577
rect 24095 4545 24121 4551
rect 2479 4521 2505 4527
rect 2479 4489 2505 4495
rect 10823 4521 10849 4527
rect 10823 4489 10849 4495
rect 14519 4521 14545 4527
rect 14519 4489 14545 4495
rect 14799 4521 14825 4527
rect 14799 4489 14825 4495
rect 20511 4521 20537 4527
rect 20511 4489 20537 4495
rect 23815 4521 23841 4527
rect 23815 4489 23841 4495
rect 26223 4521 26249 4527
rect 26223 4489 26249 4495
rect 26391 4521 26417 4527
rect 29577 4495 29583 4521
rect 29609 4495 29615 4521
rect 31089 4495 31095 4521
rect 31121 4495 31127 4521
rect 26391 4489 26417 4495
rect 2759 4465 2785 4471
rect 2759 4433 2785 4439
rect 26671 4465 26697 4471
rect 30249 4439 30255 4465
rect 30281 4439 30287 4465
rect 31425 4439 31431 4465
rect 31457 4439 31463 4465
rect 26671 4433 26697 4439
rect 1639 4409 1665 4415
rect 1639 4377 1665 4383
rect 1751 4409 1777 4415
rect 1751 4377 1777 4383
rect 8527 4409 8553 4415
rect 8527 4377 8553 4383
rect 8639 4409 8665 4415
rect 8639 4377 8665 4383
rect 27959 4409 27985 4415
rect 27959 4377 27985 4383
rect 28127 4409 28153 4415
rect 28127 4377 28153 4383
rect 28575 4409 28601 4415
rect 28575 4377 28601 4383
rect 336 4325 31864 4342
rect 336 4299 2233 4325
rect 2259 4299 2285 4325
rect 2311 4299 2337 4325
rect 2363 4299 12233 4325
rect 12259 4299 12285 4325
rect 12311 4299 12337 4325
rect 12363 4299 22233 4325
rect 22259 4299 22285 4325
rect 22311 4299 22337 4325
rect 22363 4299 31864 4325
rect 336 4282 31864 4299
rect 2255 4185 2281 4191
rect 2255 4153 2281 4159
rect 2367 4185 2393 4191
rect 2367 4153 2393 4159
rect 21967 4185 21993 4191
rect 21967 4153 21993 4159
rect 22079 4185 22105 4191
rect 22079 4153 22105 4159
rect 28239 4185 28265 4191
rect 30137 4159 30143 4185
rect 30169 4159 30175 4185
rect 30529 4159 30535 4185
rect 30561 4159 30567 4185
rect 28239 4153 28265 4159
rect 6231 4129 6257 4135
rect 6231 4097 6257 4103
rect 27959 4129 27985 4135
rect 27959 4097 27985 4103
rect 28463 4129 28489 4135
rect 28463 4097 28489 4103
rect 28743 4129 28769 4135
rect 28743 4097 28769 4103
rect 28911 4129 28937 4135
rect 28911 4097 28937 4103
rect 29191 4129 29217 4135
rect 29353 4103 29359 4129
rect 29385 4103 29391 4129
rect 30921 4103 30927 4129
rect 30953 4103 30959 4129
rect 29191 4097 29217 4103
rect 2647 4073 2673 4079
rect 2647 4041 2673 4047
rect 6063 4073 6089 4079
rect 6063 4041 6089 4047
rect 6511 4073 6537 4079
rect 27735 4073 27761 4079
rect 21737 4047 21743 4073
rect 21769 4047 21775 4073
rect 6511 4041 6537 4047
rect 27735 4041 27761 4047
rect 29863 4073 29889 4079
rect 29863 4041 29889 4047
rect 31431 4017 31457 4023
rect 31431 3985 31457 3991
rect 336 3933 31864 3950
rect 336 3907 1903 3933
rect 1929 3907 1955 3933
rect 1981 3907 2007 3933
rect 2033 3907 11903 3933
rect 11929 3907 11955 3933
rect 11981 3907 12007 3933
rect 12033 3907 21903 3933
rect 21929 3907 21955 3933
rect 21981 3907 22007 3933
rect 22033 3907 31864 3933
rect 336 3890 31864 3907
rect 31543 3849 31569 3855
rect 31543 3817 31569 3823
rect 17263 3793 17289 3799
rect 21239 3793 21265 3799
rect 7401 3767 7407 3793
rect 7433 3767 7439 3793
rect 17649 3767 17655 3793
rect 17681 3767 17687 3793
rect 17263 3761 17289 3767
rect 21239 3761 21265 3767
rect 28351 3793 28377 3799
rect 30759 3793 30785 3799
rect 29129 3767 29135 3793
rect 29161 3767 29167 3793
rect 29577 3767 29583 3793
rect 29609 3767 29615 3793
rect 28351 3761 28377 3767
rect 30759 3761 30785 3767
rect 17431 3737 17457 3743
rect 17431 3705 17457 3711
rect 21127 3737 21153 3743
rect 21127 3705 21153 3711
rect 28799 3737 28825 3743
rect 29409 3711 29415 3737
rect 29441 3711 29447 3737
rect 31145 3711 31151 3737
rect 31177 3711 31183 3737
rect 28799 3705 28825 3711
rect 7743 3681 7769 3687
rect 7743 3649 7769 3655
rect 20847 3681 20873 3687
rect 30249 3655 30255 3681
rect 30281 3655 30287 3681
rect 20847 3649 20873 3655
rect 7631 3625 7657 3631
rect 7631 3593 7657 3599
rect 28631 3625 28657 3631
rect 28631 3593 28657 3599
rect 28911 3625 28937 3631
rect 28911 3593 28937 3599
rect 336 3541 31864 3558
rect 336 3515 2233 3541
rect 2259 3515 2285 3541
rect 2311 3515 2337 3541
rect 2363 3515 12233 3541
rect 12259 3515 12285 3541
rect 12311 3515 12337 3541
rect 12363 3515 22233 3541
rect 22259 3515 22285 3541
rect 22311 3515 22337 3541
rect 22363 3515 31864 3541
rect 336 3498 31864 3515
rect 30921 3375 30927 3401
rect 30953 3375 30959 3401
rect 8751 3345 8777 3351
rect 8751 3313 8777 3319
rect 9031 3345 9057 3351
rect 9031 3313 9057 3319
rect 15359 3345 15385 3351
rect 15359 3313 15385 3319
rect 18439 3345 18465 3351
rect 18439 3313 18465 3319
rect 18551 3345 18577 3351
rect 18551 3313 18577 3319
rect 23479 3345 23505 3351
rect 23479 3313 23505 3319
rect 23759 3345 23785 3351
rect 23759 3313 23785 3319
rect 25215 3345 25241 3351
rect 25215 3313 25241 3319
rect 25495 3345 25521 3351
rect 25495 3313 25521 3319
rect 29135 3345 29161 3351
rect 29135 3313 29161 3319
rect 29247 3345 29273 3351
rect 29247 3313 29273 3319
rect 29695 3345 29721 3351
rect 29695 3313 29721 3319
rect 29975 3345 30001 3351
rect 30137 3319 30143 3345
rect 30169 3319 30175 3345
rect 29975 3313 30001 3319
rect 9199 3289 9225 3295
rect 15527 3289 15553 3295
rect 15129 3263 15135 3289
rect 15161 3263 15167 3289
rect 9199 3257 9225 3263
rect 15527 3257 15553 3263
rect 18159 3289 18185 3295
rect 18159 3257 18185 3263
rect 23367 3289 23393 3295
rect 23367 3257 23393 3263
rect 25047 3289 25073 3295
rect 25047 3257 25073 3263
rect 28911 3289 28937 3295
rect 28911 3257 28937 3263
rect 29023 3289 29049 3295
rect 31431 3289 31457 3295
rect 29465 3263 29471 3289
rect 29497 3263 29503 3289
rect 29023 3257 29049 3263
rect 31431 3257 31457 3263
rect 30647 3233 30673 3239
rect 30647 3201 30673 3207
rect 336 3149 31864 3166
rect 336 3123 1903 3149
rect 1929 3123 1955 3149
rect 1981 3123 2007 3149
rect 2033 3123 11903 3149
rect 11929 3123 11955 3149
rect 11981 3123 12007 3149
rect 12033 3123 21903 3149
rect 21929 3123 21955 3149
rect 21981 3123 22007 3149
rect 22033 3123 31864 3149
rect 336 3106 31864 3123
rect 30759 3065 30785 3071
rect 30759 3033 30785 3039
rect 31543 3065 31569 3071
rect 31543 3033 31569 3039
rect 1359 3009 1385 3015
rect 4439 3009 4465 3015
rect 4097 2983 4103 3009
rect 4129 2983 4135 3009
rect 1359 2977 1385 2983
rect 4439 2977 4465 2983
rect 13287 3009 13313 3015
rect 13287 2977 13313 2983
rect 13679 3009 13705 3015
rect 13679 2977 13705 2983
rect 14799 3009 14825 3015
rect 14799 2977 14825 2983
rect 21295 3009 21321 3015
rect 21295 2977 21321 2983
rect 28967 3009 28993 3015
rect 28967 2977 28993 2983
rect 29639 3009 29665 3015
rect 29639 2977 29665 2983
rect 1247 2953 1273 2959
rect 1247 2921 1273 2927
rect 4327 2953 4353 2959
rect 4327 2921 4353 2927
rect 13567 2953 13593 2959
rect 30249 2927 30255 2953
rect 30281 2927 30287 2953
rect 31089 2927 31095 2953
rect 31121 2927 31127 2953
rect 13567 2921 13593 2927
rect 967 2897 993 2903
rect 967 2865 993 2871
rect 15079 2897 15105 2903
rect 15079 2865 15105 2871
rect 15191 2897 15217 2903
rect 15191 2865 15217 2871
rect 22359 2897 22385 2903
rect 22359 2865 22385 2871
rect 21855 2841 21881 2847
rect 21855 2809 21881 2815
rect 22079 2841 22105 2847
rect 22079 2809 22105 2815
rect 28519 2841 28545 2847
rect 28519 2809 28545 2815
rect 28687 2841 28713 2847
rect 28687 2809 28713 2815
rect 29191 2841 29217 2847
rect 29191 2809 29217 2815
rect 29359 2841 29385 2847
rect 29359 2809 29385 2815
rect 336 2757 31864 2774
rect 336 2731 2233 2757
rect 2259 2731 2285 2757
rect 2311 2731 2337 2757
rect 2363 2731 12233 2757
rect 12259 2731 12285 2757
rect 12311 2731 12337 2757
rect 12363 2731 22233 2757
rect 22259 2731 22285 2757
rect 22311 2731 22337 2757
rect 22363 2731 31864 2757
rect 336 2714 31864 2731
rect 8639 2673 8665 2679
rect 8639 2641 8665 2647
rect 8807 2673 8833 2679
rect 8807 2641 8833 2647
rect 9647 2673 9673 2679
rect 9647 2641 9673 2647
rect 9815 2673 9841 2679
rect 9815 2641 9841 2647
rect 10935 2673 10961 2679
rect 10935 2641 10961 2647
rect 11103 2673 11129 2679
rect 11103 2641 11129 2647
rect 12559 2673 12585 2679
rect 12559 2641 12585 2647
rect 12727 2673 12753 2679
rect 12727 2641 12753 2647
rect 14799 2673 14825 2679
rect 14799 2641 14825 2647
rect 14911 2673 14937 2679
rect 14911 2641 14937 2647
rect 19895 2673 19921 2679
rect 19895 2641 19921 2647
rect 20175 2673 20201 2679
rect 20175 2641 20201 2647
rect 21183 2673 21209 2679
rect 21183 2641 21209 2647
rect 21351 2673 21377 2679
rect 21351 2641 21377 2647
rect 21463 2673 21489 2679
rect 21463 2641 21489 2647
rect 967 2617 993 2623
rect 967 2585 993 2591
rect 9367 2617 9393 2623
rect 9367 2585 9393 2591
rect 10655 2617 10681 2623
rect 10655 2585 10681 2591
rect 12279 2617 12305 2623
rect 12279 2585 12305 2591
rect 14519 2617 14545 2623
rect 14519 2585 14545 2591
rect 20455 2617 20481 2623
rect 20455 2585 20481 2591
rect 20903 2617 20929 2623
rect 20903 2585 20929 2591
rect 25439 2617 25465 2623
rect 25439 2585 25465 2591
rect 29191 2617 29217 2623
rect 30137 2591 30143 2617
rect 30169 2591 30175 2617
rect 30529 2591 30535 2617
rect 30561 2591 30567 2617
rect 31313 2591 31319 2617
rect 31345 2591 31351 2617
rect 29191 2585 29217 2591
rect 1247 2561 1273 2567
rect 1247 2529 1273 2535
rect 1415 2561 1441 2567
rect 1415 2529 1441 2535
rect 21743 2561 21769 2567
rect 21743 2529 21769 2535
rect 24991 2561 25017 2567
rect 24991 2529 25017 2535
rect 25159 2561 25185 2567
rect 25159 2529 25185 2535
rect 28183 2561 28209 2567
rect 28183 2529 28209 2535
rect 28351 2561 28377 2567
rect 28351 2529 28377 2535
rect 28631 2561 28657 2567
rect 28631 2529 28657 2535
rect 28743 2561 28769 2567
rect 28743 2529 28769 2535
rect 28911 2561 28937 2567
rect 28911 2529 28937 2535
rect 29583 2561 29609 2567
rect 29583 2529 29609 2535
rect 29695 2561 29721 2567
rect 29695 2529 29721 2535
rect 29975 2561 30001 2567
rect 30921 2535 30927 2561
rect 30953 2535 30959 2561
rect 29975 2529 30001 2535
rect 8409 2479 8415 2505
rect 8441 2479 8447 2505
rect 336 2365 31864 2382
rect 336 2339 1903 2365
rect 1929 2339 1955 2365
rect 1981 2339 2007 2365
rect 2033 2339 11903 2365
rect 11929 2339 11955 2365
rect 11981 2339 12007 2365
rect 12033 2339 21903 2365
rect 21929 2339 21955 2365
rect 21981 2339 22007 2365
rect 22033 2339 31864 2365
rect 336 2322 31864 2339
rect 31543 2281 31569 2287
rect 31543 2249 31569 2255
rect 911 2225 937 2231
rect 911 2193 937 2199
rect 8247 2225 8273 2231
rect 8247 2193 8273 2199
rect 21015 2225 21041 2231
rect 21015 2193 21041 2199
rect 21407 2225 21433 2231
rect 21407 2193 21433 2199
rect 24655 2225 24681 2231
rect 27841 2199 27847 2225
rect 27873 2199 27879 2225
rect 24655 2193 24681 2199
rect 21295 2169 21321 2175
rect 21295 2137 21321 2143
rect 24543 2169 24569 2175
rect 30305 2143 30311 2169
rect 30337 2143 30343 2169
rect 31145 2143 31151 2169
rect 31177 2143 31183 2169
rect 24543 2137 24569 2143
rect 24263 2113 24289 2119
rect 30641 2087 30647 2113
rect 30673 2087 30679 2113
rect 24263 2081 24289 2087
rect 1191 2057 1217 2063
rect 1191 2025 1217 2031
rect 1303 2057 1329 2063
rect 1303 2025 1329 2031
rect 8527 2057 8553 2063
rect 8527 2025 8553 2031
rect 8639 2057 8665 2063
rect 8639 2025 8665 2031
rect 28071 2057 28097 2063
rect 28071 2025 28097 2031
rect 28239 2057 28265 2063
rect 28239 2025 28265 2031
rect 336 1973 31864 1990
rect 336 1947 2233 1973
rect 2259 1947 2285 1973
rect 2311 1947 2337 1973
rect 2363 1947 12233 1973
rect 12259 1947 12285 1973
rect 12311 1947 12337 1973
rect 12363 1947 22233 1973
rect 22259 1947 22285 1973
rect 22311 1947 22337 1973
rect 22363 1947 31864 1973
rect 336 1930 31864 1947
rect 2479 1889 2505 1895
rect 2479 1857 2505 1863
rect 2591 1889 2617 1895
rect 2591 1857 2617 1863
rect 8639 1889 8665 1895
rect 8639 1857 8665 1863
rect 8807 1889 8833 1895
rect 8807 1857 8833 1863
rect 12279 1889 12305 1895
rect 12279 1857 12305 1863
rect 20399 1889 20425 1895
rect 20399 1857 20425 1863
rect 20511 1889 20537 1895
rect 20511 1857 20537 1863
rect 23535 1889 23561 1895
rect 23535 1857 23561 1863
rect 23703 1889 23729 1895
rect 23703 1857 23729 1863
rect 25271 1889 25297 1895
rect 25271 1857 25297 1863
rect 25383 1889 25409 1895
rect 25383 1857 25409 1863
rect 29527 1889 29553 1895
rect 29527 1857 29553 1863
rect 29695 1889 29721 1895
rect 29695 1857 29721 1863
rect 2871 1833 2897 1839
rect 2871 1801 2897 1807
rect 8359 1833 8385 1839
rect 8359 1801 8385 1807
rect 11999 1833 12025 1839
rect 11999 1801 12025 1807
rect 22023 1833 22049 1839
rect 22023 1801 22049 1807
rect 22191 1833 22217 1839
rect 22191 1801 22217 1807
rect 22471 1833 22497 1839
rect 22471 1801 22497 1807
rect 23255 1833 23281 1839
rect 23255 1801 23281 1807
rect 24991 1833 25017 1839
rect 30921 1807 30927 1833
rect 30953 1807 30959 1833
rect 24991 1801 25017 1807
rect 1303 1777 1329 1783
rect 1303 1745 1329 1751
rect 1471 1777 1497 1783
rect 1471 1745 1497 1751
rect 29975 1777 30001 1783
rect 30137 1751 30143 1777
rect 30169 1751 30175 1777
rect 29975 1745 30001 1751
rect 29247 1721 29273 1727
rect 1073 1695 1079 1721
rect 1105 1695 1111 1721
rect 11769 1695 11775 1721
rect 11801 1695 11807 1721
rect 20169 1695 20175 1721
rect 20201 1695 20207 1721
rect 29247 1689 29273 1695
rect 30647 1721 30673 1727
rect 30647 1689 30673 1695
rect 31431 1721 31457 1727
rect 31431 1689 31457 1695
rect 336 1581 31864 1598
rect 336 1555 1903 1581
rect 1929 1555 1955 1581
rect 1981 1555 2007 1581
rect 2033 1555 11903 1581
rect 11929 1555 11955 1581
rect 11981 1555 12007 1581
rect 12033 1555 21903 1581
rect 21929 1555 21955 1581
rect 21981 1555 22007 1581
rect 22033 1555 31864 1581
rect 336 1538 31864 1555
rect 31543 1497 31569 1503
rect 31543 1465 31569 1471
rect 26049 1415 26055 1441
rect 26081 1415 26087 1441
rect 29639 1385 29665 1391
rect 29409 1359 29415 1385
rect 29441 1359 29447 1385
rect 31089 1359 31095 1385
rect 31121 1359 31127 1385
rect 29639 1353 29665 1359
rect 29191 1329 29217 1335
rect 30249 1303 30255 1329
rect 30281 1303 30287 1329
rect 30641 1303 30647 1329
rect 30673 1303 30679 1329
rect 29191 1297 29217 1303
rect 26279 1273 26305 1279
rect 26279 1241 26305 1247
rect 26447 1273 26473 1279
rect 26447 1241 26473 1247
rect 28799 1273 28825 1279
rect 28799 1241 28825 1247
rect 28911 1273 28937 1279
rect 28911 1241 28937 1247
rect 336 1189 31864 1206
rect 336 1163 2233 1189
rect 2259 1163 2285 1189
rect 2311 1163 2337 1189
rect 2363 1163 12233 1189
rect 12259 1163 12285 1189
rect 12311 1163 12337 1189
rect 12363 1163 22233 1189
rect 22259 1163 22285 1189
rect 22311 1163 22337 1189
rect 22363 1163 31864 1189
rect 336 1146 31864 1163
rect 1247 1105 1273 1111
rect 1247 1073 1273 1079
rect 1415 1105 1441 1111
rect 1415 1073 1441 1079
rect 7631 1105 7657 1111
rect 7631 1073 7657 1079
rect 8079 1105 8105 1111
rect 8079 1073 8105 1079
rect 8359 1105 8385 1111
rect 8359 1073 8385 1079
rect 11439 1105 11465 1111
rect 11439 1073 11465 1079
rect 11607 1105 11633 1111
rect 11607 1073 11633 1079
rect 15079 1105 15105 1111
rect 15079 1073 15105 1079
rect 15247 1105 15273 1111
rect 18439 1105 18465 1111
rect 15409 1079 15415 1105
rect 15441 1079 15447 1105
rect 15247 1073 15273 1079
rect 18439 1073 18465 1079
rect 18607 1105 18633 1111
rect 18607 1073 18633 1079
rect 19055 1105 19081 1111
rect 19055 1073 19081 1079
rect 19223 1105 19249 1111
rect 19223 1073 19249 1079
rect 19727 1105 19753 1111
rect 19727 1073 19753 1079
rect 19895 1105 19921 1111
rect 19895 1073 19921 1079
rect 20903 1105 20929 1111
rect 20903 1073 20929 1079
rect 21351 1105 21377 1111
rect 21351 1073 21377 1079
rect 22919 1105 22945 1111
rect 22919 1073 22945 1079
rect 23087 1105 23113 1111
rect 23087 1073 23113 1079
rect 6119 1049 6145 1055
rect 6119 1017 6145 1023
rect 6231 1049 6257 1055
rect 6231 1017 6257 1023
rect 6511 1049 6537 1055
rect 6511 1017 6537 1023
rect 7351 1049 7377 1055
rect 7351 1017 7377 1023
rect 7799 1049 7825 1055
rect 7799 1017 7825 1023
rect 11159 1049 11185 1055
rect 11159 1017 11185 1023
rect 16199 1049 16225 1055
rect 16199 1017 16225 1023
rect 16647 1049 16673 1055
rect 16647 1017 16673 1023
rect 17655 1049 17681 1055
rect 17655 1017 17681 1023
rect 18159 1049 18185 1055
rect 18159 1017 18185 1023
rect 20623 1049 20649 1055
rect 20623 1017 20649 1023
rect 21071 1049 21097 1055
rect 21071 1017 21097 1023
rect 21519 1049 21545 1055
rect 21519 1017 21545 1023
rect 24319 1049 24345 1055
rect 24319 1017 24345 1023
rect 24879 1049 24905 1055
rect 24879 1017 24905 1023
rect 25439 1049 25465 1055
rect 25439 1017 25465 1023
rect 28799 1049 28825 1055
rect 28799 1017 28825 1023
rect 29247 1049 29273 1055
rect 30137 1023 30143 1049
rect 30169 1023 30175 1049
rect 29247 1017 29273 1023
rect 4383 993 4409 999
rect 4383 961 4409 967
rect 4551 993 4577 999
rect 5279 993 5305 999
rect 17935 993 17961 999
rect 5049 967 5055 993
rect 5081 967 5087 993
rect 16417 967 16423 993
rect 16449 967 16455 993
rect 4551 961 4577 967
rect 5279 961 5305 967
rect 17935 961 17961 967
rect 19447 993 19473 999
rect 19447 961 19473 967
rect 21799 993 21825 999
rect 21799 961 21825 967
rect 21967 993 21993 999
rect 21967 961 21993 967
rect 24039 993 24065 999
rect 24039 961 24065 967
rect 24599 993 24625 999
rect 24599 961 24625 967
rect 25159 993 25185 999
rect 25159 961 25185 967
rect 28519 993 28545 999
rect 28519 961 28545 967
rect 28967 993 28993 999
rect 28967 961 28993 967
rect 29695 993 29721 999
rect 29695 961 29721 967
rect 29975 993 30001 999
rect 30921 967 30927 993
rect 30953 967 30959 993
rect 29975 961 30001 967
rect 4831 937 4857 943
rect 1017 911 1023 937
rect 1049 911 1055 937
rect 4831 905 4857 911
rect 18775 937 18801 943
rect 23759 937 23785 943
rect 22689 911 22695 937
rect 22721 911 22727 937
rect 18775 905 18801 911
rect 23759 905 23785 911
rect 24431 937 24457 943
rect 24431 905 24457 911
rect 24991 937 25017 943
rect 24991 905 25017 911
rect 28351 937 28377 943
rect 28351 905 28377 911
rect 29583 937 29609 943
rect 29583 905 29609 911
rect 31431 937 31457 943
rect 31431 905 31457 911
rect 30647 881 30673 887
rect 30647 849 30673 855
rect 336 797 31864 814
rect 336 771 1903 797
rect 1929 771 1955 797
rect 1981 771 2007 797
rect 2033 771 11903 797
rect 11929 771 11955 797
rect 11981 771 12007 797
rect 12033 771 21903 797
rect 21929 771 21955 797
rect 21981 771 22007 797
rect 22033 771 31864 797
rect 336 754 31864 771
rect 31543 713 31569 719
rect 31543 681 31569 687
rect 5279 657 5305 663
rect 5279 625 5305 631
rect 7799 657 7825 663
rect 7799 625 7825 631
rect 18103 657 18129 663
rect 18103 625 18129 631
rect 21071 657 21097 663
rect 21071 625 21097 631
rect 21519 657 21545 663
rect 21519 625 21545 631
rect 28855 657 28881 663
rect 28855 625 28881 631
rect 29807 657 29833 663
rect 29807 625 29833 631
rect 30591 657 30617 663
rect 30591 625 30617 631
rect 29297 575 29303 601
rect 29329 575 29335 601
rect 30081 575 30087 601
rect 30113 575 30119 601
rect 31089 575 31095 601
rect 31121 575 31127 601
rect 911 545 937 551
rect 911 513 937 519
rect 4999 545 5025 551
rect 4999 513 5025 519
rect 1191 489 1217 495
rect 1191 457 1217 463
rect 1303 489 1329 495
rect 1303 457 1329 463
rect 4775 489 4801 495
rect 4775 457 4801 463
rect 4831 489 4857 495
rect 4831 457 4857 463
rect 336 405 31864 422
rect 336 379 2233 405
rect 2259 379 2285 405
rect 2311 379 2337 405
rect 2363 379 12233 405
rect 12259 379 12285 405
rect 12311 379 12337 405
rect 12363 379 22233 405
rect 22259 379 22285 405
rect 22311 379 22337 405
rect 22363 379 31864 405
rect 336 362 31864 379
<< via1 >>
rect 2233 6651 2259 6677
rect 2285 6651 2311 6677
rect 2337 6651 2363 6677
rect 12233 6651 12259 6677
rect 12285 6651 12311 6677
rect 12337 6651 12363 6677
rect 22233 6651 22259 6677
rect 22285 6651 22311 6677
rect 22337 6651 22363 6677
rect 1863 6567 1889 6593
rect 2983 6567 3009 6593
rect 3767 6567 3793 6593
rect 4887 6567 4913 6593
rect 5671 6567 5697 6593
rect 8695 6567 8721 6593
rect 9479 6567 9505 6593
rect 10599 6567 10625 6593
rect 11383 6567 11409 6593
rect 12503 6567 12529 6593
rect 13287 6567 13313 6593
rect 25439 6567 25465 6593
rect 26055 6567 26081 6593
rect 27455 6567 27481 6593
rect 28239 6567 28265 6593
rect 31263 6567 31289 6593
rect 7463 6511 7489 6537
rect 30255 6511 30281 6537
rect 855 6455 881 6481
rect 2143 6455 2169 6481
rect 3207 6455 3233 6481
rect 3991 6455 4017 6481
rect 5167 6455 5193 6481
rect 5951 6455 5977 6481
rect 6455 6455 6481 6481
rect 7855 6455 7881 6481
rect 8975 6455 9001 6481
rect 9759 6455 9785 6481
rect 10879 6455 10905 6481
rect 11663 6455 11689 6481
rect 12727 6455 12753 6481
rect 13567 6455 13593 6481
rect 14463 6455 14489 6481
rect 25607 6455 25633 6481
rect 25775 6455 25801 6481
rect 27175 6455 27201 6481
rect 27959 6455 27985 6481
rect 29079 6455 29105 6481
rect 29863 6455 29889 6481
rect 30983 6455 31009 6481
rect 1247 6399 1273 6425
rect 6959 6399 6985 6425
rect 13959 6399 13985 6425
rect 29415 6399 29441 6425
rect 1903 6259 1929 6285
rect 1955 6259 1981 6285
rect 2007 6259 2033 6285
rect 11903 6259 11929 6285
rect 11955 6259 11981 6285
rect 12007 6259 12033 6285
rect 21903 6259 21929 6285
rect 21955 6259 21981 6285
rect 22007 6259 22033 6285
rect 3487 6175 3513 6201
rect 4271 6175 4297 6201
rect 5055 6175 5081 6201
rect 5839 6175 5865 6201
rect 8191 6175 8217 6201
rect 8975 6175 9001 6201
rect 9927 6175 9953 6201
rect 11215 6175 11241 6201
rect 11999 6175 12025 6201
rect 12559 6175 12585 6201
rect 26279 6175 26305 6201
rect 27063 6175 27089 6201
rect 27847 6175 27873 6201
rect 28631 6175 28657 6201
rect 1807 6119 1833 6145
rect 7519 6119 7545 6145
rect 13455 6119 13481 6145
rect 14911 6119 14937 6145
rect 15191 6119 15217 6145
rect 15583 6119 15609 6145
rect 17487 6119 17513 6145
rect 30311 6119 30337 6145
rect 31095 6119 31121 6145
rect 6063 6063 6089 6089
rect 9199 6063 9225 6089
rect 9423 6063 9449 6089
rect 13735 6063 13761 6089
rect 15471 6063 15497 6089
rect 17599 6063 17625 6089
rect 20679 6063 20705 6089
rect 26055 6063 26081 6089
rect 26783 6063 26809 6089
rect 2199 6007 2225 6033
rect 3767 6007 3793 6033
rect 4551 6007 4577 6033
rect 5335 6007 5361 6033
rect 7071 6007 7097 6033
rect 8471 6007 8497 6033
rect 11495 6007 11521 6033
rect 12279 6007 12305 6033
rect 13063 6007 13089 6033
rect 17879 6007 17905 6033
rect 20287 6007 20313 6033
rect 20399 6007 20425 6033
rect 21799 6007 21825 6033
rect 27567 6007 27593 6033
rect 28351 6007 28377 6033
rect 29583 6007 29609 6033
rect 29919 6007 29945 6033
rect 30703 6007 30729 6033
rect 14519 5951 14545 5977
rect 14631 5951 14657 5977
rect 21407 5951 21433 5977
rect 21519 5951 21545 5977
rect 29135 5951 29161 5977
rect 29303 5951 29329 5977
rect 2233 5867 2259 5893
rect 2285 5867 2311 5893
rect 2337 5867 2363 5893
rect 12233 5867 12259 5893
rect 12285 5867 12311 5893
rect 12337 5867 12363 5893
rect 22233 5867 22259 5893
rect 22285 5867 22311 5893
rect 22337 5867 22363 5893
rect 2311 5783 2337 5809
rect 3879 5783 3905 5809
rect 5447 5783 5473 5809
rect 9311 5783 9337 5809
rect 10151 5783 10177 5809
rect 26503 5783 26529 5809
rect 27287 5783 27313 5809
rect 28239 5783 28265 5809
rect 29023 5783 29049 5809
rect 29807 5783 29833 5809
rect 30591 5783 30617 5809
rect 10431 5727 10457 5753
rect 23087 5727 23113 5753
rect 1191 5671 1217 5697
rect 2591 5671 2617 5697
rect 3263 5671 3289 5697
rect 4159 5671 4185 5697
rect 5727 5671 5753 5697
rect 6511 5671 6537 5697
rect 6735 5671 6761 5697
rect 7463 5671 7489 5697
rect 9031 5671 9057 5697
rect 11159 5671 11185 5697
rect 11999 5671 12025 5697
rect 13623 5671 13649 5697
rect 14015 5671 14041 5697
rect 23367 5671 23393 5697
rect 26223 5671 26249 5697
rect 27007 5671 27033 5697
rect 28015 5671 28041 5697
rect 28743 5671 28769 5697
rect 29527 5671 29553 5697
rect 30367 5671 30393 5697
rect 31319 5671 31345 5697
rect 967 5615 993 5641
rect 1359 5615 1385 5641
rect 3039 5615 3065 5641
rect 6175 5615 6201 5641
rect 7183 5615 7209 5641
rect 7967 5615 7993 5641
rect 10711 5615 10737 5641
rect 11551 5615 11577 5641
rect 13119 5615 13145 5641
rect 13847 5615 13873 5641
rect 14239 5615 14265 5641
rect 23479 5615 23505 5641
rect 31095 5615 31121 5641
rect 31487 5615 31513 5641
rect 1903 5475 1929 5501
rect 1955 5475 1981 5501
rect 2007 5475 2033 5501
rect 11903 5475 11929 5501
rect 11955 5475 11981 5501
rect 12007 5475 12033 5501
rect 21903 5475 21929 5501
rect 21955 5475 21981 5501
rect 22007 5475 22033 5501
rect 4047 5391 4073 5417
rect 4831 5391 4857 5417
rect 5615 5391 5641 5417
rect 7183 5391 7209 5417
rect 8135 5391 8161 5417
rect 8919 5391 8945 5417
rect 9535 5391 9561 5417
rect 11103 5391 11129 5417
rect 11999 5391 12025 5417
rect 3431 5335 3457 5361
rect 10767 5335 10793 5361
rect 27679 5335 27705 5361
rect 28575 5335 28601 5361
rect 29415 5335 29441 5361
rect 30759 5335 30785 5361
rect 3655 5279 3681 5305
rect 4551 5279 4577 5305
rect 5335 5279 5361 5305
rect 8639 5279 8665 5305
rect 9983 5279 10009 5305
rect 11607 5279 11633 5305
rect 21575 5279 21601 5305
rect 29023 5279 29049 5305
rect 30311 5279 30337 5305
rect 31151 5279 31177 5305
rect 6119 5223 6145 5249
rect 6399 5223 6425 5249
rect 6791 5223 6817 5249
rect 7687 5223 7713 5249
rect 7855 5223 7881 5249
rect 12503 5223 12529 5249
rect 21799 5223 21825 5249
rect 28071 5223 28097 5249
rect 28239 5223 28265 5249
rect 31431 5223 31457 5249
rect 6511 5167 6537 5193
rect 10375 5167 10401 5193
rect 10487 5167 10513 5193
rect 21407 5167 21433 5193
rect 2233 5083 2259 5109
rect 2285 5083 2311 5109
rect 2337 5083 2363 5109
rect 12233 5083 12259 5109
rect 12285 5083 12311 5109
rect 12337 5083 12363 5109
rect 22233 5083 22259 5109
rect 22285 5083 22311 5109
rect 22337 5083 22363 5109
rect 3767 4999 3793 5025
rect 3879 4999 3905 5025
rect 4159 4943 4185 4969
rect 30143 4943 30169 4969
rect 30535 4943 30561 4969
rect 5783 4887 5809 4913
rect 7519 4887 7545 4913
rect 27959 4887 27985 4913
rect 28687 4887 28713 4913
rect 29415 4887 29441 4913
rect 30983 4887 31009 4913
rect 5279 4831 5305 4857
rect 7071 4831 7097 4857
rect 27735 4831 27761 4857
rect 28239 4831 28265 4857
rect 28407 4831 28433 4857
rect 28967 4831 28993 4857
rect 29863 4831 29889 4857
rect 31375 4831 31401 4857
rect 1903 4691 1929 4717
rect 1955 4691 1981 4717
rect 2007 4691 2033 4717
rect 11903 4691 11929 4717
rect 11955 4691 11981 4717
rect 12007 4691 12033 4717
rect 21903 4691 21929 4717
rect 21955 4691 21981 4717
rect 22007 4691 22033 4717
rect 29359 4607 29385 4633
rect 30759 4607 30785 4633
rect 1415 4551 1441 4577
rect 2199 4551 2225 4577
rect 8919 4551 8945 4577
rect 10711 4551 10737 4577
rect 11103 4551 11129 4577
rect 14911 4551 14937 4577
rect 20231 4551 20257 4577
rect 20623 4551 20649 4577
rect 23703 4551 23729 4577
rect 24095 4551 24121 4577
rect 28351 4551 28377 4577
rect 28799 4551 28825 4577
rect 2479 4495 2505 4521
rect 10823 4495 10849 4521
rect 14519 4495 14545 4521
rect 14799 4495 14825 4521
rect 20511 4495 20537 4521
rect 23815 4495 23841 4521
rect 26223 4495 26249 4521
rect 26391 4495 26417 4521
rect 29583 4495 29609 4521
rect 31095 4495 31121 4521
rect 2759 4439 2785 4465
rect 26671 4439 26697 4465
rect 30255 4439 30281 4465
rect 31431 4439 31457 4465
rect 1639 4383 1665 4409
rect 1751 4383 1777 4409
rect 8527 4383 8553 4409
rect 8639 4383 8665 4409
rect 27959 4383 27985 4409
rect 28127 4383 28153 4409
rect 28575 4383 28601 4409
rect 2233 4299 2259 4325
rect 2285 4299 2311 4325
rect 2337 4299 2363 4325
rect 12233 4299 12259 4325
rect 12285 4299 12311 4325
rect 12337 4299 12363 4325
rect 22233 4299 22259 4325
rect 22285 4299 22311 4325
rect 22337 4299 22363 4325
rect 2255 4159 2281 4185
rect 2367 4159 2393 4185
rect 21967 4159 21993 4185
rect 22079 4159 22105 4185
rect 28239 4159 28265 4185
rect 30143 4159 30169 4185
rect 30535 4159 30561 4185
rect 6231 4103 6257 4129
rect 27959 4103 27985 4129
rect 28463 4103 28489 4129
rect 28743 4103 28769 4129
rect 28911 4103 28937 4129
rect 29191 4103 29217 4129
rect 29359 4103 29385 4129
rect 30927 4103 30953 4129
rect 2647 4047 2673 4073
rect 6063 4047 6089 4073
rect 6511 4047 6537 4073
rect 21743 4047 21769 4073
rect 27735 4047 27761 4073
rect 29863 4047 29889 4073
rect 31431 3991 31457 4017
rect 1903 3907 1929 3933
rect 1955 3907 1981 3933
rect 2007 3907 2033 3933
rect 11903 3907 11929 3933
rect 11955 3907 11981 3933
rect 12007 3907 12033 3933
rect 21903 3907 21929 3933
rect 21955 3907 21981 3933
rect 22007 3907 22033 3933
rect 31543 3823 31569 3849
rect 7407 3767 7433 3793
rect 17263 3767 17289 3793
rect 17655 3767 17681 3793
rect 21239 3767 21265 3793
rect 28351 3767 28377 3793
rect 29135 3767 29161 3793
rect 29583 3767 29609 3793
rect 30759 3767 30785 3793
rect 17431 3711 17457 3737
rect 21127 3711 21153 3737
rect 28799 3711 28825 3737
rect 29415 3711 29441 3737
rect 31151 3711 31177 3737
rect 7743 3655 7769 3681
rect 20847 3655 20873 3681
rect 30255 3655 30281 3681
rect 7631 3599 7657 3625
rect 28631 3599 28657 3625
rect 28911 3599 28937 3625
rect 2233 3515 2259 3541
rect 2285 3515 2311 3541
rect 2337 3515 2363 3541
rect 12233 3515 12259 3541
rect 12285 3515 12311 3541
rect 12337 3515 12363 3541
rect 22233 3515 22259 3541
rect 22285 3515 22311 3541
rect 22337 3515 22363 3541
rect 30927 3375 30953 3401
rect 8751 3319 8777 3345
rect 9031 3319 9057 3345
rect 15359 3319 15385 3345
rect 18439 3319 18465 3345
rect 18551 3319 18577 3345
rect 23479 3319 23505 3345
rect 23759 3319 23785 3345
rect 25215 3319 25241 3345
rect 25495 3319 25521 3345
rect 29135 3319 29161 3345
rect 29247 3319 29273 3345
rect 29695 3319 29721 3345
rect 29975 3319 30001 3345
rect 30143 3319 30169 3345
rect 9199 3263 9225 3289
rect 15135 3263 15161 3289
rect 15527 3263 15553 3289
rect 18159 3263 18185 3289
rect 23367 3263 23393 3289
rect 25047 3263 25073 3289
rect 28911 3263 28937 3289
rect 29023 3263 29049 3289
rect 29471 3263 29497 3289
rect 31431 3263 31457 3289
rect 30647 3207 30673 3233
rect 1903 3123 1929 3149
rect 1955 3123 1981 3149
rect 2007 3123 2033 3149
rect 11903 3123 11929 3149
rect 11955 3123 11981 3149
rect 12007 3123 12033 3149
rect 21903 3123 21929 3149
rect 21955 3123 21981 3149
rect 22007 3123 22033 3149
rect 30759 3039 30785 3065
rect 31543 3039 31569 3065
rect 1359 2983 1385 3009
rect 4103 2983 4129 3009
rect 4439 2983 4465 3009
rect 13287 2983 13313 3009
rect 13679 2983 13705 3009
rect 14799 2983 14825 3009
rect 21295 2983 21321 3009
rect 28967 2983 28993 3009
rect 29639 2983 29665 3009
rect 1247 2927 1273 2953
rect 4327 2927 4353 2953
rect 13567 2927 13593 2953
rect 30255 2927 30281 2953
rect 31095 2927 31121 2953
rect 967 2871 993 2897
rect 15079 2871 15105 2897
rect 15191 2871 15217 2897
rect 22359 2871 22385 2897
rect 21855 2815 21881 2841
rect 22079 2815 22105 2841
rect 28519 2815 28545 2841
rect 28687 2815 28713 2841
rect 29191 2815 29217 2841
rect 29359 2815 29385 2841
rect 2233 2731 2259 2757
rect 2285 2731 2311 2757
rect 2337 2731 2363 2757
rect 12233 2731 12259 2757
rect 12285 2731 12311 2757
rect 12337 2731 12363 2757
rect 22233 2731 22259 2757
rect 22285 2731 22311 2757
rect 22337 2731 22363 2757
rect 8639 2647 8665 2673
rect 8807 2647 8833 2673
rect 9647 2647 9673 2673
rect 9815 2647 9841 2673
rect 10935 2647 10961 2673
rect 11103 2647 11129 2673
rect 12559 2647 12585 2673
rect 12727 2647 12753 2673
rect 14799 2647 14825 2673
rect 14911 2647 14937 2673
rect 19895 2647 19921 2673
rect 20175 2647 20201 2673
rect 21183 2647 21209 2673
rect 21351 2647 21377 2673
rect 21463 2647 21489 2673
rect 967 2591 993 2617
rect 9367 2591 9393 2617
rect 10655 2591 10681 2617
rect 12279 2591 12305 2617
rect 14519 2591 14545 2617
rect 20455 2591 20481 2617
rect 20903 2591 20929 2617
rect 25439 2591 25465 2617
rect 29191 2591 29217 2617
rect 30143 2591 30169 2617
rect 30535 2591 30561 2617
rect 31319 2591 31345 2617
rect 1247 2535 1273 2561
rect 1415 2535 1441 2561
rect 21743 2535 21769 2561
rect 24991 2535 25017 2561
rect 25159 2535 25185 2561
rect 28183 2535 28209 2561
rect 28351 2535 28377 2561
rect 28631 2535 28657 2561
rect 28743 2535 28769 2561
rect 28911 2535 28937 2561
rect 29583 2535 29609 2561
rect 29695 2535 29721 2561
rect 29975 2535 30001 2561
rect 30927 2535 30953 2561
rect 8415 2479 8441 2505
rect 1903 2339 1929 2365
rect 1955 2339 1981 2365
rect 2007 2339 2033 2365
rect 11903 2339 11929 2365
rect 11955 2339 11981 2365
rect 12007 2339 12033 2365
rect 21903 2339 21929 2365
rect 21955 2339 21981 2365
rect 22007 2339 22033 2365
rect 31543 2255 31569 2281
rect 911 2199 937 2225
rect 8247 2199 8273 2225
rect 21015 2199 21041 2225
rect 21407 2199 21433 2225
rect 24655 2199 24681 2225
rect 27847 2199 27873 2225
rect 21295 2143 21321 2169
rect 24543 2143 24569 2169
rect 30311 2143 30337 2169
rect 31151 2143 31177 2169
rect 24263 2087 24289 2113
rect 30647 2087 30673 2113
rect 1191 2031 1217 2057
rect 1303 2031 1329 2057
rect 8527 2031 8553 2057
rect 8639 2031 8665 2057
rect 28071 2031 28097 2057
rect 28239 2031 28265 2057
rect 2233 1947 2259 1973
rect 2285 1947 2311 1973
rect 2337 1947 2363 1973
rect 12233 1947 12259 1973
rect 12285 1947 12311 1973
rect 12337 1947 12363 1973
rect 22233 1947 22259 1973
rect 22285 1947 22311 1973
rect 22337 1947 22363 1973
rect 2479 1863 2505 1889
rect 2591 1863 2617 1889
rect 8639 1863 8665 1889
rect 8807 1863 8833 1889
rect 12279 1863 12305 1889
rect 20399 1863 20425 1889
rect 20511 1863 20537 1889
rect 23535 1863 23561 1889
rect 23703 1863 23729 1889
rect 25271 1863 25297 1889
rect 25383 1863 25409 1889
rect 29527 1863 29553 1889
rect 29695 1863 29721 1889
rect 2871 1807 2897 1833
rect 8359 1807 8385 1833
rect 11999 1807 12025 1833
rect 22023 1807 22049 1833
rect 22191 1807 22217 1833
rect 22471 1807 22497 1833
rect 23255 1807 23281 1833
rect 24991 1807 25017 1833
rect 30927 1807 30953 1833
rect 1303 1751 1329 1777
rect 1471 1751 1497 1777
rect 29975 1751 30001 1777
rect 30143 1751 30169 1777
rect 1079 1695 1105 1721
rect 11775 1695 11801 1721
rect 20175 1695 20201 1721
rect 29247 1695 29273 1721
rect 30647 1695 30673 1721
rect 31431 1695 31457 1721
rect 1903 1555 1929 1581
rect 1955 1555 1981 1581
rect 2007 1555 2033 1581
rect 11903 1555 11929 1581
rect 11955 1555 11981 1581
rect 12007 1555 12033 1581
rect 21903 1555 21929 1581
rect 21955 1555 21981 1581
rect 22007 1555 22033 1581
rect 31543 1471 31569 1497
rect 26055 1415 26081 1441
rect 29415 1359 29441 1385
rect 29639 1359 29665 1385
rect 31095 1359 31121 1385
rect 29191 1303 29217 1329
rect 30255 1303 30281 1329
rect 30647 1303 30673 1329
rect 26279 1247 26305 1273
rect 26447 1247 26473 1273
rect 28799 1247 28825 1273
rect 28911 1247 28937 1273
rect 2233 1163 2259 1189
rect 2285 1163 2311 1189
rect 2337 1163 2363 1189
rect 12233 1163 12259 1189
rect 12285 1163 12311 1189
rect 12337 1163 12363 1189
rect 22233 1163 22259 1189
rect 22285 1163 22311 1189
rect 22337 1163 22363 1189
rect 1247 1079 1273 1105
rect 1415 1079 1441 1105
rect 7631 1079 7657 1105
rect 8079 1079 8105 1105
rect 8359 1079 8385 1105
rect 11439 1079 11465 1105
rect 11607 1079 11633 1105
rect 15079 1079 15105 1105
rect 15247 1079 15273 1105
rect 15415 1079 15441 1105
rect 18439 1079 18465 1105
rect 18607 1079 18633 1105
rect 19055 1079 19081 1105
rect 19223 1079 19249 1105
rect 19727 1079 19753 1105
rect 19895 1079 19921 1105
rect 20903 1079 20929 1105
rect 21351 1079 21377 1105
rect 22919 1079 22945 1105
rect 23087 1079 23113 1105
rect 6119 1023 6145 1049
rect 6231 1023 6257 1049
rect 6511 1023 6537 1049
rect 7351 1023 7377 1049
rect 7799 1023 7825 1049
rect 11159 1023 11185 1049
rect 16199 1023 16225 1049
rect 16647 1023 16673 1049
rect 17655 1023 17681 1049
rect 18159 1023 18185 1049
rect 20623 1023 20649 1049
rect 21071 1023 21097 1049
rect 21519 1023 21545 1049
rect 24319 1023 24345 1049
rect 24879 1023 24905 1049
rect 25439 1023 25465 1049
rect 28799 1023 28825 1049
rect 29247 1023 29273 1049
rect 30143 1023 30169 1049
rect 4383 967 4409 993
rect 4551 967 4577 993
rect 5055 967 5081 993
rect 5279 967 5305 993
rect 16423 967 16449 993
rect 17935 967 17961 993
rect 19447 967 19473 993
rect 21799 967 21825 993
rect 21967 967 21993 993
rect 24039 967 24065 993
rect 24599 967 24625 993
rect 25159 967 25185 993
rect 28519 967 28545 993
rect 28967 967 28993 993
rect 29695 967 29721 993
rect 29975 967 30001 993
rect 30927 967 30953 993
rect 1023 911 1049 937
rect 4831 911 4857 937
rect 18775 911 18801 937
rect 22695 911 22721 937
rect 23759 911 23785 937
rect 24431 911 24457 937
rect 24991 911 25017 937
rect 28351 911 28377 937
rect 29583 911 29609 937
rect 31431 911 31457 937
rect 30647 855 30673 881
rect 1903 771 1929 797
rect 1955 771 1981 797
rect 2007 771 2033 797
rect 11903 771 11929 797
rect 11955 771 11981 797
rect 12007 771 12033 797
rect 21903 771 21929 797
rect 21955 771 21981 797
rect 22007 771 22033 797
rect 31543 687 31569 713
rect 5279 631 5305 657
rect 7799 631 7825 657
rect 18103 631 18129 657
rect 21071 631 21097 657
rect 21519 631 21545 657
rect 28855 631 28881 657
rect 29807 631 29833 657
rect 30591 631 30617 657
rect 29303 575 29329 601
rect 30087 575 30113 601
rect 31095 575 31121 601
rect 911 519 937 545
rect 4999 519 5025 545
rect 1191 463 1217 489
rect 1303 463 1329 489
rect 4775 463 4801 489
rect 4831 463 4857 489
rect 2233 379 2259 405
rect 2285 379 2311 405
rect 2337 379 2363 405
rect 12233 379 12259 405
rect 12285 379 12311 405
rect 12337 379 12363 405
rect 22233 379 22259 405
rect 22285 379 22311 405
rect 22337 379 22363 405
<< metal2 >>
rect 2128 7056 2184 7112
rect 2352 7056 2408 7112
rect 2576 7056 2632 7112
rect 2800 7056 2856 7112
rect 3024 7056 3080 7112
rect 3248 7056 3304 7112
rect 3472 7056 3528 7112
rect 3696 7056 3752 7112
rect 3920 7056 3976 7112
rect 4144 7056 4200 7112
rect 4368 7056 4424 7112
rect 4592 7056 4648 7112
rect 4816 7056 4872 7112
rect 5040 7056 5096 7112
rect 5264 7056 5320 7112
rect 5488 7056 5544 7112
rect 5712 7056 5768 7112
rect 5936 7056 5992 7112
rect 6160 7056 6216 7112
rect 6384 7056 6440 7112
rect 6608 7056 6664 7112
rect 6832 7056 6888 7112
rect 7056 7056 7112 7112
rect 7280 7056 7336 7112
rect 7504 7056 7560 7112
rect 7728 7056 7784 7112
rect 7952 7056 8008 7112
rect 8176 7056 8232 7112
rect 8400 7056 8456 7112
rect 8624 7056 8680 7112
rect 8848 7056 8904 7112
rect 9072 7056 9128 7112
rect 9296 7056 9352 7112
rect 9520 7056 9576 7112
rect 9744 7056 9800 7112
rect 9968 7056 10024 7112
rect 10192 7056 10248 7112
rect 10416 7056 10472 7112
rect 10640 7056 10696 7112
rect 10864 7056 10920 7112
rect 11088 7056 11144 7112
rect 11312 7056 11368 7112
rect 11536 7056 11592 7112
rect 11760 7056 11816 7112
rect 11984 7056 12040 7112
rect 12208 7056 12264 7112
rect 12432 7056 12488 7112
rect 12656 7056 12712 7112
rect 12880 7056 12936 7112
rect 13104 7056 13160 7112
rect 13328 7056 13384 7112
rect 13552 7056 13608 7112
rect 13776 7056 13832 7112
rect 14000 7056 14056 7112
rect 14224 7056 14280 7112
rect 14448 7056 14504 7112
rect 14672 7056 14728 7112
rect 14896 7056 14952 7112
rect 15120 7056 15176 7112
rect 15344 7056 15400 7112
rect 15568 7056 15624 7112
rect 15792 7056 15848 7112
rect 16016 7056 16072 7112
rect 16240 7056 16296 7112
rect 16464 7056 16520 7112
rect 16688 7056 16744 7112
rect 16912 7056 16968 7112
rect 17136 7056 17192 7112
rect 17360 7056 17416 7112
rect 17584 7056 17640 7112
rect 17808 7056 17864 7112
rect 18032 7056 18088 7112
rect 18256 7056 18312 7112
rect 18480 7056 18536 7112
rect 18704 7056 18760 7112
rect 18928 7056 18984 7112
rect 19152 7056 19208 7112
rect 19376 7056 19432 7112
rect 19600 7056 19656 7112
rect 19824 7056 19880 7112
rect 20048 7056 20104 7112
rect 20272 7056 20328 7112
rect 20496 7056 20552 7112
rect 20720 7056 20776 7112
rect 20944 7056 21000 7112
rect 21168 7056 21224 7112
rect 21392 7056 21448 7112
rect 21616 7056 21672 7112
rect 21840 7056 21896 7112
rect 22064 7056 22120 7112
rect 22288 7056 22344 7112
rect 22512 7056 22568 7112
rect 22736 7056 22792 7112
rect 22960 7056 23016 7112
rect 23184 7056 23240 7112
rect 23408 7056 23464 7112
rect 23632 7056 23688 7112
rect 23856 7056 23912 7112
rect 24080 7056 24136 7112
rect 24304 7056 24360 7112
rect 24528 7056 24584 7112
rect 24752 7056 24808 7112
rect 24976 7056 25032 7112
rect 25200 7056 25256 7112
rect 25424 7056 25480 7112
rect 25648 7056 25704 7112
rect 25872 7056 25928 7112
rect 26096 7056 26152 7112
rect 26320 7056 26376 7112
rect 26544 7056 26600 7112
rect 26768 7056 26824 7112
rect 26992 7056 27048 7112
rect 27216 7056 27272 7112
rect 27440 7056 27496 7112
rect 27664 7056 27720 7112
rect 27888 7056 27944 7112
rect 28112 7056 28168 7112
rect 28336 7056 28392 7112
rect 28560 7056 28616 7112
rect 28784 7056 28840 7112
rect 29008 7056 29064 7112
rect 29232 7056 29288 7112
rect 29456 7056 29512 7112
rect 29680 7056 29736 7112
rect 29904 7056 29960 7112
rect 126 6986 154 6991
rect 126 4130 154 6958
rect 1862 6818 1890 6823
rect 1806 6762 1834 6767
rect 1246 6594 1274 6599
rect 854 6481 882 6487
rect 854 6455 855 6481
rect 881 6455 882 6481
rect 126 4097 154 4102
rect 182 6314 210 6319
rect 182 3738 210 6286
rect 798 6090 826 6095
rect 798 5754 826 6062
rect 798 5721 826 5726
rect 854 4214 882 6455
rect 1078 6426 1106 6431
rect 966 5642 994 5647
rect 966 5595 994 5614
rect 854 4186 1050 4214
rect 182 3705 210 3710
rect 462 4074 490 4079
rect 462 1050 490 4046
rect 966 2898 994 2903
rect 966 2851 994 2870
rect 910 2618 938 2623
rect 910 2225 938 2590
rect 966 2618 994 2623
rect 1022 2618 1050 4186
rect 966 2617 1050 2618
rect 966 2591 967 2617
rect 993 2591 1050 2617
rect 966 2590 1050 2591
rect 966 2585 994 2590
rect 910 2199 911 2225
rect 937 2199 938 2225
rect 910 2193 938 2199
rect 1078 1721 1106 6398
rect 1246 6425 1274 6566
rect 1246 6399 1247 6425
rect 1273 6399 1274 6425
rect 1246 6393 1274 6399
rect 1806 6145 1834 6734
rect 1862 6593 1890 6790
rect 1862 6567 1863 6593
rect 1889 6567 1890 6593
rect 1862 6561 1890 6567
rect 2086 6706 2114 6711
rect 1902 6286 2034 6291
rect 1930 6258 1954 6286
rect 1982 6258 2006 6286
rect 1902 6253 2034 6258
rect 1806 6119 1807 6145
rect 1833 6119 1834 6145
rect 1806 6113 1834 6119
rect 1190 5697 1218 5703
rect 1190 5671 1191 5697
rect 1217 5671 1218 5697
rect 1190 5642 1218 5671
rect 1358 5642 1386 5647
rect 1190 5641 1386 5642
rect 1190 5615 1359 5641
rect 1385 5615 1386 5641
rect 1190 5614 1386 5615
rect 1246 5418 1274 5423
rect 1246 3794 1274 5390
rect 1358 5418 1386 5614
rect 1902 5502 2034 5507
rect 1930 5474 1954 5502
rect 1982 5474 2006 5502
rect 1902 5469 2034 5474
rect 1358 5385 1386 5390
rect 1902 4718 2034 4723
rect 1930 4690 1954 4718
rect 1982 4690 2006 4718
rect 1902 4685 2034 4690
rect 1414 4578 1442 4583
rect 1414 4531 1442 4550
rect 1638 4410 1666 4415
rect 1638 4363 1666 4382
rect 1750 4410 1778 4415
rect 1750 4363 1778 4382
rect 2086 4298 2114 6678
rect 2142 6594 2170 7056
rect 2366 6762 2394 7056
rect 2366 6729 2394 6734
rect 2232 6678 2364 6683
rect 2260 6650 2284 6678
rect 2312 6650 2336 6678
rect 2232 6645 2364 6650
rect 2142 6561 2170 6566
rect 2142 6481 2170 6487
rect 2142 6455 2143 6481
rect 2169 6455 2170 6481
rect 2142 5698 2170 6455
rect 2198 6033 2226 6039
rect 2198 6007 2199 6033
rect 2225 6007 2226 6033
rect 2198 5978 2226 6007
rect 2198 5945 2226 5950
rect 2534 6034 2562 6039
rect 2232 5894 2364 5899
rect 2260 5866 2284 5894
rect 2312 5866 2336 5894
rect 2232 5861 2364 5866
rect 2310 5810 2338 5815
rect 2310 5763 2338 5782
rect 2478 5698 2506 5703
rect 2534 5698 2562 6006
rect 2590 5810 2618 7056
rect 2814 6818 2842 7056
rect 2814 6785 2842 6790
rect 2982 6650 3010 6655
rect 2982 6593 3010 6622
rect 2982 6567 2983 6593
rect 3009 6567 3010 6593
rect 2982 6561 3010 6567
rect 2590 5777 2618 5782
rect 2142 5670 2226 5698
rect 2142 5586 2170 5591
rect 2142 4578 2170 5558
rect 2198 5530 2226 5670
rect 2506 5670 2562 5698
rect 2590 5697 2618 5703
rect 2590 5671 2591 5697
rect 2617 5671 2618 5697
rect 2478 5665 2506 5670
rect 2198 5497 2226 5502
rect 2232 5110 2364 5115
rect 2260 5082 2284 5110
rect 2312 5082 2336 5110
rect 2232 5077 2364 5082
rect 2590 5082 2618 5671
rect 3038 5641 3066 7056
rect 3262 6594 3290 7056
rect 3486 6650 3514 7056
rect 3486 6617 3514 6622
rect 3262 6566 3458 6594
rect 3038 5615 3039 5641
rect 3065 5615 3066 5641
rect 3038 5609 3066 5615
rect 3206 6481 3234 6487
rect 3206 6455 3207 6481
rect 3233 6455 3234 6481
rect 2590 5049 2618 5054
rect 3150 5586 3178 5591
rect 2198 4578 2226 4583
rect 2142 4577 2226 4578
rect 2142 4551 2199 4577
rect 2225 4551 2226 4577
rect 2142 4550 2226 4551
rect 2198 4522 2226 4550
rect 2198 4489 2226 4494
rect 2478 4522 2506 4527
rect 2478 4475 2506 4494
rect 2758 4466 2786 4471
rect 2758 4419 2786 4438
rect 2232 4326 2364 4331
rect 2260 4298 2284 4326
rect 2312 4298 2336 4326
rect 2086 4270 2170 4298
rect 2232 4293 2364 4298
rect 2142 4186 2170 4270
rect 2254 4186 2282 4191
rect 2366 4186 2394 4191
rect 2142 4185 2394 4186
rect 2142 4159 2255 4185
rect 2281 4159 2367 4185
rect 2393 4159 2394 4185
rect 2142 4158 2394 4159
rect 2254 4153 2282 4158
rect 2366 4153 2394 4158
rect 2646 4073 2674 4079
rect 2646 4047 2647 4073
rect 2673 4047 2674 4073
rect 2646 3962 2674 4047
rect 1902 3934 2034 3939
rect 1930 3906 1954 3934
rect 1982 3906 2006 3934
rect 2646 3929 2674 3934
rect 1902 3901 2034 3906
rect 1246 3761 1274 3766
rect 2232 3542 2364 3547
rect 2260 3514 2284 3542
rect 2312 3514 2336 3542
rect 2232 3509 2364 3514
rect 1358 3346 1386 3351
rect 1358 3010 1386 3318
rect 1902 3150 2034 3155
rect 1930 3122 1954 3150
rect 1982 3122 2006 3150
rect 1902 3117 2034 3122
rect 1246 3009 1386 3010
rect 1246 2983 1359 3009
rect 1385 2983 1386 3009
rect 1246 2982 1386 2983
rect 1246 2953 1274 2982
rect 1358 2977 1386 2982
rect 1246 2927 1247 2953
rect 1273 2927 1274 2953
rect 1246 2921 1274 2927
rect 2232 2758 2364 2763
rect 2260 2730 2284 2758
rect 2312 2730 2336 2758
rect 2232 2725 2364 2730
rect 3150 2618 3178 5558
rect 3206 2618 3234 6455
rect 3262 5697 3290 5703
rect 3262 5671 3263 5697
rect 3289 5671 3290 5697
rect 3262 4298 3290 5671
rect 3430 5361 3458 6566
rect 3486 6202 3514 6207
rect 3710 6202 3738 7056
rect 3766 6650 3794 6655
rect 3766 6593 3794 6622
rect 3766 6567 3767 6593
rect 3793 6567 3794 6593
rect 3766 6561 3794 6567
rect 3934 6594 3962 7056
rect 3934 6566 4074 6594
rect 3486 6201 3738 6202
rect 3486 6175 3487 6201
rect 3513 6175 3738 6201
rect 3486 6174 3738 6175
rect 3990 6481 4018 6487
rect 3990 6455 3991 6481
rect 4017 6455 4018 6481
rect 3486 6169 3514 6174
rect 3766 6034 3794 6039
rect 3766 6033 3962 6034
rect 3766 6007 3767 6033
rect 3793 6007 3962 6033
rect 3766 6006 3962 6007
rect 3766 6001 3794 6006
rect 3878 5810 3906 5815
rect 3878 5763 3906 5782
rect 3430 5335 3431 5361
rect 3457 5335 3458 5361
rect 3430 5329 3458 5335
rect 3654 5305 3682 5311
rect 3654 5279 3655 5305
rect 3681 5279 3682 5305
rect 3318 5250 3346 5255
rect 3318 4802 3346 5222
rect 3318 4769 3346 4774
rect 3262 4265 3290 4270
rect 3654 3906 3682 5279
rect 3710 5194 3738 5199
rect 3710 5026 3738 5166
rect 3766 5026 3794 5031
rect 3878 5026 3906 5031
rect 3710 5025 3906 5026
rect 3710 4999 3767 5025
rect 3793 4999 3879 5025
rect 3905 4999 3906 5025
rect 3710 4998 3906 4999
rect 3766 4993 3794 4998
rect 3878 4993 3906 4998
rect 3654 3873 3682 3878
rect 3262 2618 3290 2623
rect 3206 2590 3262 2618
rect 3150 2585 3178 2590
rect 3262 2585 3290 2590
rect 1246 2562 1274 2567
rect 1246 2515 1274 2534
rect 1414 2562 1442 2567
rect 1414 2515 1442 2534
rect 1902 2366 2034 2371
rect 1930 2338 1954 2366
rect 1982 2338 2006 2366
rect 1902 2333 2034 2338
rect 2478 2114 2506 2119
rect 1190 2058 1218 2063
rect 1190 2011 1218 2030
rect 1302 2058 1330 2063
rect 1302 2011 1330 2030
rect 2232 1974 2364 1979
rect 2260 1946 2284 1974
rect 2312 1946 2336 1974
rect 2232 1941 2364 1946
rect 2478 1890 2506 2086
rect 2870 2002 2898 2007
rect 2590 1890 2618 1895
rect 2478 1889 2618 1890
rect 2478 1863 2479 1889
rect 2505 1863 2591 1889
rect 2617 1863 2618 1889
rect 2478 1862 2618 1863
rect 2478 1857 2506 1862
rect 2590 1857 2618 1862
rect 2870 1833 2898 1974
rect 2870 1807 2871 1833
rect 2897 1807 2898 1833
rect 2870 1801 2898 1807
rect 1302 1778 1330 1783
rect 1302 1731 1330 1750
rect 1470 1778 1498 1783
rect 1470 1731 1498 1750
rect 1078 1695 1079 1721
rect 1105 1695 1106 1721
rect 1078 1689 1106 1695
rect 1526 1722 1554 1727
rect 1414 1330 1442 1335
rect 1246 1106 1274 1111
rect 1414 1106 1442 1302
rect 1246 1105 1442 1106
rect 1246 1079 1247 1105
rect 1273 1079 1415 1105
rect 1441 1079 1442 1105
rect 1246 1078 1442 1079
rect 1246 1073 1274 1078
rect 1414 1073 1442 1078
rect 462 1017 490 1022
rect 1022 938 1050 943
rect 1022 891 1050 910
rect 1526 882 1554 1694
rect 1902 1582 2034 1587
rect 1930 1554 1954 1582
rect 1982 1554 2006 1582
rect 1902 1549 2034 1554
rect 2232 1190 2364 1195
rect 2260 1162 2284 1190
rect 2312 1162 2336 1190
rect 2232 1157 2364 1162
rect 3934 1106 3962 6006
rect 3990 4186 4018 6455
rect 4046 5417 4074 6566
rect 4046 5391 4047 5417
rect 4073 5391 4074 5417
rect 4046 5385 4074 5391
rect 4102 5866 4130 5871
rect 3990 4153 4018 4158
rect 4102 3009 4130 5838
rect 4158 5810 4186 7056
rect 4382 6650 4410 7056
rect 4382 6617 4410 6622
rect 4270 6202 4298 6207
rect 4270 6155 4298 6174
rect 4550 6033 4578 6039
rect 4550 6007 4551 6033
rect 4577 6007 4578 6033
rect 4550 5922 4578 6007
rect 4550 5889 4578 5894
rect 4158 5777 4186 5782
rect 4158 5698 4186 5703
rect 4158 5651 4186 5670
rect 4606 5418 4634 7056
rect 4830 6202 4858 7056
rect 4886 6762 4914 6767
rect 4886 6593 4914 6734
rect 4886 6567 4887 6593
rect 4913 6567 4914 6593
rect 4886 6561 4914 6567
rect 5054 6314 5082 7056
rect 5166 6481 5194 6487
rect 5166 6455 5167 6481
rect 5193 6455 5194 6481
rect 5166 6314 5194 6455
rect 5054 6286 5138 6314
rect 4830 6169 4858 6174
rect 5054 6202 5082 6207
rect 5054 6155 5082 6174
rect 4830 5418 4858 5423
rect 4606 5417 4858 5418
rect 4606 5391 4831 5417
rect 4857 5391 4858 5417
rect 4606 5390 4858 5391
rect 4830 5385 4858 5390
rect 4550 5362 4578 5367
rect 4550 5305 4578 5334
rect 4550 5279 4551 5305
rect 4577 5279 4578 5305
rect 4550 5273 4578 5279
rect 4942 5082 4970 5087
rect 4158 5026 4186 5031
rect 4158 4969 4186 4998
rect 4158 4943 4159 4969
rect 4185 4943 4186 4969
rect 4158 4937 4186 4943
rect 4438 3010 4466 3015
rect 4102 2983 4103 3009
rect 4129 2983 4130 3009
rect 4102 2977 4130 2983
rect 4326 2982 4438 3010
rect 4326 2953 4354 2982
rect 4438 2963 4466 2982
rect 4326 2927 4327 2953
rect 4353 2927 4354 2953
rect 4326 2921 4354 2927
rect 4942 2730 4970 5054
rect 5110 4858 5138 6286
rect 5166 6281 5194 6286
rect 5278 6202 5306 7056
rect 5278 6169 5306 6174
rect 5502 6146 5530 7056
rect 5670 6650 5698 6655
rect 5670 6593 5698 6622
rect 5670 6567 5671 6593
rect 5697 6567 5698 6593
rect 5670 6561 5698 6567
rect 5502 6118 5642 6146
rect 5334 6034 5362 6039
rect 5334 6033 5418 6034
rect 5334 6007 5335 6033
rect 5361 6007 5418 6033
rect 5334 6006 5418 6007
rect 5334 6001 5362 6006
rect 5334 5306 5362 5311
rect 5334 5259 5362 5278
rect 5278 4858 5306 4863
rect 5110 4857 5306 4858
rect 5110 4831 5279 4857
rect 5305 4831 5306 4857
rect 5110 4830 5306 4831
rect 5278 4825 5306 4830
rect 5054 4746 5082 4751
rect 4942 2697 4970 2702
rect 4998 3906 5026 3911
rect 4158 2674 4186 2679
rect 4158 2338 4186 2646
rect 4998 2506 5026 3878
rect 5054 3626 5082 4718
rect 5390 4074 5418 6006
rect 5446 5810 5474 5815
rect 5446 5763 5474 5782
rect 5614 5417 5642 6118
rect 5726 5810 5754 7056
rect 5950 6762 5978 7056
rect 5950 6729 5978 6734
rect 5950 6482 5978 6487
rect 5950 6435 5978 6454
rect 5838 6202 5866 6207
rect 5838 6155 5866 6174
rect 6062 6089 6090 6095
rect 6062 6063 6063 6089
rect 6089 6063 6090 6089
rect 5726 5777 5754 5782
rect 5838 6034 5866 6039
rect 5614 5391 5615 5417
rect 5641 5391 5642 5417
rect 5614 5385 5642 5391
rect 5726 5697 5754 5703
rect 5726 5671 5727 5697
rect 5753 5671 5754 5697
rect 5390 4041 5418 4046
rect 5670 4298 5698 4303
rect 5054 3593 5082 3598
rect 4998 2473 5026 2478
rect 4158 2305 4186 2310
rect 5670 1890 5698 4270
rect 5726 3178 5754 5671
rect 5838 5474 5866 6006
rect 5838 5441 5866 5446
rect 6006 5418 6034 5423
rect 5950 5362 5978 5367
rect 5894 4970 5922 4975
rect 5782 4913 5810 4919
rect 5782 4887 5783 4913
rect 5809 4887 5810 4913
rect 5782 4858 5810 4887
rect 5782 4825 5810 4830
rect 5894 4018 5922 4942
rect 5894 3985 5922 3990
rect 5726 3145 5754 3150
rect 5894 3122 5922 3127
rect 5894 2562 5922 3094
rect 5894 2529 5922 2534
rect 5950 2226 5978 5334
rect 6006 5026 6034 5390
rect 6006 4993 6034 4998
rect 6062 4186 6090 6063
rect 6174 5641 6202 7056
rect 6398 6202 6426 7056
rect 6566 6986 6594 6991
rect 6454 6481 6482 6487
rect 6454 6455 6455 6481
rect 6481 6455 6482 6481
rect 6454 6426 6482 6455
rect 6454 6393 6482 6398
rect 6398 6169 6426 6174
rect 6286 5978 6314 5983
rect 6174 5615 6175 5641
rect 6201 5615 6202 5641
rect 6174 5609 6202 5615
rect 6230 5698 6258 5703
rect 6118 5249 6146 5255
rect 6118 5223 6119 5249
rect 6145 5223 6146 5249
rect 6118 5082 6146 5223
rect 6118 5049 6146 5054
rect 6230 4522 6258 5670
rect 6230 4489 6258 4494
rect 6006 4158 6090 4186
rect 6006 2842 6034 4158
rect 6230 4129 6258 4135
rect 6230 4103 6231 4129
rect 6257 4103 6258 4129
rect 6062 4074 6090 4079
rect 6230 4074 6258 4103
rect 6062 4073 6258 4074
rect 6062 4047 6063 4073
rect 6089 4047 6258 4073
rect 6062 4046 6258 4047
rect 6062 2954 6090 4046
rect 6062 2921 6090 2926
rect 6006 2809 6034 2814
rect 5950 2193 5978 2198
rect 5670 1857 5698 1862
rect 3934 1073 3962 1078
rect 6118 1050 6146 1055
rect 6118 1003 6146 1022
rect 6230 1050 6258 1055
rect 6230 1003 6258 1022
rect 4382 994 4410 999
rect 4382 947 4410 966
rect 4550 994 4578 999
rect 4550 947 4578 966
rect 5054 993 5082 999
rect 5054 967 5055 993
rect 5081 967 5082 993
rect 4830 938 4858 943
rect 4830 937 4914 938
rect 4830 911 4831 937
rect 4857 911 4914 937
rect 4830 910 4914 911
rect 4830 905 4858 910
rect 1470 854 1554 882
rect 910 546 938 551
rect 910 499 938 518
rect 1190 490 1218 495
rect 1190 443 1218 462
rect 1302 490 1330 495
rect 1302 443 1330 462
rect 1470 56 1498 854
rect 1902 798 2034 803
rect 1930 770 1954 798
rect 1982 770 2006 798
rect 1902 765 2034 770
rect 4382 770 4410 775
rect 2232 406 2364 411
rect 2260 378 2284 406
rect 2312 378 2336 406
rect 2232 373 2364 378
rect 2926 154 2954 159
rect 2926 56 2954 126
rect 4382 56 4410 742
rect 4774 546 4802 551
rect 4774 489 4802 518
rect 4774 463 4775 489
rect 4801 463 4802 489
rect 1456 0 1512 56
rect 2912 0 2968 56
rect 4368 0 4424 56
rect 4774 42 4802 463
rect 4830 489 4858 495
rect 4830 463 4831 489
rect 4857 463 4858 489
rect 4830 266 4858 463
rect 4830 233 4858 238
rect 4886 210 4914 910
rect 4998 546 5026 551
rect 4998 499 5026 518
rect 5054 266 5082 967
rect 5278 994 5306 999
rect 5278 947 5306 966
rect 5838 826 5866 831
rect 5278 658 5306 663
rect 5278 611 5306 630
rect 5054 233 5082 238
rect 4886 177 4914 182
rect 5838 56 5866 798
rect 6286 770 6314 5950
rect 6510 5697 6538 5703
rect 6510 5671 6511 5697
rect 6537 5671 6538 5697
rect 6342 5306 6370 5311
rect 6342 3066 6370 5278
rect 6510 5306 6538 5671
rect 6510 5273 6538 5278
rect 6398 5250 6426 5255
rect 6426 5222 6482 5250
rect 6398 5203 6426 5222
rect 6454 5194 6482 5222
rect 6510 5194 6538 5199
rect 6454 5193 6538 5194
rect 6454 5167 6511 5193
rect 6537 5167 6538 5193
rect 6454 5166 6538 5167
rect 6510 5161 6538 5166
rect 6342 3033 6370 3038
rect 6510 4073 6538 4079
rect 6510 4047 6511 4073
rect 6537 4047 6538 4073
rect 6510 2562 6538 4047
rect 6566 3010 6594 6958
rect 6622 6650 6650 7056
rect 6622 6617 6650 6622
rect 6678 6986 6706 6991
rect 6678 6426 6706 6958
rect 6846 6874 6874 7056
rect 6846 6846 7042 6874
rect 6622 6398 6706 6426
rect 6958 6762 6986 6767
rect 6958 6425 6986 6734
rect 6958 6399 6959 6425
rect 6985 6399 6986 6425
rect 6622 3122 6650 6398
rect 6958 6393 6986 6399
rect 6678 6314 6706 6319
rect 6678 5082 6706 6286
rect 6902 6090 6930 6095
rect 6734 5697 6762 5703
rect 6734 5671 6735 5697
rect 6761 5671 6762 5697
rect 6734 5586 6762 5671
rect 6734 5553 6762 5558
rect 6790 5249 6818 5255
rect 6790 5223 6791 5249
rect 6817 5223 6818 5249
rect 6678 5054 6762 5082
rect 6734 3906 6762 5054
rect 6678 3878 6762 3906
rect 6678 3570 6706 3878
rect 6734 3794 6762 3799
rect 6734 3682 6762 3766
rect 6734 3649 6762 3654
rect 6734 3570 6762 3575
rect 6678 3542 6734 3570
rect 6734 3537 6762 3542
rect 6622 3089 6650 3094
rect 6790 3122 6818 5223
rect 6902 4578 6930 6062
rect 7014 4858 7042 6846
rect 7070 6146 7098 7056
rect 7294 6314 7322 7056
rect 7518 6762 7546 7056
rect 7518 6729 7546 6734
rect 7462 6538 7490 6543
rect 7462 6491 7490 6510
rect 7182 6286 7322 6314
rect 7350 6482 7378 6487
rect 7070 6118 7154 6146
rect 7070 6033 7098 6039
rect 7070 6007 7071 6033
rect 7097 6007 7098 6033
rect 7070 4970 7098 6007
rect 7126 5418 7154 6118
rect 7182 5641 7210 6286
rect 7182 5615 7183 5641
rect 7209 5615 7210 5641
rect 7182 5609 7210 5615
rect 7238 5810 7266 5815
rect 7182 5418 7210 5423
rect 7126 5417 7210 5418
rect 7126 5391 7183 5417
rect 7209 5391 7210 5417
rect 7126 5390 7210 5391
rect 7182 5385 7210 5390
rect 7070 4942 7154 4970
rect 7070 4858 7098 4863
rect 7014 4857 7098 4858
rect 7014 4831 7071 4857
rect 7097 4831 7098 4857
rect 7014 4830 7098 4831
rect 7070 4825 7098 4830
rect 7126 4690 7154 4942
rect 6902 4545 6930 4550
rect 6958 4662 7154 4690
rect 6958 3850 6986 4662
rect 7182 4634 7210 4639
rect 6790 3089 6818 3094
rect 6846 3822 6986 3850
rect 7070 4578 7098 4583
rect 6566 2977 6594 2982
rect 6510 2529 6538 2534
rect 6678 1778 6706 1783
rect 6510 1274 6538 1279
rect 6510 1049 6538 1246
rect 6510 1023 6511 1049
rect 6537 1023 6538 1049
rect 6510 1017 6538 1023
rect 6286 737 6314 742
rect 6678 322 6706 1750
rect 6846 434 6874 3822
rect 7014 3682 7042 3687
rect 6902 3626 6930 3631
rect 6902 826 6930 3598
rect 7014 1442 7042 3654
rect 7070 2898 7098 4550
rect 7182 2954 7210 4606
rect 7238 3626 7266 5782
rect 7238 3593 7266 3598
rect 7294 5082 7322 5087
rect 7182 2921 7210 2926
rect 7070 2865 7098 2870
rect 7014 1409 7042 1414
rect 7070 2450 7098 2455
rect 7070 1386 7098 2422
rect 7070 1353 7098 1358
rect 7126 2114 7154 2119
rect 7126 1330 7154 2086
rect 7126 1297 7154 1302
rect 7182 1834 7210 1839
rect 6902 793 6930 798
rect 7182 770 7210 1806
rect 7294 1694 7322 5054
rect 7350 3458 7378 6454
rect 7518 6482 7546 6487
rect 7518 6145 7546 6454
rect 7518 6119 7519 6145
rect 7545 6119 7546 6145
rect 7518 6113 7546 6119
rect 7406 5698 7434 5703
rect 7406 3793 7434 5670
rect 7462 5697 7490 5703
rect 7462 5671 7463 5697
rect 7489 5671 7490 5697
rect 7462 4578 7490 5671
rect 7742 5418 7770 7056
rect 7854 6482 7882 6487
rect 7966 6482 7994 7056
rect 7854 6481 7938 6482
rect 7854 6455 7855 6481
rect 7881 6455 7938 6481
rect 7854 6454 7938 6455
rect 7854 6449 7882 6454
rect 7742 5385 7770 5390
rect 7686 5250 7714 5255
rect 7686 5203 7714 5222
rect 7854 5249 7882 5255
rect 7854 5223 7855 5249
rect 7881 5223 7882 5249
rect 7518 4914 7546 4919
rect 7518 4867 7546 4886
rect 7462 4545 7490 4550
rect 7686 4578 7714 4583
rect 7406 3767 7407 3793
rect 7433 3767 7434 3793
rect 7406 3761 7434 3767
rect 7462 4410 7490 4415
rect 7350 3425 7378 3430
rect 7462 2058 7490 4382
rect 7518 3962 7546 3967
rect 7546 3934 7602 3962
rect 7518 3929 7546 3934
rect 7574 2674 7602 3934
rect 7630 3626 7658 3631
rect 7630 3579 7658 3598
rect 7574 2641 7602 2646
rect 7686 2394 7714 4550
rect 7742 3682 7770 3687
rect 7742 3681 7826 3682
rect 7742 3655 7743 3681
rect 7769 3655 7826 3681
rect 7742 3654 7826 3655
rect 7742 3649 7770 3654
rect 7798 3626 7826 3654
rect 7798 3402 7826 3598
rect 7798 3369 7826 3374
rect 7462 2025 7490 2030
rect 7574 2366 7714 2394
rect 7798 2730 7826 2735
rect 7574 1778 7602 2366
rect 7518 1750 7602 1778
rect 7630 2282 7658 2287
rect 7294 1666 7378 1694
rect 7350 1330 7378 1666
rect 7350 1297 7378 1302
rect 7350 1106 7378 1111
rect 7350 1049 7378 1078
rect 7350 1023 7351 1049
rect 7377 1023 7378 1049
rect 7350 1017 7378 1023
rect 7182 737 7210 742
rect 7518 546 7546 1750
rect 7574 1666 7602 1671
rect 7574 826 7602 1638
rect 7630 1554 7658 2254
rect 7630 1521 7658 1526
rect 7686 2170 7714 2175
rect 7630 1106 7658 1111
rect 7686 1106 7714 2142
rect 7630 1105 7770 1106
rect 7630 1079 7631 1105
rect 7657 1079 7770 1105
rect 7630 1078 7770 1079
rect 7630 1073 7658 1078
rect 7574 793 7602 798
rect 7742 658 7770 1078
rect 7798 1049 7826 2702
rect 7854 2058 7882 5223
rect 7910 3346 7938 6454
rect 7966 6449 7994 6454
rect 8190 6370 8218 7056
rect 8414 6538 8442 7056
rect 8414 6505 8442 6510
rect 7966 6342 8218 6370
rect 7966 5641 7994 6342
rect 8190 6202 8218 6207
rect 8190 6155 8218 6174
rect 8638 6202 8666 7056
rect 8694 6650 8722 6655
rect 8694 6593 8722 6622
rect 8694 6567 8695 6593
rect 8721 6567 8722 6593
rect 8694 6561 8722 6567
rect 8638 6169 8666 6174
rect 8470 6034 8498 6039
rect 8470 5987 8498 6006
rect 8750 5922 8778 5927
rect 7966 5615 7967 5641
rect 7993 5615 7994 5641
rect 7966 5609 7994 5615
rect 8638 5642 8666 5647
rect 8134 5418 8162 5423
rect 8134 5371 8162 5390
rect 8638 5305 8666 5614
rect 8750 5642 8778 5894
rect 8750 5609 8778 5614
rect 8862 5418 8890 7056
rect 9086 6538 9114 7056
rect 9086 6510 9226 6538
rect 8974 6482 9002 6487
rect 8974 6481 9170 6482
rect 8974 6455 8975 6481
rect 9001 6455 9170 6481
rect 8974 6454 9170 6455
rect 8974 6449 9002 6454
rect 8974 6202 9002 6207
rect 8974 6155 9002 6174
rect 9030 5698 9058 5703
rect 9030 5651 9058 5670
rect 8918 5418 8946 5423
rect 8862 5417 8946 5418
rect 8862 5391 8919 5417
rect 8945 5391 8946 5417
rect 8862 5390 8946 5391
rect 8918 5385 8946 5390
rect 8638 5279 8639 5305
rect 8665 5279 8666 5305
rect 8638 5273 8666 5279
rect 8246 5250 8274 5255
rect 7910 3313 7938 3318
rect 7966 3626 7994 3631
rect 7854 2030 7938 2058
rect 7798 1023 7799 1049
rect 7825 1023 7826 1049
rect 7798 1017 7826 1023
rect 7854 1946 7882 1951
rect 7854 714 7882 1918
rect 7910 938 7938 2030
rect 7910 905 7938 910
rect 7854 681 7882 686
rect 7798 658 7826 663
rect 7742 657 7826 658
rect 7742 631 7799 657
rect 7825 631 7826 657
rect 7742 630 7826 631
rect 7798 625 7826 630
rect 7518 513 7546 518
rect 6846 401 6874 406
rect 6678 289 6706 294
rect 7294 154 7322 159
rect 7294 56 7322 126
rect 7966 98 7994 3598
rect 8022 3570 8050 3575
rect 8022 546 8050 3542
rect 8246 2225 8274 5222
rect 8918 4690 8946 4695
rect 8918 4577 8946 4662
rect 8918 4551 8919 4577
rect 8945 4551 8946 4577
rect 8918 4545 8946 4551
rect 8526 4410 8554 4415
rect 8638 4410 8666 4415
rect 8526 4409 8666 4410
rect 8526 4383 8527 4409
rect 8553 4383 8639 4409
rect 8665 4383 8666 4409
rect 8526 4382 8666 4383
rect 8526 3234 8554 4382
rect 8638 4377 8666 4382
rect 8806 3794 8834 3799
rect 8526 3201 8554 3206
rect 8582 3458 8610 3463
rect 8414 2506 8442 2511
rect 8414 2459 8442 2478
rect 8246 2199 8247 2225
rect 8273 2199 8274 2225
rect 8246 2193 8274 2199
rect 8470 2282 8498 2287
rect 8414 2002 8442 2007
rect 8358 1834 8386 1839
rect 8358 1787 8386 1806
rect 8414 1498 8442 1974
rect 8414 1465 8442 1470
rect 8414 1162 8442 1167
rect 8078 1106 8106 1111
rect 8078 1059 8106 1078
rect 8358 1106 8386 1111
rect 8358 1059 8386 1078
rect 8414 714 8442 1134
rect 8414 681 8442 686
rect 8470 658 8498 2254
rect 8526 2058 8554 2063
rect 8526 2011 8554 2030
rect 8582 1162 8610 3430
rect 8750 3346 8778 3351
rect 8750 3299 8778 3318
rect 8638 2674 8666 2679
rect 8806 2674 8834 3766
rect 8638 2673 8834 2674
rect 8638 2647 8639 2673
rect 8665 2647 8807 2673
rect 8833 2647 8834 2673
rect 8638 2646 8834 2647
rect 8638 2641 8666 2646
rect 8806 2641 8834 2646
rect 8974 3738 9002 3743
rect 8638 2058 8666 2063
rect 8638 2011 8666 2030
rect 8638 1890 8666 1895
rect 8638 1843 8666 1862
rect 8806 1890 8834 1895
rect 8806 1843 8834 1862
rect 8974 1778 9002 3710
rect 9030 3345 9058 3351
rect 9030 3319 9031 3345
rect 9057 3319 9058 3345
rect 9030 3010 9058 3319
rect 9030 2977 9058 2982
rect 9142 2786 9170 6454
rect 9198 6202 9226 6510
rect 9198 6174 9282 6202
rect 9198 6089 9226 6095
rect 9198 6063 9199 6089
rect 9225 6063 9226 6089
rect 9198 4186 9226 6063
rect 9254 5810 9282 6174
rect 9310 5922 9338 7056
rect 9478 6594 9506 6599
rect 9478 6547 9506 6566
rect 9534 6202 9562 7056
rect 9758 6650 9786 7056
rect 9870 6930 9898 6935
rect 9758 6617 9786 6622
rect 9814 6874 9842 6879
rect 9534 6169 9562 6174
rect 9646 6538 9674 6543
rect 9422 6090 9450 6095
rect 9422 6043 9450 6062
rect 9590 6034 9618 6039
rect 9310 5894 9562 5922
rect 9310 5810 9338 5815
rect 9254 5809 9338 5810
rect 9254 5783 9311 5809
rect 9337 5783 9338 5809
rect 9254 5782 9338 5783
rect 9310 5777 9338 5782
rect 9366 5754 9394 5759
rect 9310 5530 9338 5535
rect 9198 4153 9226 4158
rect 9254 4298 9282 4303
rect 9254 4074 9282 4270
rect 9254 4041 9282 4046
rect 9310 3906 9338 5502
rect 9366 5026 9394 5726
rect 9366 4993 9394 4998
rect 9422 5698 9450 5703
rect 9310 3873 9338 3878
rect 9366 4074 9394 4079
rect 9366 3626 9394 4046
rect 9422 3738 9450 5670
rect 9534 5417 9562 5894
rect 9534 5391 9535 5417
rect 9561 5391 9562 5417
rect 9534 5385 9562 5391
rect 9422 3705 9450 3710
rect 9366 3593 9394 3598
rect 9198 3289 9226 3295
rect 9198 3263 9199 3289
rect 9225 3263 9226 3289
rect 9198 3010 9226 3263
rect 9198 2977 9226 2982
rect 9254 3290 9282 3295
rect 9142 2753 9170 2758
rect 9254 2562 9282 3262
rect 9366 2618 9394 2623
rect 9366 2571 9394 2590
rect 9590 2618 9618 6006
rect 9646 5362 9674 6510
rect 9758 6482 9786 6487
rect 9758 6435 9786 6454
rect 9646 5329 9674 5334
rect 9702 6426 9730 6431
rect 9702 4410 9730 6398
rect 9702 4377 9730 4382
rect 9814 4354 9842 6846
rect 9814 4321 9842 4326
rect 9814 3458 9842 3463
rect 9646 2674 9674 2679
rect 9814 2674 9842 3430
rect 9646 2673 9842 2674
rect 9646 2647 9647 2673
rect 9673 2647 9815 2673
rect 9841 2647 9842 2673
rect 9646 2646 9842 2647
rect 9646 2641 9674 2646
rect 9814 2641 9842 2646
rect 9590 2585 9618 2590
rect 9254 2529 9282 2534
rect 9870 1890 9898 6902
rect 9926 6202 9954 6207
rect 9982 6202 10010 7056
rect 9926 6201 10010 6202
rect 9926 6175 9927 6201
rect 9953 6175 10010 6201
rect 9926 6174 10010 6175
rect 9926 6169 9954 6174
rect 10150 5810 10178 5815
rect 10206 5810 10234 7056
rect 10430 6594 10458 7056
rect 10430 6561 10458 6566
rect 10598 6594 10626 6599
rect 10598 6547 10626 6566
rect 10150 5809 10234 5810
rect 10150 5783 10151 5809
rect 10177 5783 10234 5809
rect 10150 5782 10234 5783
rect 10430 6034 10458 6039
rect 10150 5777 10178 5782
rect 10430 5753 10458 6006
rect 10430 5727 10431 5753
rect 10457 5727 10458 5753
rect 10430 5721 10458 5727
rect 10654 5642 10682 7056
rect 10878 6594 10906 7056
rect 10822 6566 10906 6594
rect 11102 6594 11130 7056
rect 10710 5642 10738 5647
rect 10654 5641 10738 5642
rect 10654 5615 10711 5641
rect 10737 5615 10738 5641
rect 10654 5614 10738 5615
rect 10710 5609 10738 5614
rect 10822 5418 10850 6566
rect 11102 6561 11130 6566
rect 10822 5385 10850 5390
rect 10878 6481 10906 6487
rect 10878 6455 10879 6481
rect 10905 6455 10906 6481
rect 10766 5362 10794 5367
rect 10766 5315 10794 5334
rect 9982 5305 10010 5311
rect 9982 5279 9983 5305
rect 10009 5279 10010 5305
rect 9926 2954 9954 2959
rect 9926 1946 9954 2926
rect 9982 2730 10010 5279
rect 10374 5194 10402 5199
rect 10486 5194 10514 5199
rect 10374 5193 10514 5194
rect 10374 5167 10375 5193
rect 10401 5167 10487 5193
rect 10513 5167 10514 5193
rect 10374 5166 10514 5167
rect 10206 4410 10234 4415
rect 9982 2697 10010 2702
rect 10094 2954 10122 2959
rect 10094 2394 10122 2926
rect 10094 2361 10122 2366
rect 10038 1946 10066 1951
rect 9926 1918 10038 1946
rect 10038 1913 10066 1918
rect 9870 1857 9898 1862
rect 8974 1745 9002 1750
rect 8582 1129 8610 1134
rect 8750 1722 8778 1727
rect 8470 625 8498 630
rect 8022 513 8050 518
rect 7966 65 7994 70
rect 8750 56 8778 1694
rect 10206 1554 10234 4382
rect 10374 3514 10402 5166
rect 10486 5161 10514 5166
rect 10542 5138 10570 5143
rect 10374 3481 10402 3486
rect 10430 4354 10458 4359
rect 10430 2338 10458 4326
rect 10430 2305 10458 2310
rect 10486 3906 10514 3911
rect 10486 1666 10514 3878
rect 10486 1633 10514 1638
rect 10206 1521 10234 1526
rect 10206 770 10234 775
rect 10206 56 10234 742
rect 10542 266 10570 5110
rect 10878 5026 10906 6455
rect 10878 4993 10906 4998
rect 10934 6370 10962 6375
rect 10710 4746 10738 4751
rect 10710 4578 10738 4718
rect 10710 4577 10850 4578
rect 10710 4551 10711 4577
rect 10737 4551 10850 4577
rect 10710 4550 10850 4551
rect 10710 4545 10738 4550
rect 10822 4521 10850 4550
rect 10822 4495 10823 4521
rect 10849 4495 10850 4521
rect 10822 4489 10850 4495
rect 10822 3850 10850 3855
rect 10654 2618 10682 2623
rect 10654 2571 10682 2590
rect 10822 2338 10850 3822
rect 10934 2674 10962 6342
rect 11158 6202 11186 6207
rect 11158 5697 11186 6174
rect 11214 6202 11242 6207
rect 11326 6202 11354 7056
rect 11382 6594 11410 6599
rect 11382 6547 11410 6566
rect 11214 6201 11354 6202
rect 11214 6175 11215 6201
rect 11241 6175 11354 6201
rect 11214 6174 11354 6175
rect 11214 6169 11242 6174
rect 11158 5671 11159 5697
rect 11185 5671 11186 5697
rect 11158 5665 11186 5671
rect 11494 6033 11522 6039
rect 11494 6007 11495 6033
rect 11521 6007 11522 6033
rect 11102 5418 11130 5423
rect 11102 5371 11130 5390
rect 11438 5250 11466 5255
rect 11102 4914 11130 4919
rect 11102 4577 11130 4886
rect 11102 4551 11103 4577
rect 11129 4551 11130 4577
rect 11102 4545 11130 4551
rect 11438 4578 11466 5222
rect 11494 5138 11522 6007
rect 11550 5641 11578 7056
rect 11662 6482 11690 6487
rect 11662 6481 11746 6482
rect 11662 6455 11663 6481
rect 11689 6455 11746 6481
rect 11662 6454 11746 6455
rect 11662 6449 11690 6454
rect 11550 5615 11551 5641
rect 11577 5615 11578 5641
rect 11550 5609 11578 5615
rect 11606 6090 11634 6095
rect 11606 5305 11634 6062
rect 11606 5279 11607 5305
rect 11633 5279 11634 5305
rect 11606 5273 11634 5279
rect 11718 5194 11746 6454
rect 11774 5474 11802 7056
rect 11998 6594 12026 7056
rect 12222 6762 12250 7056
rect 11998 6561 12026 6566
rect 12166 6734 12250 6762
rect 11902 6286 12034 6291
rect 11930 6258 11954 6286
rect 11982 6258 12006 6286
rect 11902 6253 12034 6258
rect 11998 6202 12026 6207
rect 12166 6202 12194 6734
rect 12232 6678 12364 6683
rect 12260 6650 12284 6678
rect 12312 6650 12336 6678
rect 12232 6645 12364 6650
rect 11998 6201 12194 6202
rect 11998 6175 11999 6201
rect 12025 6175 12194 6201
rect 11998 6174 12194 6175
rect 12222 6258 12250 6263
rect 11998 6169 12026 6174
rect 12222 6146 12250 6230
rect 12446 6202 12474 7056
rect 12670 6706 12698 7056
rect 12502 6678 12698 6706
rect 12502 6593 12530 6678
rect 12502 6567 12503 6593
rect 12529 6567 12530 6593
rect 12502 6561 12530 6567
rect 12726 6481 12754 6487
rect 12726 6455 12727 6481
rect 12753 6455 12754 6481
rect 12558 6202 12586 6207
rect 12446 6201 12586 6202
rect 12446 6175 12559 6201
rect 12585 6175 12586 6201
rect 12446 6174 12586 6175
rect 12558 6169 12586 6174
rect 12166 6118 12250 6146
rect 11998 5697 12026 5703
rect 11998 5671 11999 5697
rect 12025 5671 12026 5697
rect 11998 5586 12026 5671
rect 11998 5553 12026 5558
rect 11902 5502 12034 5507
rect 11930 5474 11954 5502
rect 11982 5474 12006 5502
rect 11774 5446 11858 5474
rect 11902 5469 12034 5474
rect 11830 5418 11858 5446
rect 11998 5418 12026 5423
rect 11830 5417 12026 5418
rect 11830 5391 11999 5417
rect 12025 5391 12026 5417
rect 11830 5390 12026 5391
rect 11998 5385 12026 5390
rect 11718 5166 11802 5194
rect 11494 5110 11746 5138
rect 11438 4545 11466 4550
rect 10934 2627 10962 2646
rect 10990 4242 11018 4247
rect 10822 2305 10850 2310
rect 10878 2562 10906 2567
rect 10878 1722 10906 2534
rect 10878 1689 10906 1694
rect 10990 826 11018 4214
rect 11662 4186 11690 4191
rect 11606 3402 11634 3407
rect 11102 2674 11130 2679
rect 11102 2627 11130 2646
rect 11158 1666 11186 1671
rect 11158 1049 11186 1638
rect 11158 1023 11159 1049
rect 11185 1023 11186 1049
rect 11158 1017 11186 1023
rect 11326 1442 11354 1447
rect 11326 882 11354 1414
rect 11438 1106 11466 1111
rect 11606 1106 11634 3374
rect 11662 3290 11690 4158
rect 11662 3257 11690 3262
rect 11662 2506 11690 2511
rect 11662 2170 11690 2478
rect 11662 2137 11690 2142
rect 11718 1666 11746 5110
rect 11774 4970 11802 5166
rect 11774 4937 11802 4942
rect 11902 4718 12034 4723
rect 11930 4690 11954 4718
rect 11982 4690 12006 4718
rect 11902 4685 12034 4690
rect 12110 4690 12138 4695
rect 12110 4354 12138 4662
rect 12110 4321 12138 4326
rect 11902 3934 12034 3939
rect 11930 3906 11954 3934
rect 11982 3906 12006 3934
rect 11902 3901 12034 3906
rect 12110 3906 12138 3911
rect 11902 3150 12034 3155
rect 11930 3122 11954 3150
rect 11982 3122 12006 3150
rect 11902 3117 12034 3122
rect 12110 2954 12138 3878
rect 12166 3402 12194 6118
rect 12278 6034 12306 6039
rect 12278 6033 12586 6034
rect 12278 6007 12279 6033
rect 12305 6007 12586 6033
rect 12278 6006 12586 6007
rect 12278 6001 12306 6006
rect 12502 5922 12530 5927
rect 12232 5894 12364 5899
rect 12260 5866 12284 5894
rect 12312 5866 12336 5894
rect 12232 5861 12364 5866
rect 12502 5418 12530 5894
rect 12502 5385 12530 5390
rect 12502 5249 12530 5255
rect 12502 5223 12503 5249
rect 12529 5223 12530 5249
rect 12232 5110 12364 5115
rect 12260 5082 12284 5110
rect 12312 5082 12336 5110
rect 12232 5077 12364 5082
rect 12502 5082 12530 5223
rect 12502 5049 12530 5054
rect 12502 4410 12530 4415
rect 12232 4326 12364 4331
rect 12260 4298 12284 4326
rect 12312 4298 12336 4326
rect 12232 4293 12364 4298
rect 12232 3542 12364 3547
rect 12260 3514 12284 3542
rect 12312 3514 12336 3542
rect 12232 3509 12364 3514
rect 12166 3369 12194 3374
rect 12110 2921 12138 2926
rect 12166 3066 12194 3071
rect 12166 2618 12194 3038
rect 12502 2954 12530 4382
rect 12558 3962 12586 6006
rect 12726 5362 12754 6455
rect 12894 5642 12922 7056
rect 13118 6146 13146 7056
rect 13286 6594 13314 6599
rect 13342 6594 13370 7056
rect 13566 6762 13594 7056
rect 13566 6729 13594 6734
rect 13286 6593 13370 6594
rect 13286 6567 13287 6593
rect 13313 6567 13370 6593
rect 13286 6566 13370 6567
rect 13510 6706 13538 6711
rect 13286 6561 13314 6566
rect 13118 6113 13146 6118
rect 13454 6146 13482 6151
rect 13454 6099 13482 6118
rect 13062 6034 13090 6039
rect 13062 6033 13202 6034
rect 13062 6007 13063 6033
rect 13089 6007 13202 6033
rect 13062 6006 13202 6007
rect 13062 6001 13090 6006
rect 13118 5642 13146 5647
rect 12894 5641 13146 5642
rect 12894 5615 13119 5641
rect 13145 5615 13146 5641
rect 12894 5614 13146 5615
rect 13118 5609 13146 5614
rect 13118 5530 13146 5535
rect 12726 5334 12810 5362
rect 12558 3929 12586 3934
rect 12614 5138 12642 5143
rect 12558 3738 12586 3743
rect 12614 3738 12642 5110
rect 12726 4746 12754 4751
rect 12726 4130 12754 4718
rect 12726 4097 12754 4102
rect 12586 3710 12642 3738
rect 12558 3705 12586 3710
rect 12502 2921 12530 2926
rect 12232 2758 12364 2763
rect 12260 2730 12284 2758
rect 12312 2730 12336 2758
rect 12232 2725 12364 2730
rect 12558 2674 12586 2679
rect 12558 2627 12586 2646
rect 12726 2674 12754 2679
rect 12726 2627 12754 2646
rect 12278 2618 12306 2623
rect 12166 2617 12306 2618
rect 12166 2591 12279 2617
rect 12305 2591 12306 2617
rect 12166 2590 12306 2591
rect 12278 2585 12306 2590
rect 12446 2562 12474 2567
rect 11902 2366 12034 2371
rect 11830 2338 11858 2343
rect 11930 2338 11954 2366
rect 11982 2338 12006 2366
rect 11902 2333 12034 2338
rect 12110 2338 12138 2343
rect 11774 2226 11802 2231
rect 11830 2226 11858 2310
rect 11886 2226 11914 2231
rect 11830 2198 11886 2226
rect 11774 1721 11802 2198
rect 11886 2193 11914 2198
rect 11942 2114 11970 2119
rect 11942 1834 11970 2086
rect 12110 2002 12138 2310
rect 12110 1969 12138 1974
rect 12166 2114 12194 2119
rect 12166 1946 12194 2086
rect 12232 1974 12364 1979
rect 12260 1946 12284 1974
rect 12312 1946 12336 1974
rect 12232 1941 12364 1946
rect 12166 1913 12194 1918
rect 12278 1890 12306 1895
rect 12446 1890 12474 2534
rect 12782 1946 12810 5334
rect 13006 4018 13034 4023
rect 13006 2786 13034 3990
rect 13006 2753 13034 2758
rect 12782 1913 12810 1918
rect 12950 2226 12978 2231
rect 12222 1889 12474 1890
rect 12222 1863 12279 1889
rect 12305 1863 12474 1889
rect 12222 1862 12474 1863
rect 11942 1801 11970 1806
rect 11998 1834 12026 1839
rect 12222 1834 12250 1862
rect 12278 1857 12306 1862
rect 11998 1833 12250 1834
rect 11998 1807 11999 1833
rect 12025 1807 12250 1833
rect 11998 1806 12250 1807
rect 11998 1801 12026 1806
rect 11774 1695 11775 1721
rect 11801 1695 11802 1721
rect 11774 1689 11802 1695
rect 12894 1778 12922 1783
rect 12950 1778 12978 2198
rect 13118 1890 13146 5502
rect 13174 4578 13202 6006
rect 13342 5866 13370 5871
rect 13342 4690 13370 5838
rect 13510 5810 13538 6678
rect 13510 5777 13538 5782
rect 13566 6481 13594 6487
rect 13566 6455 13567 6481
rect 13593 6455 13594 6481
rect 13510 5642 13538 5647
rect 13454 5530 13482 5535
rect 13342 4657 13370 4662
rect 13398 4858 13426 4863
rect 13174 4545 13202 4550
rect 13230 4354 13258 4359
rect 13174 2954 13202 2959
rect 13174 2450 13202 2926
rect 13174 2417 13202 2422
rect 13230 2282 13258 4326
rect 13398 3570 13426 4830
rect 13398 3537 13426 3542
rect 13286 3290 13314 3295
rect 13286 3009 13314 3262
rect 13286 2983 13287 3009
rect 13313 2983 13314 3009
rect 13286 2977 13314 2983
rect 13398 2954 13426 2959
rect 13230 2249 13258 2254
rect 13286 2394 13314 2399
rect 13118 1857 13146 1862
rect 13118 1778 13146 1783
rect 12950 1750 13118 1778
rect 11718 1633 11746 1638
rect 12894 1666 12922 1750
rect 13118 1745 13146 1750
rect 12894 1633 12922 1638
rect 11830 1610 11858 1615
rect 11830 1386 11858 1582
rect 11902 1582 12034 1587
rect 11930 1554 11954 1582
rect 11982 1554 12006 1582
rect 11902 1549 12034 1554
rect 13006 1554 13034 1559
rect 11830 1353 11858 1358
rect 12232 1190 12364 1195
rect 11438 1105 11634 1106
rect 11438 1079 11439 1105
rect 11465 1079 11607 1105
rect 11633 1079 11634 1105
rect 11438 1078 11634 1079
rect 11438 1073 11466 1078
rect 11606 1073 11634 1078
rect 12166 1162 12194 1167
rect 12260 1162 12284 1190
rect 12312 1162 12336 1190
rect 12232 1157 12364 1162
rect 12166 1050 12194 1134
rect 12166 1017 12194 1022
rect 13006 994 13034 1526
rect 13286 1498 13314 2366
rect 13398 2114 13426 2926
rect 13454 2674 13482 5502
rect 13510 4410 13538 5614
rect 13510 4377 13538 4382
rect 13566 4214 13594 6455
rect 13790 6258 13818 7056
rect 13958 6762 13986 6767
rect 13958 6425 13986 6734
rect 13958 6399 13959 6425
rect 13985 6399 13986 6425
rect 13958 6393 13986 6399
rect 14014 6314 14042 7056
rect 14238 7042 14266 7056
rect 14238 7009 14266 7014
rect 14462 6986 14490 7056
rect 14462 6953 14490 6958
rect 14574 6594 14602 6599
rect 14462 6481 14490 6487
rect 14462 6455 14463 6481
rect 14489 6455 14490 6481
rect 14014 6286 14154 6314
rect 13790 6225 13818 6230
rect 14070 6202 14098 6207
rect 13734 6089 13762 6095
rect 13734 6063 13735 6089
rect 13761 6063 13762 6089
rect 13622 5698 13650 5703
rect 13622 5651 13650 5670
rect 13734 5138 13762 6063
rect 13790 6090 13818 6095
rect 13790 5810 13818 6062
rect 13790 5777 13818 5782
rect 14014 5697 14042 5703
rect 14014 5671 14015 5697
rect 14041 5671 14042 5697
rect 13734 5105 13762 5110
rect 13846 5642 13874 5647
rect 14014 5642 14042 5671
rect 13846 5641 14042 5642
rect 13846 5615 13847 5641
rect 13873 5615 14042 5641
rect 13846 5614 14042 5615
rect 13566 4186 13818 4214
rect 13734 3850 13762 3855
rect 13510 3402 13538 3407
rect 13510 2898 13538 3374
rect 13678 3010 13706 3015
rect 13566 2982 13678 3010
rect 13566 2953 13594 2982
rect 13678 2963 13706 2982
rect 13566 2927 13567 2953
rect 13593 2927 13594 2953
rect 13566 2921 13594 2927
rect 13510 2865 13538 2870
rect 13622 2898 13650 2903
rect 13454 2641 13482 2646
rect 13398 2081 13426 2086
rect 13566 2282 13594 2287
rect 13286 1465 13314 1470
rect 13454 2058 13482 2063
rect 13006 961 13034 966
rect 11326 849 11354 854
rect 11830 938 11858 943
rect 10990 793 11018 798
rect 11830 770 11858 910
rect 13454 826 13482 2030
rect 11902 798 12034 803
rect 11930 770 11954 798
rect 11982 770 12006 798
rect 13454 793 13482 798
rect 13510 1442 13538 1447
rect 11902 765 12034 770
rect 11830 737 11858 742
rect 10542 233 10570 238
rect 11662 658 11690 663
rect 11662 56 11690 630
rect 13510 546 13538 1414
rect 13566 602 13594 2254
rect 13566 569 13594 574
rect 13510 513 13538 518
rect 12232 406 12364 411
rect 12260 378 12284 406
rect 12312 378 12336 406
rect 12232 373 12364 378
rect 13118 322 13146 327
rect 13118 56 13146 294
rect 13622 154 13650 2870
rect 13734 1722 13762 3822
rect 13734 1689 13762 1694
rect 13790 1162 13818 4186
rect 13846 4074 13874 5614
rect 14070 4970 14098 6174
rect 13846 4041 13874 4046
rect 13958 4942 14098 4970
rect 13902 4018 13930 4023
rect 13902 2394 13930 3990
rect 13902 2361 13930 2366
rect 13958 2114 13986 4942
rect 14014 4746 14042 4751
rect 14014 3458 14042 4718
rect 14014 3425 14042 3430
rect 14070 3962 14098 3967
rect 13958 2081 13986 2086
rect 14070 2058 14098 3934
rect 14070 2025 14098 2030
rect 13958 1778 13986 1783
rect 13958 1610 13986 1750
rect 13958 1577 13986 1582
rect 13790 1129 13818 1134
rect 14126 1106 14154 6286
rect 14462 6146 14490 6455
rect 14462 6113 14490 6118
rect 14294 6034 14322 6039
rect 14238 5642 14266 5647
rect 14238 5595 14266 5614
rect 14294 5586 14322 6006
rect 14518 5978 14546 5983
rect 14518 5931 14546 5950
rect 14294 5553 14322 5558
rect 14406 5922 14434 5927
rect 14406 5474 14434 5894
rect 14574 5866 14602 6566
rect 14630 5978 14658 5983
rect 14630 5931 14658 5950
rect 14294 5446 14434 5474
rect 14518 5838 14602 5866
rect 14182 5026 14210 5031
rect 14182 4186 14210 4998
rect 14182 4153 14210 4158
rect 14238 4242 14266 4247
rect 14238 2562 14266 4214
rect 14294 3626 14322 5446
rect 14518 5418 14546 5838
rect 14686 5530 14714 7056
rect 14910 6650 14938 7056
rect 14910 6617 14938 6622
rect 14910 6538 14938 6543
rect 14910 6145 14938 6510
rect 15134 6314 15162 7056
rect 14910 6119 14911 6145
rect 14937 6119 14938 6145
rect 14910 6113 14938 6119
rect 14966 6286 15162 6314
rect 14686 5497 14714 5502
rect 14350 5390 14546 5418
rect 14574 5418 14602 5423
rect 14350 3850 14378 5390
rect 14350 3817 14378 3822
rect 14406 4858 14434 4863
rect 14294 3593 14322 3598
rect 14350 3738 14378 3743
rect 14350 2618 14378 3710
rect 14350 2585 14378 2590
rect 14238 2529 14266 2534
rect 14406 2338 14434 4830
rect 14518 4522 14546 4527
rect 14518 4475 14546 4494
rect 14462 3962 14490 3967
rect 14462 2898 14490 3934
rect 14462 2865 14490 2870
rect 14518 2618 14546 2623
rect 14518 2571 14546 2590
rect 14406 2305 14434 2310
rect 14126 1073 14154 1078
rect 14182 1946 14210 1951
rect 14182 994 14210 1918
rect 14182 961 14210 966
rect 14294 1946 14322 1951
rect 14294 938 14322 1918
rect 14294 905 14322 910
rect 14350 1834 14378 1839
rect 14350 602 14378 1806
rect 14574 1778 14602 5390
rect 14966 5306 14994 6286
rect 14910 5278 14994 5306
rect 15022 6202 15050 6207
rect 14742 4634 14770 4639
rect 14686 4522 14714 4527
rect 14574 1745 14602 1750
rect 14630 1890 14658 1895
rect 14630 1498 14658 1862
rect 14630 1465 14658 1470
rect 14406 882 14434 887
rect 14406 770 14434 854
rect 14406 737 14434 742
rect 14686 658 14714 4494
rect 14742 3010 14770 4606
rect 14910 4578 14938 5278
rect 14798 4577 14938 4578
rect 14798 4551 14911 4577
rect 14937 4551 14938 4577
rect 14798 4550 14938 4551
rect 14798 4521 14826 4550
rect 14910 4545 14938 4550
rect 14966 5138 14994 5143
rect 14798 4495 14799 4521
rect 14825 4495 14826 4521
rect 14798 4489 14826 4495
rect 14910 3458 14938 3463
rect 14798 3010 14826 3015
rect 14742 3009 14826 3010
rect 14742 2983 14799 3009
rect 14825 2983 14826 3009
rect 14742 2982 14826 2983
rect 14798 2977 14826 2982
rect 14798 2674 14826 2679
rect 14910 2674 14938 3430
rect 14798 2673 14938 2674
rect 14798 2647 14799 2673
rect 14825 2647 14911 2673
rect 14937 2647 14938 2673
rect 14798 2646 14938 2647
rect 14798 2641 14826 2646
rect 14910 2641 14938 2646
rect 14966 994 14994 5110
rect 15022 2282 15050 6174
rect 15190 6146 15218 6151
rect 15190 6099 15218 6118
rect 15302 6146 15330 6151
rect 15246 6034 15274 6039
rect 15190 5978 15218 5983
rect 15190 4970 15218 5950
rect 15190 4937 15218 4942
rect 15246 4522 15274 6006
rect 15246 4489 15274 4494
rect 15134 4242 15162 4247
rect 15302 4214 15330 6118
rect 15078 4186 15162 4214
rect 15246 4186 15330 4214
rect 15078 4153 15106 4158
rect 15134 3289 15162 3295
rect 15134 3263 15135 3289
rect 15161 3263 15162 3289
rect 15078 2898 15106 2903
rect 15078 2851 15106 2870
rect 15134 2730 15162 3263
rect 15190 2898 15218 2903
rect 15246 2898 15274 4186
rect 15358 3738 15386 7056
rect 15582 6594 15610 7056
rect 15582 6561 15610 6566
rect 15414 6370 15442 6375
rect 15414 5978 15442 6342
rect 15582 6370 15610 6375
rect 15582 6146 15610 6342
rect 15470 6145 15610 6146
rect 15470 6119 15583 6145
rect 15609 6119 15610 6145
rect 15470 6118 15610 6119
rect 15470 6089 15498 6118
rect 15582 6113 15610 6118
rect 15470 6063 15471 6089
rect 15497 6063 15498 6089
rect 15470 6057 15498 6063
rect 15414 5950 15778 5978
rect 15582 5866 15610 5871
rect 15358 3705 15386 3710
rect 15470 4914 15498 4919
rect 15358 3345 15386 3351
rect 15358 3319 15359 3345
rect 15385 3319 15386 3345
rect 15358 3290 15386 3319
rect 15358 3257 15386 3262
rect 15246 2870 15386 2898
rect 15190 2851 15218 2870
rect 15134 2697 15162 2702
rect 15022 2249 15050 2254
rect 15078 2562 15106 2567
rect 15078 1106 15106 2534
rect 15190 2562 15218 2567
rect 15134 2282 15162 2287
rect 15134 1442 15162 2254
rect 15190 1666 15218 2534
rect 15190 1633 15218 1638
rect 15134 1409 15162 1414
rect 15246 1106 15274 1111
rect 15078 1105 15274 1106
rect 15078 1079 15079 1105
rect 15105 1079 15247 1105
rect 15273 1079 15274 1105
rect 15078 1078 15274 1079
rect 15078 1073 15106 1078
rect 15246 1073 15274 1078
rect 14966 961 14994 966
rect 14686 625 14714 630
rect 14350 569 14378 574
rect 15358 490 15386 2870
rect 15414 2786 15442 2791
rect 15414 2506 15442 2758
rect 15414 2473 15442 2478
rect 15470 2394 15498 4886
rect 15582 4914 15610 5838
rect 15582 4881 15610 4886
rect 15638 5698 15666 5703
rect 15582 3850 15610 3855
rect 15526 3290 15554 3295
rect 15526 3243 15554 3262
rect 15470 2361 15498 2366
rect 15582 2170 15610 3822
rect 15582 2137 15610 2142
rect 15414 1274 15442 1279
rect 15414 1105 15442 1246
rect 15414 1079 15415 1105
rect 15441 1079 15442 1105
rect 15414 1073 15442 1079
rect 15638 1106 15666 5670
rect 15694 4298 15722 4303
rect 15694 3122 15722 4270
rect 15750 4214 15778 5950
rect 15806 5922 15834 7056
rect 15862 6426 15890 6431
rect 15862 6314 15890 6398
rect 15862 6281 15890 6286
rect 15918 5922 15946 5927
rect 15806 5889 15834 5894
rect 15862 5894 15918 5922
rect 15862 4858 15890 5894
rect 15918 5889 15946 5894
rect 15862 4825 15890 4830
rect 15918 5250 15946 5255
rect 15750 4186 15834 4214
rect 15806 4130 15834 4186
rect 15806 4097 15834 4102
rect 15694 3089 15722 3094
rect 15918 2618 15946 5222
rect 16030 3794 16058 7056
rect 16254 6930 16282 7056
rect 16254 6897 16282 6902
rect 16310 6986 16338 6991
rect 16254 6426 16282 6431
rect 16254 6090 16282 6398
rect 16254 6057 16282 6062
rect 16310 5978 16338 6958
rect 16254 5950 16338 5978
rect 16366 6090 16394 6095
rect 16030 3761 16058 3766
rect 16086 5082 16114 5087
rect 16086 2954 16114 5054
rect 16086 2921 16114 2926
rect 16142 4970 16170 4975
rect 15918 2585 15946 2590
rect 16142 2282 16170 4942
rect 16254 4214 16282 5950
rect 16310 5642 16338 5647
rect 16310 5362 16338 5614
rect 16310 5329 16338 5334
rect 16254 4186 16338 4214
rect 16142 2249 16170 2254
rect 15638 1073 15666 1078
rect 16198 1050 16226 1055
rect 16310 1050 16338 4186
rect 16366 3010 16394 6062
rect 16478 5978 16506 7056
rect 16478 5945 16506 5950
rect 16590 6650 16618 6655
rect 16590 3794 16618 6622
rect 16646 5306 16674 5311
rect 16646 3906 16674 5278
rect 16646 3873 16674 3878
rect 16590 3761 16618 3766
rect 16702 3458 16730 7056
rect 16926 6594 16954 7056
rect 16926 6561 16954 6566
rect 17150 6482 17178 7056
rect 17150 6449 17178 6454
rect 16814 6314 16842 6319
rect 16814 5866 16842 6286
rect 17206 6202 17234 6207
rect 17094 6034 17122 6039
rect 16758 5838 16842 5866
rect 16982 5922 17010 5927
rect 16758 4746 16786 5838
rect 16758 4713 16786 4718
rect 16926 4858 16954 4863
rect 16926 3850 16954 4830
rect 16926 3817 16954 3822
rect 16702 3425 16730 3430
rect 16366 2977 16394 2982
rect 16758 3402 16786 3407
rect 16758 2506 16786 3374
rect 16982 3402 17010 5894
rect 17038 5754 17066 5759
rect 17038 5530 17066 5726
rect 17038 5497 17066 5502
rect 16982 3369 17010 3374
rect 17038 4242 17066 4247
rect 16758 2473 16786 2478
rect 17038 2338 17066 4214
rect 17094 3738 17122 6006
rect 17150 5866 17178 5871
rect 17150 5754 17178 5838
rect 17150 5721 17178 5726
rect 17150 4802 17178 4807
rect 17150 4074 17178 4774
rect 17150 4041 17178 4046
rect 17094 3705 17122 3710
rect 17206 2674 17234 6174
rect 17318 6202 17346 6207
rect 17262 5866 17290 5871
rect 17262 3962 17290 5838
rect 17318 5250 17346 6174
rect 17374 5922 17402 7056
rect 17598 6818 17626 7056
rect 17598 6785 17626 6790
rect 17486 6706 17514 6711
rect 17374 5889 17402 5894
rect 17430 6258 17458 6263
rect 17318 5222 17402 5250
rect 17318 5138 17346 5143
rect 17318 5026 17346 5110
rect 17318 4993 17346 4998
rect 17374 4970 17402 5222
rect 17430 5026 17458 6230
rect 17486 6146 17514 6678
rect 17486 6145 17626 6146
rect 17486 6119 17487 6145
rect 17513 6119 17626 6145
rect 17486 6118 17626 6119
rect 17486 6113 17514 6118
rect 17598 6089 17626 6118
rect 17598 6063 17599 6089
rect 17625 6063 17626 6089
rect 17598 6057 17626 6063
rect 17598 5978 17626 5983
rect 17430 4993 17458 4998
rect 17486 5642 17514 5647
rect 17374 4937 17402 4942
rect 17262 3929 17290 3934
rect 17262 3794 17290 3799
rect 17290 3766 17458 3794
rect 17262 3747 17290 3766
rect 17430 3737 17458 3766
rect 17430 3711 17431 3737
rect 17457 3711 17458 3737
rect 17430 3705 17458 3711
rect 17262 3402 17290 3407
rect 17262 2786 17290 3374
rect 17486 3178 17514 5614
rect 17542 5194 17570 5199
rect 17542 4802 17570 5166
rect 17542 4769 17570 4774
rect 17598 3850 17626 5950
rect 17598 3817 17626 3822
rect 17654 3793 17682 3799
rect 17654 3767 17655 3793
rect 17681 3767 17682 3793
rect 17654 3682 17682 3767
rect 17822 3794 17850 7056
rect 17878 6033 17906 6039
rect 17878 6007 17879 6033
rect 17905 6007 17906 6033
rect 17878 5698 17906 6007
rect 17878 5665 17906 5670
rect 17990 5922 18018 5927
rect 17822 3761 17850 3766
rect 17878 4298 17906 4303
rect 17654 3649 17682 3654
rect 17486 3145 17514 3150
rect 17262 2753 17290 2758
rect 17206 2641 17234 2646
rect 17038 2305 17066 2310
rect 17374 2618 17402 2623
rect 17374 2282 17402 2590
rect 17878 2562 17906 4270
rect 17934 3794 17962 3799
rect 17934 3626 17962 3766
rect 17934 3593 17962 3598
rect 17990 3178 18018 5894
rect 18046 4522 18074 7056
rect 18270 6874 18298 7056
rect 18270 6841 18298 6846
rect 18270 6594 18298 6599
rect 18046 4489 18074 4494
rect 18214 5082 18242 5087
rect 17990 3145 18018 3150
rect 18046 4410 18074 4415
rect 18046 3066 18074 4382
rect 18214 3794 18242 5054
rect 18270 4410 18298 6566
rect 18494 6538 18522 7056
rect 18494 6510 18690 6538
rect 18550 6426 18578 6431
rect 18270 4377 18298 4382
rect 18326 5418 18354 5423
rect 18214 3761 18242 3766
rect 18270 4298 18298 4303
rect 18046 3033 18074 3038
rect 18158 3289 18186 3295
rect 18158 3263 18159 3289
rect 18185 3263 18186 3289
rect 18158 2842 18186 3263
rect 18158 2809 18186 2814
rect 17374 2249 17402 2254
rect 17822 2534 17906 2562
rect 18158 2618 18186 2623
rect 17094 1778 17122 1783
rect 17094 1610 17122 1750
rect 17094 1577 17122 1582
rect 17486 1666 17514 1671
rect 16646 1050 16674 1055
rect 16310 1049 16674 1050
rect 16310 1023 16647 1049
rect 16673 1023 16674 1049
rect 16310 1022 16674 1023
rect 16198 1003 16226 1022
rect 16422 993 16450 1022
rect 16646 1017 16674 1022
rect 17486 1050 17514 1638
rect 17486 1017 17514 1022
rect 17654 1162 17682 1167
rect 17654 1049 17682 1134
rect 17654 1023 17655 1049
rect 17681 1023 17682 1049
rect 17654 1017 17682 1023
rect 16422 967 16423 993
rect 16449 967 16450 993
rect 16422 961 16450 967
rect 17822 882 17850 2534
rect 18158 1330 18186 2590
rect 18158 1297 18186 1302
rect 18214 1946 18242 1951
rect 17822 849 17850 854
rect 17878 1162 17906 1167
rect 15358 457 15386 462
rect 17878 322 17906 1134
rect 18158 1106 18186 1111
rect 18158 1049 18186 1078
rect 18158 1023 18159 1049
rect 18185 1023 18186 1049
rect 18158 1017 18186 1023
rect 17934 993 17962 999
rect 17934 967 17935 993
rect 17961 967 17962 993
rect 17934 770 17962 967
rect 17934 737 17962 742
rect 18102 770 18130 775
rect 18102 657 18130 742
rect 18102 631 18103 657
rect 18129 631 18130 657
rect 18102 625 18130 631
rect 18214 378 18242 1918
rect 18270 1610 18298 4270
rect 18326 3010 18354 5390
rect 18494 5082 18522 5087
rect 18494 4410 18522 5054
rect 18382 4382 18522 4410
rect 18382 4074 18410 4382
rect 18550 4354 18578 6398
rect 18494 4326 18578 4354
rect 18382 4041 18410 4046
rect 18438 4186 18466 4191
rect 18382 3682 18410 3687
rect 18382 3234 18410 3654
rect 18438 3570 18466 4158
rect 18494 4074 18522 4326
rect 18662 4242 18690 6510
rect 18718 6090 18746 7056
rect 18718 6057 18746 6062
rect 18494 4041 18522 4046
rect 18550 4214 18690 4242
rect 18438 3537 18466 3542
rect 18438 3346 18466 3351
rect 18550 3346 18578 4214
rect 18438 3345 18578 3346
rect 18438 3319 18439 3345
rect 18465 3319 18551 3345
rect 18577 3319 18578 3345
rect 18438 3318 18578 3319
rect 18438 3313 18466 3318
rect 18550 3313 18578 3318
rect 18774 3290 18802 3295
rect 18942 3290 18970 7056
rect 19166 6314 19194 7056
rect 19390 6426 19418 7056
rect 19166 6281 19194 6286
rect 19278 6398 19418 6426
rect 19054 5922 19082 5927
rect 18802 3262 18970 3290
rect 18998 3402 19026 3407
rect 18774 3257 18802 3262
rect 18998 3234 19026 3374
rect 18382 3206 18746 3234
rect 18326 2977 18354 2982
rect 18494 2898 18522 2903
rect 18270 1577 18298 1582
rect 18326 2674 18354 2679
rect 18326 1330 18354 2646
rect 18382 2338 18410 2343
rect 18382 1610 18410 2310
rect 18494 1890 18522 2870
rect 18382 1577 18410 1582
rect 18438 1862 18522 1890
rect 18606 2674 18634 2679
rect 18326 1297 18354 1302
rect 18438 1218 18466 1862
rect 18494 1778 18522 1783
rect 18494 1498 18522 1750
rect 18494 1465 18522 1470
rect 18438 1185 18466 1190
rect 18270 1106 18298 1111
rect 18270 826 18298 1078
rect 18438 1106 18466 1111
rect 18606 1106 18634 2646
rect 18438 1105 18634 1106
rect 18438 1079 18439 1105
rect 18465 1079 18607 1105
rect 18633 1079 18634 1105
rect 18438 1078 18634 1079
rect 18438 1073 18466 1078
rect 18606 1073 18634 1078
rect 18662 2450 18690 2455
rect 18270 793 18298 798
rect 18662 602 18690 2422
rect 18662 569 18690 574
rect 18718 490 18746 3206
rect 18998 3201 19026 3206
rect 19054 3122 19082 5894
rect 19278 5530 19306 6398
rect 19614 5754 19642 7056
rect 19614 5721 19642 5726
rect 19670 6874 19698 6879
rect 19278 5497 19306 5502
rect 19334 5418 19362 5423
rect 19334 5026 19362 5390
rect 19334 4993 19362 4998
rect 19558 5138 19586 5143
rect 19390 4970 19418 4975
rect 19390 4690 19418 4942
rect 19390 4657 19418 4662
rect 19278 4354 19306 4359
rect 19278 4186 19306 4326
rect 19278 4153 19306 4158
rect 19222 3850 19250 3855
rect 19054 3089 19082 3094
rect 19166 3122 19194 3127
rect 19166 1890 19194 3094
rect 19222 2842 19250 3822
rect 19334 3850 19362 3855
rect 19278 3794 19306 3799
rect 19278 3234 19306 3766
rect 19278 3201 19306 3206
rect 19334 3122 19362 3822
rect 19222 2809 19250 2814
rect 19278 3094 19362 3122
rect 19166 1857 19194 1862
rect 19222 2450 19250 2455
rect 18886 1722 18914 1727
rect 18886 1274 18914 1694
rect 18886 1241 18914 1246
rect 19054 1106 19082 1111
rect 19222 1106 19250 2422
rect 19054 1105 19250 1106
rect 19054 1079 19055 1105
rect 19081 1079 19223 1105
rect 19249 1079 19250 1105
rect 19054 1078 19250 1079
rect 19054 1073 19082 1078
rect 19222 1073 19250 1078
rect 18774 938 18802 943
rect 18774 891 18802 910
rect 18718 457 18746 462
rect 18942 826 18970 831
rect 18214 345 18242 350
rect 17878 289 17906 294
rect 17486 266 17514 271
rect 13622 121 13650 126
rect 14574 154 14602 159
rect 14574 56 14602 126
rect 16030 98 16058 103
rect 16030 56 16058 70
rect 17486 56 17514 238
rect 18942 56 18970 798
rect 19278 658 19306 3094
rect 19278 625 19306 630
rect 19334 2730 19362 2735
rect 19334 546 19362 2702
rect 19558 2618 19586 5110
rect 19558 2585 19586 2590
rect 19446 994 19474 999
rect 19446 947 19474 966
rect 19670 770 19698 6846
rect 19838 5642 19866 7056
rect 19838 5609 19866 5614
rect 20006 5978 20034 5983
rect 20006 3570 20034 5950
rect 20062 4858 20090 7056
rect 20286 6146 20314 7056
rect 20286 6113 20314 6118
rect 20342 6650 20370 6655
rect 20286 6034 20314 6039
rect 20286 5987 20314 6006
rect 20342 5922 20370 6622
rect 20398 6034 20426 6039
rect 20398 5987 20426 6006
rect 20342 5894 20426 5922
rect 20062 4825 20090 4830
rect 20174 5642 20202 5647
rect 20174 3850 20202 5614
rect 20230 4578 20258 4583
rect 20230 4531 20258 4550
rect 20174 3817 20202 3822
rect 20006 3537 20034 3542
rect 19894 3458 19922 3463
rect 19894 2730 19922 3430
rect 20006 3458 20034 3463
rect 20006 2954 20034 3430
rect 20006 2921 20034 2926
rect 19894 2673 19922 2702
rect 19894 2647 19895 2673
rect 19921 2647 19922 2673
rect 19894 2641 19922 2647
rect 20174 2730 20202 2735
rect 20174 2673 20202 2702
rect 20174 2647 20175 2673
rect 20201 2647 20202 2673
rect 20174 2641 20202 2647
rect 20398 2506 20426 5894
rect 20510 5642 20538 7056
rect 20678 6090 20706 6095
rect 20678 6043 20706 6062
rect 20734 5922 20762 7056
rect 20846 6482 20874 6487
rect 20734 5889 20762 5894
rect 20790 6426 20818 6431
rect 20510 5609 20538 5614
rect 20790 5306 20818 6398
rect 20678 5278 20818 5306
rect 20454 4802 20482 4807
rect 20454 2617 20482 4774
rect 20622 4578 20650 4583
rect 20510 4550 20622 4578
rect 20510 4521 20538 4550
rect 20622 4531 20650 4550
rect 20510 4495 20511 4521
rect 20537 4495 20538 4521
rect 20510 4489 20538 4495
rect 20678 2674 20706 5278
rect 20678 2641 20706 2646
rect 20734 4690 20762 4695
rect 20454 2591 20455 2617
rect 20481 2591 20482 2617
rect 20454 2585 20482 2591
rect 20398 2473 20426 2478
rect 20510 2282 20538 2287
rect 20174 2058 20202 2063
rect 19894 2002 19922 2007
rect 19726 1106 19754 1111
rect 19894 1106 19922 1974
rect 20174 1721 20202 2030
rect 20174 1695 20175 1721
rect 20201 1695 20202 1721
rect 20174 1689 20202 1695
rect 20230 1890 20258 1895
rect 20230 1666 20258 1862
rect 20398 1890 20426 1895
rect 20510 1890 20538 2254
rect 20398 1889 20538 1890
rect 20398 1863 20399 1889
rect 20425 1863 20511 1889
rect 20537 1863 20538 1889
rect 20398 1862 20538 1863
rect 20398 1857 20426 1862
rect 20510 1857 20538 1862
rect 20230 1633 20258 1638
rect 20622 1834 20650 1839
rect 19726 1105 19922 1106
rect 19726 1079 19727 1105
rect 19753 1079 19895 1105
rect 19921 1079 19922 1105
rect 19726 1078 19922 1079
rect 19726 1073 19754 1078
rect 19894 1073 19922 1078
rect 20398 1330 20426 1335
rect 19838 938 19866 943
rect 19838 826 19866 910
rect 19838 793 19866 798
rect 19670 737 19698 742
rect 20174 714 20202 719
rect 20174 602 20202 686
rect 20174 569 20202 574
rect 19334 513 19362 518
rect 20398 56 20426 1302
rect 20622 1049 20650 1806
rect 20622 1023 20623 1049
rect 20649 1023 20650 1049
rect 20622 1017 20650 1023
rect 20734 882 20762 4662
rect 20846 4214 20874 6454
rect 20790 4186 20874 4214
rect 20902 4298 20930 4303
rect 20790 3290 20818 4186
rect 20902 3850 20930 4270
rect 20958 3962 20986 7056
rect 21070 6762 21098 6767
rect 21014 5194 21042 5199
rect 21014 4634 21042 5166
rect 21014 4601 21042 4606
rect 20958 3929 20986 3934
rect 21014 4018 21042 4023
rect 21014 3850 21042 3990
rect 20902 3817 20930 3822
rect 20958 3822 21042 3850
rect 20958 3794 20986 3822
rect 20958 3761 20986 3766
rect 21014 3738 21042 3743
rect 20790 3257 20818 3262
rect 20846 3681 20874 3687
rect 20846 3655 20847 3681
rect 20873 3655 20874 3681
rect 20846 2114 20874 3655
rect 20958 3346 20986 3351
rect 20958 2674 20986 3318
rect 20958 2641 20986 2646
rect 20902 2618 20930 2623
rect 20902 2571 20930 2590
rect 21014 2225 21042 3710
rect 21014 2199 21015 2225
rect 21041 2199 21042 2225
rect 21014 2193 21042 2199
rect 20846 2081 20874 2086
rect 21014 2114 21042 2119
rect 21014 1946 21042 2086
rect 21070 2002 21098 6734
rect 21126 5642 21154 5647
rect 21126 4018 21154 5614
rect 21126 3985 21154 3990
rect 21126 3794 21154 3799
rect 21126 3737 21154 3766
rect 21126 3711 21127 3737
rect 21153 3711 21154 3737
rect 21126 3705 21154 3711
rect 21182 3178 21210 7056
rect 21406 6818 21434 7056
rect 21630 6986 21658 7056
rect 21630 6953 21658 6958
rect 21350 6790 21434 6818
rect 21350 4214 21378 6790
rect 21854 6370 21882 7056
rect 22078 6874 22106 7056
rect 22078 6841 22106 6846
rect 22302 6762 22330 7056
rect 22302 6729 22330 6734
rect 22232 6678 22364 6683
rect 22260 6650 22284 6678
rect 22312 6650 22336 6678
rect 22232 6645 22364 6650
rect 22526 6426 22554 7056
rect 22526 6393 22554 6398
rect 22638 6930 22666 6935
rect 21854 6337 21882 6342
rect 21902 6286 22034 6291
rect 21930 6258 21954 6286
rect 21982 6258 22006 6286
rect 21902 6253 22034 6258
rect 21798 6034 21826 6039
rect 21798 5987 21826 6006
rect 21406 5978 21434 5983
rect 21406 5931 21434 5950
rect 21518 5978 21546 5983
rect 21518 5931 21546 5950
rect 22582 5922 22610 5927
rect 22232 5894 22364 5899
rect 22260 5866 22284 5894
rect 22312 5866 22336 5894
rect 22232 5861 22364 5866
rect 22414 5586 22442 5591
rect 21902 5502 22034 5507
rect 21930 5474 21954 5502
rect 21982 5474 22006 5502
rect 21902 5469 22034 5474
rect 21574 5305 21602 5311
rect 21574 5279 21575 5305
rect 21601 5279 21602 5305
rect 21406 5194 21434 5199
rect 21574 5194 21602 5279
rect 21798 5250 21826 5255
rect 21798 5203 21826 5222
rect 21406 5193 21602 5194
rect 21406 5167 21407 5193
rect 21433 5167 21602 5193
rect 21406 5166 21602 5167
rect 21406 5161 21434 5166
rect 21294 4186 21378 4214
rect 21238 3794 21266 3799
rect 21238 3747 21266 3766
rect 21294 3458 21322 4186
rect 21294 3425 21322 3430
rect 21182 3150 21266 3178
rect 21182 2730 21210 2735
rect 21182 2673 21210 2702
rect 21182 2647 21183 2673
rect 21209 2647 21210 2673
rect 21182 2641 21210 2647
rect 21070 1969 21098 1974
rect 21014 1913 21042 1918
rect 20790 1834 20818 1839
rect 20790 1162 20818 1806
rect 21070 1778 21098 1783
rect 20790 1129 20818 1134
rect 20902 1274 20930 1279
rect 20902 1106 20930 1246
rect 20902 1105 21042 1106
rect 20902 1079 20903 1105
rect 20929 1079 21042 1105
rect 20902 1078 21042 1079
rect 20902 1073 20930 1078
rect 20734 849 20762 854
rect 21014 658 21042 1078
rect 21070 1049 21098 1750
rect 21238 1106 21266 3150
rect 21462 3066 21490 3071
rect 21294 3010 21322 3015
rect 21294 2730 21322 2982
rect 21294 2697 21322 2702
rect 21350 2842 21378 2847
rect 21350 2674 21378 2814
rect 21462 2842 21490 3038
rect 21462 2809 21490 2814
rect 21462 2674 21490 2679
rect 21350 2673 21490 2674
rect 21350 2647 21351 2673
rect 21377 2647 21463 2673
rect 21489 2647 21490 2673
rect 21350 2646 21490 2647
rect 21350 2641 21378 2646
rect 21462 2641 21490 2646
rect 21406 2226 21434 2231
rect 21294 2198 21406 2226
rect 21294 2169 21322 2198
rect 21406 2179 21434 2198
rect 21294 2143 21295 2169
rect 21321 2143 21322 2169
rect 21294 2137 21322 2143
rect 21518 1610 21546 1615
rect 21238 1073 21266 1078
rect 21350 1106 21378 1111
rect 21350 1059 21378 1078
rect 21462 1106 21490 1111
rect 21070 1023 21071 1049
rect 21097 1023 21098 1049
rect 21070 1017 21098 1023
rect 21070 658 21098 663
rect 21014 657 21098 658
rect 21014 631 21071 657
rect 21097 631 21098 657
rect 21014 630 21098 631
rect 21462 658 21490 1078
rect 21518 1049 21546 1582
rect 21518 1023 21519 1049
rect 21545 1023 21546 1049
rect 21518 1017 21546 1023
rect 21518 658 21546 663
rect 21462 657 21546 658
rect 21462 631 21519 657
rect 21545 631 21546 657
rect 21462 630 21546 631
rect 21070 625 21098 630
rect 21518 625 21546 630
rect 21574 378 21602 5166
rect 22232 5110 22364 5115
rect 22260 5082 22284 5110
rect 22312 5082 22336 5110
rect 22232 5077 22364 5082
rect 22414 5082 22442 5558
rect 22414 5049 22442 5054
rect 21902 4718 22034 4723
rect 21930 4690 21954 4718
rect 21982 4690 22006 4718
rect 21902 4685 22034 4690
rect 22582 4578 22610 5894
rect 22582 4545 22610 4550
rect 22232 4326 22364 4331
rect 22260 4298 22284 4326
rect 22312 4298 22336 4326
rect 22232 4293 22364 4298
rect 22414 4298 22442 4303
rect 22414 4214 22442 4270
rect 21966 4186 21994 4191
rect 22078 4186 22442 4214
rect 21966 4185 22106 4186
rect 21966 4159 21967 4185
rect 21993 4159 22079 4185
rect 22105 4159 22106 4185
rect 21966 4158 22106 4159
rect 21966 4153 21994 4158
rect 22078 4153 22106 4158
rect 21742 4073 21770 4079
rect 21742 4047 21743 4073
rect 21769 4047 21770 4073
rect 21742 4018 21770 4047
rect 21742 3985 21770 3990
rect 21902 3934 22034 3939
rect 21930 3906 21954 3934
rect 21982 3906 22006 3934
rect 21902 3901 22034 3906
rect 22232 3542 22364 3547
rect 22260 3514 22284 3542
rect 22312 3514 22336 3542
rect 22232 3509 22364 3514
rect 21798 3206 22106 3234
rect 21798 3178 21826 3206
rect 22078 3178 22106 3206
rect 21798 3145 21826 3150
rect 21902 3150 22034 3155
rect 21930 3122 21954 3150
rect 21982 3122 22006 3150
rect 22078 3145 22106 3150
rect 21902 3117 22034 3122
rect 22638 3010 22666 6902
rect 22638 2977 22666 2982
rect 21854 2898 21882 2903
rect 21854 2842 21882 2870
rect 22134 2898 22162 2903
rect 22078 2842 22106 2847
rect 21854 2841 22106 2842
rect 21854 2815 21855 2841
rect 21881 2815 22079 2841
rect 22105 2815 22106 2841
rect 21854 2814 22106 2815
rect 21854 2809 21882 2814
rect 22078 2809 22106 2814
rect 21742 2562 21770 2567
rect 21742 2515 21770 2534
rect 21902 2366 22034 2371
rect 21930 2338 21954 2366
rect 21982 2338 22006 2366
rect 21902 2333 22034 2338
rect 22022 1834 22050 1839
rect 22022 1787 22050 1806
rect 21902 1582 22034 1587
rect 21930 1554 21954 1582
rect 21982 1554 22006 1582
rect 21902 1549 22034 1554
rect 21798 994 21826 999
rect 21798 947 21826 966
rect 21966 994 21994 999
rect 21966 947 21994 966
rect 21902 798 22034 803
rect 21930 770 21954 798
rect 21982 770 22006 798
rect 21902 765 22034 770
rect 22134 714 22162 2870
rect 22358 2898 22386 2903
rect 22358 2897 22442 2898
rect 22358 2871 22359 2897
rect 22385 2871 22442 2897
rect 22358 2870 22442 2871
rect 22358 2865 22386 2870
rect 22232 2758 22364 2763
rect 22260 2730 22284 2758
rect 22312 2730 22336 2758
rect 22232 2725 22364 2730
rect 22414 2562 22442 2870
rect 22414 2529 22442 2534
rect 22750 2450 22778 7056
rect 22974 5922 23002 7056
rect 22974 5889 23002 5894
rect 22750 2417 22778 2422
rect 22806 5754 22834 5759
rect 22694 2394 22722 2399
rect 22358 2338 22386 2343
rect 22358 2114 22386 2310
rect 22638 2170 22666 2175
rect 22358 2081 22386 2086
rect 22470 2114 22498 2119
rect 22232 1974 22364 1979
rect 22260 1946 22284 1974
rect 22312 1946 22336 1974
rect 22232 1941 22364 1946
rect 22190 1834 22218 1839
rect 22190 1787 22218 1806
rect 22470 1833 22498 2086
rect 22470 1807 22471 1833
rect 22497 1807 22498 1833
rect 22470 1801 22498 1807
rect 22638 1610 22666 2142
rect 22638 1577 22666 1582
rect 22694 1274 22722 2366
rect 22694 1241 22722 1246
rect 22232 1190 22364 1195
rect 22260 1162 22284 1190
rect 22312 1162 22336 1190
rect 22232 1157 22364 1162
rect 22694 938 22722 943
rect 22806 938 22834 5726
rect 23086 5754 23114 5759
rect 23086 5707 23114 5726
rect 23142 5026 23170 5031
rect 23142 3010 23170 4998
rect 23198 3794 23226 7056
rect 23254 6818 23282 6823
rect 23254 5642 23282 6790
rect 23254 5609 23282 5614
rect 23310 5922 23338 5927
rect 23310 5362 23338 5894
rect 23366 5697 23394 5703
rect 23366 5671 23367 5697
rect 23393 5671 23394 5697
rect 23366 5586 23394 5671
rect 23366 5553 23394 5558
rect 23310 5329 23338 5334
rect 23422 4214 23450 7056
rect 23646 6930 23674 7056
rect 23646 6897 23674 6902
rect 23478 5641 23506 5647
rect 23478 5615 23479 5641
rect 23505 5615 23506 5641
rect 23478 5586 23506 5615
rect 23478 5362 23506 5558
rect 23478 5329 23506 5334
rect 23198 3761 23226 3766
rect 23310 4186 23450 4214
rect 23646 5138 23674 5143
rect 23646 4186 23674 5110
rect 23702 4634 23730 4639
rect 23702 4578 23730 4606
rect 23702 4577 23842 4578
rect 23702 4551 23703 4577
rect 23729 4551 23842 4577
rect 23702 4550 23842 4551
rect 23702 4545 23730 4550
rect 23814 4521 23842 4550
rect 23814 4495 23815 4521
rect 23841 4495 23842 4521
rect 23814 4489 23842 4495
rect 23142 2977 23170 2982
rect 22694 937 22834 938
rect 22694 911 22695 937
rect 22721 911 22834 937
rect 22694 910 22834 911
rect 22862 2674 22890 2679
rect 22694 905 22722 910
rect 21574 345 21602 350
rect 21854 686 22162 714
rect 22694 714 22722 719
rect 21854 56 21882 686
rect 22694 434 22722 686
rect 22232 406 22364 411
rect 22260 378 22284 406
rect 22312 378 22336 406
rect 22694 401 22722 406
rect 22232 373 22364 378
rect 22862 378 22890 2646
rect 22974 2618 23002 2623
rect 22974 1274 23002 2590
rect 23254 2506 23282 2511
rect 23254 1833 23282 2478
rect 23310 2226 23338 4186
rect 23646 4153 23674 4158
rect 23478 3345 23506 3351
rect 23478 3319 23479 3345
rect 23505 3319 23506 3345
rect 23366 3290 23394 3295
rect 23478 3290 23506 3319
rect 23758 3346 23786 3351
rect 23758 3299 23786 3318
rect 23394 3262 23506 3290
rect 23366 3243 23394 3262
rect 23478 2842 23506 2847
rect 23310 2193 23338 2198
rect 23366 2730 23394 2735
rect 23254 1807 23255 1833
rect 23281 1807 23282 1833
rect 23254 1801 23282 1807
rect 22974 1241 23002 1246
rect 22918 1106 22946 1111
rect 22918 1059 22946 1078
rect 23086 1106 23114 1111
rect 23086 1059 23114 1078
rect 23366 1050 23394 2702
rect 23478 2002 23506 2814
rect 23478 1969 23506 1974
rect 23702 2226 23730 2231
rect 23534 1890 23562 1895
rect 23702 1890 23730 2198
rect 23534 1889 23730 1890
rect 23534 1863 23535 1889
rect 23561 1863 23703 1889
rect 23729 1863 23730 1889
rect 23534 1862 23730 1863
rect 23534 1857 23562 1862
rect 23702 1857 23730 1862
rect 23478 1778 23506 1783
rect 23478 1498 23506 1750
rect 23478 1465 23506 1470
rect 23366 1017 23394 1022
rect 23422 1218 23450 1223
rect 23422 546 23450 1190
rect 23870 1162 23898 7056
rect 24094 5642 24122 7056
rect 24318 5642 24346 7056
rect 24542 6650 24570 7056
rect 24038 5614 24122 5642
rect 24150 5614 24346 5642
rect 24486 6622 24570 6650
rect 24038 4214 24066 5614
rect 24094 5026 24122 5031
rect 24094 4577 24122 4998
rect 24094 4551 24095 4577
rect 24121 4551 24122 4577
rect 24094 4545 24122 4551
rect 23982 4186 24066 4214
rect 23982 2394 24010 4186
rect 23982 2361 24010 2366
rect 23870 1129 23898 1134
rect 24038 993 24066 999
rect 24038 967 24039 993
rect 24065 967 24066 993
rect 23422 513 23450 518
rect 23478 938 23506 943
rect 22862 345 22890 350
rect 23310 490 23338 495
rect 23310 56 23338 462
rect 23478 98 23506 910
rect 23758 938 23786 943
rect 24038 938 24066 967
rect 24150 994 24178 5614
rect 24262 5418 24290 5423
rect 24150 961 24178 966
rect 24206 4298 24234 4303
rect 23758 937 24066 938
rect 23758 911 23759 937
rect 23785 911 24066 937
rect 23758 910 24066 911
rect 23758 154 23786 910
rect 24206 490 24234 4270
rect 24262 3570 24290 5390
rect 24262 3537 24290 3542
rect 24318 5194 24346 5199
rect 24318 2450 24346 5166
rect 24318 2417 24346 2422
rect 24262 2113 24290 2119
rect 24262 2087 24263 2113
rect 24289 2087 24290 2113
rect 24262 1610 24290 2087
rect 24262 1577 24290 1582
rect 24318 1554 24346 1559
rect 24318 1049 24346 1526
rect 24486 1106 24514 6622
rect 24766 4214 24794 7056
rect 24542 4186 24794 4214
rect 24878 5082 24906 5087
rect 24542 2226 24570 4186
rect 24766 2282 24794 2287
rect 24654 2226 24682 2231
rect 24542 2225 24682 2226
rect 24542 2199 24655 2225
rect 24681 2199 24682 2225
rect 24542 2198 24682 2199
rect 24542 2169 24570 2198
rect 24654 2193 24682 2198
rect 24542 2143 24543 2169
rect 24569 2143 24570 2169
rect 24542 2137 24570 2143
rect 24486 1073 24514 1078
rect 24318 1023 24319 1049
rect 24345 1023 24346 1049
rect 24318 1017 24346 1023
rect 24598 993 24626 999
rect 24598 967 24599 993
rect 24625 967 24626 993
rect 24430 938 24458 943
rect 24430 891 24458 910
rect 24598 938 24626 967
rect 24598 905 24626 910
rect 24206 457 24234 462
rect 23758 121 23786 126
rect 23478 65 23506 70
rect 24766 56 24794 2254
rect 24878 1834 24906 5054
rect 24990 4214 25018 7056
rect 24934 4186 25018 4214
rect 25214 4214 25242 7056
rect 25438 6593 25466 7056
rect 25438 6567 25439 6593
rect 25465 6567 25466 6593
rect 25438 6561 25466 6567
rect 25662 6594 25690 7056
rect 25662 6561 25690 6566
rect 25606 6481 25634 6487
rect 25606 6455 25607 6481
rect 25633 6455 25634 6481
rect 25550 5362 25578 5367
rect 25214 4186 25298 4214
rect 24934 2226 24962 4186
rect 25214 3345 25242 3351
rect 25214 3319 25215 3345
rect 25241 3319 25242 3345
rect 25046 3290 25074 3295
rect 25214 3290 25242 3319
rect 25046 3289 25242 3290
rect 25046 3263 25047 3289
rect 25073 3263 25242 3289
rect 25046 3262 25242 3263
rect 25046 2898 25074 3262
rect 25046 2865 25074 2870
rect 24990 2562 25018 2567
rect 25158 2562 25186 2567
rect 24990 2561 25186 2562
rect 24990 2535 24991 2561
rect 25017 2535 25159 2561
rect 25185 2535 25186 2561
rect 24990 2534 25186 2535
rect 24990 2529 25018 2534
rect 24934 2193 24962 2198
rect 24990 1834 25018 1839
rect 24878 1833 25018 1834
rect 24878 1807 24991 1833
rect 25017 1807 25018 1833
rect 24878 1806 25018 1807
rect 24990 1801 25018 1806
rect 25046 1330 25074 2534
rect 25158 2529 25186 2534
rect 25270 1890 25298 4186
rect 25494 3346 25522 3351
rect 25494 3299 25522 3318
rect 25438 2618 25466 2623
rect 25438 2571 25466 2590
rect 25438 2394 25466 2399
rect 25382 1890 25410 1895
rect 25270 1889 25410 1890
rect 25270 1863 25271 1889
rect 25297 1863 25383 1889
rect 25409 1863 25410 1889
rect 25270 1862 25410 1863
rect 25270 1857 25298 1862
rect 25382 1857 25410 1862
rect 25046 1297 25074 1302
rect 24878 1050 24906 1055
rect 24878 1003 24906 1022
rect 25438 1049 25466 2366
rect 25438 1023 25439 1049
rect 25465 1023 25466 1049
rect 25438 1017 25466 1023
rect 25158 993 25186 999
rect 25158 967 25159 993
rect 25185 967 25186 993
rect 24990 938 25018 943
rect 25158 938 25186 967
rect 24990 937 25186 938
rect 24990 911 24991 937
rect 25017 911 25186 937
rect 24990 910 25186 911
rect 24878 826 24906 831
rect 24878 602 24906 798
rect 24878 569 24906 574
rect 24990 266 25018 910
rect 25550 546 25578 5334
rect 25606 1666 25634 6455
rect 25774 6481 25802 6487
rect 25774 6455 25775 6481
rect 25801 6455 25802 6481
rect 25774 5922 25802 6455
rect 25886 6202 25914 7056
rect 26054 6594 26082 6599
rect 26054 6547 26082 6566
rect 25886 6169 25914 6174
rect 26054 6482 26082 6487
rect 26054 6089 26082 6454
rect 26054 6063 26055 6089
rect 26081 6063 26082 6089
rect 26054 6057 26082 6063
rect 25774 5889 25802 5894
rect 26110 5810 26138 7056
rect 26334 6538 26362 7056
rect 26558 6762 26586 7056
rect 26558 6729 26586 6734
rect 26334 6505 26362 6510
rect 26558 6426 26586 6431
rect 26278 6202 26306 6207
rect 26278 6155 26306 6174
rect 26502 5810 26530 5815
rect 26110 5809 26530 5810
rect 26110 5783 26503 5809
rect 26529 5783 26530 5809
rect 26110 5782 26530 5783
rect 26502 5777 26530 5782
rect 26558 5754 26586 6398
rect 26558 5721 26586 5726
rect 26614 6370 26642 6375
rect 26782 6370 26810 7056
rect 26782 6342 26866 6370
rect 26222 5698 26250 5703
rect 26222 5651 26250 5670
rect 26054 5642 26082 5647
rect 25718 5362 25746 5367
rect 25718 5138 25746 5334
rect 25718 5105 25746 5110
rect 25998 4410 26026 4415
rect 25998 3850 26026 4382
rect 25998 3817 26026 3822
rect 25998 2338 26026 2343
rect 26054 2338 26082 5614
rect 26222 4522 26250 4527
rect 26222 4475 26250 4494
rect 26390 4522 26418 4527
rect 26390 4475 26418 4494
rect 26614 4214 26642 6342
rect 26670 6146 26698 6151
rect 26670 4578 26698 6118
rect 26782 6090 26810 6095
rect 26782 6043 26810 6062
rect 26838 5810 26866 6342
rect 27006 6202 27034 7056
rect 27230 6594 27258 7056
rect 27454 6874 27482 7056
rect 27454 6841 27482 6846
rect 27230 6561 27258 6566
rect 27454 6762 27482 6767
rect 27454 6593 27482 6734
rect 27454 6567 27455 6593
rect 27481 6567 27482 6593
rect 27454 6561 27482 6567
rect 27006 6169 27034 6174
rect 27062 6538 27090 6543
rect 27062 6201 27090 6510
rect 27062 6175 27063 6201
rect 27089 6175 27090 6201
rect 27062 6169 27090 6175
rect 27174 6481 27202 6487
rect 27174 6455 27175 6481
rect 27201 6455 27202 6481
rect 27174 6034 27202 6455
rect 27678 6482 27706 7056
rect 27902 6762 27930 7056
rect 27902 6729 27930 6734
rect 27958 6482 27986 6487
rect 27678 6449 27706 6454
rect 27902 6481 27986 6482
rect 27902 6455 27959 6481
rect 27985 6455 27986 6481
rect 27902 6454 27986 6455
rect 27846 6202 27874 6207
rect 27846 6155 27874 6174
rect 27174 6001 27202 6006
rect 27566 6033 27594 6039
rect 27566 6007 27567 6033
rect 27593 6007 27594 6033
rect 26838 5777 26866 5782
rect 27286 5810 27314 5815
rect 27286 5763 27314 5782
rect 27006 5697 27034 5703
rect 27006 5671 27007 5697
rect 27033 5671 27034 5697
rect 27006 5250 27034 5671
rect 27006 5217 27034 5222
rect 26670 4545 26698 4550
rect 27118 5026 27146 5031
rect 26670 4466 26698 4471
rect 26670 4419 26698 4438
rect 26446 4186 26642 4214
rect 26446 3346 26474 4186
rect 26446 3313 26474 3318
rect 27118 2618 27146 4998
rect 27118 2585 27146 2590
rect 26026 2310 26082 2338
rect 26334 2562 26362 2567
rect 25998 2305 26026 2310
rect 25606 1633 25634 1638
rect 26110 1778 26138 1783
rect 26054 1498 26082 1503
rect 26054 1441 26082 1470
rect 26054 1415 26055 1441
rect 26081 1415 26082 1441
rect 26054 1409 26082 1415
rect 26110 770 26138 1750
rect 26110 737 26138 742
rect 26166 1442 26194 1447
rect 26166 658 26194 1414
rect 26278 1274 26306 1279
rect 26278 1227 26306 1246
rect 26166 625 26194 630
rect 25550 513 25578 518
rect 24990 233 25018 238
rect 26222 490 26250 495
rect 26222 56 26250 462
rect 26334 434 26362 2534
rect 27566 2506 27594 6007
rect 27678 5530 27706 5535
rect 27678 5361 27706 5502
rect 27678 5335 27679 5361
rect 27705 5335 27706 5361
rect 27678 5329 27706 5335
rect 27734 4858 27762 4863
rect 27734 4811 27762 4830
rect 27734 4073 27762 4079
rect 27734 4047 27735 4073
rect 27761 4047 27762 4073
rect 27734 3962 27762 4047
rect 27734 3929 27762 3934
rect 27566 2473 27594 2478
rect 27846 2226 27874 2231
rect 27846 2179 27874 2198
rect 27902 2114 27930 6454
rect 27958 6449 27986 6454
rect 28126 6146 28154 7056
rect 28238 6594 28266 6599
rect 28238 6547 28266 6566
rect 28126 6113 28154 6118
rect 28238 6482 28266 6487
rect 28238 5809 28266 6454
rect 28350 6314 28378 7056
rect 28574 6538 28602 7056
rect 28574 6505 28602 6510
rect 28630 6874 28658 6879
rect 28350 6281 28378 6286
rect 28630 6201 28658 6846
rect 28630 6175 28631 6201
rect 28657 6175 28658 6201
rect 28630 6169 28658 6175
rect 28574 6146 28602 6151
rect 28350 6034 28378 6039
rect 28238 5783 28239 5809
rect 28265 5783 28266 5809
rect 28238 5777 28266 5783
rect 28294 6033 28378 6034
rect 28294 6007 28351 6033
rect 28377 6007 28378 6033
rect 28294 6006 28378 6007
rect 28014 5697 28042 5703
rect 28014 5671 28015 5697
rect 28041 5671 28042 5697
rect 27958 4913 27986 4919
rect 27958 4887 27959 4913
rect 27985 4887 27986 4913
rect 27958 4858 27986 4887
rect 27958 4825 27986 4830
rect 27958 4409 27986 4415
rect 27958 4383 27959 4409
rect 27985 4383 27986 4409
rect 27958 4354 27986 4383
rect 27958 4321 27986 4326
rect 27958 4129 27986 4135
rect 27958 4103 27959 4129
rect 27985 4103 27986 4129
rect 27958 3962 27986 4103
rect 27958 3929 27986 3934
rect 27902 2081 27930 2086
rect 26446 1274 26474 1279
rect 26446 1227 26474 1246
rect 28014 1050 28042 5671
rect 28070 5250 28098 5255
rect 28070 5203 28098 5222
rect 28238 5249 28266 5255
rect 28238 5223 28239 5249
rect 28265 5223 28266 5249
rect 28238 5082 28266 5223
rect 28238 5049 28266 5054
rect 28238 4857 28266 4863
rect 28238 4831 28239 4857
rect 28265 4831 28266 4857
rect 28238 4466 28266 4831
rect 28238 4433 28266 4438
rect 28126 4409 28154 4415
rect 28126 4383 28127 4409
rect 28153 4383 28154 4409
rect 28126 4354 28154 4383
rect 28126 4321 28154 4326
rect 28238 4186 28266 4191
rect 28238 4139 28266 4158
rect 28294 2954 28322 6006
rect 28350 6001 28378 6006
rect 28462 5474 28490 5479
rect 28406 4857 28434 4863
rect 28406 4831 28407 4857
rect 28433 4831 28434 4857
rect 28350 4578 28378 4583
rect 28350 4531 28378 4550
rect 28406 4410 28434 4831
rect 28406 4377 28434 4382
rect 28462 4129 28490 5446
rect 28574 5361 28602 6118
rect 28798 6146 28826 7056
rect 29022 6482 29050 7056
rect 29022 6449 29050 6454
rect 29078 6481 29106 6487
rect 29078 6455 29079 6481
rect 29105 6455 29106 6481
rect 28798 6113 28826 6118
rect 29022 6314 29050 6319
rect 29022 5809 29050 6286
rect 29022 5783 29023 5809
rect 29049 5783 29050 5809
rect 29022 5777 29050 5783
rect 28574 5335 28575 5361
rect 28601 5335 28602 5361
rect 28574 5329 28602 5335
rect 28630 5698 28658 5703
rect 28574 4410 28602 4415
rect 28574 4363 28602 4382
rect 28462 4103 28463 4129
rect 28489 4103 28490 4129
rect 28350 3794 28378 3799
rect 28462 3794 28490 4103
rect 28630 4018 28658 5670
rect 28742 5697 28770 5703
rect 28742 5671 28743 5697
rect 28769 5671 28770 5697
rect 28742 5026 28770 5671
rect 29022 5306 29050 5311
rect 29022 5259 29050 5278
rect 29078 5194 29106 6455
rect 29246 6258 29274 7056
rect 29414 6762 29442 6767
rect 29414 6425 29442 6734
rect 29470 6594 29498 7056
rect 29470 6561 29498 6566
rect 29414 6399 29415 6425
rect 29441 6399 29442 6425
rect 29414 6393 29442 6399
rect 29246 6225 29274 6230
rect 29414 6146 29442 6151
rect 29134 5978 29162 5983
rect 29302 5978 29330 5983
rect 29134 5977 29330 5978
rect 29134 5951 29135 5977
rect 29161 5951 29303 5977
rect 29329 5951 29330 5977
rect 29134 5950 29330 5951
rect 29134 5866 29162 5950
rect 29302 5945 29330 5950
rect 29134 5833 29162 5838
rect 29414 5361 29442 6118
rect 29694 6146 29722 7056
rect 29862 6481 29890 6487
rect 29862 6455 29863 6481
rect 29889 6455 29890 6481
rect 29806 6370 29834 6375
rect 29862 6370 29890 6455
rect 29834 6342 29890 6370
rect 29918 6370 29946 7056
rect 30422 6986 30450 6991
rect 30254 6538 30282 6543
rect 30254 6491 30282 6510
rect 29806 6337 29834 6342
rect 29918 6337 29946 6342
rect 30310 6482 30338 6487
rect 29694 6113 29722 6118
rect 29806 6258 29834 6263
rect 29582 6033 29610 6039
rect 29582 6007 29583 6033
rect 29609 6007 29610 6033
rect 29526 5698 29554 5703
rect 29526 5651 29554 5670
rect 29414 5335 29415 5361
rect 29441 5335 29442 5361
rect 29414 5329 29442 5335
rect 29470 5418 29498 5423
rect 28742 4993 28770 4998
rect 29022 5166 29106 5194
rect 28686 4914 28714 4919
rect 28686 4913 28826 4914
rect 28686 4887 28687 4913
rect 28713 4887 28826 4913
rect 28686 4886 28826 4887
rect 28686 4881 28714 4886
rect 28798 4577 28826 4886
rect 28966 4858 28994 4863
rect 28966 4811 28994 4830
rect 28798 4551 28799 4577
rect 28825 4551 28826 4577
rect 28798 4545 28826 4551
rect 28742 4130 28770 4135
rect 28742 4083 28770 4102
rect 28910 4129 28938 4135
rect 28910 4103 28911 4129
rect 28937 4103 28938 4129
rect 28630 3985 28658 3990
rect 28350 3793 28490 3794
rect 28350 3767 28351 3793
rect 28377 3767 28490 3793
rect 28350 3766 28490 3767
rect 28350 3761 28378 3766
rect 28798 3738 28826 3743
rect 28910 3738 28938 4103
rect 28826 3710 28938 3738
rect 28798 3691 28826 3710
rect 28630 3626 28658 3631
rect 28630 3579 28658 3598
rect 28910 3626 28938 3631
rect 28910 3579 28938 3598
rect 28238 2926 28322 2954
rect 28742 3514 28770 3519
rect 28182 2562 28210 2567
rect 28182 2515 28210 2534
rect 28238 2170 28266 2926
rect 28182 2142 28266 2170
rect 28294 2842 28322 2847
rect 28070 2058 28098 2063
rect 28070 2011 28098 2030
rect 28182 1722 28210 2142
rect 28238 2058 28266 2063
rect 28238 2011 28266 2030
rect 28182 1689 28210 1694
rect 28014 1017 28042 1022
rect 28294 714 28322 2814
rect 28518 2842 28546 2847
rect 28518 2795 28546 2814
rect 28686 2842 28714 2847
rect 28686 2795 28714 2814
rect 28742 2674 28770 3486
rect 29022 3402 29050 5166
rect 29078 5026 29106 5031
rect 29078 3514 29106 4998
rect 29414 4914 29442 4919
rect 29414 4867 29442 4886
rect 29358 4802 29386 4807
rect 29358 4633 29386 4774
rect 29358 4607 29359 4633
rect 29385 4607 29386 4633
rect 29358 4601 29386 4607
rect 29134 4242 29162 4247
rect 29134 3793 29162 4214
rect 29190 4130 29218 4135
rect 29358 4130 29386 4135
rect 29190 4129 29386 4130
rect 29190 4103 29191 4129
rect 29217 4103 29359 4129
rect 29385 4103 29386 4129
rect 29190 4102 29386 4103
rect 29190 4097 29218 4102
rect 29358 4097 29386 4102
rect 29134 3767 29135 3793
rect 29161 3767 29162 3793
rect 29134 3761 29162 3767
rect 29414 3737 29442 3743
rect 29414 3711 29415 3737
rect 29441 3711 29442 3737
rect 29078 3481 29106 3486
rect 29134 3570 29162 3575
rect 29022 3374 29106 3402
rect 28910 3289 28938 3295
rect 28910 3263 28911 3289
rect 28937 3263 28938 3289
rect 28910 3234 28938 3263
rect 28910 3201 28938 3206
rect 28966 3290 28994 3295
rect 28966 3009 28994 3262
rect 29022 3289 29050 3295
rect 29022 3263 29023 3289
rect 29049 3263 29050 3289
rect 29022 3178 29050 3263
rect 29022 3145 29050 3150
rect 28966 2983 28967 3009
rect 28993 2983 28994 3009
rect 28966 2977 28994 2983
rect 28686 2646 28770 2674
rect 28350 2562 28378 2567
rect 28350 2515 28378 2534
rect 28630 2562 28658 2567
rect 28630 2515 28658 2534
rect 28686 1498 28714 2646
rect 28742 2562 28770 2567
rect 28910 2562 28938 2567
rect 28742 2561 28938 2562
rect 28742 2535 28743 2561
rect 28769 2535 28911 2561
rect 28937 2535 28938 2561
rect 28742 2534 28938 2535
rect 28742 2450 28770 2534
rect 28910 2529 28938 2534
rect 28742 2417 28770 2422
rect 29078 2394 29106 3374
rect 29134 3345 29162 3542
rect 29414 3570 29442 3711
rect 29414 3537 29442 3542
rect 29302 3458 29330 3463
rect 29134 3319 29135 3345
rect 29161 3319 29162 3345
rect 29134 3313 29162 3319
rect 29246 3345 29274 3351
rect 29246 3319 29247 3345
rect 29273 3319 29274 3345
rect 29246 3178 29274 3319
rect 29246 3145 29274 3150
rect 29134 3010 29162 3015
rect 29134 2506 29162 2982
rect 29302 2954 29330 3430
rect 29470 3289 29498 5390
rect 29526 5250 29554 5255
rect 29526 4214 29554 5222
rect 29582 4521 29610 6007
rect 29806 5809 29834 6230
rect 30310 6145 30338 6454
rect 30310 6119 30311 6145
rect 30337 6119 30338 6145
rect 30310 6113 30338 6119
rect 29806 5783 29807 5809
rect 29833 5783 29834 5809
rect 29806 5777 29834 5783
rect 29918 6033 29946 6039
rect 29918 6007 29919 6033
rect 29945 6007 29946 6033
rect 29862 4858 29890 4863
rect 29862 4811 29890 4830
rect 29582 4495 29583 4521
rect 29609 4495 29610 4521
rect 29582 4489 29610 4495
rect 29526 4186 29610 4214
rect 29582 3793 29610 4186
rect 29862 4130 29890 4135
rect 29862 4073 29890 4102
rect 29862 4047 29863 4073
rect 29889 4047 29890 4073
rect 29862 4041 29890 4047
rect 29582 3767 29583 3793
rect 29609 3767 29610 3793
rect 29582 3761 29610 3767
rect 29470 3263 29471 3289
rect 29497 3263 29498 3289
rect 29470 3257 29498 3263
rect 29694 3345 29722 3351
rect 29694 3319 29695 3345
rect 29721 3319 29722 3345
rect 29694 3234 29722 3319
rect 29694 3201 29722 3206
rect 29638 3010 29666 3015
rect 29638 2963 29666 2982
rect 29302 2921 29330 2926
rect 29190 2842 29218 2847
rect 29358 2842 29386 2847
rect 29190 2841 29386 2842
rect 29190 2815 29191 2841
rect 29217 2815 29359 2841
rect 29385 2815 29386 2841
rect 29190 2814 29386 2815
rect 29190 2730 29218 2814
rect 29358 2809 29386 2814
rect 29190 2697 29218 2702
rect 29190 2618 29218 2623
rect 29190 2571 29218 2590
rect 29134 2473 29162 2478
rect 29582 2562 29610 2567
rect 29694 2562 29722 2567
rect 29582 2561 29722 2562
rect 29582 2535 29583 2561
rect 29609 2535 29695 2561
rect 29721 2535 29722 2561
rect 29582 2534 29722 2535
rect 29078 2361 29106 2366
rect 29526 1890 29554 1895
rect 29526 1843 29554 1862
rect 29582 1778 29610 2534
rect 29694 2529 29722 2534
rect 29918 1946 29946 6007
rect 30366 5697 30394 5703
rect 30366 5671 30367 5697
rect 30393 5671 30394 5697
rect 30310 5305 30338 5311
rect 30310 5279 30311 5305
rect 30337 5279 30338 5305
rect 30142 4970 30170 4975
rect 30142 4923 30170 4942
rect 30142 4466 30170 4471
rect 30142 4185 30170 4438
rect 30142 4159 30143 4185
rect 30169 4159 30170 4185
rect 30142 4153 30170 4159
rect 30254 4465 30282 4471
rect 30254 4439 30255 4465
rect 30281 4439 30282 4465
rect 30254 4186 30282 4439
rect 30254 4153 30282 4158
rect 30254 3682 30282 3687
rect 30254 3635 30282 3654
rect 30254 3402 30282 3407
rect 29974 3346 30002 3351
rect 29974 3299 30002 3318
rect 30142 3345 30170 3351
rect 30142 3319 30143 3345
rect 30169 3319 30170 3345
rect 30142 3122 30170 3319
rect 30142 3089 30170 3094
rect 30254 2953 30282 3374
rect 30310 3290 30338 5279
rect 30310 3257 30338 3262
rect 30254 2927 30255 2953
rect 30281 2927 30282 2953
rect 30254 2921 30282 2927
rect 30142 2618 30170 2623
rect 30142 2571 30170 2590
rect 29974 2562 30002 2567
rect 29974 2515 30002 2534
rect 30366 2226 30394 5671
rect 30422 5530 30450 6958
rect 32102 6762 32130 6767
rect 31262 6594 31290 6599
rect 31262 6547 31290 6566
rect 31542 6538 31570 6543
rect 30982 6481 31010 6487
rect 30982 6455 30983 6481
rect 31009 6455 31010 6481
rect 30982 6426 31010 6455
rect 30982 6393 31010 6398
rect 30590 6370 30618 6375
rect 30590 5809 30618 6342
rect 31094 6146 31122 6151
rect 31094 6099 31122 6118
rect 30590 5783 30591 5809
rect 30617 5783 30618 5809
rect 30590 5777 30618 5783
rect 30702 6033 30730 6039
rect 30702 6007 30703 6033
rect 30729 6007 30730 6033
rect 30422 5497 30450 5502
rect 30702 5026 30730 6007
rect 31206 5866 31234 5871
rect 31094 5641 31122 5647
rect 31094 5615 31095 5641
rect 31121 5615 31122 5641
rect 30758 5361 30786 5367
rect 30758 5335 30759 5361
rect 30785 5335 30786 5361
rect 30758 5082 30786 5335
rect 30758 5049 30786 5054
rect 30702 4993 30730 4998
rect 30534 4970 30562 4975
rect 30534 4923 30562 4942
rect 30982 4913 31010 4919
rect 30982 4887 30983 4913
rect 31009 4887 31010 4913
rect 30758 4634 30786 4639
rect 30758 4587 30786 4606
rect 30534 4186 30562 4191
rect 30534 4139 30562 4158
rect 30926 4130 30954 4135
rect 30870 4129 30954 4130
rect 30870 4103 30927 4129
rect 30953 4103 30954 4129
rect 30870 4102 30954 4103
rect 30758 3793 30786 3799
rect 30758 3767 30759 3793
rect 30785 3767 30786 3793
rect 30758 3402 30786 3767
rect 30758 3369 30786 3374
rect 30646 3233 30674 3239
rect 30646 3207 30647 3233
rect 30673 3207 30674 3233
rect 30646 2954 30674 3207
rect 30758 3066 30786 3071
rect 30758 3019 30786 3038
rect 30870 3010 30898 4102
rect 30926 4097 30954 4102
rect 30926 3458 30954 3463
rect 30926 3401 30954 3430
rect 30926 3375 30927 3401
rect 30953 3375 30954 3401
rect 30926 3369 30954 3375
rect 30982 3346 31010 4887
rect 31094 4521 31122 5615
rect 31150 5362 31178 5367
rect 31150 5305 31178 5334
rect 31150 5279 31151 5305
rect 31177 5279 31178 5305
rect 31150 5273 31178 5279
rect 31150 5194 31178 5199
rect 31150 4970 31178 5166
rect 31150 4937 31178 4942
rect 31094 4495 31095 4521
rect 31121 4495 31122 4521
rect 31094 4489 31122 4495
rect 31206 4186 31234 5838
rect 31318 5697 31346 5703
rect 31318 5671 31319 5697
rect 31345 5671 31346 5697
rect 31318 5642 31346 5671
rect 31318 5609 31346 5614
rect 31486 5642 31514 5647
rect 31486 5595 31514 5614
rect 31318 5418 31346 5423
rect 31318 4634 31346 5390
rect 31430 5249 31458 5255
rect 31430 5223 31431 5249
rect 31457 5223 31458 5249
rect 31318 4601 31346 4606
rect 31374 4857 31402 4863
rect 31374 4831 31375 4857
rect 31401 4831 31402 4857
rect 31374 4522 31402 4831
rect 31430 4746 31458 5223
rect 31542 4914 31570 6510
rect 31822 6314 31850 6319
rect 31710 6090 31738 6095
rect 31542 4881 31570 4886
rect 31598 5642 31626 5647
rect 31598 4858 31626 5614
rect 31598 4825 31626 4830
rect 31710 4802 31738 6062
rect 31710 4769 31738 4774
rect 31430 4713 31458 4718
rect 31374 4489 31402 4494
rect 31430 4465 31458 4471
rect 31430 4439 31431 4465
rect 31457 4439 31458 4465
rect 31430 4298 31458 4439
rect 31430 4265 31458 4270
rect 31206 4153 31234 4158
rect 31822 4130 31850 6286
rect 31822 4097 31850 4102
rect 31542 4074 31570 4079
rect 31430 4017 31458 4023
rect 31430 3991 31431 4017
rect 31457 3991 31458 4017
rect 31430 3850 31458 3991
rect 31430 3817 31458 3822
rect 31542 3849 31570 4046
rect 31542 3823 31543 3849
rect 31569 3823 31570 3849
rect 31542 3817 31570 3823
rect 31150 3738 31178 3743
rect 31150 3737 31234 3738
rect 31150 3711 31151 3737
rect 31177 3711 31234 3737
rect 31150 3710 31234 3711
rect 31150 3705 31178 3710
rect 30982 3313 31010 3318
rect 30870 2977 30898 2982
rect 30646 2921 30674 2926
rect 31094 2953 31122 2959
rect 31094 2927 31095 2953
rect 31121 2927 31122 2953
rect 30534 2618 30562 2623
rect 30534 2571 30562 2590
rect 30926 2562 30954 2567
rect 30926 2515 30954 2534
rect 31094 2506 31122 2927
rect 31094 2473 31122 2478
rect 31150 2674 31178 2679
rect 30366 2193 30394 2198
rect 29918 1913 29946 1918
rect 30310 2169 30338 2175
rect 30310 2143 30311 2169
rect 30337 2143 30338 2169
rect 29694 1890 29722 1895
rect 29694 1843 29722 1862
rect 29526 1750 29610 1778
rect 29974 1778 30002 1783
rect 30142 1778 30170 1783
rect 29974 1777 30170 1778
rect 29974 1751 29975 1777
rect 30001 1751 30143 1777
rect 30169 1751 30170 1777
rect 29974 1750 30170 1751
rect 28686 1465 28714 1470
rect 29246 1721 29274 1727
rect 29246 1695 29247 1721
rect 29273 1695 29274 1721
rect 29246 1386 29274 1695
rect 29246 1353 29274 1358
rect 29414 1386 29442 1391
rect 29414 1339 29442 1358
rect 29190 1330 29218 1335
rect 29190 1283 29218 1302
rect 28798 1274 28826 1279
rect 28910 1274 28938 1279
rect 28798 1273 28938 1274
rect 28798 1247 28799 1273
rect 28825 1247 28911 1273
rect 28937 1247 28938 1273
rect 28798 1246 28938 1247
rect 28798 1218 28826 1246
rect 28910 1241 28938 1246
rect 29134 1274 29162 1279
rect 28798 1185 28826 1190
rect 28798 1050 28826 1055
rect 28798 1003 28826 1022
rect 28518 993 28546 999
rect 28518 967 28519 993
rect 28545 967 28546 993
rect 28294 681 28322 686
rect 28350 938 28378 943
rect 28518 938 28546 967
rect 28350 937 28546 938
rect 28350 911 28351 937
rect 28377 911 28546 937
rect 28350 910 28546 911
rect 28966 993 28994 999
rect 28966 967 28967 993
rect 28993 967 28994 993
rect 26334 401 26362 406
rect 27678 546 27706 551
rect 27678 56 27706 518
rect 28350 378 28378 910
rect 28854 770 28882 775
rect 28966 770 28994 967
rect 28882 742 28994 770
rect 28854 657 28882 742
rect 28854 631 28855 657
rect 28881 631 28882 657
rect 28854 625 28882 631
rect 28350 345 28378 350
rect 29134 56 29162 1246
rect 29246 1106 29274 1111
rect 29246 1049 29274 1078
rect 29246 1023 29247 1049
rect 29273 1023 29274 1049
rect 29246 1017 29274 1023
rect 29302 658 29330 663
rect 29302 601 29330 630
rect 29302 575 29303 601
rect 29329 575 29330 601
rect 29302 569 29330 575
rect 29526 322 29554 1750
rect 29974 1745 30002 1750
rect 30142 1745 30170 1750
rect 29638 1386 29666 1391
rect 29638 1339 29666 1358
rect 30086 1330 30114 1335
rect 29694 993 29722 999
rect 29694 967 29695 993
rect 29721 967 29722 993
rect 29582 938 29610 943
rect 29694 938 29722 967
rect 29974 994 30002 999
rect 29974 947 30002 966
rect 29582 937 29722 938
rect 29582 911 29583 937
rect 29609 911 29722 937
rect 29582 910 29722 911
rect 29582 826 29610 910
rect 29582 793 29610 798
rect 29526 289 29554 294
rect 29806 657 29834 663
rect 29806 631 29807 657
rect 29833 631 29834 657
rect 29806 266 29834 631
rect 30086 601 30114 1302
rect 30254 1329 30282 1335
rect 30254 1303 30255 1329
rect 30281 1303 30282 1329
rect 30142 1050 30170 1055
rect 30142 1003 30170 1022
rect 30086 575 30087 601
rect 30113 575 30114 601
rect 30086 569 30114 575
rect 30254 602 30282 1303
rect 30310 1106 30338 2143
rect 31150 2169 31178 2646
rect 31150 2143 31151 2169
rect 31177 2143 31178 2169
rect 31150 2137 31178 2143
rect 30646 2113 30674 2119
rect 30646 2087 30647 2113
rect 30673 2087 30674 2113
rect 30310 1073 30338 1078
rect 30534 2058 30562 2063
rect 30254 569 30282 574
rect 30534 378 30562 2030
rect 30646 1834 30674 2087
rect 30646 1801 30674 1806
rect 30926 2002 30954 2007
rect 30926 1833 30954 1974
rect 30926 1807 30927 1833
rect 30953 1807 30954 1833
rect 30926 1801 30954 1807
rect 30646 1722 30674 1727
rect 30646 1675 30674 1694
rect 31206 1554 31234 3710
rect 31430 3626 31458 3631
rect 31430 3289 31458 3598
rect 31430 3263 31431 3289
rect 31457 3263 31458 3289
rect 31430 3257 31458 3263
rect 31542 3178 31570 3183
rect 31542 3065 31570 3150
rect 31542 3039 31543 3065
rect 31569 3039 31570 3065
rect 31542 3033 31570 3039
rect 32102 3066 32130 6734
rect 32102 3033 32130 3038
rect 31318 2730 31346 2735
rect 31262 2618 31290 2623
rect 31262 2282 31290 2590
rect 31318 2617 31346 2702
rect 31318 2591 31319 2617
rect 31345 2591 31346 2617
rect 31318 2585 31346 2591
rect 31262 2249 31290 2254
rect 31542 2506 31570 2511
rect 31542 2281 31570 2478
rect 31542 2255 31543 2281
rect 31569 2255 31570 2281
rect 31542 2249 31570 2255
rect 31430 2058 31458 2063
rect 31206 1521 31234 1526
rect 31318 1722 31346 1727
rect 31094 1386 31122 1391
rect 31094 1339 31122 1358
rect 31318 1386 31346 1694
rect 31430 1721 31458 2030
rect 31430 1695 31431 1721
rect 31457 1695 31458 1721
rect 31430 1689 31458 1695
rect 31542 1610 31570 1615
rect 31542 1497 31570 1582
rect 31542 1471 31543 1497
rect 31569 1471 31570 1497
rect 31542 1465 31570 1471
rect 31318 1353 31346 1358
rect 30646 1330 30674 1335
rect 30646 1283 30674 1302
rect 31374 1330 31402 1335
rect 30926 994 30954 999
rect 30926 947 30954 966
rect 30646 882 30674 887
rect 30646 835 30674 854
rect 30590 657 30618 663
rect 30590 631 30591 657
rect 30617 631 30618 657
rect 30590 490 30618 631
rect 30590 457 30618 462
rect 31094 601 31122 607
rect 31094 575 31095 601
rect 31121 575 31122 601
rect 30534 350 30618 378
rect 29806 233 29834 238
rect 30590 56 30618 350
rect 31094 210 31122 575
rect 31094 177 31122 182
rect 4774 9 4802 14
rect 5824 0 5880 56
rect 7280 0 7336 56
rect 8736 0 8792 56
rect 10192 0 10248 56
rect 11648 0 11704 56
rect 13104 0 13160 56
rect 14560 0 14616 56
rect 16016 0 16072 56
rect 17472 0 17528 56
rect 18928 0 18984 56
rect 20384 0 20440 56
rect 21840 0 21896 56
rect 23296 0 23352 56
rect 24752 0 24808 56
rect 26208 0 26264 56
rect 27664 0 27720 56
rect 29120 0 29176 56
rect 30576 0 30632 56
rect 31374 42 31402 1302
rect 31430 1162 31458 1167
rect 31430 937 31458 1134
rect 31430 911 31431 937
rect 31457 911 31458 937
rect 31430 905 31458 911
rect 31542 938 31570 943
rect 31542 713 31570 910
rect 31542 687 31543 713
rect 31569 687 31570 713
rect 31542 681 31570 687
rect 31374 9 31402 14
<< via2 >>
rect 126 6958 154 6986
rect 1862 6790 1890 6818
rect 1806 6734 1834 6762
rect 1246 6566 1274 6594
rect 126 4102 154 4130
rect 182 6286 210 6314
rect 798 6062 826 6090
rect 798 5726 826 5754
rect 1078 6398 1106 6426
rect 966 5641 994 5642
rect 966 5615 967 5641
rect 967 5615 993 5641
rect 993 5615 994 5641
rect 966 5614 994 5615
rect 182 3710 210 3738
rect 462 4046 490 4074
rect 966 2897 994 2898
rect 966 2871 967 2897
rect 967 2871 993 2897
rect 993 2871 994 2897
rect 966 2870 994 2871
rect 910 2590 938 2618
rect 2086 6678 2114 6706
rect 1902 6285 1930 6286
rect 1902 6259 1903 6285
rect 1903 6259 1929 6285
rect 1929 6259 1930 6285
rect 1902 6258 1930 6259
rect 1954 6285 1982 6286
rect 1954 6259 1955 6285
rect 1955 6259 1981 6285
rect 1981 6259 1982 6285
rect 1954 6258 1982 6259
rect 2006 6285 2034 6286
rect 2006 6259 2007 6285
rect 2007 6259 2033 6285
rect 2033 6259 2034 6285
rect 2006 6258 2034 6259
rect 1246 5390 1274 5418
rect 1902 5501 1930 5502
rect 1902 5475 1903 5501
rect 1903 5475 1929 5501
rect 1929 5475 1930 5501
rect 1902 5474 1930 5475
rect 1954 5501 1982 5502
rect 1954 5475 1955 5501
rect 1955 5475 1981 5501
rect 1981 5475 1982 5501
rect 1954 5474 1982 5475
rect 2006 5501 2034 5502
rect 2006 5475 2007 5501
rect 2007 5475 2033 5501
rect 2033 5475 2034 5501
rect 2006 5474 2034 5475
rect 1358 5390 1386 5418
rect 1902 4717 1930 4718
rect 1902 4691 1903 4717
rect 1903 4691 1929 4717
rect 1929 4691 1930 4717
rect 1902 4690 1930 4691
rect 1954 4717 1982 4718
rect 1954 4691 1955 4717
rect 1955 4691 1981 4717
rect 1981 4691 1982 4717
rect 1954 4690 1982 4691
rect 2006 4717 2034 4718
rect 2006 4691 2007 4717
rect 2007 4691 2033 4717
rect 2033 4691 2034 4717
rect 2006 4690 2034 4691
rect 1414 4577 1442 4578
rect 1414 4551 1415 4577
rect 1415 4551 1441 4577
rect 1441 4551 1442 4577
rect 1414 4550 1442 4551
rect 1638 4409 1666 4410
rect 1638 4383 1639 4409
rect 1639 4383 1665 4409
rect 1665 4383 1666 4409
rect 1638 4382 1666 4383
rect 1750 4409 1778 4410
rect 1750 4383 1751 4409
rect 1751 4383 1777 4409
rect 1777 4383 1778 4409
rect 1750 4382 1778 4383
rect 2366 6734 2394 6762
rect 2232 6677 2260 6678
rect 2232 6651 2233 6677
rect 2233 6651 2259 6677
rect 2259 6651 2260 6677
rect 2232 6650 2260 6651
rect 2284 6677 2312 6678
rect 2284 6651 2285 6677
rect 2285 6651 2311 6677
rect 2311 6651 2312 6677
rect 2284 6650 2312 6651
rect 2336 6677 2364 6678
rect 2336 6651 2337 6677
rect 2337 6651 2363 6677
rect 2363 6651 2364 6677
rect 2336 6650 2364 6651
rect 2142 6566 2170 6594
rect 2198 5950 2226 5978
rect 2534 6006 2562 6034
rect 2232 5893 2260 5894
rect 2232 5867 2233 5893
rect 2233 5867 2259 5893
rect 2259 5867 2260 5893
rect 2232 5866 2260 5867
rect 2284 5893 2312 5894
rect 2284 5867 2285 5893
rect 2285 5867 2311 5893
rect 2311 5867 2312 5893
rect 2284 5866 2312 5867
rect 2336 5893 2364 5894
rect 2336 5867 2337 5893
rect 2337 5867 2363 5893
rect 2363 5867 2364 5893
rect 2336 5866 2364 5867
rect 2310 5809 2338 5810
rect 2310 5783 2311 5809
rect 2311 5783 2337 5809
rect 2337 5783 2338 5809
rect 2310 5782 2338 5783
rect 2814 6790 2842 6818
rect 2982 6622 3010 6650
rect 2590 5782 2618 5810
rect 2142 5558 2170 5586
rect 2478 5670 2506 5698
rect 2198 5502 2226 5530
rect 2232 5109 2260 5110
rect 2232 5083 2233 5109
rect 2233 5083 2259 5109
rect 2259 5083 2260 5109
rect 2232 5082 2260 5083
rect 2284 5109 2312 5110
rect 2284 5083 2285 5109
rect 2285 5083 2311 5109
rect 2311 5083 2312 5109
rect 2284 5082 2312 5083
rect 2336 5109 2364 5110
rect 2336 5083 2337 5109
rect 2337 5083 2363 5109
rect 2363 5083 2364 5109
rect 2336 5082 2364 5083
rect 3486 6622 3514 6650
rect 2590 5054 2618 5082
rect 3150 5558 3178 5586
rect 2198 4494 2226 4522
rect 2478 4521 2506 4522
rect 2478 4495 2479 4521
rect 2479 4495 2505 4521
rect 2505 4495 2506 4521
rect 2478 4494 2506 4495
rect 2758 4465 2786 4466
rect 2758 4439 2759 4465
rect 2759 4439 2785 4465
rect 2785 4439 2786 4465
rect 2758 4438 2786 4439
rect 2232 4325 2260 4326
rect 2232 4299 2233 4325
rect 2233 4299 2259 4325
rect 2259 4299 2260 4325
rect 2232 4298 2260 4299
rect 2284 4325 2312 4326
rect 2284 4299 2285 4325
rect 2285 4299 2311 4325
rect 2311 4299 2312 4325
rect 2284 4298 2312 4299
rect 2336 4325 2364 4326
rect 2336 4299 2337 4325
rect 2337 4299 2363 4325
rect 2363 4299 2364 4325
rect 2336 4298 2364 4299
rect 1902 3933 1930 3934
rect 1902 3907 1903 3933
rect 1903 3907 1929 3933
rect 1929 3907 1930 3933
rect 1902 3906 1930 3907
rect 1954 3933 1982 3934
rect 1954 3907 1955 3933
rect 1955 3907 1981 3933
rect 1981 3907 1982 3933
rect 1954 3906 1982 3907
rect 2006 3933 2034 3934
rect 2006 3907 2007 3933
rect 2007 3907 2033 3933
rect 2033 3907 2034 3933
rect 2646 3934 2674 3962
rect 2006 3906 2034 3907
rect 1246 3766 1274 3794
rect 2232 3541 2260 3542
rect 2232 3515 2233 3541
rect 2233 3515 2259 3541
rect 2259 3515 2260 3541
rect 2232 3514 2260 3515
rect 2284 3541 2312 3542
rect 2284 3515 2285 3541
rect 2285 3515 2311 3541
rect 2311 3515 2312 3541
rect 2284 3514 2312 3515
rect 2336 3541 2364 3542
rect 2336 3515 2337 3541
rect 2337 3515 2363 3541
rect 2363 3515 2364 3541
rect 2336 3514 2364 3515
rect 1358 3318 1386 3346
rect 1902 3149 1930 3150
rect 1902 3123 1903 3149
rect 1903 3123 1929 3149
rect 1929 3123 1930 3149
rect 1902 3122 1930 3123
rect 1954 3149 1982 3150
rect 1954 3123 1955 3149
rect 1955 3123 1981 3149
rect 1981 3123 1982 3149
rect 1954 3122 1982 3123
rect 2006 3149 2034 3150
rect 2006 3123 2007 3149
rect 2007 3123 2033 3149
rect 2033 3123 2034 3149
rect 2006 3122 2034 3123
rect 2232 2757 2260 2758
rect 2232 2731 2233 2757
rect 2233 2731 2259 2757
rect 2259 2731 2260 2757
rect 2232 2730 2260 2731
rect 2284 2757 2312 2758
rect 2284 2731 2285 2757
rect 2285 2731 2311 2757
rect 2311 2731 2312 2757
rect 2284 2730 2312 2731
rect 2336 2757 2364 2758
rect 2336 2731 2337 2757
rect 2337 2731 2363 2757
rect 2363 2731 2364 2757
rect 2336 2730 2364 2731
rect 3150 2590 3178 2618
rect 3766 6622 3794 6650
rect 3878 5809 3906 5810
rect 3878 5783 3879 5809
rect 3879 5783 3905 5809
rect 3905 5783 3906 5809
rect 3878 5782 3906 5783
rect 3318 5222 3346 5250
rect 3318 4774 3346 4802
rect 3262 4270 3290 4298
rect 3710 5166 3738 5194
rect 3654 3878 3682 3906
rect 3262 2590 3290 2618
rect 1246 2561 1274 2562
rect 1246 2535 1247 2561
rect 1247 2535 1273 2561
rect 1273 2535 1274 2561
rect 1246 2534 1274 2535
rect 1414 2561 1442 2562
rect 1414 2535 1415 2561
rect 1415 2535 1441 2561
rect 1441 2535 1442 2561
rect 1414 2534 1442 2535
rect 1902 2365 1930 2366
rect 1902 2339 1903 2365
rect 1903 2339 1929 2365
rect 1929 2339 1930 2365
rect 1902 2338 1930 2339
rect 1954 2365 1982 2366
rect 1954 2339 1955 2365
rect 1955 2339 1981 2365
rect 1981 2339 1982 2365
rect 1954 2338 1982 2339
rect 2006 2365 2034 2366
rect 2006 2339 2007 2365
rect 2007 2339 2033 2365
rect 2033 2339 2034 2365
rect 2006 2338 2034 2339
rect 2478 2086 2506 2114
rect 1190 2057 1218 2058
rect 1190 2031 1191 2057
rect 1191 2031 1217 2057
rect 1217 2031 1218 2057
rect 1190 2030 1218 2031
rect 1302 2057 1330 2058
rect 1302 2031 1303 2057
rect 1303 2031 1329 2057
rect 1329 2031 1330 2057
rect 1302 2030 1330 2031
rect 2232 1973 2260 1974
rect 2232 1947 2233 1973
rect 2233 1947 2259 1973
rect 2259 1947 2260 1973
rect 2232 1946 2260 1947
rect 2284 1973 2312 1974
rect 2284 1947 2285 1973
rect 2285 1947 2311 1973
rect 2311 1947 2312 1973
rect 2284 1946 2312 1947
rect 2336 1973 2364 1974
rect 2336 1947 2337 1973
rect 2337 1947 2363 1973
rect 2363 1947 2364 1973
rect 2336 1946 2364 1947
rect 2870 1974 2898 2002
rect 1302 1777 1330 1778
rect 1302 1751 1303 1777
rect 1303 1751 1329 1777
rect 1329 1751 1330 1777
rect 1302 1750 1330 1751
rect 1470 1777 1498 1778
rect 1470 1751 1471 1777
rect 1471 1751 1497 1777
rect 1497 1751 1498 1777
rect 1470 1750 1498 1751
rect 1526 1694 1554 1722
rect 1414 1302 1442 1330
rect 462 1022 490 1050
rect 1022 937 1050 938
rect 1022 911 1023 937
rect 1023 911 1049 937
rect 1049 911 1050 937
rect 1022 910 1050 911
rect 1902 1581 1930 1582
rect 1902 1555 1903 1581
rect 1903 1555 1929 1581
rect 1929 1555 1930 1581
rect 1902 1554 1930 1555
rect 1954 1581 1982 1582
rect 1954 1555 1955 1581
rect 1955 1555 1981 1581
rect 1981 1555 1982 1581
rect 1954 1554 1982 1555
rect 2006 1581 2034 1582
rect 2006 1555 2007 1581
rect 2007 1555 2033 1581
rect 2033 1555 2034 1581
rect 2006 1554 2034 1555
rect 2232 1189 2260 1190
rect 2232 1163 2233 1189
rect 2233 1163 2259 1189
rect 2259 1163 2260 1189
rect 2232 1162 2260 1163
rect 2284 1189 2312 1190
rect 2284 1163 2285 1189
rect 2285 1163 2311 1189
rect 2311 1163 2312 1189
rect 2284 1162 2312 1163
rect 2336 1189 2364 1190
rect 2336 1163 2337 1189
rect 2337 1163 2363 1189
rect 2363 1163 2364 1189
rect 2336 1162 2364 1163
rect 4102 5838 4130 5866
rect 3990 4158 4018 4186
rect 4382 6622 4410 6650
rect 4270 6201 4298 6202
rect 4270 6175 4271 6201
rect 4271 6175 4297 6201
rect 4297 6175 4298 6201
rect 4270 6174 4298 6175
rect 4550 5894 4578 5922
rect 4158 5782 4186 5810
rect 4158 5697 4186 5698
rect 4158 5671 4159 5697
rect 4159 5671 4185 5697
rect 4185 5671 4186 5697
rect 4158 5670 4186 5671
rect 4886 6734 4914 6762
rect 4830 6174 4858 6202
rect 5054 6201 5082 6202
rect 5054 6175 5055 6201
rect 5055 6175 5081 6201
rect 5081 6175 5082 6201
rect 5054 6174 5082 6175
rect 4550 5334 4578 5362
rect 4942 5054 4970 5082
rect 4158 4998 4186 5026
rect 4438 3009 4466 3010
rect 4438 2983 4439 3009
rect 4439 2983 4465 3009
rect 4465 2983 4466 3009
rect 4438 2982 4466 2983
rect 5166 6286 5194 6314
rect 5278 6174 5306 6202
rect 5670 6622 5698 6650
rect 5334 5305 5362 5306
rect 5334 5279 5335 5305
rect 5335 5279 5361 5305
rect 5361 5279 5362 5305
rect 5334 5278 5362 5279
rect 5054 4718 5082 4746
rect 4942 2702 4970 2730
rect 4998 3878 5026 3906
rect 4158 2646 4186 2674
rect 5446 5809 5474 5810
rect 5446 5783 5447 5809
rect 5447 5783 5473 5809
rect 5473 5783 5474 5809
rect 5446 5782 5474 5783
rect 5950 6734 5978 6762
rect 5950 6481 5978 6482
rect 5950 6455 5951 6481
rect 5951 6455 5977 6481
rect 5977 6455 5978 6481
rect 5950 6454 5978 6455
rect 5838 6201 5866 6202
rect 5838 6175 5839 6201
rect 5839 6175 5865 6201
rect 5865 6175 5866 6201
rect 5838 6174 5866 6175
rect 5726 5782 5754 5810
rect 5838 6006 5866 6034
rect 5390 4046 5418 4074
rect 5670 4270 5698 4298
rect 5054 3598 5082 3626
rect 4998 2478 5026 2506
rect 4158 2310 4186 2338
rect 5838 5446 5866 5474
rect 6006 5390 6034 5418
rect 5950 5334 5978 5362
rect 5894 4942 5922 4970
rect 5782 4830 5810 4858
rect 5894 3990 5922 4018
rect 5726 3150 5754 3178
rect 5894 3094 5922 3122
rect 5894 2534 5922 2562
rect 6006 4998 6034 5026
rect 6566 6958 6594 6986
rect 6454 6398 6482 6426
rect 6398 6174 6426 6202
rect 6286 5950 6314 5978
rect 6230 5670 6258 5698
rect 6118 5054 6146 5082
rect 6230 4494 6258 4522
rect 6062 2926 6090 2954
rect 6006 2814 6034 2842
rect 5950 2198 5978 2226
rect 5670 1862 5698 1890
rect 3934 1078 3962 1106
rect 6118 1049 6146 1050
rect 6118 1023 6119 1049
rect 6119 1023 6145 1049
rect 6145 1023 6146 1049
rect 6118 1022 6146 1023
rect 6230 1049 6258 1050
rect 6230 1023 6231 1049
rect 6231 1023 6257 1049
rect 6257 1023 6258 1049
rect 6230 1022 6258 1023
rect 4382 993 4410 994
rect 4382 967 4383 993
rect 4383 967 4409 993
rect 4409 967 4410 993
rect 4382 966 4410 967
rect 4550 993 4578 994
rect 4550 967 4551 993
rect 4551 967 4577 993
rect 4577 967 4578 993
rect 4550 966 4578 967
rect 910 545 938 546
rect 910 519 911 545
rect 911 519 937 545
rect 937 519 938 545
rect 910 518 938 519
rect 1190 489 1218 490
rect 1190 463 1191 489
rect 1191 463 1217 489
rect 1217 463 1218 489
rect 1190 462 1218 463
rect 1302 489 1330 490
rect 1302 463 1303 489
rect 1303 463 1329 489
rect 1329 463 1330 489
rect 1302 462 1330 463
rect 1902 797 1930 798
rect 1902 771 1903 797
rect 1903 771 1929 797
rect 1929 771 1930 797
rect 1902 770 1930 771
rect 1954 797 1982 798
rect 1954 771 1955 797
rect 1955 771 1981 797
rect 1981 771 1982 797
rect 1954 770 1982 771
rect 2006 797 2034 798
rect 2006 771 2007 797
rect 2007 771 2033 797
rect 2033 771 2034 797
rect 2006 770 2034 771
rect 4382 742 4410 770
rect 2232 405 2260 406
rect 2232 379 2233 405
rect 2233 379 2259 405
rect 2259 379 2260 405
rect 2232 378 2260 379
rect 2284 405 2312 406
rect 2284 379 2285 405
rect 2285 379 2311 405
rect 2311 379 2312 405
rect 2284 378 2312 379
rect 2336 405 2364 406
rect 2336 379 2337 405
rect 2337 379 2363 405
rect 2363 379 2364 405
rect 2336 378 2364 379
rect 2926 126 2954 154
rect 4774 518 4802 546
rect 4830 238 4858 266
rect 4998 545 5026 546
rect 4998 519 4999 545
rect 4999 519 5025 545
rect 5025 519 5026 545
rect 4998 518 5026 519
rect 5278 993 5306 994
rect 5278 967 5279 993
rect 5279 967 5305 993
rect 5305 967 5306 993
rect 5278 966 5306 967
rect 5838 798 5866 826
rect 5278 657 5306 658
rect 5278 631 5279 657
rect 5279 631 5305 657
rect 5305 631 5306 657
rect 5278 630 5306 631
rect 5054 238 5082 266
rect 4886 182 4914 210
rect 6342 5278 6370 5306
rect 6510 5278 6538 5306
rect 6398 5249 6426 5250
rect 6398 5223 6399 5249
rect 6399 5223 6425 5249
rect 6425 5223 6426 5249
rect 6398 5222 6426 5223
rect 6342 3038 6370 3066
rect 6622 6622 6650 6650
rect 6678 6958 6706 6986
rect 6958 6734 6986 6762
rect 6678 6286 6706 6314
rect 6902 6062 6930 6090
rect 6734 5558 6762 5586
rect 6734 3766 6762 3794
rect 6734 3654 6762 3682
rect 6734 3542 6762 3570
rect 6622 3094 6650 3122
rect 7518 6734 7546 6762
rect 7462 6537 7490 6538
rect 7462 6511 7463 6537
rect 7463 6511 7489 6537
rect 7489 6511 7490 6537
rect 7462 6510 7490 6511
rect 7350 6454 7378 6482
rect 7238 5782 7266 5810
rect 6902 4550 6930 4578
rect 7182 4606 7210 4634
rect 6790 3094 6818 3122
rect 7070 4550 7098 4578
rect 6566 2982 6594 3010
rect 6510 2534 6538 2562
rect 6678 1750 6706 1778
rect 6510 1246 6538 1274
rect 6286 742 6314 770
rect 7014 3654 7042 3682
rect 6902 3598 6930 3626
rect 7238 3598 7266 3626
rect 7294 5054 7322 5082
rect 7182 2926 7210 2954
rect 7070 2870 7098 2898
rect 7014 1414 7042 1442
rect 7070 2422 7098 2450
rect 7070 1358 7098 1386
rect 7126 2086 7154 2114
rect 7126 1302 7154 1330
rect 7182 1806 7210 1834
rect 6902 798 6930 826
rect 7518 6454 7546 6482
rect 7406 5670 7434 5698
rect 7742 5390 7770 5418
rect 7686 5249 7714 5250
rect 7686 5223 7687 5249
rect 7687 5223 7713 5249
rect 7713 5223 7714 5249
rect 7686 5222 7714 5223
rect 7518 4913 7546 4914
rect 7518 4887 7519 4913
rect 7519 4887 7545 4913
rect 7545 4887 7546 4913
rect 7518 4886 7546 4887
rect 7462 4550 7490 4578
rect 7686 4550 7714 4578
rect 7462 4382 7490 4410
rect 7350 3430 7378 3458
rect 7518 3934 7546 3962
rect 7630 3625 7658 3626
rect 7630 3599 7631 3625
rect 7631 3599 7657 3625
rect 7657 3599 7658 3625
rect 7630 3598 7658 3599
rect 7574 2646 7602 2674
rect 7798 3598 7826 3626
rect 7798 3374 7826 3402
rect 7462 2030 7490 2058
rect 7798 2702 7826 2730
rect 7630 2254 7658 2282
rect 7350 1302 7378 1330
rect 7350 1078 7378 1106
rect 7182 742 7210 770
rect 7574 1638 7602 1666
rect 7630 1526 7658 1554
rect 7686 2142 7714 2170
rect 7574 798 7602 826
rect 7966 6454 7994 6482
rect 8414 6510 8442 6538
rect 8190 6201 8218 6202
rect 8190 6175 8191 6201
rect 8191 6175 8217 6201
rect 8217 6175 8218 6201
rect 8190 6174 8218 6175
rect 8694 6622 8722 6650
rect 8638 6174 8666 6202
rect 8470 6033 8498 6034
rect 8470 6007 8471 6033
rect 8471 6007 8497 6033
rect 8497 6007 8498 6033
rect 8470 6006 8498 6007
rect 8750 5894 8778 5922
rect 8638 5614 8666 5642
rect 8134 5417 8162 5418
rect 8134 5391 8135 5417
rect 8135 5391 8161 5417
rect 8161 5391 8162 5417
rect 8134 5390 8162 5391
rect 8750 5614 8778 5642
rect 8974 6201 9002 6202
rect 8974 6175 8975 6201
rect 8975 6175 9001 6201
rect 9001 6175 9002 6201
rect 8974 6174 9002 6175
rect 9030 5697 9058 5698
rect 9030 5671 9031 5697
rect 9031 5671 9057 5697
rect 9057 5671 9058 5697
rect 9030 5670 9058 5671
rect 8246 5222 8274 5250
rect 7910 3318 7938 3346
rect 7966 3598 7994 3626
rect 7854 1918 7882 1946
rect 7910 910 7938 938
rect 7854 686 7882 714
rect 7518 518 7546 546
rect 6846 406 6874 434
rect 6678 294 6706 322
rect 7294 126 7322 154
rect 8022 3542 8050 3570
rect 8918 4662 8946 4690
rect 8806 3766 8834 3794
rect 8526 3206 8554 3234
rect 8582 3430 8610 3458
rect 8414 2505 8442 2506
rect 8414 2479 8415 2505
rect 8415 2479 8441 2505
rect 8441 2479 8442 2505
rect 8414 2478 8442 2479
rect 8470 2254 8498 2282
rect 8414 1974 8442 2002
rect 8358 1833 8386 1834
rect 8358 1807 8359 1833
rect 8359 1807 8385 1833
rect 8385 1807 8386 1833
rect 8358 1806 8386 1807
rect 8414 1470 8442 1498
rect 8414 1134 8442 1162
rect 8078 1105 8106 1106
rect 8078 1079 8079 1105
rect 8079 1079 8105 1105
rect 8105 1079 8106 1105
rect 8078 1078 8106 1079
rect 8358 1105 8386 1106
rect 8358 1079 8359 1105
rect 8359 1079 8385 1105
rect 8385 1079 8386 1105
rect 8358 1078 8386 1079
rect 8414 686 8442 714
rect 8526 2057 8554 2058
rect 8526 2031 8527 2057
rect 8527 2031 8553 2057
rect 8553 2031 8554 2057
rect 8526 2030 8554 2031
rect 8750 3345 8778 3346
rect 8750 3319 8751 3345
rect 8751 3319 8777 3345
rect 8777 3319 8778 3345
rect 8750 3318 8778 3319
rect 8974 3710 9002 3738
rect 8638 2057 8666 2058
rect 8638 2031 8639 2057
rect 8639 2031 8665 2057
rect 8665 2031 8666 2057
rect 8638 2030 8666 2031
rect 8638 1889 8666 1890
rect 8638 1863 8639 1889
rect 8639 1863 8665 1889
rect 8665 1863 8666 1889
rect 8638 1862 8666 1863
rect 8806 1889 8834 1890
rect 8806 1863 8807 1889
rect 8807 1863 8833 1889
rect 8833 1863 8834 1889
rect 8806 1862 8834 1863
rect 9030 2982 9058 3010
rect 9478 6593 9506 6594
rect 9478 6567 9479 6593
rect 9479 6567 9505 6593
rect 9505 6567 9506 6593
rect 9478 6566 9506 6567
rect 9870 6902 9898 6930
rect 9758 6622 9786 6650
rect 9814 6846 9842 6874
rect 9534 6174 9562 6202
rect 9646 6510 9674 6538
rect 9422 6089 9450 6090
rect 9422 6063 9423 6089
rect 9423 6063 9449 6089
rect 9449 6063 9450 6089
rect 9422 6062 9450 6063
rect 9590 6006 9618 6034
rect 9366 5726 9394 5754
rect 9310 5502 9338 5530
rect 9198 4158 9226 4186
rect 9254 4270 9282 4298
rect 9254 4046 9282 4074
rect 9366 4998 9394 5026
rect 9422 5670 9450 5698
rect 9310 3878 9338 3906
rect 9366 4046 9394 4074
rect 9422 3710 9450 3738
rect 9366 3598 9394 3626
rect 9198 2982 9226 3010
rect 9254 3262 9282 3290
rect 9142 2758 9170 2786
rect 9366 2617 9394 2618
rect 9366 2591 9367 2617
rect 9367 2591 9393 2617
rect 9393 2591 9394 2617
rect 9366 2590 9394 2591
rect 9758 6481 9786 6482
rect 9758 6455 9759 6481
rect 9759 6455 9785 6481
rect 9785 6455 9786 6481
rect 9758 6454 9786 6455
rect 9646 5334 9674 5362
rect 9702 6398 9730 6426
rect 9702 4382 9730 4410
rect 9814 4326 9842 4354
rect 9814 3430 9842 3458
rect 9590 2590 9618 2618
rect 9254 2534 9282 2562
rect 10430 6566 10458 6594
rect 10598 6593 10626 6594
rect 10598 6567 10599 6593
rect 10599 6567 10625 6593
rect 10625 6567 10626 6593
rect 10598 6566 10626 6567
rect 10430 6006 10458 6034
rect 11102 6566 11130 6594
rect 10822 5390 10850 5418
rect 10766 5361 10794 5362
rect 10766 5335 10767 5361
rect 10767 5335 10793 5361
rect 10793 5335 10794 5361
rect 10766 5334 10794 5335
rect 9926 2926 9954 2954
rect 10206 4382 10234 4410
rect 9982 2702 10010 2730
rect 10094 2926 10122 2954
rect 10094 2366 10122 2394
rect 10038 1918 10066 1946
rect 9870 1862 9898 1890
rect 8974 1750 9002 1778
rect 8582 1134 8610 1162
rect 8750 1694 8778 1722
rect 8470 630 8498 658
rect 8022 518 8050 546
rect 7966 70 7994 98
rect 10542 5110 10570 5138
rect 10374 3486 10402 3514
rect 10430 4326 10458 4354
rect 10430 2310 10458 2338
rect 10486 3878 10514 3906
rect 10486 1638 10514 1666
rect 10206 1526 10234 1554
rect 10206 742 10234 770
rect 10878 4998 10906 5026
rect 10934 6342 10962 6370
rect 10710 4718 10738 4746
rect 10822 3822 10850 3850
rect 10654 2617 10682 2618
rect 10654 2591 10655 2617
rect 10655 2591 10681 2617
rect 10681 2591 10682 2617
rect 10654 2590 10682 2591
rect 11158 6174 11186 6202
rect 11382 6593 11410 6594
rect 11382 6567 11383 6593
rect 11383 6567 11409 6593
rect 11409 6567 11410 6593
rect 11382 6566 11410 6567
rect 11102 5417 11130 5418
rect 11102 5391 11103 5417
rect 11103 5391 11129 5417
rect 11129 5391 11130 5417
rect 11102 5390 11130 5391
rect 11438 5222 11466 5250
rect 11102 4886 11130 4914
rect 11606 6062 11634 6090
rect 11998 6566 12026 6594
rect 11902 6285 11930 6286
rect 11902 6259 11903 6285
rect 11903 6259 11929 6285
rect 11929 6259 11930 6285
rect 11902 6258 11930 6259
rect 11954 6285 11982 6286
rect 11954 6259 11955 6285
rect 11955 6259 11981 6285
rect 11981 6259 11982 6285
rect 11954 6258 11982 6259
rect 12006 6285 12034 6286
rect 12006 6259 12007 6285
rect 12007 6259 12033 6285
rect 12033 6259 12034 6285
rect 12006 6258 12034 6259
rect 12232 6677 12260 6678
rect 12232 6651 12233 6677
rect 12233 6651 12259 6677
rect 12259 6651 12260 6677
rect 12232 6650 12260 6651
rect 12284 6677 12312 6678
rect 12284 6651 12285 6677
rect 12285 6651 12311 6677
rect 12311 6651 12312 6677
rect 12284 6650 12312 6651
rect 12336 6677 12364 6678
rect 12336 6651 12337 6677
rect 12337 6651 12363 6677
rect 12363 6651 12364 6677
rect 12336 6650 12364 6651
rect 12222 6230 12250 6258
rect 11998 5558 12026 5586
rect 11902 5501 11930 5502
rect 11902 5475 11903 5501
rect 11903 5475 11929 5501
rect 11929 5475 11930 5501
rect 11902 5474 11930 5475
rect 11954 5501 11982 5502
rect 11954 5475 11955 5501
rect 11955 5475 11981 5501
rect 11981 5475 11982 5501
rect 11954 5474 11982 5475
rect 12006 5501 12034 5502
rect 12006 5475 12007 5501
rect 12007 5475 12033 5501
rect 12033 5475 12034 5501
rect 12006 5474 12034 5475
rect 11438 4550 11466 4578
rect 10934 2673 10962 2674
rect 10934 2647 10935 2673
rect 10935 2647 10961 2673
rect 10961 2647 10962 2673
rect 10934 2646 10962 2647
rect 10990 4214 11018 4242
rect 10822 2310 10850 2338
rect 10878 2534 10906 2562
rect 10878 1694 10906 1722
rect 11662 4158 11690 4186
rect 11606 3374 11634 3402
rect 11102 2673 11130 2674
rect 11102 2647 11103 2673
rect 11103 2647 11129 2673
rect 11129 2647 11130 2673
rect 11102 2646 11130 2647
rect 11158 1638 11186 1666
rect 11326 1414 11354 1442
rect 11662 3262 11690 3290
rect 11662 2478 11690 2506
rect 11662 2142 11690 2170
rect 11774 4942 11802 4970
rect 11902 4717 11930 4718
rect 11902 4691 11903 4717
rect 11903 4691 11929 4717
rect 11929 4691 11930 4717
rect 11902 4690 11930 4691
rect 11954 4717 11982 4718
rect 11954 4691 11955 4717
rect 11955 4691 11981 4717
rect 11981 4691 11982 4717
rect 11954 4690 11982 4691
rect 12006 4717 12034 4718
rect 12006 4691 12007 4717
rect 12007 4691 12033 4717
rect 12033 4691 12034 4717
rect 12006 4690 12034 4691
rect 12110 4662 12138 4690
rect 12110 4326 12138 4354
rect 11902 3933 11930 3934
rect 11902 3907 11903 3933
rect 11903 3907 11929 3933
rect 11929 3907 11930 3933
rect 11902 3906 11930 3907
rect 11954 3933 11982 3934
rect 11954 3907 11955 3933
rect 11955 3907 11981 3933
rect 11981 3907 11982 3933
rect 11954 3906 11982 3907
rect 12006 3933 12034 3934
rect 12006 3907 12007 3933
rect 12007 3907 12033 3933
rect 12033 3907 12034 3933
rect 12006 3906 12034 3907
rect 12110 3878 12138 3906
rect 11902 3149 11930 3150
rect 11902 3123 11903 3149
rect 11903 3123 11929 3149
rect 11929 3123 11930 3149
rect 11902 3122 11930 3123
rect 11954 3149 11982 3150
rect 11954 3123 11955 3149
rect 11955 3123 11981 3149
rect 11981 3123 11982 3149
rect 11954 3122 11982 3123
rect 12006 3149 12034 3150
rect 12006 3123 12007 3149
rect 12007 3123 12033 3149
rect 12033 3123 12034 3149
rect 12006 3122 12034 3123
rect 12232 5893 12260 5894
rect 12232 5867 12233 5893
rect 12233 5867 12259 5893
rect 12259 5867 12260 5893
rect 12232 5866 12260 5867
rect 12284 5893 12312 5894
rect 12284 5867 12285 5893
rect 12285 5867 12311 5893
rect 12311 5867 12312 5893
rect 12284 5866 12312 5867
rect 12336 5893 12364 5894
rect 12336 5867 12337 5893
rect 12337 5867 12363 5893
rect 12363 5867 12364 5893
rect 12336 5866 12364 5867
rect 12502 5894 12530 5922
rect 12502 5390 12530 5418
rect 12232 5109 12260 5110
rect 12232 5083 12233 5109
rect 12233 5083 12259 5109
rect 12259 5083 12260 5109
rect 12232 5082 12260 5083
rect 12284 5109 12312 5110
rect 12284 5083 12285 5109
rect 12285 5083 12311 5109
rect 12311 5083 12312 5109
rect 12284 5082 12312 5083
rect 12336 5109 12364 5110
rect 12336 5083 12337 5109
rect 12337 5083 12363 5109
rect 12363 5083 12364 5109
rect 12336 5082 12364 5083
rect 12502 5054 12530 5082
rect 12502 4382 12530 4410
rect 12232 4325 12260 4326
rect 12232 4299 12233 4325
rect 12233 4299 12259 4325
rect 12259 4299 12260 4325
rect 12232 4298 12260 4299
rect 12284 4325 12312 4326
rect 12284 4299 12285 4325
rect 12285 4299 12311 4325
rect 12311 4299 12312 4325
rect 12284 4298 12312 4299
rect 12336 4325 12364 4326
rect 12336 4299 12337 4325
rect 12337 4299 12363 4325
rect 12363 4299 12364 4325
rect 12336 4298 12364 4299
rect 12232 3541 12260 3542
rect 12232 3515 12233 3541
rect 12233 3515 12259 3541
rect 12259 3515 12260 3541
rect 12232 3514 12260 3515
rect 12284 3541 12312 3542
rect 12284 3515 12285 3541
rect 12285 3515 12311 3541
rect 12311 3515 12312 3541
rect 12284 3514 12312 3515
rect 12336 3541 12364 3542
rect 12336 3515 12337 3541
rect 12337 3515 12363 3541
rect 12363 3515 12364 3541
rect 12336 3514 12364 3515
rect 12166 3374 12194 3402
rect 12110 2926 12138 2954
rect 12166 3038 12194 3066
rect 13566 6734 13594 6762
rect 13510 6678 13538 6706
rect 13118 6118 13146 6146
rect 13454 6145 13482 6146
rect 13454 6119 13455 6145
rect 13455 6119 13481 6145
rect 13481 6119 13482 6145
rect 13454 6118 13482 6119
rect 13118 5502 13146 5530
rect 12558 3934 12586 3962
rect 12614 5110 12642 5138
rect 12726 4718 12754 4746
rect 12726 4102 12754 4130
rect 12558 3710 12586 3738
rect 12502 2926 12530 2954
rect 12232 2757 12260 2758
rect 12232 2731 12233 2757
rect 12233 2731 12259 2757
rect 12259 2731 12260 2757
rect 12232 2730 12260 2731
rect 12284 2757 12312 2758
rect 12284 2731 12285 2757
rect 12285 2731 12311 2757
rect 12311 2731 12312 2757
rect 12284 2730 12312 2731
rect 12336 2757 12364 2758
rect 12336 2731 12337 2757
rect 12337 2731 12363 2757
rect 12363 2731 12364 2757
rect 12336 2730 12364 2731
rect 12558 2673 12586 2674
rect 12558 2647 12559 2673
rect 12559 2647 12585 2673
rect 12585 2647 12586 2673
rect 12558 2646 12586 2647
rect 12726 2673 12754 2674
rect 12726 2647 12727 2673
rect 12727 2647 12753 2673
rect 12753 2647 12754 2673
rect 12726 2646 12754 2647
rect 12446 2534 12474 2562
rect 11902 2365 11930 2366
rect 11830 2310 11858 2338
rect 11902 2339 11903 2365
rect 11903 2339 11929 2365
rect 11929 2339 11930 2365
rect 11902 2338 11930 2339
rect 11954 2365 11982 2366
rect 11954 2339 11955 2365
rect 11955 2339 11981 2365
rect 11981 2339 11982 2365
rect 11954 2338 11982 2339
rect 12006 2365 12034 2366
rect 12006 2339 12007 2365
rect 12007 2339 12033 2365
rect 12033 2339 12034 2365
rect 12006 2338 12034 2339
rect 11774 2198 11802 2226
rect 12110 2310 12138 2338
rect 11886 2198 11914 2226
rect 11942 2086 11970 2114
rect 12110 1974 12138 2002
rect 12166 2086 12194 2114
rect 12166 1918 12194 1946
rect 12232 1973 12260 1974
rect 12232 1947 12233 1973
rect 12233 1947 12259 1973
rect 12259 1947 12260 1973
rect 12232 1946 12260 1947
rect 12284 1973 12312 1974
rect 12284 1947 12285 1973
rect 12285 1947 12311 1973
rect 12311 1947 12312 1973
rect 12284 1946 12312 1947
rect 12336 1973 12364 1974
rect 12336 1947 12337 1973
rect 12337 1947 12363 1973
rect 12363 1947 12364 1973
rect 12336 1946 12364 1947
rect 13006 3990 13034 4018
rect 13006 2758 13034 2786
rect 12782 1918 12810 1946
rect 12950 2198 12978 2226
rect 11942 1806 11970 1834
rect 12894 1750 12922 1778
rect 13342 5838 13370 5866
rect 13510 5782 13538 5810
rect 13510 5614 13538 5642
rect 13454 5502 13482 5530
rect 13342 4662 13370 4690
rect 13398 4830 13426 4858
rect 13174 4550 13202 4578
rect 13230 4326 13258 4354
rect 13174 2926 13202 2954
rect 13174 2422 13202 2450
rect 13398 3542 13426 3570
rect 13286 3262 13314 3290
rect 13398 2926 13426 2954
rect 13230 2254 13258 2282
rect 13286 2366 13314 2394
rect 13118 1862 13146 1890
rect 13118 1750 13146 1778
rect 11718 1638 11746 1666
rect 12894 1638 12922 1666
rect 11830 1582 11858 1610
rect 11902 1581 11930 1582
rect 11902 1555 11903 1581
rect 11903 1555 11929 1581
rect 11929 1555 11930 1581
rect 11902 1554 11930 1555
rect 11954 1581 11982 1582
rect 11954 1555 11955 1581
rect 11955 1555 11981 1581
rect 11981 1555 11982 1581
rect 11954 1554 11982 1555
rect 12006 1581 12034 1582
rect 12006 1555 12007 1581
rect 12007 1555 12033 1581
rect 12033 1555 12034 1581
rect 12006 1554 12034 1555
rect 11830 1358 11858 1386
rect 13006 1526 13034 1554
rect 12232 1189 12260 1190
rect 12166 1134 12194 1162
rect 12232 1163 12233 1189
rect 12233 1163 12259 1189
rect 12259 1163 12260 1189
rect 12232 1162 12260 1163
rect 12284 1189 12312 1190
rect 12284 1163 12285 1189
rect 12285 1163 12311 1189
rect 12311 1163 12312 1189
rect 12284 1162 12312 1163
rect 12336 1189 12364 1190
rect 12336 1163 12337 1189
rect 12337 1163 12363 1189
rect 12363 1163 12364 1189
rect 12336 1162 12364 1163
rect 12166 1022 12194 1050
rect 13510 4382 13538 4410
rect 13958 6734 13986 6762
rect 14238 7014 14266 7042
rect 14462 6958 14490 6986
rect 14574 6566 14602 6594
rect 13790 6230 13818 6258
rect 14070 6174 14098 6202
rect 13622 5697 13650 5698
rect 13622 5671 13623 5697
rect 13623 5671 13649 5697
rect 13649 5671 13650 5697
rect 13622 5670 13650 5671
rect 13790 6062 13818 6090
rect 13790 5782 13818 5810
rect 13734 5110 13762 5138
rect 13734 3822 13762 3850
rect 13510 3374 13538 3402
rect 13678 3009 13706 3010
rect 13678 2983 13679 3009
rect 13679 2983 13705 3009
rect 13705 2983 13706 3009
rect 13678 2982 13706 2983
rect 13510 2870 13538 2898
rect 13622 2870 13650 2898
rect 13454 2646 13482 2674
rect 13398 2086 13426 2114
rect 13566 2254 13594 2282
rect 13286 1470 13314 1498
rect 13454 2030 13482 2058
rect 13006 966 13034 994
rect 11326 854 11354 882
rect 11830 910 11858 938
rect 10990 798 11018 826
rect 11830 742 11858 770
rect 11902 797 11930 798
rect 11902 771 11903 797
rect 11903 771 11929 797
rect 11929 771 11930 797
rect 11902 770 11930 771
rect 11954 797 11982 798
rect 11954 771 11955 797
rect 11955 771 11981 797
rect 11981 771 11982 797
rect 11954 770 11982 771
rect 12006 797 12034 798
rect 12006 771 12007 797
rect 12007 771 12033 797
rect 12033 771 12034 797
rect 13454 798 13482 826
rect 13510 1414 13538 1442
rect 12006 770 12034 771
rect 10542 238 10570 266
rect 11662 630 11690 658
rect 13566 574 13594 602
rect 13510 518 13538 546
rect 12232 405 12260 406
rect 12232 379 12233 405
rect 12233 379 12259 405
rect 12259 379 12260 405
rect 12232 378 12260 379
rect 12284 405 12312 406
rect 12284 379 12285 405
rect 12285 379 12311 405
rect 12311 379 12312 405
rect 12284 378 12312 379
rect 12336 405 12364 406
rect 12336 379 12337 405
rect 12337 379 12363 405
rect 12363 379 12364 405
rect 12336 378 12364 379
rect 13118 294 13146 322
rect 13734 1694 13762 1722
rect 13846 4046 13874 4074
rect 13902 3990 13930 4018
rect 13902 2366 13930 2394
rect 14014 4718 14042 4746
rect 14014 3430 14042 3458
rect 14070 3934 14098 3962
rect 13958 2086 13986 2114
rect 14070 2030 14098 2058
rect 13958 1750 13986 1778
rect 13958 1582 13986 1610
rect 13790 1134 13818 1162
rect 14462 6118 14490 6146
rect 14294 6006 14322 6034
rect 14238 5641 14266 5642
rect 14238 5615 14239 5641
rect 14239 5615 14265 5641
rect 14265 5615 14266 5641
rect 14238 5614 14266 5615
rect 14518 5977 14546 5978
rect 14518 5951 14519 5977
rect 14519 5951 14545 5977
rect 14545 5951 14546 5977
rect 14518 5950 14546 5951
rect 14294 5558 14322 5586
rect 14406 5894 14434 5922
rect 14630 5977 14658 5978
rect 14630 5951 14631 5977
rect 14631 5951 14657 5977
rect 14657 5951 14658 5977
rect 14630 5950 14658 5951
rect 14182 4998 14210 5026
rect 14182 4158 14210 4186
rect 14238 4214 14266 4242
rect 14910 6622 14938 6650
rect 14910 6510 14938 6538
rect 14686 5502 14714 5530
rect 14574 5390 14602 5418
rect 14350 3822 14378 3850
rect 14406 4830 14434 4858
rect 14294 3598 14322 3626
rect 14350 3710 14378 3738
rect 14350 2590 14378 2618
rect 14238 2534 14266 2562
rect 14518 4521 14546 4522
rect 14518 4495 14519 4521
rect 14519 4495 14545 4521
rect 14545 4495 14546 4521
rect 14518 4494 14546 4495
rect 14462 3934 14490 3962
rect 14462 2870 14490 2898
rect 14518 2617 14546 2618
rect 14518 2591 14519 2617
rect 14519 2591 14545 2617
rect 14545 2591 14546 2617
rect 14518 2590 14546 2591
rect 14406 2310 14434 2338
rect 14126 1078 14154 1106
rect 14182 1918 14210 1946
rect 14182 966 14210 994
rect 14294 1918 14322 1946
rect 14294 910 14322 938
rect 14350 1806 14378 1834
rect 15022 6174 15050 6202
rect 14742 4606 14770 4634
rect 14686 4494 14714 4522
rect 14574 1750 14602 1778
rect 14630 1862 14658 1890
rect 14630 1470 14658 1498
rect 14406 854 14434 882
rect 14406 742 14434 770
rect 14966 5110 14994 5138
rect 14910 3430 14938 3458
rect 15190 6145 15218 6146
rect 15190 6119 15191 6145
rect 15191 6119 15217 6145
rect 15217 6119 15218 6145
rect 15190 6118 15218 6119
rect 15302 6118 15330 6146
rect 15246 6006 15274 6034
rect 15190 5950 15218 5978
rect 15190 4942 15218 4970
rect 15246 4494 15274 4522
rect 15134 4214 15162 4242
rect 15078 4158 15106 4186
rect 15078 2897 15106 2898
rect 15078 2871 15079 2897
rect 15079 2871 15105 2897
rect 15105 2871 15106 2897
rect 15078 2870 15106 2871
rect 15190 2897 15218 2898
rect 15190 2871 15191 2897
rect 15191 2871 15217 2897
rect 15217 2871 15218 2897
rect 15190 2870 15218 2871
rect 15582 6566 15610 6594
rect 15414 6342 15442 6370
rect 15582 6342 15610 6370
rect 15582 5838 15610 5866
rect 15358 3710 15386 3738
rect 15470 4886 15498 4914
rect 15358 3262 15386 3290
rect 15134 2702 15162 2730
rect 15022 2254 15050 2282
rect 15078 2534 15106 2562
rect 15190 2534 15218 2562
rect 15134 2254 15162 2282
rect 15190 1638 15218 1666
rect 15134 1414 15162 1442
rect 14966 966 14994 994
rect 14686 630 14714 658
rect 14350 574 14378 602
rect 15414 2758 15442 2786
rect 15414 2478 15442 2506
rect 15582 4886 15610 4914
rect 15638 5670 15666 5698
rect 15582 3822 15610 3850
rect 15526 3289 15554 3290
rect 15526 3263 15527 3289
rect 15527 3263 15553 3289
rect 15553 3263 15554 3289
rect 15526 3262 15554 3263
rect 15470 2366 15498 2394
rect 15582 2142 15610 2170
rect 15414 1246 15442 1274
rect 15694 4270 15722 4298
rect 15862 6398 15890 6426
rect 15862 6286 15890 6314
rect 15806 5894 15834 5922
rect 15918 5894 15946 5922
rect 15862 4830 15890 4858
rect 15918 5222 15946 5250
rect 15806 4102 15834 4130
rect 15694 3094 15722 3122
rect 16254 6902 16282 6930
rect 16310 6958 16338 6986
rect 16254 6398 16282 6426
rect 16254 6062 16282 6090
rect 16366 6062 16394 6090
rect 16030 3766 16058 3794
rect 16086 5054 16114 5082
rect 16086 2926 16114 2954
rect 16142 4942 16170 4970
rect 15918 2590 15946 2618
rect 16310 5614 16338 5642
rect 16310 5334 16338 5362
rect 16142 2254 16170 2282
rect 15638 1078 15666 1106
rect 16198 1049 16226 1050
rect 16198 1023 16199 1049
rect 16199 1023 16225 1049
rect 16225 1023 16226 1049
rect 16198 1022 16226 1023
rect 16478 5950 16506 5978
rect 16590 6622 16618 6650
rect 16646 5278 16674 5306
rect 16646 3878 16674 3906
rect 16590 3766 16618 3794
rect 16926 6566 16954 6594
rect 17150 6454 17178 6482
rect 16814 6286 16842 6314
rect 17206 6174 17234 6202
rect 17094 6006 17122 6034
rect 16982 5894 17010 5922
rect 16758 4718 16786 4746
rect 16926 4830 16954 4858
rect 16926 3822 16954 3850
rect 16702 3430 16730 3458
rect 16366 2982 16394 3010
rect 16758 3374 16786 3402
rect 17038 5726 17066 5754
rect 17038 5502 17066 5530
rect 16982 3374 17010 3402
rect 17038 4214 17066 4242
rect 16758 2478 16786 2506
rect 17150 5838 17178 5866
rect 17150 5726 17178 5754
rect 17150 4774 17178 4802
rect 17150 4046 17178 4074
rect 17094 3710 17122 3738
rect 17318 6174 17346 6202
rect 17262 5838 17290 5866
rect 17598 6790 17626 6818
rect 17486 6678 17514 6706
rect 17374 5894 17402 5922
rect 17430 6230 17458 6258
rect 17318 5110 17346 5138
rect 17318 4998 17346 5026
rect 17598 5950 17626 5978
rect 17430 4998 17458 5026
rect 17486 5614 17514 5642
rect 17374 4942 17402 4970
rect 17262 3934 17290 3962
rect 17262 3793 17290 3794
rect 17262 3767 17263 3793
rect 17263 3767 17289 3793
rect 17289 3767 17290 3793
rect 17262 3766 17290 3767
rect 17262 3374 17290 3402
rect 17542 5166 17570 5194
rect 17542 4774 17570 4802
rect 17598 3822 17626 3850
rect 17878 5670 17906 5698
rect 17990 5894 18018 5922
rect 17822 3766 17850 3794
rect 17878 4270 17906 4298
rect 17654 3654 17682 3682
rect 17486 3150 17514 3178
rect 17262 2758 17290 2786
rect 17206 2646 17234 2674
rect 17038 2310 17066 2338
rect 17374 2590 17402 2618
rect 17934 3766 17962 3794
rect 17934 3598 17962 3626
rect 18270 6846 18298 6874
rect 18270 6566 18298 6594
rect 18046 4494 18074 4522
rect 18214 5054 18242 5082
rect 17990 3150 18018 3178
rect 18046 4382 18074 4410
rect 18550 6398 18578 6426
rect 18270 4382 18298 4410
rect 18326 5390 18354 5418
rect 18214 3766 18242 3794
rect 18270 4270 18298 4298
rect 18046 3038 18074 3066
rect 18158 2814 18186 2842
rect 17374 2254 17402 2282
rect 18158 2590 18186 2618
rect 17094 1750 17122 1778
rect 17094 1582 17122 1610
rect 17486 1638 17514 1666
rect 17486 1022 17514 1050
rect 17654 1134 17682 1162
rect 18158 1302 18186 1330
rect 18214 1918 18242 1946
rect 17822 854 17850 882
rect 17878 1134 17906 1162
rect 15358 462 15386 490
rect 18158 1078 18186 1106
rect 17934 742 17962 770
rect 18102 742 18130 770
rect 18494 5054 18522 5082
rect 18382 4046 18410 4074
rect 18438 4158 18466 4186
rect 18382 3654 18410 3682
rect 18718 6062 18746 6090
rect 18494 4046 18522 4074
rect 18438 3542 18466 3570
rect 19166 6286 19194 6314
rect 19054 5894 19082 5922
rect 18774 3262 18802 3290
rect 18998 3374 19026 3402
rect 18326 2982 18354 3010
rect 18494 2870 18522 2898
rect 18270 1582 18298 1610
rect 18326 2646 18354 2674
rect 18382 2310 18410 2338
rect 18382 1582 18410 1610
rect 18606 2646 18634 2674
rect 18326 1302 18354 1330
rect 18494 1750 18522 1778
rect 18494 1470 18522 1498
rect 18438 1190 18466 1218
rect 18270 1078 18298 1106
rect 18662 2422 18690 2450
rect 18270 798 18298 826
rect 18662 574 18690 602
rect 18998 3206 19026 3234
rect 19614 5726 19642 5754
rect 19670 6846 19698 6874
rect 19278 5502 19306 5530
rect 19334 5390 19362 5418
rect 19334 4998 19362 5026
rect 19558 5110 19586 5138
rect 19390 4942 19418 4970
rect 19390 4662 19418 4690
rect 19278 4326 19306 4354
rect 19278 4158 19306 4186
rect 19222 3822 19250 3850
rect 19054 3094 19082 3122
rect 19166 3094 19194 3122
rect 19334 3822 19362 3850
rect 19278 3766 19306 3794
rect 19278 3206 19306 3234
rect 19222 2814 19250 2842
rect 19166 1862 19194 1890
rect 19222 2422 19250 2450
rect 18886 1694 18914 1722
rect 18886 1246 18914 1274
rect 18774 937 18802 938
rect 18774 911 18775 937
rect 18775 911 18801 937
rect 18801 911 18802 937
rect 18774 910 18802 911
rect 18718 462 18746 490
rect 18942 798 18970 826
rect 18214 350 18242 378
rect 17878 294 17906 322
rect 17486 238 17514 266
rect 13622 126 13650 154
rect 14574 126 14602 154
rect 16030 70 16058 98
rect 19278 630 19306 658
rect 19334 2702 19362 2730
rect 19558 2590 19586 2618
rect 19446 993 19474 994
rect 19446 967 19447 993
rect 19447 967 19473 993
rect 19473 967 19474 993
rect 19446 966 19474 967
rect 19838 5614 19866 5642
rect 20006 5950 20034 5978
rect 20286 6118 20314 6146
rect 20342 6622 20370 6650
rect 20286 6033 20314 6034
rect 20286 6007 20287 6033
rect 20287 6007 20313 6033
rect 20313 6007 20314 6033
rect 20286 6006 20314 6007
rect 20398 6033 20426 6034
rect 20398 6007 20399 6033
rect 20399 6007 20425 6033
rect 20425 6007 20426 6033
rect 20398 6006 20426 6007
rect 20062 4830 20090 4858
rect 20174 5614 20202 5642
rect 20230 4577 20258 4578
rect 20230 4551 20231 4577
rect 20231 4551 20257 4577
rect 20257 4551 20258 4577
rect 20230 4550 20258 4551
rect 20174 3822 20202 3850
rect 20006 3542 20034 3570
rect 19894 3430 19922 3458
rect 20006 3430 20034 3458
rect 20006 2926 20034 2954
rect 19894 2702 19922 2730
rect 20174 2702 20202 2730
rect 20678 6089 20706 6090
rect 20678 6063 20679 6089
rect 20679 6063 20705 6089
rect 20705 6063 20706 6089
rect 20678 6062 20706 6063
rect 20846 6454 20874 6482
rect 20734 5894 20762 5922
rect 20790 6398 20818 6426
rect 20510 5614 20538 5642
rect 20454 4774 20482 4802
rect 20622 4577 20650 4578
rect 20622 4551 20623 4577
rect 20623 4551 20649 4577
rect 20649 4551 20650 4577
rect 20622 4550 20650 4551
rect 20678 2646 20706 2674
rect 20734 4662 20762 4690
rect 20398 2478 20426 2506
rect 20510 2254 20538 2282
rect 20174 2030 20202 2058
rect 19894 1974 19922 2002
rect 20230 1862 20258 1890
rect 20230 1638 20258 1666
rect 20622 1806 20650 1834
rect 20398 1302 20426 1330
rect 19838 910 19866 938
rect 19838 798 19866 826
rect 19670 742 19698 770
rect 20174 686 20202 714
rect 20174 574 20202 602
rect 19334 518 19362 546
rect 20902 4270 20930 4298
rect 21070 6734 21098 6762
rect 21014 5166 21042 5194
rect 21014 4606 21042 4634
rect 20958 3934 20986 3962
rect 21014 3990 21042 4018
rect 20902 3822 20930 3850
rect 20958 3766 20986 3794
rect 21014 3710 21042 3738
rect 20790 3262 20818 3290
rect 20958 3318 20986 3346
rect 20958 2646 20986 2674
rect 20902 2617 20930 2618
rect 20902 2591 20903 2617
rect 20903 2591 20929 2617
rect 20929 2591 20930 2617
rect 20902 2590 20930 2591
rect 20846 2086 20874 2114
rect 21014 2086 21042 2114
rect 21126 5614 21154 5642
rect 21126 3990 21154 4018
rect 21126 3766 21154 3794
rect 21630 6958 21658 6986
rect 22078 6846 22106 6874
rect 22302 6734 22330 6762
rect 22232 6677 22260 6678
rect 22232 6651 22233 6677
rect 22233 6651 22259 6677
rect 22259 6651 22260 6677
rect 22232 6650 22260 6651
rect 22284 6677 22312 6678
rect 22284 6651 22285 6677
rect 22285 6651 22311 6677
rect 22311 6651 22312 6677
rect 22284 6650 22312 6651
rect 22336 6677 22364 6678
rect 22336 6651 22337 6677
rect 22337 6651 22363 6677
rect 22363 6651 22364 6677
rect 22336 6650 22364 6651
rect 22526 6398 22554 6426
rect 22638 6902 22666 6930
rect 21854 6342 21882 6370
rect 21902 6285 21930 6286
rect 21902 6259 21903 6285
rect 21903 6259 21929 6285
rect 21929 6259 21930 6285
rect 21902 6258 21930 6259
rect 21954 6285 21982 6286
rect 21954 6259 21955 6285
rect 21955 6259 21981 6285
rect 21981 6259 21982 6285
rect 21954 6258 21982 6259
rect 22006 6285 22034 6286
rect 22006 6259 22007 6285
rect 22007 6259 22033 6285
rect 22033 6259 22034 6285
rect 22006 6258 22034 6259
rect 21798 6033 21826 6034
rect 21798 6007 21799 6033
rect 21799 6007 21825 6033
rect 21825 6007 21826 6033
rect 21798 6006 21826 6007
rect 21406 5977 21434 5978
rect 21406 5951 21407 5977
rect 21407 5951 21433 5977
rect 21433 5951 21434 5977
rect 21406 5950 21434 5951
rect 21518 5977 21546 5978
rect 21518 5951 21519 5977
rect 21519 5951 21545 5977
rect 21545 5951 21546 5977
rect 21518 5950 21546 5951
rect 22232 5893 22260 5894
rect 22232 5867 22233 5893
rect 22233 5867 22259 5893
rect 22259 5867 22260 5893
rect 22232 5866 22260 5867
rect 22284 5893 22312 5894
rect 22284 5867 22285 5893
rect 22285 5867 22311 5893
rect 22311 5867 22312 5893
rect 22284 5866 22312 5867
rect 22336 5893 22364 5894
rect 22336 5867 22337 5893
rect 22337 5867 22363 5893
rect 22363 5867 22364 5893
rect 22336 5866 22364 5867
rect 22582 5894 22610 5922
rect 22414 5558 22442 5586
rect 21902 5501 21930 5502
rect 21902 5475 21903 5501
rect 21903 5475 21929 5501
rect 21929 5475 21930 5501
rect 21902 5474 21930 5475
rect 21954 5501 21982 5502
rect 21954 5475 21955 5501
rect 21955 5475 21981 5501
rect 21981 5475 21982 5501
rect 21954 5474 21982 5475
rect 22006 5501 22034 5502
rect 22006 5475 22007 5501
rect 22007 5475 22033 5501
rect 22033 5475 22034 5501
rect 22006 5474 22034 5475
rect 21798 5249 21826 5250
rect 21798 5223 21799 5249
rect 21799 5223 21825 5249
rect 21825 5223 21826 5249
rect 21798 5222 21826 5223
rect 21238 3793 21266 3794
rect 21238 3767 21239 3793
rect 21239 3767 21265 3793
rect 21265 3767 21266 3793
rect 21238 3766 21266 3767
rect 21294 3430 21322 3458
rect 21182 2702 21210 2730
rect 21070 1974 21098 2002
rect 21014 1918 21042 1946
rect 20790 1806 20818 1834
rect 21070 1750 21098 1778
rect 20790 1134 20818 1162
rect 20902 1246 20930 1274
rect 20734 854 20762 882
rect 21462 3038 21490 3066
rect 21294 3009 21322 3010
rect 21294 2983 21295 3009
rect 21295 2983 21321 3009
rect 21321 2983 21322 3009
rect 21294 2982 21322 2983
rect 21294 2702 21322 2730
rect 21350 2814 21378 2842
rect 21462 2814 21490 2842
rect 21406 2225 21434 2226
rect 21406 2199 21407 2225
rect 21407 2199 21433 2225
rect 21433 2199 21434 2225
rect 21406 2198 21434 2199
rect 21518 1582 21546 1610
rect 21238 1078 21266 1106
rect 21350 1105 21378 1106
rect 21350 1079 21351 1105
rect 21351 1079 21377 1105
rect 21377 1079 21378 1105
rect 21350 1078 21378 1079
rect 21462 1078 21490 1106
rect 22232 5109 22260 5110
rect 22232 5083 22233 5109
rect 22233 5083 22259 5109
rect 22259 5083 22260 5109
rect 22232 5082 22260 5083
rect 22284 5109 22312 5110
rect 22284 5083 22285 5109
rect 22285 5083 22311 5109
rect 22311 5083 22312 5109
rect 22284 5082 22312 5083
rect 22336 5109 22364 5110
rect 22336 5083 22337 5109
rect 22337 5083 22363 5109
rect 22363 5083 22364 5109
rect 22336 5082 22364 5083
rect 22414 5054 22442 5082
rect 21902 4717 21930 4718
rect 21902 4691 21903 4717
rect 21903 4691 21929 4717
rect 21929 4691 21930 4717
rect 21902 4690 21930 4691
rect 21954 4717 21982 4718
rect 21954 4691 21955 4717
rect 21955 4691 21981 4717
rect 21981 4691 21982 4717
rect 21954 4690 21982 4691
rect 22006 4717 22034 4718
rect 22006 4691 22007 4717
rect 22007 4691 22033 4717
rect 22033 4691 22034 4717
rect 22006 4690 22034 4691
rect 22582 4550 22610 4578
rect 22232 4325 22260 4326
rect 22232 4299 22233 4325
rect 22233 4299 22259 4325
rect 22259 4299 22260 4325
rect 22232 4298 22260 4299
rect 22284 4325 22312 4326
rect 22284 4299 22285 4325
rect 22285 4299 22311 4325
rect 22311 4299 22312 4325
rect 22284 4298 22312 4299
rect 22336 4325 22364 4326
rect 22336 4299 22337 4325
rect 22337 4299 22363 4325
rect 22363 4299 22364 4325
rect 22336 4298 22364 4299
rect 22414 4270 22442 4298
rect 21742 3990 21770 4018
rect 21902 3933 21930 3934
rect 21902 3907 21903 3933
rect 21903 3907 21929 3933
rect 21929 3907 21930 3933
rect 21902 3906 21930 3907
rect 21954 3933 21982 3934
rect 21954 3907 21955 3933
rect 21955 3907 21981 3933
rect 21981 3907 21982 3933
rect 21954 3906 21982 3907
rect 22006 3933 22034 3934
rect 22006 3907 22007 3933
rect 22007 3907 22033 3933
rect 22033 3907 22034 3933
rect 22006 3906 22034 3907
rect 22232 3541 22260 3542
rect 22232 3515 22233 3541
rect 22233 3515 22259 3541
rect 22259 3515 22260 3541
rect 22232 3514 22260 3515
rect 22284 3541 22312 3542
rect 22284 3515 22285 3541
rect 22285 3515 22311 3541
rect 22311 3515 22312 3541
rect 22284 3514 22312 3515
rect 22336 3541 22364 3542
rect 22336 3515 22337 3541
rect 22337 3515 22363 3541
rect 22363 3515 22364 3541
rect 22336 3514 22364 3515
rect 21798 3150 21826 3178
rect 21902 3149 21930 3150
rect 21902 3123 21903 3149
rect 21903 3123 21929 3149
rect 21929 3123 21930 3149
rect 21902 3122 21930 3123
rect 21954 3149 21982 3150
rect 21954 3123 21955 3149
rect 21955 3123 21981 3149
rect 21981 3123 21982 3149
rect 21954 3122 21982 3123
rect 22006 3149 22034 3150
rect 22006 3123 22007 3149
rect 22007 3123 22033 3149
rect 22033 3123 22034 3149
rect 22078 3150 22106 3178
rect 22006 3122 22034 3123
rect 22638 2982 22666 3010
rect 21854 2870 21882 2898
rect 22134 2870 22162 2898
rect 21742 2561 21770 2562
rect 21742 2535 21743 2561
rect 21743 2535 21769 2561
rect 21769 2535 21770 2561
rect 21742 2534 21770 2535
rect 21902 2365 21930 2366
rect 21902 2339 21903 2365
rect 21903 2339 21929 2365
rect 21929 2339 21930 2365
rect 21902 2338 21930 2339
rect 21954 2365 21982 2366
rect 21954 2339 21955 2365
rect 21955 2339 21981 2365
rect 21981 2339 21982 2365
rect 21954 2338 21982 2339
rect 22006 2365 22034 2366
rect 22006 2339 22007 2365
rect 22007 2339 22033 2365
rect 22033 2339 22034 2365
rect 22006 2338 22034 2339
rect 22022 1833 22050 1834
rect 22022 1807 22023 1833
rect 22023 1807 22049 1833
rect 22049 1807 22050 1833
rect 22022 1806 22050 1807
rect 21902 1581 21930 1582
rect 21902 1555 21903 1581
rect 21903 1555 21929 1581
rect 21929 1555 21930 1581
rect 21902 1554 21930 1555
rect 21954 1581 21982 1582
rect 21954 1555 21955 1581
rect 21955 1555 21981 1581
rect 21981 1555 21982 1581
rect 21954 1554 21982 1555
rect 22006 1581 22034 1582
rect 22006 1555 22007 1581
rect 22007 1555 22033 1581
rect 22033 1555 22034 1581
rect 22006 1554 22034 1555
rect 21798 993 21826 994
rect 21798 967 21799 993
rect 21799 967 21825 993
rect 21825 967 21826 993
rect 21798 966 21826 967
rect 21966 993 21994 994
rect 21966 967 21967 993
rect 21967 967 21993 993
rect 21993 967 21994 993
rect 21966 966 21994 967
rect 21902 797 21930 798
rect 21902 771 21903 797
rect 21903 771 21929 797
rect 21929 771 21930 797
rect 21902 770 21930 771
rect 21954 797 21982 798
rect 21954 771 21955 797
rect 21955 771 21981 797
rect 21981 771 21982 797
rect 21954 770 21982 771
rect 22006 797 22034 798
rect 22006 771 22007 797
rect 22007 771 22033 797
rect 22033 771 22034 797
rect 22006 770 22034 771
rect 22232 2757 22260 2758
rect 22232 2731 22233 2757
rect 22233 2731 22259 2757
rect 22259 2731 22260 2757
rect 22232 2730 22260 2731
rect 22284 2757 22312 2758
rect 22284 2731 22285 2757
rect 22285 2731 22311 2757
rect 22311 2731 22312 2757
rect 22284 2730 22312 2731
rect 22336 2757 22364 2758
rect 22336 2731 22337 2757
rect 22337 2731 22363 2757
rect 22363 2731 22364 2757
rect 22336 2730 22364 2731
rect 22414 2534 22442 2562
rect 22974 5894 23002 5922
rect 22750 2422 22778 2450
rect 22806 5726 22834 5754
rect 22694 2366 22722 2394
rect 22358 2310 22386 2338
rect 22638 2142 22666 2170
rect 22358 2086 22386 2114
rect 22470 2086 22498 2114
rect 22232 1973 22260 1974
rect 22232 1947 22233 1973
rect 22233 1947 22259 1973
rect 22259 1947 22260 1973
rect 22232 1946 22260 1947
rect 22284 1973 22312 1974
rect 22284 1947 22285 1973
rect 22285 1947 22311 1973
rect 22311 1947 22312 1973
rect 22284 1946 22312 1947
rect 22336 1973 22364 1974
rect 22336 1947 22337 1973
rect 22337 1947 22363 1973
rect 22363 1947 22364 1973
rect 22336 1946 22364 1947
rect 22190 1833 22218 1834
rect 22190 1807 22191 1833
rect 22191 1807 22217 1833
rect 22217 1807 22218 1833
rect 22190 1806 22218 1807
rect 22638 1582 22666 1610
rect 22694 1246 22722 1274
rect 22232 1189 22260 1190
rect 22232 1163 22233 1189
rect 22233 1163 22259 1189
rect 22259 1163 22260 1189
rect 22232 1162 22260 1163
rect 22284 1189 22312 1190
rect 22284 1163 22285 1189
rect 22285 1163 22311 1189
rect 22311 1163 22312 1189
rect 22284 1162 22312 1163
rect 22336 1189 22364 1190
rect 22336 1163 22337 1189
rect 22337 1163 22363 1189
rect 22363 1163 22364 1189
rect 22336 1162 22364 1163
rect 23086 5753 23114 5754
rect 23086 5727 23087 5753
rect 23087 5727 23113 5753
rect 23113 5727 23114 5753
rect 23086 5726 23114 5727
rect 23142 4998 23170 5026
rect 23254 6790 23282 6818
rect 23254 5614 23282 5642
rect 23310 5894 23338 5922
rect 23366 5558 23394 5586
rect 23310 5334 23338 5362
rect 23646 6902 23674 6930
rect 23478 5558 23506 5586
rect 23478 5334 23506 5362
rect 23198 3766 23226 3794
rect 23646 5110 23674 5138
rect 23702 4606 23730 4634
rect 23142 2982 23170 3010
rect 22862 2646 22890 2674
rect 21574 350 21602 378
rect 22694 686 22722 714
rect 22232 405 22260 406
rect 22232 379 22233 405
rect 22233 379 22259 405
rect 22259 379 22260 405
rect 22232 378 22260 379
rect 22284 405 22312 406
rect 22284 379 22285 405
rect 22285 379 22311 405
rect 22311 379 22312 405
rect 22284 378 22312 379
rect 22336 405 22364 406
rect 22336 379 22337 405
rect 22337 379 22363 405
rect 22363 379 22364 405
rect 22694 406 22722 434
rect 22336 378 22364 379
rect 22974 2590 23002 2618
rect 23254 2478 23282 2506
rect 23646 4158 23674 4186
rect 23758 3345 23786 3346
rect 23758 3319 23759 3345
rect 23759 3319 23785 3345
rect 23785 3319 23786 3345
rect 23758 3318 23786 3319
rect 23366 3289 23394 3290
rect 23366 3263 23367 3289
rect 23367 3263 23393 3289
rect 23393 3263 23394 3289
rect 23366 3262 23394 3263
rect 23478 2814 23506 2842
rect 23310 2198 23338 2226
rect 23366 2702 23394 2730
rect 22974 1246 23002 1274
rect 22918 1105 22946 1106
rect 22918 1079 22919 1105
rect 22919 1079 22945 1105
rect 22945 1079 22946 1105
rect 22918 1078 22946 1079
rect 23086 1105 23114 1106
rect 23086 1079 23087 1105
rect 23087 1079 23113 1105
rect 23113 1079 23114 1105
rect 23086 1078 23114 1079
rect 23478 1974 23506 2002
rect 23702 2198 23730 2226
rect 23478 1750 23506 1778
rect 23478 1470 23506 1498
rect 23366 1022 23394 1050
rect 23422 1190 23450 1218
rect 24094 4998 24122 5026
rect 23982 2366 24010 2394
rect 23870 1134 23898 1162
rect 23422 518 23450 546
rect 23478 910 23506 938
rect 22862 350 22890 378
rect 23310 462 23338 490
rect 24262 5390 24290 5418
rect 24150 966 24178 994
rect 24206 4270 24234 4298
rect 24262 3542 24290 3570
rect 24318 5166 24346 5194
rect 24318 2422 24346 2450
rect 24262 1582 24290 1610
rect 24318 1526 24346 1554
rect 24878 5054 24906 5082
rect 24766 2254 24794 2282
rect 24486 1078 24514 1106
rect 24430 937 24458 938
rect 24430 911 24431 937
rect 24431 911 24457 937
rect 24457 911 24458 937
rect 24430 910 24458 911
rect 24598 910 24626 938
rect 24206 462 24234 490
rect 23758 126 23786 154
rect 23478 70 23506 98
rect 25662 6566 25690 6594
rect 25550 5334 25578 5362
rect 25046 2870 25074 2898
rect 24934 2198 24962 2226
rect 25494 3345 25522 3346
rect 25494 3319 25495 3345
rect 25495 3319 25521 3345
rect 25521 3319 25522 3345
rect 25494 3318 25522 3319
rect 25438 2617 25466 2618
rect 25438 2591 25439 2617
rect 25439 2591 25465 2617
rect 25465 2591 25466 2617
rect 25438 2590 25466 2591
rect 25438 2366 25466 2394
rect 25046 1302 25074 1330
rect 24878 1049 24906 1050
rect 24878 1023 24879 1049
rect 24879 1023 24905 1049
rect 24905 1023 24906 1049
rect 24878 1022 24906 1023
rect 24878 798 24906 826
rect 24878 574 24906 602
rect 26054 6593 26082 6594
rect 26054 6567 26055 6593
rect 26055 6567 26081 6593
rect 26081 6567 26082 6593
rect 26054 6566 26082 6567
rect 25886 6174 25914 6202
rect 26054 6454 26082 6482
rect 25774 5894 25802 5922
rect 26558 6734 26586 6762
rect 26334 6510 26362 6538
rect 26558 6398 26586 6426
rect 26278 6201 26306 6202
rect 26278 6175 26279 6201
rect 26279 6175 26305 6201
rect 26305 6175 26306 6201
rect 26278 6174 26306 6175
rect 26558 5726 26586 5754
rect 26614 6342 26642 6370
rect 26222 5697 26250 5698
rect 26222 5671 26223 5697
rect 26223 5671 26249 5697
rect 26249 5671 26250 5697
rect 26222 5670 26250 5671
rect 26054 5614 26082 5642
rect 25718 5334 25746 5362
rect 25718 5110 25746 5138
rect 25998 4382 26026 4410
rect 25998 3822 26026 3850
rect 26222 4521 26250 4522
rect 26222 4495 26223 4521
rect 26223 4495 26249 4521
rect 26249 4495 26250 4521
rect 26222 4494 26250 4495
rect 26390 4521 26418 4522
rect 26390 4495 26391 4521
rect 26391 4495 26417 4521
rect 26417 4495 26418 4521
rect 26390 4494 26418 4495
rect 26670 6118 26698 6146
rect 26782 6089 26810 6090
rect 26782 6063 26783 6089
rect 26783 6063 26809 6089
rect 26809 6063 26810 6089
rect 26782 6062 26810 6063
rect 27454 6846 27482 6874
rect 27230 6566 27258 6594
rect 27454 6734 27482 6762
rect 27006 6174 27034 6202
rect 27062 6510 27090 6538
rect 27902 6734 27930 6762
rect 27678 6454 27706 6482
rect 27846 6201 27874 6202
rect 27846 6175 27847 6201
rect 27847 6175 27873 6201
rect 27873 6175 27874 6201
rect 27846 6174 27874 6175
rect 27174 6006 27202 6034
rect 26838 5782 26866 5810
rect 27286 5809 27314 5810
rect 27286 5783 27287 5809
rect 27287 5783 27313 5809
rect 27313 5783 27314 5809
rect 27286 5782 27314 5783
rect 27006 5222 27034 5250
rect 26670 4550 26698 4578
rect 27118 4998 27146 5026
rect 26670 4465 26698 4466
rect 26670 4439 26671 4465
rect 26671 4439 26697 4465
rect 26697 4439 26698 4465
rect 26670 4438 26698 4439
rect 26446 3318 26474 3346
rect 27118 2590 27146 2618
rect 25998 2310 26026 2338
rect 26334 2534 26362 2562
rect 25606 1638 25634 1666
rect 26110 1750 26138 1778
rect 26054 1470 26082 1498
rect 26110 742 26138 770
rect 26166 1414 26194 1442
rect 26278 1273 26306 1274
rect 26278 1247 26279 1273
rect 26279 1247 26305 1273
rect 26305 1247 26306 1273
rect 26278 1246 26306 1247
rect 26166 630 26194 658
rect 25550 518 25578 546
rect 24990 238 25018 266
rect 26222 462 26250 490
rect 27678 5502 27706 5530
rect 27734 4857 27762 4858
rect 27734 4831 27735 4857
rect 27735 4831 27761 4857
rect 27761 4831 27762 4857
rect 27734 4830 27762 4831
rect 27734 3934 27762 3962
rect 27566 2478 27594 2506
rect 27846 2225 27874 2226
rect 27846 2199 27847 2225
rect 27847 2199 27873 2225
rect 27873 2199 27874 2225
rect 27846 2198 27874 2199
rect 28238 6593 28266 6594
rect 28238 6567 28239 6593
rect 28239 6567 28265 6593
rect 28265 6567 28266 6593
rect 28238 6566 28266 6567
rect 28126 6118 28154 6146
rect 28238 6454 28266 6482
rect 28574 6510 28602 6538
rect 28630 6846 28658 6874
rect 28350 6286 28378 6314
rect 28574 6118 28602 6146
rect 27958 4830 27986 4858
rect 27958 4326 27986 4354
rect 27958 3934 27986 3962
rect 27902 2086 27930 2114
rect 26446 1273 26474 1274
rect 26446 1247 26447 1273
rect 26447 1247 26473 1273
rect 26473 1247 26474 1273
rect 26446 1246 26474 1247
rect 28070 5249 28098 5250
rect 28070 5223 28071 5249
rect 28071 5223 28097 5249
rect 28097 5223 28098 5249
rect 28070 5222 28098 5223
rect 28238 5054 28266 5082
rect 28238 4438 28266 4466
rect 28126 4326 28154 4354
rect 28238 4185 28266 4186
rect 28238 4159 28239 4185
rect 28239 4159 28265 4185
rect 28265 4159 28266 4185
rect 28238 4158 28266 4159
rect 28462 5446 28490 5474
rect 28350 4577 28378 4578
rect 28350 4551 28351 4577
rect 28351 4551 28377 4577
rect 28377 4551 28378 4577
rect 28350 4550 28378 4551
rect 28406 4382 28434 4410
rect 29022 6454 29050 6482
rect 28798 6118 28826 6146
rect 29022 6286 29050 6314
rect 28630 5670 28658 5698
rect 28574 4409 28602 4410
rect 28574 4383 28575 4409
rect 28575 4383 28601 4409
rect 28601 4383 28602 4409
rect 28574 4382 28602 4383
rect 29022 5305 29050 5306
rect 29022 5279 29023 5305
rect 29023 5279 29049 5305
rect 29049 5279 29050 5305
rect 29022 5278 29050 5279
rect 29414 6734 29442 6762
rect 29470 6566 29498 6594
rect 29246 6230 29274 6258
rect 29414 6118 29442 6146
rect 29134 5838 29162 5866
rect 29806 6342 29834 6370
rect 30422 6958 30450 6986
rect 30254 6537 30282 6538
rect 30254 6511 30255 6537
rect 30255 6511 30281 6537
rect 30281 6511 30282 6537
rect 30254 6510 30282 6511
rect 29918 6342 29946 6370
rect 30310 6454 30338 6482
rect 29694 6118 29722 6146
rect 29806 6230 29834 6258
rect 29526 5697 29554 5698
rect 29526 5671 29527 5697
rect 29527 5671 29553 5697
rect 29553 5671 29554 5697
rect 29526 5670 29554 5671
rect 29470 5390 29498 5418
rect 28742 4998 28770 5026
rect 28966 4857 28994 4858
rect 28966 4831 28967 4857
rect 28967 4831 28993 4857
rect 28993 4831 28994 4857
rect 28966 4830 28994 4831
rect 28742 4129 28770 4130
rect 28742 4103 28743 4129
rect 28743 4103 28769 4129
rect 28769 4103 28770 4129
rect 28742 4102 28770 4103
rect 28630 3990 28658 4018
rect 28798 3737 28826 3738
rect 28798 3711 28799 3737
rect 28799 3711 28825 3737
rect 28825 3711 28826 3737
rect 28798 3710 28826 3711
rect 28630 3625 28658 3626
rect 28630 3599 28631 3625
rect 28631 3599 28657 3625
rect 28657 3599 28658 3625
rect 28630 3598 28658 3599
rect 28910 3625 28938 3626
rect 28910 3599 28911 3625
rect 28911 3599 28937 3625
rect 28937 3599 28938 3625
rect 28910 3598 28938 3599
rect 28742 3486 28770 3514
rect 28182 2561 28210 2562
rect 28182 2535 28183 2561
rect 28183 2535 28209 2561
rect 28209 2535 28210 2561
rect 28182 2534 28210 2535
rect 28294 2814 28322 2842
rect 28070 2057 28098 2058
rect 28070 2031 28071 2057
rect 28071 2031 28097 2057
rect 28097 2031 28098 2057
rect 28070 2030 28098 2031
rect 28238 2057 28266 2058
rect 28238 2031 28239 2057
rect 28239 2031 28265 2057
rect 28265 2031 28266 2057
rect 28238 2030 28266 2031
rect 28182 1694 28210 1722
rect 28014 1022 28042 1050
rect 28518 2841 28546 2842
rect 28518 2815 28519 2841
rect 28519 2815 28545 2841
rect 28545 2815 28546 2841
rect 28518 2814 28546 2815
rect 28686 2841 28714 2842
rect 28686 2815 28687 2841
rect 28687 2815 28713 2841
rect 28713 2815 28714 2841
rect 28686 2814 28714 2815
rect 29078 4998 29106 5026
rect 29414 4913 29442 4914
rect 29414 4887 29415 4913
rect 29415 4887 29441 4913
rect 29441 4887 29442 4913
rect 29414 4886 29442 4887
rect 29358 4774 29386 4802
rect 29134 4214 29162 4242
rect 29078 3486 29106 3514
rect 29134 3542 29162 3570
rect 28910 3206 28938 3234
rect 28966 3262 28994 3290
rect 29022 3150 29050 3178
rect 28350 2561 28378 2562
rect 28350 2535 28351 2561
rect 28351 2535 28377 2561
rect 28377 2535 28378 2561
rect 28350 2534 28378 2535
rect 28630 2561 28658 2562
rect 28630 2535 28631 2561
rect 28631 2535 28657 2561
rect 28657 2535 28658 2561
rect 28630 2534 28658 2535
rect 28742 2422 28770 2450
rect 29414 3542 29442 3570
rect 29302 3430 29330 3458
rect 29246 3150 29274 3178
rect 29134 2982 29162 3010
rect 29526 5222 29554 5250
rect 29862 4857 29890 4858
rect 29862 4831 29863 4857
rect 29863 4831 29889 4857
rect 29889 4831 29890 4857
rect 29862 4830 29890 4831
rect 29862 4102 29890 4130
rect 29694 3206 29722 3234
rect 29638 3009 29666 3010
rect 29638 2983 29639 3009
rect 29639 2983 29665 3009
rect 29665 2983 29666 3009
rect 29638 2982 29666 2983
rect 29302 2926 29330 2954
rect 29190 2702 29218 2730
rect 29190 2617 29218 2618
rect 29190 2591 29191 2617
rect 29191 2591 29217 2617
rect 29217 2591 29218 2617
rect 29190 2590 29218 2591
rect 29134 2478 29162 2506
rect 29078 2366 29106 2394
rect 29526 1889 29554 1890
rect 29526 1863 29527 1889
rect 29527 1863 29553 1889
rect 29553 1863 29554 1889
rect 29526 1862 29554 1863
rect 30142 4969 30170 4970
rect 30142 4943 30143 4969
rect 30143 4943 30169 4969
rect 30169 4943 30170 4969
rect 30142 4942 30170 4943
rect 30142 4438 30170 4466
rect 30254 4158 30282 4186
rect 30254 3681 30282 3682
rect 30254 3655 30255 3681
rect 30255 3655 30281 3681
rect 30281 3655 30282 3681
rect 30254 3654 30282 3655
rect 30254 3374 30282 3402
rect 29974 3345 30002 3346
rect 29974 3319 29975 3345
rect 29975 3319 30001 3345
rect 30001 3319 30002 3345
rect 29974 3318 30002 3319
rect 30142 3094 30170 3122
rect 30310 3262 30338 3290
rect 30142 2617 30170 2618
rect 30142 2591 30143 2617
rect 30143 2591 30169 2617
rect 30169 2591 30170 2617
rect 30142 2590 30170 2591
rect 29974 2561 30002 2562
rect 29974 2535 29975 2561
rect 29975 2535 30001 2561
rect 30001 2535 30002 2561
rect 29974 2534 30002 2535
rect 32102 6734 32130 6762
rect 31262 6593 31290 6594
rect 31262 6567 31263 6593
rect 31263 6567 31289 6593
rect 31289 6567 31290 6593
rect 31262 6566 31290 6567
rect 31542 6510 31570 6538
rect 30982 6398 31010 6426
rect 30590 6342 30618 6370
rect 31094 6145 31122 6146
rect 31094 6119 31095 6145
rect 31095 6119 31121 6145
rect 31121 6119 31122 6145
rect 31094 6118 31122 6119
rect 30422 5502 30450 5530
rect 31206 5838 31234 5866
rect 30758 5054 30786 5082
rect 30702 4998 30730 5026
rect 30534 4969 30562 4970
rect 30534 4943 30535 4969
rect 30535 4943 30561 4969
rect 30561 4943 30562 4969
rect 30534 4942 30562 4943
rect 30758 4633 30786 4634
rect 30758 4607 30759 4633
rect 30759 4607 30785 4633
rect 30785 4607 30786 4633
rect 30758 4606 30786 4607
rect 30534 4185 30562 4186
rect 30534 4159 30535 4185
rect 30535 4159 30561 4185
rect 30561 4159 30562 4185
rect 30534 4158 30562 4159
rect 30758 3374 30786 3402
rect 30758 3065 30786 3066
rect 30758 3039 30759 3065
rect 30759 3039 30785 3065
rect 30785 3039 30786 3065
rect 30758 3038 30786 3039
rect 30926 3430 30954 3458
rect 31150 5334 31178 5362
rect 31150 5166 31178 5194
rect 31150 4942 31178 4970
rect 31318 5614 31346 5642
rect 31486 5641 31514 5642
rect 31486 5615 31487 5641
rect 31487 5615 31513 5641
rect 31513 5615 31514 5641
rect 31486 5614 31514 5615
rect 31318 5390 31346 5418
rect 31318 4606 31346 4634
rect 31822 6286 31850 6314
rect 31710 6062 31738 6090
rect 31542 4886 31570 4914
rect 31598 5614 31626 5642
rect 31598 4830 31626 4858
rect 31710 4774 31738 4802
rect 31430 4718 31458 4746
rect 31374 4494 31402 4522
rect 31430 4270 31458 4298
rect 31206 4158 31234 4186
rect 31822 4102 31850 4130
rect 31542 4046 31570 4074
rect 31430 3822 31458 3850
rect 30982 3318 31010 3346
rect 30870 2982 30898 3010
rect 30646 2926 30674 2954
rect 30534 2617 30562 2618
rect 30534 2591 30535 2617
rect 30535 2591 30561 2617
rect 30561 2591 30562 2617
rect 30534 2590 30562 2591
rect 30926 2561 30954 2562
rect 30926 2535 30927 2561
rect 30927 2535 30953 2561
rect 30953 2535 30954 2561
rect 30926 2534 30954 2535
rect 31094 2478 31122 2506
rect 31150 2646 31178 2674
rect 30366 2198 30394 2226
rect 29918 1918 29946 1946
rect 29694 1889 29722 1890
rect 29694 1863 29695 1889
rect 29695 1863 29721 1889
rect 29721 1863 29722 1889
rect 29694 1862 29722 1863
rect 28686 1470 28714 1498
rect 29246 1358 29274 1386
rect 29414 1385 29442 1386
rect 29414 1359 29415 1385
rect 29415 1359 29441 1385
rect 29441 1359 29442 1385
rect 29414 1358 29442 1359
rect 29190 1329 29218 1330
rect 29190 1303 29191 1329
rect 29191 1303 29217 1329
rect 29217 1303 29218 1329
rect 29190 1302 29218 1303
rect 29134 1246 29162 1274
rect 28798 1190 28826 1218
rect 28798 1049 28826 1050
rect 28798 1023 28799 1049
rect 28799 1023 28825 1049
rect 28825 1023 28826 1049
rect 28798 1022 28826 1023
rect 28294 686 28322 714
rect 26334 406 26362 434
rect 27678 518 27706 546
rect 28854 742 28882 770
rect 28350 350 28378 378
rect 29246 1078 29274 1106
rect 29302 630 29330 658
rect 29638 1385 29666 1386
rect 29638 1359 29639 1385
rect 29639 1359 29665 1385
rect 29665 1359 29666 1385
rect 29638 1358 29666 1359
rect 30086 1302 30114 1330
rect 29974 993 30002 994
rect 29974 967 29975 993
rect 29975 967 30001 993
rect 30001 967 30002 993
rect 29974 966 30002 967
rect 29582 798 29610 826
rect 29526 294 29554 322
rect 30142 1049 30170 1050
rect 30142 1023 30143 1049
rect 30143 1023 30169 1049
rect 30169 1023 30170 1049
rect 30142 1022 30170 1023
rect 30310 1078 30338 1106
rect 30534 2030 30562 2058
rect 30254 574 30282 602
rect 30646 1806 30674 1834
rect 30926 1974 30954 2002
rect 30646 1721 30674 1722
rect 30646 1695 30647 1721
rect 30647 1695 30673 1721
rect 30673 1695 30674 1721
rect 30646 1694 30674 1695
rect 31430 3598 31458 3626
rect 31542 3150 31570 3178
rect 32102 3038 32130 3066
rect 31318 2702 31346 2730
rect 31262 2590 31290 2618
rect 31262 2254 31290 2282
rect 31542 2478 31570 2506
rect 31430 2030 31458 2058
rect 31206 1526 31234 1554
rect 31318 1694 31346 1722
rect 31094 1385 31122 1386
rect 31094 1359 31095 1385
rect 31095 1359 31121 1385
rect 31121 1359 31122 1385
rect 31094 1358 31122 1359
rect 31542 1582 31570 1610
rect 31318 1358 31346 1386
rect 30646 1329 30674 1330
rect 30646 1303 30647 1329
rect 30647 1303 30673 1329
rect 30673 1303 30674 1329
rect 30646 1302 30674 1303
rect 31374 1302 31402 1330
rect 30926 993 30954 994
rect 30926 967 30927 993
rect 30927 967 30953 993
rect 30953 967 30954 993
rect 30926 966 30954 967
rect 30646 881 30674 882
rect 30646 855 30647 881
rect 30647 855 30673 881
rect 30673 855 30674 881
rect 30646 854 30674 855
rect 30590 462 30618 490
rect 29806 238 29834 266
rect 31094 182 31122 210
rect 4774 14 4802 42
rect 31430 1134 31458 1162
rect 31542 910 31570 938
rect 31374 14 31402 42
<< metal3 >>
rect 6566 7014 14238 7042
rect 14266 7014 14271 7042
rect 0 6986 56 7000
rect 6566 6986 6594 7014
rect 32144 6986 32200 7000
rect 0 6958 126 6986
rect 154 6958 159 6986
rect 6561 6958 6566 6986
rect 6594 6958 6599 6986
rect 6673 6958 6678 6986
rect 6706 6958 14462 6986
rect 14490 6958 14495 6986
rect 16305 6958 16310 6986
rect 16338 6958 21630 6986
rect 21658 6958 21663 6986
rect 30417 6958 30422 6986
rect 30450 6958 32200 6986
rect 0 6944 56 6958
rect 32144 6944 32200 6958
rect 9865 6902 9870 6930
rect 9898 6902 16254 6930
rect 16282 6902 16287 6930
rect 22633 6902 22638 6930
rect 22666 6902 23646 6930
rect 23674 6902 23679 6930
rect 9809 6846 9814 6874
rect 9842 6846 18270 6874
rect 18298 6846 18303 6874
rect 19665 6846 19670 6874
rect 19698 6846 22078 6874
rect 22106 6846 22111 6874
rect 27449 6846 27454 6874
rect 27482 6846 28630 6874
rect 28658 6846 28663 6874
rect 1857 6790 1862 6818
rect 1890 6790 2814 6818
rect 2842 6790 2847 6818
rect 17593 6790 17598 6818
rect 17626 6790 23254 6818
rect 23282 6790 23287 6818
rect 0 6762 56 6776
rect 32144 6762 32200 6776
rect 0 6734 1694 6762
rect 1801 6734 1806 6762
rect 1834 6734 2366 6762
rect 2394 6734 2399 6762
rect 4881 6734 4886 6762
rect 4914 6734 5950 6762
rect 5978 6734 5983 6762
rect 6953 6734 6958 6762
rect 6986 6734 7518 6762
rect 7546 6734 7551 6762
rect 13561 6734 13566 6762
rect 13594 6734 13958 6762
rect 13986 6734 13991 6762
rect 21065 6734 21070 6762
rect 21098 6734 22302 6762
rect 22330 6734 22335 6762
rect 26553 6734 26558 6762
rect 26586 6734 27454 6762
rect 27482 6734 27487 6762
rect 27897 6734 27902 6762
rect 27930 6734 29414 6762
rect 29442 6734 29447 6762
rect 32097 6734 32102 6762
rect 32130 6734 32200 6762
rect 0 6720 56 6734
rect 1666 6706 1694 6734
rect 32144 6720 32200 6734
rect 1666 6678 2086 6706
rect 2114 6678 2119 6706
rect 13505 6678 13510 6706
rect 13538 6678 17486 6706
rect 17514 6678 17519 6706
rect 2227 6650 2232 6678
rect 2260 6650 2284 6678
rect 2312 6650 2336 6678
rect 2364 6650 2369 6678
rect 12227 6650 12232 6678
rect 12260 6650 12284 6678
rect 12312 6650 12336 6678
rect 12364 6650 12369 6678
rect 22227 6650 22232 6678
rect 22260 6650 22284 6678
rect 22312 6650 22336 6678
rect 22364 6650 22369 6678
rect 2977 6622 2982 6650
rect 3010 6622 3486 6650
rect 3514 6622 3519 6650
rect 3761 6622 3766 6650
rect 3794 6622 4382 6650
rect 4410 6622 4415 6650
rect 5665 6622 5670 6650
rect 5698 6622 6622 6650
rect 6650 6622 6655 6650
rect 8689 6622 8694 6650
rect 8722 6622 9758 6650
rect 9786 6622 9791 6650
rect 14905 6622 14910 6650
rect 14938 6622 16590 6650
rect 16618 6622 16623 6650
rect 16814 6622 20342 6650
rect 20370 6622 20375 6650
rect 1241 6566 1246 6594
rect 1274 6566 2142 6594
rect 2170 6566 2175 6594
rect 2590 6566 8554 6594
rect 9473 6566 9478 6594
rect 9506 6566 10430 6594
rect 10458 6566 10463 6594
rect 10593 6566 10598 6594
rect 10626 6566 11102 6594
rect 11130 6566 11135 6594
rect 11377 6566 11382 6594
rect 11410 6566 11998 6594
rect 12026 6566 12031 6594
rect 14569 6566 14574 6594
rect 14602 6566 15582 6594
rect 15610 6566 15615 6594
rect 15946 6566 16702 6594
rect 16730 6566 16735 6594
rect 0 6538 56 6552
rect 2590 6538 2618 6566
rect 8526 6538 8554 6566
rect 15946 6538 15974 6566
rect 0 6510 2618 6538
rect 7457 6510 7462 6538
rect 7490 6510 8414 6538
rect 8442 6510 8447 6538
rect 8526 6510 9646 6538
rect 9674 6510 9679 6538
rect 14905 6510 14910 6538
rect 14938 6510 15974 6538
rect 0 6496 56 6510
rect 16814 6482 16842 6622
rect 16921 6566 16926 6594
rect 16954 6566 18270 6594
rect 18298 6566 18303 6594
rect 25657 6566 25662 6594
rect 25690 6566 26054 6594
rect 26082 6566 26087 6594
rect 27225 6566 27230 6594
rect 27258 6566 28238 6594
rect 28266 6566 28271 6594
rect 29465 6566 29470 6594
rect 29498 6566 31262 6594
rect 31290 6566 31295 6594
rect 32144 6538 32200 6552
rect 16921 6510 16926 6538
rect 16954 6510 21854 6538
rect 26329 6510 26334 6538
rect 26362 6510 27062 6538
rect 27090 6510 27095 6538
rect 28569 6510 28574 6538
rect 28602 6510 30254 6538
rect 30282 6510 30287 6538
rect 31537 6510 31542 6538
rect 31570 6510 32200 6538
rect 21826 6482 21854 6510
rect 32144 6496 32200 6510
rect 5945 6454 5950 6482
rect 5978 6454 7350 6482
rect 7378 6454 7383 6482
rect 7513 6454 7518 6482
rect 7546 6454 7966 6482
rect 7994 6454 7999 6482
rect 9753 6454 9758 6482
rect 9786 6454 16842 6482
rect 17145 6454 17150 6482
rect 17178 6454 20846 6482
rect 20874 6454 20879 6482
rect 21826 6454 26054 6482
rect 26082 6454 26087 6482
rect 27673 6454 27678 6482
rect 27706 6454 28238 6482
rect 28266 6454 28271 6482
rect 29017 6454 29022 6482
rect 29050 6454 30310 6482
rect 30338 6454 30343 6482
rect 1073 6398 1078 6426
rect 1106 6398 6454 6426
rect 6482 6398 6487 6426
rect 9697 6398 9702 6426
rect 9730 6398 12194 6426
rect 13617 6398 13622 6426
rect 13650 6398 15862 6426
rect 15890 6398 15895 6426
rect 16249 6398 16254 6426
rect 16282 6398 18550 6426
rect 18578 6398 18583 6426
rect 20785 6398 20790 6426
rect 20818 6398 22526 6426
rect 22554 6398 22559 6426
rect 26553 6398 26558 6426
rect 26586 6398 30982 6426
rect 31010 6398 31015 6426
rect 12166 6370 12194 6398
rect 10929 6342 10934 6370
rect 10962 6342 12138 6370
rect 12166 6342 15414 6370
rect 15442 6342 15447 6370
rect 15577 6342 15582 6370
rect 15610 6342 21854 6370
rect 21882 6342 21887 6370
rect 26609 6342 26614 6370
rect 26642 6342 29806 6370
rect 29834 6342 29839 6370
rect 29913 6342 29918 6370
rect 29946 6342 30590 6370
rect 30618 6342 30623 6370
rect 0 6314 56 6328
rect 12110 6314 12138 6342
rect 32144 6314 32200 6328
rect 0 6286 182 6314
rect 210 6286 215 6314
rect 5161 6286 5166 6314
rect 5194 6286 6678 6314
rect 6706 6286 6711 6314
rect 12110 6286 15694 6314
rect 15722 6286 15727 6314
rect 15857 6286 15862 6314
rect 15890 6286 16702 6314
rect 16730 6286 16735 6314
rect 16809 6286 16814 6314
rect 16842 6286 19166 6314
rect 19194 6286 19199 6314
rect 28345 6286 28350 6314
rect 28378 6286 29022 6314
rect 29050 6286 29055 6314
rect 31817 6286 31822 6314
rect 31850 6286 32200 6314
rect 0 6272 56 6286
rect 1897 6258 1902 6286
rect 1930 6258 1954 6286
rect 1982 6258 2006 6286
rect 2034 6258 2039 6286
rect 11897 6258 11902 6286
rect 11930 6258 11954 6286
rect 11982 6258 12006 6286
rect 12034 6258 12039 6286
rect 21897 6258 21902 6286
rect 21930 6258 21954 6286
rect 21982 6258 22006 6286
rect 22034 6258 22039 6286
rect 32144 6272 32200 6286
rect 12217 6230 12222 6258
rect 12250 6230 13790 6258
rect 13818 6230 13823 6258
rect 14345 6230 14350 6258
rect 14378 6230 17430 6258
rect 17458 6230 17463 6258
rect 29241 6230 29246 6258
rect 29274 6230 29806 6258
rect 29834 6230 29839 6258
rect 4265 6174 4270 6202
rect 4298 6174 4830 6202
rect 4858 6174 4863 6202
rect 5049 6174 5054 6202
rect 5082 6174 5278 6202
rect 5306 6174 5311 6202
rect 5833 6174 5838 6202
rect 5866 6174 6398 6202
rect 6426 6174 6431 6202
rect 8185 6174 8190 6202
rect 8218 6174 8638 6202
rect 8666 6174 8671 6202
rect 8969 6174 8974 6202
rect 9002 6174 9534 6202
rect 9562 6174 9567 6202
rect 11153 6174 11158 6202
rect 11186 6174 14070 6202
rect 14098 6174 14103 6202
rect 15017 6174 15022 6202
rect 15050 6174 17206 6202
rect 17234 6174 17239 6202
rect 17313 6174 17318 6202
rect 17346 6174 21854 6202
rect 25881 6174 25886 6202
rect 25914 6174 26278 6202
rect 26306 6174 26311 6202
rect 27001 6174 27006 6202
rect 27034 6174 27846 6202
rect 27874 6174 27879 6202
rect 21826 6146 21854 6174
rect 13113 6118 13118 6146
rect 13146 6118 13454 6146
rect 13482 6118 13487 6146
rect 14457 6118 14462 6146
rect 14490 6118 15190 6146
rect 15218 6118 15223 6146
rect 15297 6118 15302 6146
rect 15330 6118 20286 6146
rect 20314 6118 20319 6146
rect 21826 6118 26670 6146
rect 26698 6118 26703 6146
rect 28121 6118 28126 6146
rect 28154 6118 28574 6146
rect 28602 6118 28607 6146
rect 28793 6118 28798 6146
rect 28826 6118 29414 6146
rect 29442 6118 29447 6146
rect 29689 6118 29694 6146
rect 29722 6118 31094 6146
rect 31122 6118 31127 6146
rect 0 6090 56 6104
rect 32144 6090 32200 6104
rect 0 6062 798 6090
rect 826 6062 831 6090
rect 6897 6062 6902 6090
rect 6930 6062 9422 6090
rect 9450 6062 9455 6090
rect 11601 6062 11606 6090
rect 11634 6062 13790 6090
rect 13818 6062 13823 6090
rect 14289 6062 14294 6090
rect 14322 6062 16254 6090
rect 16282 6062 16287 6090
rect 16361 6062 16366 6090
rect 16394 6062 18718 6090
rect 18746 6062 18751 6090
rect 20673 6062 20678 6090
rect 20706 6062 26782 6090
rect 26810 6062 26815 6090
rect 31705 6062 31710 6090
rect 31738 6062 32200 6090
rect 0 6048 56 6062
rect 32144 6048 32200 6062
rect 2529 6006 2534 6034
rect 2562 6006 5838 6034
rect 5866 6006 5871 6034
rect 8465 6006 8470 6034
rect 8498 6006 9590 6034
rect 9618 6006 9623 6034
rect 10425 6006 10430 6034
rect 10458 6006 14294 6034
rect 14322 6006 14327 6034
rect 15241 6006 15246 6034
rect 15274 6006 16254 6034
rect 16282 6006 16287 6034
rect 16366 6006 17094 6034
rect 17122 6006 17127 6034
rect 18942 6006 20286 6034
rect 20314 6006 20398 6034
rect 20426 6006 20431 6034
rect 21793 6006 21798 6034
rect 21826 6006 27174 6034
rect 27202 6006 27207 6034
rect 16366 5978 16394 6006
rect 2193 5950 2198 5978
rect 2226 5950 3346 5978
rect 6281 5950 6286 5978
rect 6314 5950 10094 5978
rect 0 5866 56 5880
rect 2227 5866 2232 5894
rect 2260 5866 2284 5894
rect 2312 5866 2336 5894
rect 2364 5866 2369 5894
rect 3318 5866 3346 5950
rect 4545 5894 4550 5922
rect 4578 5894 8750 5922
rect 8778 5894 8783 5922
rect 10066 5866 10094 5950
rect 12166 5950 14518 5978
rect 14546 5950 14630 5978
rect 14658 5950 14663 5978
rect 15185 5950 15190 5978
rect 15218 5950 16394 5978
rect 16473 5950 16478 5978
rect 16506 5950 17598 5978
rect 17626 5950 17631 5978
rect 12166 5866 12194 5950
rect 12497 5894 12502 5922
rect 12530 5894 14294 5922
rect 14322 5894 14327 5922
rect 14401 5894 14406 5922
rect 14434 5894 15806 5922
rect 15834 5894 15839 5922
rect 15913 5894 15918 5922
rect 15946 5894 16982 5922
rect 17010 5894 17015 5922
rect 17369 5894 17374 5922
rect 17402 5894 17990 5922
rect 18018 5894 18023 5922
rect 12227 5866 12232 5894
rect 12260 5866 12284 5894
rect 12312 5866 12336 5894
rect 12364 5866 12369 5894
rect 18942 5866 18970 6006
rect 20001 5950 20006 5978
rect 20034 5950 21406 5978
rect 21434 5950 21518 5978
rect 21546 5950 21551 5978
rect 23361 5950 23366 5978
rect 23394 5950 25914 5978
rect 19049 5894 19054 5922
rect 19082 5894 20734 5922
rect 20762 5894 20767 5922
rect 22577 5894 22582 5922
rect 22610 5894 22974 5922
rect 23002 5894 23007 5922
rect 23305 5894 23310 5922
rect 23338 5894 25774 5922
rect 25802 5894 25807 5922
rect 22227 5866 22232 5894
rect 22260 5866 22284 5894
rect 22312 5866 22336 5894
rect 22364 5866 22369 5894
rect 25886 5866 25914 5950
rect 32144 5866 32200 5880
rect 0 5838 1778 5866
rect 3318 5838 4102 5866
rect 4130 5838 4135 5866
rect 10066 5838 12194 5866
rect 13337 5838 13342 5866
rect 13370 5838 15582 5866
rect 15610 5838 15615 5866
rect 15689 5838 15694 5866
rect 15722 5838 17150 5866
rect 17178 5838 17183 5866
rect 17257 5838 17262 5866
rect 17290 5838 18970 5866
rect 25886 5838 29134 5866
rect 29162 5838 29167 5866
rect 31201 5838 31206 5866
rect 31234 5838 32200 5866
rect 0 5824 56 5838
rect 1750 5754 1778 5838
rect 32144 5824 32200 5838
rect 2305 5782 2310 5810
rect 2338 5782 2590 5810
rect 2618 5782 2623 5810
rect 3873 5782 3878 5810
rect 3906 5782 4158 5810
rect 4186 5782 4191 5810
rect 5441 5782 5446 5810
rect 5474 5782 5726 5810
rect 5754 5782 5759 5810
rect 7233 5782 7238 5810
rect 7266 5782 13510 5810
rect 13538 5782 13543 5810
rect 13785 5782 13790 5810
rect 13818 5782 21854 5810
rect 26833 5782 26838 5810
rect 26866 5782 27286 5810
rect 27314 5782 27319 5810
rect 21826 5754 21854 5782
rect 793 5726 798 5754
rect 826 5726 1694 5754
rect 1750 5726 9170 5754
rect 9361 5726 9366 5754
rect 9394 5726 17038 5754
rect 17066 5726 17071 5754
rect 17145 5726 17150 5754
rect 17178 5726 19614 5754
rect 19642 5726 19647 5754
rect 21826 5726 22806 5754
rect 22834 5726 22839 5754
rect 23081 5726 23086 5754
rect 23114 5726 26558 5754
rect 26586 5726 26591 5754
rect 1666 5698 1694 5726
rect 9142 5698 9170 5726
rect 1666 5670 2478 5698
rect 2506 5670 2511 5698
rect 4153 5670 4158 5698
rect 4186 5670 6230 5698
rect 6258 5670 6263 5698
rect 7401 5670 7406 5698
rect 7434 5670 9030 5698
rect 9058 5670 9063 5698
rect 9142 5670 9422 5698
rect 9450 5670 9455 5698
rect 10649 5670 10654 5698
rect 10682 5670 12614 5698
rect 12642 5670 12647 5698
rect 13617 5670 13622 5698
rect 13650 5670 15638 5698
rect 15666 5670 15671 5698
rect 17873 5670 17878 5698
rect 17906 5670 26222 5698
rect 26250 5670 26255 5698
rect 28625 5670 28630 5698
rect 28658 5670 29526 5698
rect 29554 5670 29559 5698
rect 0 5642 56 5656
rect 32144 5642 32200 5656
rect 0 5614 882 5642
rect 961 5614 966 5642
rect 994 5614 8638 5642
rect 8666 5614 8671 5642
rect 8745 5614 8750 5642
rect 8778 5614 13510 5642
rect 13538 5614 13543 5642
rect 14233 5614 14238 5642
rect 14266 5614 16310 5642
rect 16338 5614 16343 5642
rect 17481 5614 17486 5642
rect 17514 5614 19838 5642
rect 19866 5614 19871 5642
rect 20169 5614 20174 5642
rect 20202 5614 20510 5642
rect 20538 5614 20543 5642
rect 21121 5614 21126 5642
rect 21154 5614 22946 5642
rect 23249 5614 23254 5642
rect 23282 5614 24962 5642
rect 26049 5614 26054 5642
rect 26082 5614 31318 5642
rect 31346 5614 31486 5642
rect 31514 5614 31519 5642
rect 31593 5614 31598 5642
rect 31626 5614 32200 5642
rect 0 5600 56 5614
rect 854 5586 882 5614
rect 854 5558 2142 5586
rect 2170 5558 2175 5586
rect 3145 5558 3150 5586
rect 3178 5558 6734 5586
rect 6762 5558 6767 5586
rect 11993 5558 11998 5586
rect 12026 5558 13146 5586
rect 14289 5558 14294 5586
rect 14322 5558 22414 5586
rect 22442 5558 22447 5586
rect 13118 5530 13146 5558
rect 2193 5502 2198 5530
rect 2226 5502 9310 5530
rect 9338 5502 9343 5530
rect 13113 5502 13118 5530
rect 13146 5502 13151 5530
rect 13449 5502 13454 5530
rect 13482 5502 14686 5530
rect 14714 5502 14719 5530
rect 17033 5502 17038 5530
rect 17066 5502 19278 5530
rect 19306 5502 19311 5530
rect 1897 5474 1902 5502
rect 1930 5474 1954 5502
rect 1982 5474 2006 5502
rect 2034 5474 2039 5502
rect 11897 5474 11902 5502
rect 11930 5474 11954 5502
rect 11982 5474 12006 5502
rect 12034 5474 12039 5502
rect 21897 5474 21902 5502
rect 21930 5474 21954 5502
rect 21982 5474 22006 5502
rect 22034 5474 22039 5502
rect 22918 5474 22946 5614
rect 23361 5558 23366 5586
rect 23394 5558 23478 5586
rect 23506 5558 23511 5586
rect 24934 5474 24962 5614
rect 32144 5600 32200 5614
rect 27673 5502 27678 5530
rect 27706 5502 30422 5530
rect 30450 5502 30455 5530
rect 5833 5446 5838 5474
rect 5866 5446 11858 5474
rect 14177 5446 14182 5474
rect 14210 5446 17598 5474
rect 17626 5446 17631 5474
rect 22918 5446 24402 5474
rect 24934 5446 28462 5474
rect 28490 5446 28495 5474
rect 0 5418 56 5432
rect 11830 5418 11858 5446
rect 24374 5418 24402 5446
rect 32144 5418 32200 5432
rect 0 5390 1246 5418
rect 1274 5390 1279 5418
rect 1353 5390 1358 5418
rect 1386 5390 6006 5418
rect 6034 5390 6039 5418
rect 7737 5390 7742 5418
rect 7770 5390 8134 5418
rect 8162 5390 8167 5418
rect 10817 5390 10822 5418
rect 10850 5390 11102 5418
rect 11130 5390 11135 5418
rect 11830 5390 12502 5418
rect 12530 5390 12535 5418
rect 12609 5390 12614 5418
rect 12642 5390 14574 5418
rect 14602 5390 14607 5418
rect 16249 5390 16254 5418
rect 16282 5390 18326 5418
rect 18354 5390 18359 5418
rect 19329 5390 19334 5418
rect 19362 5390 24262 5418
rect 24290 5390 24295 5418
rect 24374 5390 29470 5418
rect 29498 5390 29503 5418
rect 31313 5390 31318 5418
rect 31346 5390 32200 5418
rect 0 5376 56 5390
rect 32144 5376 32200 5390
rect 4545 5334 4550 5362
rect 4578 5334 5950 5362
rect 5978 5334 5983 5362
rect 9641 5334 9646 5362
rect 9674 5334 10654 5362
rect 10682 5334 10687 5362
rect 10761 5334 10766 5362
rect 10794 5334 16226 5362
rect 16305 5334 16310 5362
rect 16338 5334 23310 5362
rect 23338 5334 23343 5362
rect 23473 5334 23478 5362
rect 23506 5334 25550 5362
rect 25578 5334 25583 5362
rect 25713 5334 25718 5362
rect 25746 5334 31150 5362
rect 31178 5334 31183 5362
rect 16198 5306 16226 5334
rect 5329 5278 5334 5306
rect 5362 5278 6342 5306
rect 6370 5278 6375 5306
rect 6505 5278 6510 5306
rect 6538 5278 16086 5306
rect 16114 5278 16119 5306
rect 16198 5278 16646 5306
rect 16674 5278 16679 5306
rect 18886 5278 29022 5306
rect 29050 5278 29055 5306
rect 18886 5250 18914 5278
rect 3313 5222 3318 5250
rect 3346 5222 6398 5250
rect 6426 5222 6431 5250
rect 7681 5222 7686 5250
rect 7714 5222 8246 5250
rect 8274 5222 8279 5250
rect 11433 5222 11438 5250
rect 11466 5222 14630 5250
rect 14658 5222 14663 5250
rect 15913 5222 15918 5250
rect 15946 5222 18914 5250
rect 21793 5222 21798 5250
rect 21826 5222 27006 5250
rect 27034 5222 27039 5250
rect 28065 5222 28070 5250
rect 28098 5222 29526 5250
rect 29554 5222 29559 5250
rect 0 5194 56 5208
rect 32144 5194 32200 5208
rect 0 5166 3710 5194
rect 3738 5166 3743 5194
rect 5894 5166 14238 5194
rect 14266 5166 14271 5194
rect 16081 5166 16086 5194
rect 16114 5166 17542 5194
rect 17570 5166 17575 5194
rect 21009 5166 21014 5194
rect 21042 5166 24318 5194
rect 24346 5166 24351 5194
rect 31145 5166 31150 5194
rect 31178 5166 32200 5194
rect 0 5152 56 5166
rect 2227 5082 2232 5110
rect 2260 5082 2284 5110
rect 2312 5082 2336 5110
rect 2364 5082 2369 5110
rect 2585 5054 2590 5082
rect 2618 5054 4942 5082
rect 4970 5054 4975 5082
rect 5894 5026 5922 5166
rect 32144 5152 32200 5166
rect 6729 5110 6734 5138
rect 6762 5110 10542 5138
rect 10570 5110 10575 5138
rect 12609 5110 12614 5138
rect 12642 5110 13622 5138
rect 13650 5110 13655 5138
rect 13729 5110 13734 5138
rect 13762 5110 14966 5138
rect 14994 5110 14999 5138
rect 17313 5110 17318 5138
rect 17346 5110 19558 5138
rect 19586 5110 19591 5138
rect 23641 5110 23646 5138
rect 23674 5110 25718 5138
rect 25746 5110 25751 5138
rect 12227 5082 12232 5110
rect 12260 5082 12284 5110
rect 12312 5082 12336 5110
rect 12364 5082 12369 5110
rect 22227 5082 22232 5110
rect 22260 5082 22284 5110
rect 22312 5082 22336 5110
rect 22364 5082 22369 5110
rect 6113 5054 6118 5082
rect 6146 5054 7294 5082
rect 7322 5054 7327 5082
rect 12497 5054 12502 5082
rect 12530 5054 14322 5082
rect 16081 5054 16086 5082
rect 16114 5054 18214 5082
rect 18242 5054 18247 5082
rect 18489 5054 18494 5082
rect 18522 5054 21854 5082
rect 22409 5054 22414 5082
rect 22442 5054 24878 5082
rect 24906 5054 24911 5082
rect 26894 5054 28238 5082
rect 28266 5054 28271 5082
rect 30753 5054 30758 5082
rect 30786 5054 31346 5082
rect 14294 5026 14322 5054
rect 21826 5026 21854 5054
rect 26894 5026 26922 5054
rect 4153 4998 4158 5026
rect 4186 4998 5922 5026
rect 6001 4998 6006 5026
rect 6034 4998 9366 5026
rect 9394 4998 9399 5026
rect 10873 4998 10878 5026
rect 10906 4998 14182 5026
rect 14210 4998 14215 5026
rect 14294 4998 17318 5026
rect 17346 4998 17351 5026
rect 17425 4998 17430 5026
rect 17458 4998 19334 5026
rect 19362 4998 19367 5026
rect 21826 4998 23142 5026
rect 23170 4998 23175 5026
rect 24089 4998 24094 5026
rect 24122 4998 26922 5026
rect 27113 4998 27118 5026
rect 27146 4998 28742 5026
rect 28770 4998 28775 5026
rect 29073 4998 29078 5026
rect 29106 4998 30702 5026
rect 30730 4998 30735 5026
rect 0 4970 56 4984
rect 31318 4970 31346 5054
rect 32144 4970 32200 4984
rect 0 4942 5894 4970
rect 5922 4942 5927 4970
rect 11769 4942 11774 4970
rect 11802 4942 15190 4970
rect 15218 4942 15223 4970
rect 16137 4942 16142 4970
rect 16170 4942 17374 4970
rect 17402 4942 17407 4970
rect 19385 4942 19390 4970
rect 19418 4942 30142 4970
rect 30170 4942 30175 4970
rect 30529 4942 30534 4970
rect 30562 4942 31150 4970
rect 31178 4942 31183 4970
rect 31318 4942 32200 4970
rect 0 4928 56 4942
rect 32144 4928 32200 4942
rect 7513 4886 7518 4914
rect 7546 4886 10990 4914
rect 11018 4886 11023 4914
rect 11097 4886 11102 4914
rect 11130 4886 15470 4914
rect 15498 4886 15503 4914
rect 15577 4886 15582 4914
rect 15610 4886 16646 4914
rect 16674 4886 16679 4914
rect 17593 4886 17598 4914
rect 17626 4886 29414 4914
rect 29442 4886 29447 4914
rect 29750 4886 31542 4914
rect 31570 4886 31575 4914
rect 29750 4858 29778 4886
rect 5777 4830 5782 4858
rect 5810 4830 13398 4858
rect 13426 4830 13431 4858
rect 13897 4830 13902 4858
rect 13930 4830 14294 4858
rect 14322 4830 14327 4858
rect 14401 4830 14406 4858
rect 14434 4830 15862 4858
rect 15890 4830 15895 4858
rect 16921 4830 16926 4858
rect 16954 4830 20062 4858
rect 20090 4830 20095 4858
rect 20281 4830 20286 4858
rect 20314 4830 27734 4858
rect 27762 4830 27958 4858
rect 27986 4830 27991 4858
rect 28961 4830 28966 4858
rect 28994 4830 29778 4858
rect 29857 4830 29862 4858
rect 29890 4830 31598 4858
rect 31626 4830 31631 4858
rect 1666 4774 3318 4802
rect 3346 4774 3351 4802
rect 11830 4774 17150 4802
rect 17178 4774 17183 4802
rect 17537 4774 17542 4802
rect 17570 4774 20454 4802
rect 20482 4774 20487 4802
rect 29353 4774 29358 4802
rect 29386 4774 31710 4802
rect 31738 4774 31743 4802
rect 0 4746 56 4760
rect 1666 4746 1694 4774
rect 0 4718 1694 4746
rect 5049 4718 5054 4746
rect 5082 4718 10710 4746
rect 10738 4718 10743 4746
rect 0 4704 56 4718
rect 1897 4690 1902 4718
rect 1930 4690 1954 4718
rect 1982 4690 2006 4718
rect 2034 4690 2039 4718
rect 11830 4690 11858 4774
rect 32144 4746 32200 4760
rect 12721 4718 12726 4746
rect 12754 4718 13902 4746
rect 13930 4718 13935 4746
rect 14009 4718 14014 4746
rect 14042 4718 16758 4746
rect 16786 4718 16791 4746
rect 31425 4718 31430 4746
rect 31458 4718 32200 4746
rect 11897 4690 11902 4718
rect 11930 4690 11954 4718
rect 11982 4690 12006 4718
rect 12034 4690 12039 4718
rect 21897 4690 21902 4718
rect 21930 4690 21954 4718
rect 21982 4690 22006 4718
rect 22034 4690 22039 4718
rect 32144 4704 32200 4718
rect 8913 4662 8918 4690
rect 8946 4662 11858 4690
rect 12105 4662 12110 4690
rect 12138 4662 13342 4690
rect 13370 4662 13375 4690
rect 14233 4662 14238 4690
rect 14266 4662 19390 4690
rect 19418 4662 19423 4690
rect 20729 4662 20734 4690
rect 20762 4662 21854 4690
rect 21826 4634 21854 4662
rect 1302 4606 7182 4634
rect 7210 4606 7215 4634
rect 10985 4606 10990 4634
rect 11018 4606 14742 4634
rect 14770 4606 14775 4634
rect 15129 4606 15134 4634
rect 15162 4606 21014 4634
rect 21042 4606 21047 4634
rect 21826 4606 23702 4634
rect 23730 4606 23735 4634
rect 30753 4606 30758 4634
rect 30786 4606 31318 4634
rect 31346 4606 31351 4634
rect 0 4522 56 4536
rect 1302 4522 1330 4606
rect 1409 4550 1414 4578
rect 1442 4550 6902 4578
rect 6930 4550 6935 4578
rect 7065 4550 7070 4578
rect 7098 4550 7462 4578
rect 7490 4550 7495 4578
rect 7681 4550 7686 4578
rect 7714 4550 11438 4578
rect 11466 4550 11471 4578
rect 13169 4550 13174 4578
rect 13202 4550 20230 4578
rect 20258 4550 20263 4578
rect 20617 4550 20622 4578
rect 20650 4550 22582 4578
rect 22610 4550 22615 4578
rect 26665 4550 26670 4578
rect 26698 4550 28350 4578
rect 28378 4550 28383 4578
rect 32144 4522 32200 4536
rect 0 4494 1330 4522
rect 2193 4494 2198 4522
rect 2226 4494 2478 4522
rect 2506 4494 2511 4522
rect 6225 4494 6230 4522
rect 6258 4494 14518 4522
rect 14546 4494 14551 4522
rect 14681 4494 14686 4522
rect 14714 4494 15246 4522
rect 15274 4494 15279 4522
rect 18041 4494 18046 4522
rect 18074 4494 26222 4522
rect 26250 4494 26390 4522
rect 26418 4494 26423 4522
rect 31369 4494 31374 4522
rect 31402 4494 32200 4522
rect 0 4480 56 4494
rect 32144 4480 32200 4494
rect 2753 4438 2758 4466
rect 2786 4438 14182 4466
rect 14210 4438 14215 4466
rect 14294 4438 26670 4466
rect 26698 4438 26703 4466
rect 28233 4438 28238 4466
rect 28266 4438 30142 4466
rect 30170 4438 30175 4466
rect 14294 4410 14322 4438
rect 1633 4382 1638 4410
rect 1666 4382 1750 4410
rect 1778 4382 3626 4410
rect 7457 4382 7462 4410
rect 7490 4382 9702 4410
rect 9730 4382 9735 4410
rect 10201 4382 10206 4410
rect 10234 4382 12502 4410
rect 12530 4382 12535 4410
rect 13505 4382 13510 4410
rect 13538 4382 14322 4410
rect 15409 4382 15414 4410
rect 15442 4382 18046 4410
rect 18074 4382 18079 4410
rect 18265 4382 18270 4410
rect 18298 4382 24794 4410
rect 25993 4382 25998 4410
rect 26026 4382 28406 4410
rect 28434 4382 28574 4410
rect 28602 4382 28607 4410
rect 3598 4354 3626 4382
rect 24766 4354 24794 4382
rect 3598 4326 9814 4354
rect 9842 4326 9847 4354
rect 10425 4326 10430 4354
rect 10458 4326 12110 4354
rect 12138 4326 12143 4354
rect 13225 4326 13230 4354
rect 13258 4326 15974 4354
rect 16753 4326 16758 4354
rect 16786 4326 19278 4354
rect 19306 4326 19311 4354
rect 24766 4326 27958 4354
rect 27986 4326 28126 4354
rect 28154 4326 28159 4354
rect 0 4298 56 4312
rect 2227 4298 2232 4326
rect 2260 4298 2284 4326
rect 2312 4298 2336 4326
rect 2364 4298 2369 4326
rect 12227 4298 12232 4326
rect 12260 4298 12284 4326
rect 12312 4298 12336 4326
rect 12364 4298 12369 4326
rect 15946 4298 15974 4326
rect 22227 4298 22232 4326
rect 22260 4298 22284 4326
rect 22312 4298 22336 4326
rect 22364 4298 22369 4326
rect 32144 4298 32200 4312
rect 0 4270 1694 4298
rect 3257 4270 3262 4298
rect 3290 4270 5670 4298
rect 5698 4270 5703 4298
rect 9249 4270 9254 4298
rect 9282 4270 12110 4298
rect 12138 4270 12143 4298
rect 13617 4270 13622 4298
rect 13650 4270 15694 4298
rect 15722 4270 15727 4298
rect 15946 4270 17878 4298
rect 17906 4270 17911 4298
rect 18265 4270 18270 4298
rect 18298 4270 20902 4298
rect 20930 4270 20935 4298
rect 22409 4270 22414 4298
rect 22442 4270 24206 4298
rect 24234 4270 24239 4298
rect 31425 4270 31430 4298
rect 31458 4270 32200 4298
rect 0 4256 56 4270
rect 1666 4242 1694 4270
rect 32144 4256 32200 4270
rect 1666 4214 6734 4242
rect 6762 4214 6767 4242
rect 10985 4214 10990 4242
rect 11018 4214 14238 4242
rect 14266 4214 14271 4242
rect 15129 4214 15134 4242
rect 15162 4214 17038 4242
rect 17066 4214 17071 4242
rect 18438 4214 29134 4242
rect 29162 4214 29167 4242
rect 18438 4186 18466 4214
rect 3985 4158 3990 4186
rect 4018 4158 7126 4186
rect 7154 4158 7159 4186
rect 9193 4158 9198 4186
rect 9226 4158 11662 4186
rect 11690 4158 11695 4186
rect 12105 4158 12110 4186
rect 12138 4158 12866 4186
rect 14177 4158 14182 4186
rect 14210 4158 15078 4186
rect 15106 4158 15111 4186
rect 15190 4158 17626 4186
rect 18433 4158 18438 4186
rect 18466 4158 18471 4186
rect 19273 4158 19278 4186
rect 19306 4158 23646 4186
rect 23674 4158 23679 4186
rect 28233 4158 28238 4186
rect 28266 4158 30254 4186
rect 30282 4158 30287 4186
rect 30529 4158 30534 4186
rect 30562 4158 31206 4186
rect 31234 4158 31239 4186
rect 12838 4130 12866 4158
rect 15190 4130 15218 4158
rect 17598 4130 17626 4158
rect 121 4102 126 4130
rect 154 4102 12726 4130
rect 12754 4102 12759 4130
rect 12838 4102 15218 4130
rect 15801 4102 15806 4130
rect 15834 4102 17486 4130
rect 17514 4102 17519 4130
rect 17598 4102 28742 4130
rect 28770 4102 28775 4130
rect 29857 4102 29862 4130
rect 29890 4102 31822 4130
rect 31850 4102 31855 4130
rect 0 4074 56 4088
rect 32144 4074 32200 4088
rect 0 4046 462 4074
rect 490 4046 495 4074
rect 5385 4046 5390 4074
rect 5418 4046 9254 4074
rect 9282 4046 9287 4074
rect 9361 4046 9366 4074
rect 9394 4046 13846 4074
rect 13874 4046 13879 4074
rect 14625 4046 14630 4074
rect 14658 4046 17038 4074
rect 17066 4046 17071 4074
rect 17145 4046 17150 4074
rect 17178 4046 18382 4074
rect 18410 4046 18415 4074
rect 18489 4046 18494 4074
rect 18522 4046 23366 4074
rect 23394 4046 23399 4074
rect 31537 4046 31542 4074
rect 31570 4046 32200 4074
rect 0 4032 56 4046
rect 32144 4032 32200 4046
rect 5889 3990 5894 4018
rect 5922 3990 9282 4018
rect 9254 3962 9282 3990
rect 10066 3990 13006 4018
rect 13034 3990 13039 4018
rect 13897 3990 13902 4018
rect 13930 3990 15414 4018
rect 15442 3990 15447 4018
rect 16697 3990 16702 4018
rect 16730 3990 20286 4018
rect 20314 3990 20319 4018
rect 21009 3990 21014 4018
rect 21042 3990 21126 4018
rect 21154 3990 21159 4018
rect 21737 3990 21742 4018
rect 21770 3990 28630 4018
rect 28658 3990 28663 4018
rect 10066 3962 10094 3990
rect 2641 3934 2646 3962
rect 2674 3934 7518 3962
rect 7546 3934 7551 3962
rect 9254 3934 10094 3962
rect 12553 3934 12558 3962
rect 12586 3934 14070 3962
rect 14098 3934 14103 3962
rect 14457 3934 14462 3962
rect 14490 3934 17262 3962
rect 17290 3934 17295 3962
rect 17481 3934 17486 3962
rect 17514 3934 20958 3962
rect 20986 3934 20991 3962
rect 22633 3934 22638 3962
rect 22666 3934 27734 3962
rect 27762 3934 27958 3962
rect 27986 3934 27991 3962
rect 1897 3906 1902 3934
rect 1930 3906 1954 3934
rect 1982 3906 2006 3934
rect 2034 3906 2039 3934
rect 11897 3906 11902 3934
rect 11930 3906 11954 3934
rect 11982 3906 12006 3934
rect 12034 3906 12039 3934
rect 21897 3906 21902 3934
rect 21930 3906 21954 3934
rect 21982 3906 22006 3934
rect 22034 3906 22039 3934
rect 3649 3878 3654 3906
rect 3682 3878 4998 3906
rect 5026 3878 5031 3906
rect 9305 3878 9310 3906
rect 9338 3878 10486 3906
rect 10514 3878 10519 3906
rect 12105 3878 12110 3906
rect 12138 3878 15134 3906
rect 15162 3878 15167 3906
rect 16641 3878 16646 3906
rect 16674 3878 21238 3906
rect 21266 3878 21271 3906
rect 0 3850 56 3864
rect 32144 3850 32200 3864
rect 0 3822 10822 3850
rect 10850 3822 10855 3850
rect 13729 3822 13734 3850
rect 13762 3822 14350 3850
rect 14378 3822 14383 3850
rect 15577 3822 15582 3850
rect 15610 3822 16926 3850
rect 16954 3822 16959 3850
rect 17593 3822 17598 3850
rect 17626 3822 19222 3850
rect 19250 3822 19255 3850
rect 19329 3822 19334 3850
rect 19362 3822 20174 3850
rect 20202 3822 20207 3850
rect 20897 3822 20902 3850
rect 20930 3822 25998 3850
rect 26026 3822 26031 3850
rect 31425 3822 31430 3850
rect 31458 3822 32200 3850
rect 0 3808 56 3822
rect 32144 3808 32200 3822
rect 1241 3766 1246 3794
rect 1274 3766 6734 3794
rect 6762 3766 6767 3794
rect 8801 3766 8806 3794
rect 8834 3766 16030 3794
rect 16058 3766 16063 3794
rect 16585 3766 16590 3794
rect 16618 3766 17262 3794
rect 17290 3766 17295 3794
rect 17817 3766 17822 3794
rect 17850 3766 17934 3794
rect 17962 3766 17967 3794
rect 18209 3766 18214 3794
rect 18242 3766 19278 3794
rect 19306 3766 19311 3794
rect 19385 3766 19390 3794
rect 19418 3766 20958 3794
rect 20986 3766 20991 3794
rect 21121 3766 21126 3794
rect 21154 3766 21238 3794
rect 21266 3766 23198 3794
rect 23226 3766 23231 3794
rect 177 3710 182 3738
rect 210 3710 8974 3738
rect 9002 3710 9007 3738
rect 9417 3710 9422 3738
rect 9450 3710 12558 3738
rect 12586 3710 12591 3738
rect 14345 3710 14350 3738
rect 14378 3710 15358 3738
rect 15386 3710 15391 3738
rect 17089 3710 17094 3738
rect 17122 3710 21014 3738
rect 21042 3710 21047 3738
rect 21126 3710 28798 3738
rect 28826 3710 28831 3738
rect 21126 3682 21154 3710
rect 6729 3654 6734 3682
rect 6762 3654 7014 3682
rect 7042 3654 7047 3682
rect 7121 3654 7126 3682
rect 7154 3654 17654 3682
rect 17682 3654 17687 3682
rect 17822 3654 18382 3682
rect 18410 3654 18415 3682
rect 18489 3654 18494 3682
rect 18522 3654 21154 3682
rect 21233 3654 21238 3682
rect 21266 3654 30254 3682
rect 30282 3654 30287 3682
rect 0 3626 56 3640
rect 17822 3626 17850 3654
rect 32144 3626 32200 3640
rect 0 3598 5054 3626
rect 5082 3598 5087 3626
rect 6897 3598 6902 3626
rect 6930 3598 7238 3626
rect 7266 3598 7271 3626
rect 7625 3598 7630 3626
rect 7658 3598 7798 3626
rect 7826 3598 7831 3626
rect 7961 3598 7966 3626
rect 7994 3598 9366 3626
rect 9394 3598 9399 3626
rect 11998 3598 14294 3626
rect 14322 3598 14327 3626
rect 16585 3598 16590 3626
rect 16618 3598 17850 3626
rect 17929 3598 17934 3626
rect 17962 3598 28630 3626
rect 28658 3598 28910 3626
rect 28938 3598 28943 3626
rect 31425 3598 31430 3626
rect 31458 3598 32200 3626
rect 0 3584 56 3598
rect 6729 3542 6734 3570
rect 6762 3542 8022 3570
rect 8050 3542 8055 3570
rect 2227 3514 2232 3542
rect 2260 3514 2284 3542
rect 2312 3514 2336 3542
rect 2364 3514 2369 3542
rect 11998 3514 12026 3598
rect 32144 3584 32200 3598
rect 13393 3542 13398 3570
rect 13426 3542 18438 3570
rect 18466 3542 18471 3570
rect 18545 3542 18550 3570
rect 18578 3542 20006 3570
rect 20034 3542 20039 3570
rect 24257 3542 24262 3570
rect 24290 3542 29134 3570
rect 29162 3542 29414 3570
rect 29442 3542 29447 3570
rect 12227 3514 12232 3542
rect 12260 3514 12284 3542
rect 12312 3514 12336 3542
rect 12364 3514 12369 3542
rect 22227 3514 22232 3542
rect 22260 3514 22284 3542
rect 22312 3514 22336 3542
rect 22364 3514 22369 3542
rect 4606 3486 10374 3514
rect 10402 3486 10407 3514
rect 11438 3486 12026 3514
rect 15073 3486 15078 3514
rect 15106 3486 21854 3514
rect 28737 3486 28742 3514
rect 28770 3486 29078 3514
rect 29106 3486 29111 3514
rect 0 3402 56 3416
rect 4606 3402 4634 3486
rect 11438 3458 11466 3486
rect 21826 3458 21854 3486
rect 7345 3430 7350 3458
rect 7378 3430 8582 3458
rect 8610 3430 8615 3458
rect 9809 3430 9814 3458
rect 9842 3430 11466 3458
rect 11494 3430 14014 3458
rect 14042 3430 14047 3458
rect 14905 3430 14910 3458
rect 14938 3430 16590 3458
rect 16618 3430 16623 3458
rect 16697 3430 16702 3458
rect 16730 3430 19894 3458
rect 19922 3430 19927 3458
rect 20001 3430 20006 3458
rect 20034 3430 21294 3458
rect 21322 3430 21327 3458
rect 21826 3430 27734 3458
rect 29297 3430 29302 3458
rect 29330 3430 30926 3458
rect 30954 3430 30959 3458
rect 0 3374 4634 3402
rect 7793 3374 7798 3402
rect 7826 3374 10094 3402
rect 0 3360 56 3374
rect 10066 3346 10094 3374
rect 11494 3346 11522 3430
rect 27706 3402 27734 3430
rect 32144 3402 32200 3416
rect 11601 3374 11606 3402
rect 11634 3374 12166 3402
rect 12194 3374 12199 3402
rect 13505 3374 13510 3402
rect 13538 3374 16758 3402
rect 16786 3374 16791 3402
rect 16977 3374 16982 3402
rect 17010 3374 17178 3402
rect 17257 3374 17262 3402
rect 17290 3374 18550 3402
rect 18578 3374 18583 3402
rect 18993 3374 18998 3402
rect 19026 3374 21854 3402
rect 27706 3374 30254 3402
rect 30282 3374 30287 3402
rect 30753 3374 30758 3402
rect 30786 3374 32200 3402
rect 17150 3346 17178 3374
rect 21826 3346 21854 3374
rect 32144 3360 32200 3374
rect 1353 3318 1358 3346
rect 1386 3318 1694 3346
rect 7905 3318 7910 3346
rect 7938 3318 8750 3346
rect 8778 3318 8783 3346
rect 10066 3318 11522 3346
rect 11825 3318 11830 3346
rect 11858 3318 16758 3346
rect 16786 3318 16791 3346
rect 17150 3318 20958 3346
rect 20986 3318 20991 3346
rect 21826 3318 23758 3346
rect 23786 3318 23791 3346
rect 25489 3318 25494 3346
rect 25522 3318 26446 3346
rect 26474 3318 26479 3346
rect 29969 3318 29974 3346
rect 30002 3318 30982 3346
rect 31010 3318 31015 3346
rect 1666 3290 1694 3318
rect 1666 3262 9254 3290
rect 9282 3262 9287 3290
rect 11657 3262 11662 3290
rect 11690 3262 13286 3290
rect 13314 3262 13319 3290
rect 15353 3262 15358 3290
rect 15386 3262 15526 3290
rect 15554 3262 18774 3290
rect 18802 3262 18807 3290
rect 20785 3262 20790 3290
rect 20818 3262 23366 3290
rect 23394 3262 23399 3290
rect 28961 3262 28966 3290
rect 28994 3262 30310 3290
rect 30338 3262 30343 3290
rect 1666 3206 8526 3234
rect 8554 3206 8559 3234
rect 10066 3206 18998 3234
rect 19026 3206 19031 3234
rect 19273 3206 19278 3234
rect 19306 3206 28910 3234
rect 28938 3206 29694 3234
rect 29722 3206 29727 3234
rect 0 3178 56 3192
rect 1666 3178 1694 3206
rect 10066 3178 10094 3206
rect 32144 3178 32200 3192
rect 0 3150 1694 3178
rect 5721 3150 5726 3178
rect 5754 3150 10094 3178
rect 13062 3150 17486 3178
rect 17514 3150 17519 3178
rect 17985 3150 17990 3178
rect 18018 3150 21798 3178
rect 21826 3150 21831 3178
rect 22073 3150 22078 3178
rect 22106 3150 29022 3178
rect 29050 3150 29246 3178
rect 29274 3150 29279 3178
rect 31537 3150 31542 3178
rect 31570 3150 32200 3178
rect 0 3136 56 3150
rect 1897 3122 1902 3150
rect 1930 3122 1954 3150
rect 1982 3122 2006 3150
rect 2034 3122 2039 3150
rect 11897 3122 11902 3150
rect 11930 3122 11954 3150
rect 11982 3122 12006 3150
rect 12034 3122 12039 3150
rect 5889 3094 5894 3122
rect 5922 3094 6622 3122
rect 6650 3094 6655 3122
rect 6785 3094 6790 3122
rect 6818 3094 11830 3122
rect 11858 3094 11863 3122
rect 6337 3038 6342 3066
rect 6370 3038 12166 3066
rect 12194 3038 12199 3066
rect 13062 3010 13090 3150
rect 21897 3122 21902 3150
rect 21930 3122 21954 3150
rect 21982 3122 22006 3150
rect 22034 3122 22039 3150
rect 32144 3136 32200 3150
rect 15689 3094 15694 3122
rect 15722 3094 19054 3122
rect 19082 3094 19087 3122
rect 19161 3094 19166 3122
rect 19194 3094 21854 3122
rect 22129 3094 22134 3122
rect 22162 3094 30142 3122
rect 30170 3094 30175 3122
rect 21826 3066 21854 3094
rect 18041 3038 18046 3066
rect 18074 3038 21462 3066
rect 21490 3038 21495 3066
rect 21826 3038 22638 3066
rect 22666 3038 22671 3066
rect 30753 3038 30758 3066
rect 30786 3038 32102 3066
rect 32130 3038 32135 3066
rect 4433 2982 4438 3010
rect 4466 2982 6566 3010
rect 6594 2982 6599 3010
rect 9025 2982 9030 3010
rect 9058 2982 9198 3010
rect 9226 2982 13090 3010
rect 13673 2982 13678 3010
rect 13706 2982 16366 3010
rect 16394 2982 16399 3010
rect 18321 2982 18326 3010
rect 18354 2982 21126 3010
rect 21154 2982 21159 3010
rect 21289 2982 21294 3010
rect 21322 2982 22638 3010
rect 22666 2982 22671 3010
rect 23137 2982 23142 3010
rect 23170 2982 29134 3010
rect 29162 2982 29167 3010
rect 29633 2982 29638 3010
rect 29666 2982 30870 3010
rect 30898 2982 30903 3010
rect 0 2954 56 2968
rect 32144 2954 32200 2968
rect 0 2926 6062 2954
rect 6090 2926 6095 2954
rect 7177 2926 7182 2954
rect 7210 2926 9926 2954
rect 9954 2926 9959 2954
rect 10089 2926 10094 2954
rect 10122 2926 12110 2954
rect 12138 2926 12143 2954
rect 12497 2926 12502 2954
rect 12530 2926 13174 2954
rect 13202 2926 13207 2954
rect 13393 2926 13398 2954
rect 13426 2926 16086 2954
rect 16114 2926 16119 2954
rect 18382 2926 20006 2954
rect 20034 2926 20039 2954
rect 21233 2926 21238 2954
rect 21266 2926 29302 2954
rect 29330 2926 29335 2954
rect 30641 2926 30646 2954
rect 30674 2926 32200 2954
rect 0 2912 56 2926
rect 18382 2898 18410 2926
rect 32144 2912 32200 2926
rect 961 2870 966 2898
rect 994 2870 7070 2898
rect 7098 2870 7103 2898
rect 10066 2870 13510 2898
rect 13538 2870 13543 2898
rect 13617 2870 13622 2898
rect 13650 2870 14462 2898
rect 14490 2870 14495 2898
rect 15073 2870 15078 2898
rect 15106 2870 15190 2898
rect 15218 2870 18410 2898
rect 18489 2870 18494 2898
rect 18522 2870 21014 2898
rect 21042 2870 21047 2898
rect 21121 2870 21126 2898
rect 21154 2870 21854 2898
rect 21882 2870 21887 2898
rect 22129 2870 22134 2898
rect 22162 2870 25046 2898
rect 25074 2870 25079 2898
rect 10066 2842 10094 2870
rect 6001 2814 6006 2842
rect 6034 2814 10094 2842
rect 12166 2814 18158 2842
rect 18186 2814 18191 2842
rect 19217 2814 19222 2842
rect 19250 2814 21350 2842
rect 21378 2814 21383 2842
rect 21457 2814 21462 2842
rect 21490 2814 23478 2842
rect 23506 2814 23511 2842
rect 28289 2814 28294 2842
rect 28322 2814 28518 2842
rect 28546 2814 28686 2842
rect 28714 2814 28719 2842
rect 12166 2786 12194 2814
rect 9137 2758 9142 2786
rect 9170 2758 12194 2786
rect 13001 2758 13006 2786
rect 13034 2758 15274 2786
rect 15409 2758 15414 2786
rect 15442 2758 17262 2786
rect 17290 2758 17295 2786
rect 19273 2758 19278 2786
rect 19306 2758 22134 2786
rect 22162 2758 22167 2786
rect 0 2730 56 2744
rect 2227 2730 2232 2758
rect 2260 2730 2284 2758
rect 2312 2730 2336 2758
rect 2364 2730 2369 2758
rect 12227 2730 12232 2758
rect 12260 2730 12284 2758
rect 12312 2730 12336 2758
rect 12364 2730 12369 2758
rect 15246 2730 15274 2758
rect 22227 2730 22232 2758
rect 22260 2730 22284 2758
rect 22312 2730 22336 2758
rect 22364 2730 22369 2758
rect 32144 2730 32200 2744
rect 0 2702 1694 2730
rect 4937 2702 4942 2730
rect 4970 2702 7798 2730
rect 7826 2702 7831 2730
rect 9977 2702 9982 2730
rect 10010 2702 12194 2730
rect 0 2688 56 2702
rect 1666 2674 1694 2702
rect 12166 2674 12194 2702
rect 12446 2702 15134 2730
rect 15162 2702 15167 2730
rect 15246 2702 19334 2730
rect 19362 2702 19367 2730
rect 19889 2702 19894 2730
rect 19922 2702 20174 2730
rect 20202 2702 20207 2730
rect 21177 2702 21182 2730
rect 21210 2702 21294 2730
rect 21322 2702 21327 2730
rect 23361 2702 23366 2730
rect 23394 2702 29190 2730
rect 29218 2702 29223 2730
rect 31313 2702 31318 2730
rect 31346 2702 32200 2730
rect 12446 2674 12474 2702
rect 32144 2688 32200 2702
rect 1666 2646 4158 2674
rect 4186 2646 4191 2674
rect 7569 2646 7574 2674
rect 7602 2646 10850 2674
rect 10929 2646 10934 2674
rect 10962 2646 11102 2674
rect 11130 2646 11135 2674
rect 12166 2646 12474 2674
rect 12553 2646 12558 2674
rect 12586 2646 12726 2674
rect 12754 2646 13454 2674
rect 13482 2646 13487 2674
rect 13566 2646 15078 2674
rect 15106 2646 15111 2674
rect 17201 2646 17206 2674
rect 17234 2646 18326 2674
rect 18354 2646 18359 2674
rect 18601 2646 18606 2674
rect 18634 2646 20678 2674
rect 20706 2646 20711 2674
rect 20953 2646 20958 2674
rect 20986 2646 22862 2674
rect 22890 2646 22895 2674
rect 29190 2646 31150 2674
rect 31178 2646 31183 2674
rect 10822 2618 10850 2646
rect 13566 2618 13594 2646
rect 29190 2618 29218 2646
rect 905 2590 910 2618
rect 938 2590 3150 2618
rect 3178 2590 3183 2618
rect 3257 2590 3262 2618
rect 3290 2590 9366 2618
rect 9394 2590 9399 2618
rect 9585 2590 9590 2618
rect 9618 2590 10654 2618
rect 10682 2590 10687 2618
rect 10822 2590 13594 2618
rect 13622 2590 14350 2618
rect 14378 2590 14383 2618
rect 14513 2590 14518 2618
rect 14546 2590 15918 2618
rect 15946 2590 15951 2618
rect 16641 2590 16646 2618
rect 16674 2590 17374 2618
rect 17402 2590 17407 2618
rect 18153 2590 18158 2618
rect 18186 2590 19390 2618
rect 19418 2590 19423 2618
rect 19553 2590 19558 2618
rect 19586 2590 20902 2618
rect 20930 2590 20935 2618
rect 21009 2590 21014 2618
rect 21042 2590 22974 2618
rect 23002 2590 23007 2618
rect 25433 2590 25438 2618
rect 25466 2590 27118 2618
rect 27146 2590 27151 2618
rect 29185 2590 29190 2618
rect 29218 2590 29223 2618
rect 29302 2590 30142 2618
rect 30170 2590 30175 2618
rect 30529 2590 30534 2618
rect 30562 2590 31262 2618
rect 31290 2590 31295 2618
rect 13622 2562 13650 2590
rect 29302 2562 29330 2590
rect 1241 2534 1246 2562
rect 1274 2534 1414 2562
rect 1442 2534 5894 2562
rect 5922 2534 5927 2562
rect 6505 2534 6510 2562
rect 6538 2534 8554 2562
rect 9249 2534 9254 2562
rect 9282 2534 10094 2562
rect 10873 2534 10878 2562
rect 10906 2534 11802 2562
rect 12441 2534 12446 2562
rect 12474 2534 13650 2562
rect 14233 2534 14238 2562
rect 14266 2534 15078 2562
rect 15106 2534 15111 2562
rect 15185 2534 15190 2562
rect 15218 2534 18438 2562
rect 18466 2534 18471 2562
rect 20174 2534 21742 2562
rect 21770 2534 21775 2562
rect 22409 2534 22414 2562
rect 22442 2534 24402 2562
rect 26329 2534 26334 2562
rect 26362 2534 28182 2562
rect 28210 2534 28350 2562
rect 28378 2534 28383 2562
rect 28625 2534 28630 2562
rect 28658 2534 29330 2562
rect 29969 2534 29974 2562
rect 30002 2534 30926 2562
rect 30954 2534 30959 2562
rect 0 2506 56 2520
rect 8526 2506 8554 2534
rect 10066 2506 10094 2534
rect 11774 2506 11802 2534
rect 20174 2506 20202 2534
rect 24374 2506 24402 2534
rect 32144 2506 32200 2520
rect 0 2478 4634 2506
rect 4993 2478 4998 2506
rect 5026 2478 8414 2506
rect 8442 2478 8447 2506
rect 8526 2478 9982 2506
rect 10010 2478 10015 2506
rect 10066 2478 11662 2506
rect 11690 2478 11695 2506
rect 11774 2478 15414 2506
rect 15442 2478 15447 2506
rect 16753 2478 16758 2506
rect 16786 2478 20202 2506
rect 20393 2478 20398 2506
rect 20426 2478 23254 2506
rect 23282 2478 23287 2506
rect 24374 2478 27566 2506
rect 27594 2478 27599 2506
rect 29129 2478 29134 2506
rect 29162 2478 31094 2506
rect 31122 2478 31127 2506
rect 31537 2478 31542 2506
rect 31570 2478 32200 2506
rect 0 2464 56 2478
rect 4606 2394 4634 2478
rect 32144 2464 32200 2478
rect 7065 2422 7070 2450
rect 7098 2422 13062 2450
rect 13090 2422 13095 2450
rect 13169 2422 13174 2450
rect 13202 2422 18662 2450
rect 18690 2422 18695 2450
rect 19217 2422 19222 2450
rect 19250 2422 22750 2450
rect 22778 2422 22783 2450
rect 24313 2422 24318 2450
rect 24346 2422 28742 2450
rect 28770 2422 28775 2450
rect 4606 2366 10094 2394
rect 10122 2366 10127 2394
rect 13281 2366 13286 2394
rect 13314 2366 13902 2394
rect 13930 2366 13935 2394
rect 15465 2366 15470 2394
rect 15498 2366 21238 2394
rect 21266 2366 21271 2394
rect 22689 2366 22694 2394
rect 22722 2366 23982 2394
rect 24010 2366 24015 2394
rect 25433 2366 25438 2394
rect 25466 2366 29078 2394
rect 29106 2366 29111 2394
rect 1897 2338 1902 2366
rect 1930 2338 1954 2366
rect 1982 2338 2006 2366
rect 2034 2338 2039 2366
rect 11897 2338 11902 2366
rect 11930 2338 11954 2366
rect 11982 2338 12006 2366
rect 12034 2338 12039 2366
rect 21897 2338 21902 2366
rect 21930 2338 21954 2366
rect 21982 2338 22006 2366
rect 22034 2338 22039 2366
rect 4153 2310 4158 2338
rect 4186 2310 10430 2338
rect 10458 2310 10463 2338
rect 10817 2310 10822 2338
rect 10850 2310 11830 2338
rect 11858 2310 11863 2338
rect 12105 2310 12110 2338
rect 12138 2310 14406 2338
rect 14434 2310 14439 2338
rect 17033 2310 17038 2338
rect 17066 2310 18382 2338
rect 18410 2310 18415 2338
rect 22353 2310 22358 2338
rect 22386 2310 25998 2338
rect 26026 2310 26031 2338
rect 0 2282 56 2296
rect 32144 2282 32200 2296
rect 0 2254 7630 2282
rect 7658 2254 7663 2282
rect 8465 2254 8470 2282
rect 8498 2254 13230 2282
rect 13258 2254 13263 2282
rect 13561 2254 13566 2282
rect 13594 2254 15022 2282
rect 15050 2254 15055 2282
rect 15129 2254 15134 2282
rect 15162 2254 16142 2282
rect 16170 2254 16175 2282
rect 17369 2254 17374 2282
rect 17402 2254 20174 2282
rect 20202 2254 20207 2282
rect 20505 2254 20510 2282
rect 20538 2254 24766 2282
rect 24794 2254 24799 2282
rect 31257 2254 31262 2282
rect 31290 2254 32200 2282
rect 0 2240 56 2254
rect 32144 2240 32200 2254
rect 5945 2198 5950 2226
rect 5978 2198 11774 2226
rect 11802 2198 11807 2226
rect 11881 2198 11886 2226
rect 11914 2198 12950 2226
rect 12978 2198 12983 2226
rect 13057 2198 13062 2226
rect 13090 2198 17598 2226
rect 17626 2198 17631 2226
rect 21401 2198 21406 2226
rect 21434 2198 23310 2226
rect 23338 2198 23343 2226
rect 23697 2198 23702 2226
rect 23730 2198 24934 2226
rect 24962 2198 24967 2226
rect 27841 2198 27846 2226
rect 27874 2198 30366 2226
rect 30394 2198 30399 2226
rect 7681 2142 7686 2170
rect 7714 2142 11550 2170
rect 11578 2142 11583 2170
rect 11657 2142 11662 2170
rect 11690 2142 15582 2170
rect 15610 2142 15615 2170
rect 15946 2142 22638 2170
rect 22666 2142 22671 2170
rect 15946 2114 15974 2142
rect 1078 2086 2478 2114
rect 2506 2086 2511 2114
rect 7121 2086 7126 2114
rect 7154 2086 11942 2114
rect 11970 2086 11975 2114
rect 12161 2086 12166 2114
rect 12194 2086 13398 2114
rect 13426 2086 13431 2114
rect 13953 2086 13958 2114
rect 13986 2086 15974 2114
rect 18382 2086 20846 2114
rect 20874 2086 20879 2114
rect 21009 2086 21014 2114
rect 21042 2086 22358 2114
rect 22386 2086 22391 2114
rect 22465 2086 22470 2114
rect 22498 2086 27902 2114
rect 27930 2086 27935 2114
rect 0 2058 56 2072
rect 1078 2058 1106 2086
rect 18382 2058 18410 2086
rect 32144 2058 32200 2072
rect 0 2030 1106 2058
rect 1185 2030 1190 2058
rect 1218 2030 1302 2058
rect 1330 2030 7462 2058
rect 7490 2030 7495 2058
rect 8521 2030 8526 2058
rect 8554 2030 8638 2058
rect 8666 2030 13454 2058
rect 13482 2030 13487 2058
rect 14065 2030 14070 2058
rect 14098 2030 18410 2058
rect 20169 2030 20174 2058
rect 20202 2030 23394 2058
rect 28065 2030 28070 2058
rect 28098 2030 28238 2058
rect 28266 2030 30534 2058
rect 30562 2030 30567 2058
rect 31425 2030 31430 2058
rect 31458 2030 32200 2058
rect 0 2016 56 2030
rect 2865 1974 2870 2002
rect 2898 1974 8414 2002
rect 8442 1974 8447 2002
rect 8526 1974 12110 2002
rect 12138 1974 12143 2002
rect 12558 1974 19278 2002
rect 19306 1974 19311 2002
rect 19889 1974 19894 2002
rect 19922 1974 21070 2002
rect 21098 1974 21103 2002
rect 2227 1946 2232 1974
rect 2260 1946 2284 1974
rect 2312 1946 2336 1974
rect 2364 1946 2369 1974
rect 8526 1946 8554 1974
rect 12227 1946 12232 1974
rect 12260 1946 12284 1974
rect 12312 1946 12336 1974
rect 12364 1946 12369 1974
rect 7849 1918 7854 1946
rect 7882 1918 8554 1946
rect 10033 1918 10038 1946
rect 10066 1918 12166 1946
rect 12194 1918 12199 1946
rect 12558 1890 12586 1974
rect 22227 1946 22232 1974
rect 22260 1946 22284 1974
rect 22312 1946 22336 1974
rect 22364 1946 22369 1974
rect 23366 1946 23394 2030
rect 32144 2016 32200 2030
rect 23473 1974 23478 2002
rect 23506 1974 30926 2002
rect 30954 1974 30959 2002
rect 12777 1918 12782 1946
rect 12810 1918 14182 1946
rect 14210 1918 14215 1946
rect 14289 1918 14294 1946
rect 14322 1918 18214 1946
rect 18242 1918 18247 1946
rect 18433 1918 18438 1946
rect 18466 1918 21014 1946
rect 21042 1918 21047 1946
rect 23366 1918 29918 1946
rect 29946 1918 29951 1946
rect 5665 1862 5670 1890
rect 5698 1862 7574 1890
rect 8633 1862 8638 1890
rect 8666 1862 8806 1890
rect 8834 1862 9870 1890
rect 9898 1862 9903 1890
rect 10061 1862 10066 1890
rect 10094 1862 12586 1890
rect 13113 1862 13118 1890
rect 13146 1862 14630 1890
rect 14658 1862 14663 1890
rect 17257 1862 17262 1890
rect 17290 1862 19166 1890
rect 19194 1862 19199 1890
rect 20225 1862 20230 1890
rect 20258 1862 29526 1890
rect 29554 1862 29694 1890
rect 29722 1862 29727 1890
rect 0 1834 56 1848
rect 7546 1834 7574 1862
rect 32144 1834 32200 1848
rect 0 1806 7182 1834
rect 7210 1806 7215 1834
rect 7546 1806 8358 1834
rect 8386 1806 8391 1834
rect 11937 1806 11942 1834
rect 11970 1806 14350 1834
rect 14378 1806 14383 1834
rect 14462 1806 20622 1834
rect 20650 1806 20655 1834
rect 20785 1806 20790 1834
rect 20818 1806 22022 1834
rect 22050 1806 22190 1834
rect 22218 1806 22223 1834
rect 30641 1806 30646 1834
rect 30674 1806 32200 1834
rect 0 1792 56 1806
rect 14462 1778 14490 1806
rect 32144 1792 32200 1806
rect 1297 1750 1302 1778
rect 1330 1750 1470 1778
rect 1498 1750 6678 1778
rect 6706 1750 6711 1778
rect 8969 1750 8974 1778
rect 9002 1750 12894 1778
rect 12922 1750 12927 1778
rect 13113 1750 13118 1778
rect 13146 1750 13874 1778
rect 13953 1750 13958 1778
rect 13986 1750 14490 1778
rect 14569 1750 14574 1778
rect 14602 1750 17094 1778
rect 17122 1750 17127 1778
rect 18489 1750 18494 1778
rect 18522 1750 21070 1778
rect 21098 1750 21103 1778
rect 23473 1750 23478 1778
rect 23506 1750 26110 1778
rect 26138 1750 26143 1778
rect 13846 1722 13874 1750
rect 1521 1694 1526 1722
rect 1554 1694 5026 1722
rect 8745 1694 8750 1722
rect 8778 1694 10878 1722
rect 10906 1694 10911 1722
rect 11545 1694 11550 1722
rect 11578 1694 13734 1722
rect 13762 1694 13767 1722
rect 13846 1694 15330 1722
rect 18881 1694 18886 1722
rect 18914 1694 21042 1722
rect 4998 1666 5026 1694
rect 15302 1666 15330 1694
rect 21014 1666 21042 1694
rect 21826 1694 23534 1722
rect 21826 1666 21854 1694
rect 1806 1638 4214 1666
rect 4998 1638 7574 1666
rect 7602 1638 7607 1666
rect 10481 1638 10486 1666
rect 10514 1638 11158 1666
rect 11186 1638 11191 1666
rect 11713 1638 11718 1666
rect 11746 1638 12138 1666
rect 12889 1638 12894 1666
rect 12922 1638 15190 1666
rect 15218 1638 15223 1666
rect 15302 1638 17486 1666
rect 17514 1638 17519 1666
rect 17593 1638 17598 1666
rect 17626 1638 20230 1666
rect 20258 1638 20263 1666
rect 21014 1638 21854 1666
rect 23506 1666 23534 1694
rect 27174 1694 28182 1722
rect 28210 1694 28215 1722
rect 30641 1694 30646 1722
rect 30674 1694 31318 1722
rect 31346 1694 31351 1722
rect 23506 1638 25606 1666
rect 25634 1638 25639 1666
rect 0 1610 56 1624
rect 1806 1610 1834 1638
rect 0 1582 1834 1610
rect 4186 1610 4214 1638
rect 12110 1610 12138 1638
rect 4186 1582 11830 1610
rect 11858 1582 11863 1610
rect 12110 1582 13958 1610
rect 13986 1582 13991 1610
rect 17089 1582 17094 1610
rect 17122 1582 18270 1610
rect 18298 1582 18303 1610
rect 18377 1582 18382 1610
rect 18410 1582 21518 1610
rect 21546 1582 21551 1610
rect 22633 1582 22638 1610
rect 22666 1582 24262 1610
rect 24290 1582 24295 1610
rect 0 1568 56 1582
rect 1897 1554 1902 1582
rect 1930 1554 1954 1582
rect 1982 1554 2006 1582
rect 2034 1554 2039 1582
rect 11897 1554 11902 1582
rect 11930 1554 11954 1582
rect 11982 1554 12006 1582
rect 12034 1554 12039 1582
rect 21897 1554 21902 1582
rect 21930 1554 21954 1582
rect 21982 1554 22006 1582
rect 22034 1554 22039 1582
rect 27174 1554 27202 1694
rect 32144 1610 32200 1624
rect 31537 1582 31542 1610
rect 31570 1582 32200 1610
rect 32144 1568 32200 1582
rect 7625 1526 7630 1554
rect 7658 1526 10206 1554
rect 10234 1526 10239 1554
rect 13001 1526 13006 1554
rect 13034 1526 19362 1554
rect 24313 1526 24318 1554
rect 24346 1526 27202 1554
rect 27281 1526 27286 1554
rect 27314 1526 31206 1554
rect 31234 1526 31239 1554
rect 8409 1470 8414 1498
rect 8442 1470 13286 1498
rect 13314 1470 13319 1498
rect 14625 1470 14630 1498
rect 14658 1470 18494 1498
rect 18522 1470 18527 1498
rect 19334 1442 19362 1526
rect 19441 1470 19446 1498
rect 19474 1470 23478 1498
rect 23506 1470 23511 1498
rect 26049 1470 26054 1498
rect 26082 1470 28686 1498
rect 28714 1470 28719 1498
rect 7009 1414 7014 1442
rect 7042 1414 11326 1442
rect 11354 1414 11359 1442
rect 13505 1414 13510 1442
rect 13538 1414 15134 1442
rect 15162 1414 15167 1442
rect 19334 1414 26166 1442
rect 26194 1414 26199 1442
rect 0 1386 56 1400
rect 32144 1386 32200 1400
rect 0 1358 7070 1386
rect 7098 1358 7103 1386
rect 11825 1358 11830 1386
rect 11858 1358 29246 1386
rect 29274 1358 29414 1386
rect 29442 1358 29447 1386
rect 29633 1358 29638 1386
rect 29666 1358 31094 1386
rect 31122 1358 31127 1386
rect 31313 1358 31318 1386
rect 31346 1358 32200 1386
rect 0 1344 56 1358
rect 32144 1344 32200 1358
rect 1409 1302 1414 1330
rect 1442 1302 7126 1330
rect 7154 1302 7159 1330
rect 7345 1302 7350 1330
rect 7378 1302 18158 1330
rect 18186 1302 18191 1330
rect 18321 1302 18326 1330
rect 18354 1302 19446 1330
rect 19474 1302 19479 1330
rect 20393 1302 20398 1330
rect 20426 1302 25046 1330
rect 25074 1302 25079 1330
rect 25158 1302 27286 1330
rect 27314 1302 27319 1330
rect 29185 1302 29190 1330
rect 29218 1302 30086 1330
rect 30114 1302 30119 1330
rect 30641 1302 30646 1330
rect 30674 1302 31374 1330
rect 31402 1302 31407 1330
rect 25158 1274 25186 1302
rect 6505 1246 6510 1274
rect 6538 1246 12474 1274
rect 15409 1246 15414 1274
rect 15442 1246 18886 1274
rect 18914 1246 18919 1274
rect 20897 1246 20902 1274
rect 20930 1246 22694 1274
rect 22722 1246 22727 1274
rect 22969 1246 22974 1274
rect 23002 1246 25186 1274
rect 26273 1246 26278 1274
rect 26306 1246 26446 1274
rect 26474 1246 29134 1274
rect 29162 1246 29167 1274
rect 12446 1218 12474 1246
rect 12446 1190 18438 1218
rect 18466 1190 18471 1218
rect 23417 1190 23422 1218
rect 23450 1190 28798 1218
rect 28826 1190 28831 1218
rect 0 1162 56 1176
rect 2227 1162 2232 1190
rect 2260 1162 2284 1190
rect 2312 1162 2336 1190
rect 2364 1162 2369 1190
rect 12227 1162 12232 1190
rect 12260 1162 12284 1190
rect 12312 1162 12336 1190
rect 12364 1162 12369 1190
rect 22227 1162 22232 1190
rect 22260 1162 22284 1190
rect 22312 1162 22336 1190
rect 22364 1162 22369 1190
rect 32144 1162 32200 1176
rect 0 1134 2114 1162
rect 0 1120 56 1134
rect 2086 1106 2114 1134
rect 2422 1134 8414 1162
rect 8442 1134 8447 1162
rect 8577 1134 8582 1162
rect 8610 1134 12166 1162
rect 12194 1134 12199 1162
rect 13785 1134 13790 1162
rect 13818 1134 17654 1162
rect 17682 1134 17687 1162
rect 17873 1134 17878 1162
rect 17906 1134 20790 1162
rect 20818 1134 20823 1162
rect 22806 1134 23870 1162
rect 23898 1134 23903 1162
rect 31425 1134 31430 1162
rect 31458 1134 32200 1162
rect 2422 1106 2450 1134
rect 22806 1106 22834 1134
rect 32144 1120 32200 1134
rect 2086 1078 2450 1106
rect 3929 1078 3934 1106
rect 3962 1078 7350 1106
rect 7378 1078 7383 1106
rect 8073 1078 8078 1106
rect 8106 1078 8358 1106
rect 8386 1078 14126 1106
rect 14154 1078 14159 1106
rect 15633 1078 15638 1106
rect 15666 1078 18158 1106
rect 18186 1078 18191 1106
rect 18265 1078 18270 1106
rect 18298 1078 21238 1106
rect 21266 1078 21271 1106
rect 21345 1078 21350 1106
rect 21378 1078 21462 1106
rect 21490 1078 22834 1106
rect 22913 1078 22918 1106
rect 22946 1078 23086 1106
rect 23114 1078 24486 1106
rect 24514 1078 24519 1106
rect 29241 1078 29246 1106
rect 29274 1078 30310 1106
rect 30338 1078 30343 1106
rect 457 1022 462 1050
rect 490 1022 6118 1050
rect 6146 1022 6230 1050
rect 6258 1022 6263 1050
rect 12161 1022 12166 1050
rect 12194 1022 16198 1050
rect 16226 1022 16231 1050
rect 17481 1022 17486 1050
rect 17514 1022 23366 1050
rect 23394 1022 23399 1050
rect 24873 1022 24878 1050
rect 24906 1022 28014 1050
rect 28042 1022 28047 1050
rect 28793 1022 28798 1050
rect 28826 1022 30142 1050
rect 30170 1022 30175 1050
rect 910 966 4382 994
rect 4410 966 4550 994
rect 4578 966 4583 994
rect 5273 966 5278 994
rect 5306 966 13006 994
rect 13034 966 13039 994
rect 14177 966 14182 994
rect 14210 966 14434 994
rect 14961 966 14966 994
rect 14994 966 19446 994
rect 19474 966 19479 994
rect 21793 966 21798 994
rect 21826 966 21966 994
rect 21994 966 24150 994
rect 24178 966 24183 994
rect 29969 966 29974 994
rect 30002 966 30926 994
rect 30954 966 30959 994
rect 0 938 56 952
rect 910 938 938 966
rect 14406 938 14434 966
rect 32144 938 32200 952
rect 0 910 938 938
rect 1017 910 1022 938
rect 1050 910 7910 938
rect 7938 910 7943 938
rect 11825 910 11830 938
rect 11858 910 14294 938
rect 14322 910 14327 938
rect 14406 910 18774 938
rect 18802 910 18807 938
rect 18886 910 19838 938
rect 19866 910 19871 938
rect 23473 910 23478 938
rect 23506 910 24430 938
rect 24458 910 24598 938
rect 24626 910 24631 938
rect 31537 910 31542 938
rect 31570 910 32200 938
rect 0 896 56 910
rect 18886 882 18914 910
rect 32144 896 32200 910
rect 11321 854 11326 882
rect 11354 854 14406 882
rect 14434 854 14439 882
rect 17817 854 17822 882
rect 17850 854 18914 882
rect 19334 854 20734 882
rect 20762 854 20767 882
rect 21826 854 22106 882
rect 19334 826 19362 854
rect 21826 826 21854 854
rect 5833 798 5838 826
rect 5866 798 6902 826
rect 6930 798 6935 826
rect 7569 798 7574 826
rect 7602 798 10990 826
rect 11018 798 11023 826
rect 13449 798 13454 826
rect 13482 798 18270 826
rect 18298 798 18303 826
rect 18937 798 18942 826
rect 18970 798 19362 826
rect 19833 798 19838 826
rect 19866 798 21854 826
rect 22078 826 22106 854
rect 25214 854 27734 882
rect 30641 854 30646 882
rect 30674 854 31290 882
rect 22078 798 24878 826
rect 24906 798 24911 826
rect 1897 770 1902 798
rect 1930 770 1954 798
rect 1982 770 2006 798
rect 2034 770 2039 798
rect 11897 770 11902 798
rect 11930 770 11954 798
rect 11982 770 12006 798
rect 12034 770 12039 798
rect 21897 770 21902 798
rect 21930 770 21954 798
rect 21982 770 22006 798
rect 22034 770 22039 798
rect 25214 770 25242 854
rect 27706 826 27734 854
rect 27706 798 29582 826
rect 29610 798 29615 826
rect 4377 742 4382 770
rect 4410 742 6286 770
rect 6314 742 6319 770
rect 7177 742 7182 770
rect 7210 742 10094 770
rect 10122 742 10127 770
rect 10201 742 10206 770
rect 10234 742 11830 770
rect 11858 742 11863 770
rect 14401 742 14406 770
rect 14434 742 17262 770
rect 17290 742 17295 770
rect 17929 742 17934 770
rect 17962 742 18102 770
rect 18130 742 19670 770
rect 19698 742 19703 770
rect 23702 742 25242 770
rect 26105 742 26110 770
rect 26138 742 28854 770
rect 28882 742 28887 770
rect 0 714 56 728
rect 0 686 7854 714
rect 7882 686 7887 714
rect 8409 686 8414 714
rect 8442 686 19418 714
rect 20169 686 20174 714
rect 20202 686 22694 714
rect 22722 686 22727 714
rect 0 672 56 686
rect 19390 658 19418 686
rect 23702 658 23730 742
rect 31262 714 31290 854
rect 32144 714 32200 728
rect 4186 630 5138 658
rect 5273 630 5278 658
rect 5306 630 8470 658
rect 8498 630 8503 658
rect 11657 630 11662 658
rect 11690 630 14686 658
rect 14714 630 14719 658
rect 14798 630 19278 658
rect 19306 630 19311 658
rect 19390 630 23730 658
rect 24766 686 28294 714
rect 28322 686 28327 714
rect 31262 686 32200 714
rect 4186 602 4214 630
rect 462 574 4214 602
rect 0 490 56 504
rect 462 490 490 574
rect 5110 546 5138 630
rect 14798 602 14826 630
rect 24766 602 24794 686
rect 32144 672 32200 686
rect 26161 630 26166 658
rect 26194 630 29302 658
rect 29330 630 29335 658
rect 10089 574 10094 602
rect 10122 574 13566 602
rect 13594 574 13599 602
rect 14345 574 14350 602
rect 14378 574 14826 602
rect 14905 574 14910 602
rect 14938 574 18438 602
rect 18466 574 18471 602
rect 18657 574 18662 602
rect 18690 574 20174 602
rect 20202 574 20207 602
rect 20286 574 24794 602
rect 24873 574 24878 602
rect 24906 574 30254 602
rect 30282 574 30287 602
rect 20286 546 20314 574
rect 905 518 910 546
rect 938 518 4662 546
rect 4690 518 4695 546
rect 4769 518 4774 546
rect 4802 518 4998 546
rect 5026 518 5031 546
rect 5110 518 7518 546
rect 7546 518 7551 546
rect 8017 518 8022 546
rect 8050 518 13510 546
rect 13538 518 13543 546
rect 19329 518 19334 546
rect 19362 518 20314 546
rect 20393 518 20398 546
rect 20426 518 23422 546
rect 23450 518 23455 546
rect 25545 518 25550 546
rect 25578 518 27678 546
rect 27706 518 27711 546
rect 32144 490 32200 504
rect 0 462 490 490
rect 1185 462 1190 490
rect 1218 462 1302 490
rect 1330 462 15358 490
rect 15386 462 15391 490
rect 18713 462 18718 490
rect 18746 462 20258 490
rect 0 448 56 462
rect 20230 434 20258 462
rect 21826 462 23310 490
rect 23338 462 23343 490
rect 24201 462 24206 490
rect 24234 462 26222 490
rect 26250 462 26255 490
rect 30585 462 30590 490
rect 30618 462 32200 490
rect 21826 434 21854 462
rect 32144 448 32200 462
rect 4657 406 4662 434
rect 4690 406 6846 434
rect 6874 406 6879 434
rect 20230 406 21854 434
rect 22689 406 22694 434
rect 22722 406 26334 434
rect 26362 406 26367 434
rect 2227 378 2232 406
rect 2260 378 2284 406
rect 2312 378 2336 406
rect 2364 378 2369 406
rect 12227 378 12232 406
rect 12260 378 12284 406
rect 12312 378 12336 406
rect 12364 378 12369 406
rect 22227 378 22232 406
rect 22260 378 22284 406
rect 22312 378 22336 406
rect 22364 378 22369 406
rect 12446 350 13622 378
rect 13650 350 13655 378
rect 18209 350 18214 378
rect 18242 350 21574 378
rect 21602 350 21607 378
rect 22857 350 22862 378
rect 22890 350 28350 378
rect 28378 350 28383 378
rect 12446 322 12474 350
rect 6673 294 6678 322
rect 6706 294 12474 322
rect 13113 294 13118 322
rect 13146 294 17878 322
rect 17906 294 17911 322
rect 20169 294 20174 322
rect 20202 294 29526 322
rect 29554 294 29559 322
rect 0 266 56 280
rect 32144 266 32200 280
rect 0 238 4830 266
rect 4858 238 5054 266
rect 5082 238 5087 266
rect 10537 238 10542 266
rect 10570 238 14910 266
rect 14938 238 14943 266
rect 17481 238 17486 266
rect 17514 238 24990 266
rect 25018 238 25023 266
rect 29801 238 29806 266
rect 29834 238 32200 266
rect 0 224 56 238
rect 32144 224 32200 238
rect 4881 182 4886 210
rect 4914 182 31094 210
rect 31122 182 31127 210
rect 2921 126 2926 154
rect 2954 126 4214 154
rect 7289 126 7294 154
rect 7322 126 13622 154
rect 13650 126 13655 154
rect 14569 126 14574 154
rect 14602 126 23758 154
rect 23786 126 23791 154
rect 4186 98 4214 126
rect 4186 70 7966 98
rect 7994 70 7999 98
rect 16025 70 16030 98
rect 16058 70 23478 98
rect 23506 70 23511 98
rect 0 42 56 56
rect 32144 42 32200 56
rect 0 14 4774 42
rect 4802 14 4807 42
rect 17033 14 17038 42
rect 17066 14 20398 42
rect 20426 14 20431 42
rect 31369 14 31374 42
rect 31402 14 32200 42
rect 0 0 56 14
rect 32144 0 32200 14
<< via3 >>
rect 2232 6650 2260 6678
rect 2284 6650 2312 6678
rect 2336 6650 2364 6678
rect 12232 6650 12260 6678
rect 12284 6650 12312 6678
rect 12336 6650 12364 6678
rect 22232 6650 22260 6678
rect 22284 6650 22312 6678
rect 22336 6650 22364 6678
rect 16702 6566 16730 6594
rect 16926 6510 16954 6538
rect 13622 6398 13650 6426
rect 15694 6286 15722 6314
rect 16702 6286 16730 6314
rect 1902 6258 1930 6286
rect 1954 6258 1982 6286
rect 2006 6258 2034 6286
rect 11902 6258 11930 6286
rect 11954 6258 11982 6286
rect 12006 6258 12034 6286
rect 21902 6258 21930 6286
rect 21954 6258 21982 6286
rect 22006 6258 22034 6286
rect 14350 6230 14378 6258
rect 14294 6062 14322 6090
rect 16254 6006 16282 6034
rect 2232 5866 2260 5894
rect 2284 5866 2312 5894
rect 2336 5866 2364 5894
rect 14294 5894 14322 5922
rect 12232 5866 12260 5894
rect 12284 5866 12312 5894
rect 12336 5866 12364 5894
rect 23366 5950 23394 5978
rect 22232 5866 22260 5894
rect 22284 5866 22312 5894
rect 22336 5866 22364 5894
rect 15694 5838 15722 5866
rect 10654 5670 10682 5698
rect 12614 5670 12642 5698
rect 1902 5474 1930 5502
rect 1954 5474 1982 5502
rect 2006 5474 2034 5502
rect 11902 5474 11930 5502
rect 11954 5474 11982 5502
rect 12006 5474 12034 5502
rect 21902 5474 21930 5502
rect 21954 5474 21982 5502
rect 22006 5474 22034 5502
rect 14182 5446 14210 5474
rect 17598 5446 17626 5474
rect 12614 5390 12642 5418
rect 16254 5390 16282 5418
rect 10654 5334 10682 5362
rect 16086 5278 16114 5306
rect 14630 5222 14658 5250
rect 14238 5166 14266 5194
rect 16086 5166 16114 5194
rect 2232 5082 2260 5110
rect 2284 5082 2312 5110
rect 2336 5082 2364 5110
rect 6734 5110 6762 5138
rect 13622 5110 13650 5138
rect 12232 5082 12260 5110
rect 12284 5082 12312 5110
rect 12336 5082 12364 5110
rect 22232 5082 22260 5110
rect 22284 5082 22312 5110
rect 22336 5082 22364 5110
rect 10990 4886 11018 4914
rect 16646 4886 16674 4914
rect 17598 4886 17626 4914
rect 13902 4830 13930 4858
rect 14294 4830 14322 4858
rect 20286 4830 20314 4858
rect 1902 4690 1930 4718
rect 1954 4690 1982 4718
rect 2006 4690 2034 4718
rect 13902 4718 13930 4746
rect 11902 4690 11930 4718
rect 11954 4690 11982 4718
rect 12006 4690 12034 4718
rect 21902 4690 21930 4718
rect 21954 4690 21982 4718
rect 22006 4690 22034 4718
rect 14238 4662 14266 4690
rect 10990 4606 11018 4634
rect 15134 4606 15162 4634
rect 14182 4438 14210 4466
rect 15414 4382 15442 4410
rect 16758 4326 16786 4354
rect 2232 4298 2260 4326
rect 2284 4298 2312 4326
rect 2336 4298 2364 4326
rect 12232 4298 12260 4326
rect 12284 4298 12312 4326
rect 12336 4298 12364 4326
rect 22232 4298 22260 4326
rect 22284 4298 22312 4326
rect 22336 4298 22364 4326
rect 12110 4270 12138 4298
rect 13622 4270 13650 4298
rect 6734 4214 6762 4242
rect 7126 4158 7154 4186
rect 12110 4158 12138 4186
rect 17486 4102 17514 4130
rect 14630 4046 14658 4074
rect 17038 4046 17066 4074
rect 23366 4046 23394 4074
rect 15414 3990 15442 4018
rect 16702 3990 16730 4018
rect 20286 3990 20314 4018
rect 17486 3934 17514 3962
rect 22638 3934 22666 3962
rect 1902 3906 1930 3934
rect 1954 3906 1982 3934
rect 2006 3906 2034 3934
rect 11902 3906 11930 3934
rect 11954 3906 11982 3934
rect 12006 3906 12034 3934
rect 21902 3906 21930 3934
rect 21954 3906 21982 3934
rect 22006 3906 22034 3934
rect 15134 3878 15162 3906
rect 21238 3878 21266 3906
rect 19390 3766 19418 3794
rect 7126 3654 7154 3682
rect 18494 3654 18522 3682
rect 21238 3654 21266 3682
rect 16590 3598 16618 3626
rect 2232 3514 2260 3542
rect 2284 3514 2312 3542
rect 2336 3514 2364 3542
rect 18550 3542 18578 3570
rect 12232 3514 12260 3542
rect 12284 3514 12312 3542
rect 12336 3514 12364 3542
rect 22232 3514 22260 3542
rect 22284 3514 22312 3542
rect 22336 3514 22364 3542
rect 15078 3486 15106 3514
rect 16590 3430 16618 3458
rect 18550 3374 18578 3402
rect 11830 3318 11858 3346
rect 16758 3318 16786 3346
rect 1902 3122 1930 3150
rect 1954 3122 1982 3150
rect 2006 3122 2034 3150
rect 11902 3122 11930 3150
rect 11954 3122 11982 3150
rect 12006 3122 12034 3150
rect 11830 3094 11858 3122
rect 21902 3122 21930 3150
rect 21954 3122 21982 3150
rect 22006 3122 22034 3150
rect 22134 3094 22162 3122
rect 22638 3038 22666 3066
rect 21126 2982 21154 3010
rect 21238 2926 21266 2954
rect 21014 2870 21042 2898
rect 21126 2870 21154 2898
rect 19278 2758 19306 2786
rect 22134 2758 22162 2786
rect 2232 2730 2260 2758
rect 2284 2730 2312 2758
rect 2336 2730 2364 2758
rect 12232 2730 12260 2758
rect 12284 2730 12312 2758
rect 12336 2730 12364 2758
rect 22232 2730 22260 2758
rect 22284 2730 22312 2758
rect 22336 2730 22364 2758
rect 15078 2646 15106 2674
rect 16646 2590 16674 2618
rect 19390 2590 19418 2618
rect 21014 2590 21042 2618
rect 18438 2534 18466 2562
rect 9982 2478 10010 2506
rect 13062 2422 13090 2450
rect 21238 2366 21266 2394
rect 1902 2338 1930 2366
rect 1954 2338 1982 2366
rect 2006 2338 2034 2366
rect 11902 2338 11930 2366
rect 11954 2338 11982 2366
rect 12006 2338 12034 2366
rect 21902 2338 21930 2366
rect 21954 2338 21982 2366
rect 22006 2338 22034 2366
rect 20174 2254 20202 2282
rect 13062 2198 13090 2226
rect 17598 2198 17626 2226
rect 11550 2142 11578 2170
rect 19278 1974 19306 2002
rect 2232 1946 2260 1974
rect 2284 1946 2312 1974
rect 2336 1946 2364 1974
rect 12232 1946 12260 1974
rect 12284 1946 12312 1974
rect 12336 1946 12364 1974
rect 22232 1946 22260 1974
rect 22284 1946 22312 1974
rect 22336 1946 22364 1974
rect 18438 1918 18466 1946
rect 10066 1862 10094 1890
rect 17262 1862 17290 1890
rect 11550 1694 11578 1722
rect 17598 1638 17626 1666
rect 1902 1554 1930 1582
rect 1954 1554 1982 1582
rect 2006 1554 2034 1582
rect 11902 1554 11930 1582
rect 11954 1554 11982 1582
rect 12006 1554 12034 1582
rect 21902 1554 21930 1582
rect 21954 1554 21982 1582
rect 22006 1554 22034 1582
rect 27286 1526 27314 1554
rect 19446 1470 19474 1498
rect 19446 1302 19474 1330
rect 27286 1302 27314 1330
rect 2232 1162 2260 1190
rect 2284 1162 2312 1190
rect 2336 1162 2364 1190
rect 12232 1162 12260 1190
rect 12284 1162 12312 1190
rect 12336 1162 12364 1190
rect 22232 1162 22260 1190
rect 22284 1162 22312 1190
rect 22336 1162 22364 1190
rect 1902 770 1930 798
rect 1954 770 1982 798
rect 2006 770 2034 798
rect 11902 770 11930 798
rect 11954 770 11982 798
rect 12006 770 12034 798
rect 21902 770 21930 798
rect 21954 770 21982 798
rect 22006 770 22034 798
rect 10094 742 10122 770
rect 17262 742 17290 770
rect 10094 574 10122 602
rect 14910 574 14938 602
rect 18438 574 18466 602
rect 4662 518 4690 546
rect 20398 518 20426 546
rect 4662 406 4690 434
rect 2232 378 2260 406
rect 2284 378 2312 406
rect 2336 378 2364 406
rect 12232 378 12260 406
rect 12284 378 12312 406
rect 12336 378 12364 406
rect 22232 378 22260 406
rect 22284 378 22312 406
rect 22336 378 22364 406
rect 13622 350 13650 378
rect 20174 294 20202 322
rect 14910 238 14938 266
rect 17038 14 17066 42
rect 20398 14 20426 42
<< metal4 >>
rect 1888 6286 2048 7112
rect 1888 6258 1902 6286
rect 1930 6258 1954 6286
rect 1982 6258 2006 6286
rect 2034 6258 2048 6286
rect 1888 5502 2048 6258
rect 1888 5474 1902 5502
rect 1930 5474 1954 5502
rect 1982 5474 2006 5502
rect 2034 5474 2048 5502
rect 1888 4718 2048 5474
rect 1888 4690 1902 4718
rect 1930 4690 1954 4718
rect 1982 4690 2006 4718
rect 2034 4690 2048 4718
rect 1888 3934 2048 4690
rect 1888 3906 1902 3934
rect 1930 3906 1954 3934
rect 1982 3906 2006 3934
rect 2034 3906 2048 3934
rect 1888 3150 2048 3906
rect 1888 3122 1902 3150
rect 1930 3122 1954 3150
rect 1982 3122 2006 3150
rect 2034 3122 2048 3150
rect 1888 2366 2048 3122
rect 1888 2338 1902 2366
rect 1930 2338 1954 2366
rect 1982 2338 2006 2366
rect 2034 2338 2048 2366
rect 1888 1582 2048 2338
rect 1888 1554 1902 1582
rect 1930 1554 1954 1582
rect 1982 1554 2006 1582
rect 2034 1554 2048 1582
rect 1888 798 2048 1554
rect 1888 770 1902 798
rect 1930 770 1954 798
rect 1982 770 2006 798
rect 2034 770 2048 798
rect 1888 0 2048 770
rect 2218 6678 2378 7112
rect 2218 6650 2232 6678
rect 2260 6650 2284 6678
rect 2312 6650 2336 6678
rect 2364 6650 2378 6678
rect 2218 5894 2378 6650
rect 2218 5866 2232 5894
rect 2260 5866 2284 5894
rect 2312 5866 2336 5894
rect 2364 5866 2378 5894
rect 2218 5110 2378 5866
rect 11888 6286 12048 7112
rect 11888 6258 11902 6286
rect 11930 6258 11954 6286
rect 11982 6258 12006 6286
rect 12034 6258 12048 6286
rect 10654 5698 10682 5703
rect 10654 5362 10682 5670
rect 10654 5329 10682 5334
rect 11888 5502 12048 6258
rect 11888 5474 11902 5502
rect 11930 5474 11954 5502
rect 11982 5474 12006 5502
rect 12034 5474 12048 5502
rect 2218 5082 2232 5110
rect 2260 5082 2284 5110
rect 2312 5082 2336 5110
rect 2364 5082 2378 5110
rect 2218 4326 2378 5082
rect 2218 4298 2232 4326
rect 2260 4298 2284 4326
rect 2312 4298 2336 4326
rect 2364 4298 2378 4326
rect 2218 3542 2378 4298
rect 6734 5138 6762 5143
rect 6734 4242 6762 5110
rect 10990 4914 11018 4919
rect 10990 4634 11018 4886
rect 10990 4601 11018 4606
rect 11888 4718 12048 5474
rect 11888 4690 11902 4718
rect 11930 4690 11954 4718
rect 11982 4690 12006 4718
rect 12034 4690 12048 4718
rect 6734 4209 6762 4214
rect 7126 4186 7154 4191
rect 7126 3682 7154 4158
rect 7126 3649 7154 3654
rect 11888 3934 12048 4690
rect 12218 6678 12378 7112
rect 12218 6650 12232 6678
rect 12260 6650 12284 6678
rect 12312 6650 12336 6678
rect 12364 6650 12378 6678
rect 12218 5894 12378 6650
rect 16702 6594 16730 6599
rect 16702 6539 16730 6566
rect 16926 6539 16954 6543
rect 16702 6538 16954 6539
rect 16702 6511 16926 6538
rect 16926 6505 16954 6510
rect 12218 5866 12232 5894
rect 12260 5866 12284 5894
rect 12312 5866 12336 5894
rect 12364 5866 12378 5894
rect 12218 5110 12378 5866
rect 13622 6426 13650 6431
rect 12614 5698 12642 5703
rect 12614 5418 12642 5670
rect 12614 5385 12642 5390
rect 12218 5082 12232 5110
rect 12260 5082 12284 5110
rect 12312 5082 12336 5110
rect 12364 5082 12378 5110
rect 13622 5138 13650 6398
rect 15694 6314 15722 6319
rect 14350 6258 14378 6263
rect 14294 6090 14322 6095
rect 14294 5922 14322 6062
rect 14294 5889 14322 5894
rect 13622 5105 13650 5110
rect 14182 5474 14210 5479
rect 12218 4326 12378 5082
rect 13902 4858 13930 4863
rect 13902 4746 13930 4830
rect 13902 4713 13930 4718
rect 14182 4466 14210 5446
rect 14238 5194 14266 5199
rect 14238 4690 14266 5166
rect 14350 4919 14378 6230
rect 15694 5866 15722 6286
rect 16702 6314 16730 6319
rect 15694 5833 15722 5838
rect 16254 6034 16282 6039
rect 16254 5418 16282 6006
rect 16254 5385 16282 5390
rect 16086 5306 16114 5311
rect 14294 4891 14378 4919
rect 14630 5250 14658 5255
rect 14294 4858 14322 4891
rect 14294 4825 14322 4830
rect 14238 4657 14266 4662
rect 14182 4433 14210 4438
rect 12110 4298 12138 4303
rect 12110 4186 12138 4270
rect 12110 4153 12138 4158
rect 12218 4298 12232 4326
rect 12260 4298 12284 4326
rect 12312 4298 12336 4326
rect 12364 4298 12378 4326
rect 11888 3906 11902 3934
rect 11930 3906 11954 3934
rect 11982 3906 12006 3934
rect 12034 3906 12048 3934
rect 2218 3514 2232 3542
rect 2260 3514 2284 3542
rect 2312 3514 2336 3542
rect 2364 3514 2378 3542
rect 2218 2758 2378 3514
rect 11830 3346 11858 3351
rect 11830 3122 11858 3318
rect 11830 3089 11858 3094
rect 11888 3150 12048 3906
rect 11888 3122 11902 3150
rect 11930 3122 11954 3150
rect 11982 3122 12006 3150
rect 12034 3122 12048 3150
rect 2218 2730 2232 2758
rect 2260 2730 2284 2758
rect 2312 2730 2336 2758
rect 2364 2730 2378 2758
rect 2218 1974 2378 2730
rect 2218 1946 2232 1974
rect 2260 1946 2284 1974
rect 2312 1946 2336 1974
rect 2364 1946 2378 1974
rect 2218 1190 2378 1946
rect 9982 2506 10010 2511
rect 9982 1949 10010 2478
rect 11888 2366 12048 3122
rect 11888 2338 11902 2366
rect 11930 2338 11954 2366
rect 11982 2338 12006 2366
rect 12034 2338 12048 2366
rect 11550 2170 11578 2175
rect 9982 1921 10094 1949
rect 10066 1890 10094 1921
rect 10066 1857 10094 1862
rect 11550 1722 11578 2142
rect 11550 1689 11578 1694
rect 2218 1162 2232 1190
rect 2260 1162 2284 1190
rect 2312 1162 2336 1190
rect 2364 1162 2378 1190
rect 2218 406 2378 1162
rect 11888 1582 12048 2338
rect 11888 1554 11902 1582
rect 11930 1554 11954 1582
rect 11982 1554 12006 1582
rect 12034 1554 12048 1582
rect 11888 798 12048 1554
rect 10094 770 10122 775
rect 10094 602 10122 742
rect 10094 569 10122 574
rect 11888 770 11902 798
rect 11930 770 11954 798
rect 11982 770 12006 798
rect 12034 770 12048 798
rect 2218 378 2232 406
rect 2260 378 2284 406
rect 2312 378 2336 406
rect 2364 378 2378 406
rect 4662 546 4690 551
rect 4662 434 4690 518
rect 4662 401 4690 406
rect 2218 0 2378 378
rect 11888 0 12048 770
rect 12218 3542 12378 4298
rect 12218 3514 12232 3542
rect 12260 3514 12284 3542
rect 12312 3514 12336 3542
rect 12364 3514 12378 3542
rect 12218 2758 12378 3514
rect 12218 2730 12232 2758
rect 12260 2730 12284 2758
rect 12312 2730 12336 2758
rect 12364 2730 12378 2758
rect 12218 1974 12378 2730
rect 13622 4298 13650 4303
rect 13062 2450 13090 2455
rect 13062 2226 13090 2422
rect 13062 2193 13090 2198
rect 12218 1946 12232 1974
rect 12260 1946 12284 1974
rect 12312 1946 12336 1974
rect 12364 1946 12378 1974
rect 12218 1190 12378 1946
rect 12218 1162 12232 1190
rect 12260 1162 12284 1190
rect 12312 1162 12336 1190
rect 12364 1162 12378 1190
rect 12218 406 12378 1162
rect 12218 378 12232 406
rect 12260 378 12284 406
rect 12312 378 12336 406
rect 12364 378 12378 406
rect 12218 0 12378 378
rect 13622 378 13650 4270
rect 14630 4074 14658 5222
rect 16086 5194 16114 5278
rect 16086 5161 16114 5166
rect 16646 4914 16674 4919
rect 14630 4041 14658 4046
rect 15134 4634 15162 4639
rect 15134 3906 15162 4606
rect 15414 4410 15442 4415
rect 15414 4018 15442 4382
rect 15414 3985 15442 3990
rect 15134 3873 15162 3878
rect 16590 3626 16618 3631
rect 15078 3514 15106 3519
rect 15078 2674 15106 3486
rect 16590 3458 16618 3598
rect 16590 3425 16618 3430
rect 15078 2641 15106 2646
rect 16646 2618 16674 4886
rect 16702 4018 16730 6286
rect 21888 6286 22048 7112
rect 21888 6258 21902 6286
rect 21930 6258 21954 6286
rect 21982 6258 22006 6286
rect 22034 6258 22048 6286
rect 21888 5502 22048 6258
rect 17598 5474 17626 5479
rect 17598 4914 17626 5446
rect 17598 4881 17626 4886
rect 21888 5474 21902 5502
rect 21930 5474 21954 5502
rect 21982 5474 22006 5502
rect 22034 5474 22048 5502
rect 20286 4858 20314 4863
rect 16702 3985 16730 3990
rect 16758 4354 16786 4359
rect 16758 3346 16786 4326
rect 17486 4130 17514 4135
rect 16758 3313 16786 3318
rect 17038 4074 17066 4079
rect 16646 2585 16674 2590
rect 13622 345 13650 350
rect 14910 602 14938 607
rect 14910 266 14938 574
rect 14910 233 14938 238
rect 17038 42 17066 4046
rect 17486 3962 17514 4102
rect 20286 4018 20314 4830
rect 20286 3985 20314 3990
rect 21888 4718 22048 5474
rect 21888 4690 21902 4718
rect 21930 4690 21954 4718
rect 21982 4690 22006 4718
rect 22034 4690 22048 4718
rect 17486 3929 17514 3934
rect 21888 3934 22048 4690
rect 21238 3906 21266 3911
rect 19390 3794 19418 3799
rect 18494 3682 18522 3687
rect 18494 2579 18522 3654
rect 18550 3570 18578 3575
rect 18550 3402 18578 3542
rect 18550 3369 18578 3374
rect 18438 2562 18522 2579
rect 18466 2551 18522 2562
rect 19278 2786 19306 2791
rect 18438 2529 18466 2534
rect 17598 2226 17626 2231
rect 17262 1890 17290 1895
rect 17262 770 17290 1862
rect 17598 1666 17626 2198
rect 19278 2002 19306 2758
rect 19390 2618 19418 3766
rect 21238 3682 21266 3878
rect 21238 3649 21266 3654
rect 21888 3906 21902 3934
rect 21930 3906 21954 3934
rect 21982 3906 22006 3934
rect 22034 3906 22048 3934
rect 21888 3150 22048 3906
rect 21888 3122 21902 3150
rect 21930 3122 21954 3150
rect 21982 3122 22006 3150
rect 22034 3122 22048 3150
rect 22218 6678 22378 7112
rect 22218 6650 22232 6678
rect 22260 6650 22284 6678
rect 22312 6650 22336 6678
rect 22364 6650 22378 6678
rect 22218 5894 22378 6650
rect 22218 5866 22232 5894
rect 22260 5866 22284 5894
rect 22312 5866 22336 5894
rect 22364 5866 22378 5894
rect 22218 5110 22378 5866
rect 22218 5082 22232 5110
rect 22260 5082 22284 5110
rect 22312 5082 22336 5110
rect 22364 5082 22378 5110
rect 22218 4326 22378 5082
rect 22218 4298 22232 4326
rect 22260 4298 22284 4326
rect 22312 4298 22336 4326
rect 22364 4298 22378 4326
rect 22218 3542 22378 4298
rect 23366 5978 23394 5983
rect 23366 4074 23394 5950
rect 23366 4041 23394 4046
rect 22218 3514 22232 3542
rect 22260 3514 22284 3542
rect 22312 3514 22336 3542
rect 22364 3514 22378 3542
rect 21126 3010 21154 3015
rect 19390 2585 19418 2590
rect 21014 2898 21042 2903
rect 21014 2618 21042 2870
rect 21126 2898 21154 2982
rect 21126 2865 21154 2870
rect 21238 2954 21266 2959
rect 21014 2585 21042 2590
rect 21238 2394 21266 2926
rect 21238 2361 21266 2366
rect 21888 2366 22048 3122
rect 22134 3122 22162 3127
rect 22134 2786 22162 3094
rect 22134 2753 22162 2758
rect 22218 2758 22378 3514
rect 22638 3962 22666 3967
rect 22638 3066 22666 3934
rect 22638 3033 22666 3038
rect 21888 2338 21902 2366
rect 21930 2338 21954 2366
rect 21982 2338 22006 2366
rect 22034 2338 22048 2366
rect 19278 1969 19306 1974
rect 20174 2282 20202 2287
rect 17598 1633 17626 1638
rect 18438 1946 18466 1951
rect 17262 737 17290 742
rect 18438 602 18466 1918
rect 19446 1498 19474 1503
rect 19446 1330 19474 1470
rect 19446 1297 19474 1302
rect 18438 569 18466 574
rect 20174 322 20202 2254
rect 21888 1582 22048 2338
rect 21888 1554 21902 1582
rect 21930 1554 21954 1582
rect 21982 1554 22006 1582
rect 22034 1554 22048 1582
rect 21888 798 22048 1554
rect 21888 770 21902 798
rect 21930 770 21954 798
rect 21982 770 22006 798
rect 22034 770 22048 798
rect 20174 289 20202 294
rect 20398 546 20426 551
rect 17038 9 17066 14
rect 20398 42 20426 518
rect 20398 9 20426 14
rect 21888 0 22048 770
rect 22218 2730 22232 2758
rect 22260 2730 22284 2758
rect 22312 2730 22336 2758
rect 22364 2730 22378 2758
rect 22218 1974 22378 2730
rect 22218 1946 22232 1974
rect 22260 1946 22284 1974
rect 22312 1946 22336 1974
rect 22364 1946 22378 1974
rect 22218 1190 22378 1946
rect 27286 1554 27314 1559
rect 27286 1330 27314 1526
rect 27286 1297 27314 1302
rect 22218 1162 22232 1190
rect 22260 1162 22284 1190
rect 22312 1162 22336 1190
rect 22364 1162 22378 1190
rect 22218 406 22378 1162
rect 22218 378 22232 406
rect 22260 378 22284 406
rect 22312 378 22336 406
rect 22364 378 22378 406
rect 22218 0 22378 378
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _000_
timestamp 1486834041
transform 1 0 4928 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _001_
timestamp 1486834041
transform 1 0 4928 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _002_
timestamp 1486834041
transform 1 0 28840 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _003_
timestamp 1486834041
transform 1 0 28448 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _004_
timestamp 1486834041
transform 1 0 4480 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _005_
timestamp 1486834041
transform 1 0 29624 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _006_
timestamp 1486834041
transform 1 0 29624 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _007_
timestamp 1486834041
transform 1 0 29288 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _008_
timestamp 1486834041
transform 1 0 28896 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _009_
timestamp 1486834041
transform 1 0 2520 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _010_
timestamp 1486834041
transform 1 0 28280 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _011_
timestamp 1486834041
transform 1 0 28840 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _012_
timestamp 1486834041
transform 1 0 29624 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _013_
timestamp 1486834041
transform 1 0 6160 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _014_
timestamp 1486834041
transform 1 0 8568 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _015_
timestamp 1486834041
transform 1 0 10416 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _016_
timestamp 1486834041
transform 1 0 10752 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _017_
timestamp 1486834041
transform 1 0 29288 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _018_
timestamp 1486834041
transform 1 0 6160 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _019_
timestamp 1486834041
transform -1 0 31472 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _020_
timestamp 1486834041
transform 1 0 29624 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _021_
timestamp 1486834041
transform 1 0 6440 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _022_
timestamp 1486834041
transform 1 0 28616 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _023_
timestamp 1486834041
transform 1 0 3808 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _024_
timestamp 1486834041
transform 1 0 27888 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _025_
timestamp 1486834041
transform 1 0 2408 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _026_
timestamp 1486834041
transform 1 0 27888 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _027_
timestamp 1486834041
transform 1 0 29232 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _028_
timestamp 1486834041
transform 1 0 28840 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _029_
timestamp 1486834041
transform 1 0 28504 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _030_
timestamp 1486834041
transform 1 0 2296 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _031_
timestamp 1486834041
transform 1 0 29288 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _032_
timestamp 1486834041
transform 1 0 13944 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _033_
timestamp 1486834041
transform 1 0 14560 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _034_
timestamp 1486834041
transform 1 0 17528 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _035_
timestamp 1486834041
transform 1 0 20328 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _036_
timestamp 1486834041
transform 1 0 21448 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _037_
timestamp 1486834041
transform 1 0 21448 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _038_
timestamp 1486834041
transform 1 0 22008 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _039_
timestamp 1486834041
transform 1 0 22120 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _040_
timestamp 1486834041
transform 1 0 23968 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _041_
timestamp 1486834041
transform 1 0 24528 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _042_
timestamp 1486834041
transform 1 0 25088 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _043_
timestamp 1486834041
transform 1 0 23744 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _044_
timestamp 1486834041
transform 1 0 25088 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _045_
timestamp 1486834041
transform 1 0 25144 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _046_
timestamp 1486834041
transform -1 0 14896 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _047_
timestamp 1486834041
transform -1 0 20496 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _048_
timestamp 1486834041
transform -1 0 22064 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _049_
timestamp 1486834041
transform -1 0 23464 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _050_
timestamp 1486834041
transform -1 0 26376 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _051_
timestamp 1486834041
transform -1 0 28168 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _052_
timestamp 1486834041
transform -1 0 1344 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _053_
timestamp 1486834041
transform -1 0 4424 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _054_
timestamp 1486834041
transform -1 0 8176 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _055_
timestamp 1486834041
transform -1 0 11536 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _056_
timestamp 1486834041
transform -1 0 8736 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _057_
timestamp 1486834041
transform -1 0 8736 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _058_
timestamp 1486834041
transform -1 0 9744 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _059_
timestamp 1486834041
transform -1 0 7728 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _060_
timestamp 1486834041
transform -1 0 12096 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _061_
timestamp 1486834041
transform -1 0 14896 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _062_
timestamp 1486834041
transform 1 0 17360 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _063_
timestamp 1486834041
transform -1 0 12656 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _064_
timestamp 1486834041
transform 1 0 26320 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _065_
timestamp 1486834041
transform 1 0 28840 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _066_
timestamp 1486834041
transform 1 0 28392 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _067_
timestamp 1486834041
transform 1 0 29176 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _068_
timestamp 1486834041
transform 1 0 23408 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _069_
timestamp 1486834041
transform 1 0 28056 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _070_
timestamp 1486834041
transform 1 0 20104 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _071_
timestamp 1486834041
transform 1 0 21392 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _072_
timestamp 1486834041
transform -1 0 16576 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _073_
timestamp 1486834041
transform -1 0 15176 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _074_
timestamp 1486834041
transform -1 0 8624 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _075_
timestamp 1486834041
transform -1 0 1288 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _076_
timestamp 1486834041
transform -1 0 1400 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _077_
timestamp 1486834041
transform -1 0 1344 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _078_
timestamp 1486834041
transform -1 0 1288 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _079_
timestamp 1486834041
transform -1 0 1344 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _080_
timestamp 1486834041
transform -1 0 9128 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _081_
timestamp 1486834041
transform -1 0 11032 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _082_
timestamp 1486834041
transform -1 0 1288 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _083_
timestamp 1486834041
transform -1 0 7728 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _084_
timestamp 1486834041
transform -1 0 15456 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _085_
timestamp 1486834041
transform -1 0 13664 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _086_
timestamp 1486834041
transform -1 0 18536 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _087_
timestamp 1486834041
transform -1 0 1736 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _088_
timestamp 1486834041
transform -1 0 25368 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _089_
timestamp 1486834041
transform -1 0 23632 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _090_
timestamp 1486834041
transform -1 0 24640 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _091_
timestamp 1486834041
transform -1 0 23016 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _092_
timestamp 1486834041
transform -1 0 21896 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _093_
timestamp 1486834041
transform -1 0 21000 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _094_
timestamp 1486834041
transform -1 0 21448 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _095_
timestamp 1486834041
transform -1 0 21280 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _096_
timestamp 1486834041
transform -1 0 21392 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _097_
timestamp 1486834041
transform -1 0 21224 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _098_
timestamp 1486834041
transform -1 0 20608 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _099_
timestamp 1486834041
transform -1 0 19152 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _100_
timestamp 1486834041
transform -1 0 18536 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _101_
timestamp 1486834041
transform -1 0 19824 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _102_
timestamp 1486834041
transform -1 0 18032 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _103_
timestamp 1486834041
transform -1 0 15568 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _104_
timestamp 1486834041
transform 1 0 15176 0 -1 1176
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__000__I
timestamp 1486834041
transform -1 0 4816 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__001__I
timestamp 1486834041
transform 1 0 4816 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__002__I
timestamp 1486834041
transform -1 0 28840 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__003__I
timestamp 1486834041
transform 1 0 28336 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__004__I
timestamp 1486834041
transform 1 0 4368 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__005__I
timestamp 1486834041
transform -1 0 29624 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__006__I
timestamp 1486834041
transform 1 0 29512 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__007__I
timestamp 1486834041
transform -1 0 29288 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__008__I
timestamp 1486834041
transform -1 0 28896 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__009__I
timestamp 1486834041
transform -1 0 2520 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__010__I
timestamp 1486834041
transform 1 0 28168 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__011__I
timestamp 1486834041
transform 1 0 28728 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__012__I
timestamp 1486834041
transform -1 0 29624 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__013__I
timestamp 1486834041
transform 1 0 6048 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__014__I
timestamp 1486834041
transform -1 0 8568 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__015__I
timestamp 1486834041
transform -1 0 10416 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__016__I
timestamp 1486834041
transform -1 0 10752 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__017__I
timestamp 1486834041
transform 1 0 29176 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__018__I
timestamp 1486834041
transform -1 0 6160 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__019__I
timestamp 1486834041
transform 1 0 31472 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__020__I
timestamp 1486834041
transform -1 0 28952 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__021__I
timestamp 1486834041
transform -1 0 6440 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__022__I
timestamp 1486834041
transform 1 0 28504 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__023__I
timestamp 1486834041
transform -1 0 3808 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__024__I
timestamp 1486834041
transform -1 0 27776 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__025__I
timestamp 1486834041
transform 1 0 2184 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__026__I
timestamp 1486834041
transform -1 0 27776 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__027__I
timestamp 1486834041
transform 1 0 29120 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__028__I
timestamp 1486834041
transform -1 0 28840 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__029__I
timestamp 1486834041
transform 1 0 28392 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__030__I
timestamp 1486834041
transform -1 0 2296 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__031__I
timestamp 1486834041
transform -1 0 29176 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__032__I
timestamp 1486834041
transform 1 0 13832 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__033__I
timestamp 1486834041
transform -1 0 14560 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__034__I
timestamp 1486834041
transform -1 0 17528 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__035__I
timestamp 1486834041
transform -1 0 20328 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__036__I
timestamp 1486834041
transform -1 0 21448 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__037__I
timestamp 1486834041
transform -1 0 21448 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__038__I
timestamp 1486834041
transform -1 0 21896 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__039__I
timestamp 1486834041
transform 1 0 22008 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__040__I
timestamp 1486834041
transform 1 0 23744 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__041__I
timestamp 1486834041
transform 1 0 24416 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__042__I
timestamp 1486834041
transform 1 0 24976 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__043__I
timestamp 1486834041
transform -1 0 23744 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__044__I
timestamp 1486834041
transform 1 0 24976 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__045__I
timestamp 1486834041
transform 1 0 25032 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__046__I
timestamp 1486834041
transform 1 0 14896 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__047__I
timestamp 1486834041
transform 1 0 20496 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__048__I
timestamp 1486834041
transform 1 0 22064 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__049__I
timestamp 1486834041
transform 1 0 23464 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__050__I
timestamp 1486834041
transform -1 0 26488 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__051__I
timestamp 1486834041
transform -1 0 28280 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__052__I
timestamp 1486834041
transform -1 0 1456 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__053__I
timestamp 1486834041
transform 1 0 4424 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__054__I
timestamp 1486834041
transform -1 0 8400 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__055__I
timestamp 1486834041
transform -1 0 11648 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__056__I
timestamp 1486834041
transform -1 0 8848 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__057__I
timestamp 1486834041
transform -1 0 8848 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__058__I
timestamp 1486834041
transform -1 0 9856 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__059__I
timestamp 1486834041
transform -1 0 7840 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__060__I
timestamp 1486834041
transform -1 0 12320 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__061__I
timestamp 1486834041
transform 1 0 14896 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__062__I
timestamp 1486834041
transform 1 0 17248 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__063__I
timestamp 1486834041
transform -1 0 12768 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__064__I
timestamp 1486834041
transform 1 0 26208 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__065__I
timestamp 1486834041
transform 1 0 28616 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__066__I
timestamp 1486834041
transform -1 0 28392 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__067__I
timestamp 1486834041
transform -1 0 29064 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__068__I
timestamp 1486834041
transform -1 0 23408 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__069__I
timestamp 1486834041
transform 1 0 27944 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__070__I
timestamp 1486834041
transform -1 0 19936 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__071__I
timestamp 1486834041
transform -1 0 21392 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__072__I
timestamp 1486834041
transform -1 0 16688 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__073__I
timestamp 1486834041
transform 1 0 15176 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__074__I
timestamp 1486834041
transform 1 0 8624 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__075__I
timestamp 1486834041
transform 1 0 1288 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__076__I
timestamp 1486834041
transform -1 0 1512 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__077__I
timestamp 1486834041
transform -1 0 1456 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__078__I
timestamp 1486834041
transform 1 0 1288 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__079__I
timestamp 1486834041
transform 1 0 1344 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__080__I
timestamp 1486834041
transform -1 0 9240 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__081__I
timestamp 1486834041
transform -1 0 11144 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__082__I
timestamp 1486834041
transform -1 0 1400 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__083__I
timestamp 1486834041
transform 1 0 7728 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__084__I
timestamp 1486834041
transform -1 0 15568 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__085__I
timestamp 1486834041
transform 1 0 13664 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__086__I
timestamp 1486834041
transform 1 0 18536 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__087__I
timestamp 1486834041
transform 1 0 1736 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__088__I
timestamp 1486834041
transform 1 0 25368 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__089__I
timestamp 1486834041
transform -1 0 23744 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__090__I
timestamp 1486834041
transform 1 0 24640 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__091__I
timestamp 1486834041
transform -1 0 23128 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__092__I
timestamp 1486834041
transform -1 0 22008 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__093__I
timestamp 1486834041
transform -1 0 21112 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__094__I
timestamp 1486834041
transform -1 0 21560 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__095__I
timestamp 1486834041
transform 1 0 21280 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__096__I
timestamp 1486834041
transform 1 0 21392 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__097__I
timestamp 1486834041
transform 1 0 21224 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__098__I
timestamp 1486834041
transform 1 0 20608 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__099__I
timestamp 1486834041
transform -1 0 19264 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__100__I
timestamp 1486834041
transform -1 0 18648 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__101__I
timestamp 1486834041
transform -1 0 19936 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__102__I
timestamp 1486834041
transform -1 0 18144 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__103__I
timestamp 1486834041
transform 1 0 15568 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__104__I
timestamp 1486834041
transform 1 0 15064 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2
timestamp 1486834041
transform 1 0 448 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6
timestamp 1486834041
transform 1 0 672 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8
timestamp 1486834041
transform 1 0 784 0 1 392
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19
timestamp 1486834041
transform 1 0 1400 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27
timestamp 1486834041
transform 1 0 1848 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31
timestamp 1486834041
transform 1 0 2072 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33
timestamp 1486834041
transform 1 0 2184 0 1 392
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36
timestamp 1486834041
transform 1 0 2352 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70
timestamp 1486834041
transform 1 0 4256 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_90
timestamp 1486834041
transform 1 0 5376 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_98
timestamp 1486834041
transform 1 0 5824 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_104
timestamp 1486834041
transform 1 0 6160 0 1 392
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_120
timestamp 1486834041
transform 1 0 7056 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_128
timestamp 1486834041
transform 1 0 7504 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_134
timestamp 1486834041
transform 1 0 7840 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_138
timestamp 1486834041
transform 1 0 8064 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_172
timestamp 1486834041
transform 1 0 9968 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_206
timestamp 1486834041
transform 1 0 11872 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_240
timestamp 1486834041
transform 1 0 13776 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_274
timestamp 1486834041
transform 1 0 15680 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_308
timestamp 1486834041
transform 1 0 17584 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_318
timestamp 1486834041
transform 1 0 18144 0 1 392
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_334
timestamp 1486834041
transform 1 0 19040 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_338
timestamp 1486834041
transform 1 0 19264 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_342
timestamp 1486834041
transform 1 0 19488 0 1 392
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_358
timestamp 1486834041
transform 1 0 20384 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_366
timestamp 1486834041
transform 1 0 20832 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_368
timestamp 1486834041
transform 1 0 20944 0 1 392
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_371
timestamp 1486834041
transform 1 0 21112 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_373
timestamp 1486834041
transform 1 0 21224 0 1 392
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_376
timestamp 1486834041
transform 1 0 21392 0 1 392
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_379
timestamp 1486834041
transform 1 0 21560 0 1 392
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_395
timestamp 1486834041
transform 1 0 22456 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_403
timestamp 1486834041
transform 1 0 22904 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_407
timestamp 1486834041
transform 1 0 23128 0 1 392
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_410
timestamp 1486834041
transform 1 0 23296 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_444
timestamp 1486834041
transform 1 0 25200 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_478
timestamp 1486834041
transform 1 0 27104 0 1 392
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_494
timestamp 1486834041
transform 1 0 28000 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_502
timestamp 1486834041
transform 1 0 28448 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_506
timestamp 1486834041
transform 1 0 28672 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_512
timestamp 1486834041
transform 1 0 29008 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_546
timestamp 1486834041
transform 1 0 30912 0 1 392
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_2
timestamp 1486834041
transform 1 0 448 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_20
timestamp 1486834041
transform 1 0 1456 0 -1 1176
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_52
timestamp 1486834041
transform 1 0 3248 0 -1 1176
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_68
timestamp 1486834041
transform 1 0 4144 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_90
timestamp 1486834041
transform 1 0 5376 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_98
timestamp 1486834041
transform 1 0 5824 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_112
timestamp 1486834041
transform 1 0 6608 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_120
timestamp 1486834041
transform 1 0 7056 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_144
timestamp 1486834041
transform 1 0 8400 0 -1 1176
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_176
timestamp 1486834041
transform 1 0 10192 0 -1 1176
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_202
timestamp 1486834041
transform 1 0 11648 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_212
timestamp 1486834041
transform 1 0 12208 0 -1 1176
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_244
timestamp 1486834041
transform 1 0 14000 0 -1 1176
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_260
timestamp 1486834041
transform 1 0 14896 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_262
timestamp 1486834041
transform 1 0 15008 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_271
timestamp 1486834041
transform 1 0 15512 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_279
timestamp 1486834041
transform 1 0 15960 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_292
timestamp 1486834041
transform 1 0 16688 0 -1 1176
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_316
timestamp 1486834041
transform 1 0 18032 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_327
timestamp 1486834041
transform 1 0 18648 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_338
timestamp 1486834041
transform 1 0 19264 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_352
timestamp 1486834041
transform 1 0 20048 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_360
timestamp 1486834041
transform 1 0 20496 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_387
timestamp 1486834041
transform 1 0 22008 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_395
timestamp 1486834041
transform 1 0 22456 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_407
timestamp 1486834041
transform 1 0 23128 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_415
timestamp 1486834041
transform 1 0 23576 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_417
timestamp 1486834041
transform 1 0 23688 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_450
timestamp 1486834041
transform 1 0 25536 0 -1 1176
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_482
timestamp 1486834041
transform 1 0 27328 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_492
timestamp 1486834041
transform 1 0 27888 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_518
timestamp 1486834041
transform 1 0 29344 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_520
timestamp 1486834041
transform 1 0 29456 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_2
timestamp 1486834041
transform 1 0 448 0 1 1176
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1486834041
transform 1 0 2240 0 1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_37
timestamp 1486834041
transform 1 0 2408 0 1 1176
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_101
timestamp 1486834041
transform 1 0 5992 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_107
timestamp 1486834041
transform 1 0 6328 0 1 1176
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_171
timestamp 1486834041
transform 1 0 9912 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_177
timestamp 1486834041
transform 1 0 10248 0 1 1176
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_241
timestamp 1486834041
transform 1 0 13832 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_247
timestamp 1486834041
transform 1 0 14168 0 1 1176
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_311
timestamp 1486834041
transform 1 0 17752 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_317
timestamp 1486834041
transform 1 0 18088 0 1 1176
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_381
timestamp 1486834041
transform 1 0 21672 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_387
timestamp 1486834041
transform 1 0 22008 0 1 1176
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_451
timestamp 1486834041
transform 1 0 25592 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_467
timestamp 1486834041
transform 1 0 26488 0 1 1176
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_499
timestamp 1486834041
transform 1 0 28280 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_527
timestamp 1486834041
transform 1 0 29848 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_531
timestamp 1486834041
transform 1 0 30072 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_2
timestamp 1486834041
transform 1 0 448 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_10
timestamp 1486834041
transform 1 0 896 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_21
timestamp 1486834041
transform 1 0 1512 0 -1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_47
timestamp 1486834041
transform 1 0 2968 0 -1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_63
timestamp 1486834041
transform 1 0 3864 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_67
timestamp 1486834041
transform 1 0 4088 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_69
timestamp 1486834041
transform 1 0 4200 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_72
timestamp 1486834041
transform 1 0 4368 0 -1 1960
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_136
timestamp 1486834041
transform 1 0 7952 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_152
timestamp 1486834041
transform 1 0 8848 0 -1 1960
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_184
timestamp 1486834041
transform 1 0 10640 0 -1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_200
timestamp 1486834041
transform 1 0 11536 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_214
timestamp 1486834041
transform 1 0 12320 0 -1 1960
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_278
timestamp 1486834041
transform 1 0 15904 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_282
timestamp 1486834041
transform 1 0 16128 0 -1 1960
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_346
timestamp 1486834041
transform 1 0 19712 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_362
timestamp 1486834041
transform 1 0 20608 0 -1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_378
timestamp 1486834041
transform 1 0 21504 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_386
timestamp 1486834041
transform 1 0 21952 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_397
timestamp 1486834041
transform 1 0 22568 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_405
timestamp 1486834041
transform 1 0 23016 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_407
timestamp 1486834041
transform 1 0 23128 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_418
timestamp 1486834041
transform 1 0 23744 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_422
timestamp 1486834041
transform 1 0 23968 0 -1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_438
timestamp 1486834041
transform 1 0 24864 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_449
timestamp 1486834041
transform 1 0 25480 0 -1 1960
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_481
timestamp 1486834041
transform 1 0 27272 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_489
timestamp 1486834041
transform 1 0 27720 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_492
timestamp 1486834041
transform 1 0 27888 0 -1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_508
timestamp 1486834041
transform 1 0 28784 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_512
timestamp 1486834041
transform 1 0 29008 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_514
timestamp 1486834041
transform 1 0 29120 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_517
timestamp 1486834041
transform 1 0 29288 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_2
timestamp 1486834041
transform 1 0 448 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_6
timestamp 1486834041
transform 1 0 672 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_8
timestamp 1486834041
transform 1 0 784 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_19
timestamp 1486834041
transform 1 0 1400 0 1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_37
timestamp 1486834041
transform 1 0 2408 0 1 1960
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_101
timestamp 1486834041
transform 1 0 5992 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_107
timestamp 1486834041
transform 1 0 6328 0 1 1960
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_139
timestamp 1486834041
transform 1 0 8120 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_150
timestamp 1486834041
transform 1 0 8736 0 1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_166
timestamp 1486834041
transform 1 0 9632 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_174
timestamp 1486834041
transform 1 0 10080 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_177
timestamp 1486834041
transform 1 0 10248 0 1 1960
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_241
timestamp 1486834041
transform 1 0 13832 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_247
timestamp 1486834041
transform 1 0 14168 0 1 1960
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_311
timestamp 1486834041
transform 1 0 17752 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_317
timestamp 1486834041
transform 1 0 18088 0 1 1960
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_349
timestamp 1486834041
transform 1 0 19880 0 1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_365
timestamp 1486834041
transform 1 0 20776 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_367
timestamp 1486834041
transform 1 0 20888 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_378
timestamp 1486834041
transform 1 0 21504 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_382
timestamp 1486834041
transform 1 0 21728 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_384
timestamp 1486834041
transform 1 0 21840 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_387
timestamp 1486834041
transform 1 0 22008 0 1 1960
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_419
timestamp 1486834041
transform 1 0 23800 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_423
timestamp 1486834041
transform 1 0 24024 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_425
timestamp 1486834041
transform 1 0 24136 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_436
timestamp 1486834041
transform 1 0 24752 0 1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_452
timestamp 1486834041
transform 1 0 25648 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_454
timestamp 1486834041
transform 1 0 25760 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_457
timestamp 1486834041
transform 1 0 25928 0 1 1960
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_499
timestamp 1486834041
transform 1 0 28280 0 1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_515
timestamp 1486834041
transform 1 0 29176 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_523
timestamp 1486834041
transform 1 0 29624 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_527
timestamp 1486834041
transform 1 0 29848 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_531
timestamp 1486834041
transform 1 0 30072 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_2
timestamp 1486834041
transform 1 0 448 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_20
timestamp 1486834041
transform 1 0 1456 0 -1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_52
timestamp 1486834041
transform 1 0 3248 0 -1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_68
timestamp 1486834041
transform 1 0 4144 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_72
timestamp 1486834041
transform 1 0 4368 0 -1 2744
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_136
timestamp 1486834041
transform 1 0 7952 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_152
timestamp 1486834041
transform 1 0 8848 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_170
timestamp 1486834041
transform 1 0 9856 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_178
timestamp 1486834041
transform 1 0 10304 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_182
timestamp 1486834041
transform 1 0 10528 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_193
timestamp 1486834041
transform 1 0 11144 0 -1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_209
timestamp 1486834041
transform 1 0 12040 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_222
timestamp 1486834041
transform 1 0 12768 0 -1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_238
timestamp 1486834041
transform 1 0 13664 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_246
timestamp 1486834041
transform 1 0 14112 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_250
timestamp 1486834041
transform 1 0 14336 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_262
timestamp 1486834041
transform 1 0 15008 0 -1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_278
timestamp 1486834041
transform 1 0 15904 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_282
timestamp 1486834041
transform 1 0 16128 0 -1 2744
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_346
timestamp 1486834041
transform 1 0 19712 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_352
timestamp 1486834041
transform 1 0 20048 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_361
timestamp 1486834041
transform 1 0 20552 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_365
timestamp 1486834041
transform 1 0 20776 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_384
timestamp 1486834041
transform 1 0 21840 0 -1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_416
timestamp 1486834041
transform 1 0 23632 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_422
timestamp 1486834041
transform 1 0 23968 0 -1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_438
timestamp 1486834041
transform 1 0 24864 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_450
timestamp 1486834041
transform 1 0 25536 0 -1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_482
timestamp 1486834041
transform 1 0 27328 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_492
timestamp 1486834041
transform 1 0 27888 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_496
timestamp 1486834041
transform 1 0 28112 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_517
timestamp 1486834041
transform 1 0 29288 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_2
timestamp 1486834041
transform 1 0 448 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_20
timestamp 1486834041
transform 1 0 1456 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_28
timestamp 1486834041
transform 1 0 1904 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_32
timestamp 1486834041
transform 1 0 2128 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1486834041
transform 1 0 2240 0 1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_37
timestamp 1486834041
transform 1 0 2408 0 1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_53
timestamp 1486834041
transform 1 0 3304 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_61
timestamp 1486834041
transform 1 0 3752 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_75
timestamp 1486834041
transform 1 0 4536 0 1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_91
timestamp 1486834041
transform 1 0 5432 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_99
timestamp 1486834041
transform 1 0 5880 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_103
timestamp 1486834041
transform 1 0 6104 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_107
timestamp 1486834041
transform 1 0 6328 0 1 2744
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_171
timestamp 1486834041
transform 1 0 9912 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_177
timestamp 1486834041
transform 1 0 10248 0 1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_209
timestamp 1486834041
transform 1 0 12040 0 1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_225
timestamp 1486834041
transform 1 0 12936 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_229
timestamp 1486834041
transform 1 0 13160 0 1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_240
timestamp 1486834041
transform 1 0 13776 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_244
timestamp 1486834041
transform 1 0 14000 0 1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_247
timestamp 1486834041
transform 1 0 14168 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_255
timestamp 1486834041
transform 1 0 14616 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_267
timestamp 1486834041
transform 1 0 15288 0 1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_299
timestamp 1486834041
transform 1 0 17080 0 1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_317
timestamp 1486834041
transform 1 0 18088 0 1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_349
timestamp 1486834041
transform 1 0 19880 0 1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_365
timestamp 1486834041
transform 1 0 20776 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_373
timestamp 1486834041
transform 1 0 21224 0 1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_376
timestamp 1486834041
transform 1 0 21392 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_380
timestamp 1486834041
transform 1 0 21616 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_382
timestamp 1486834041
transform 1 0 21728 0 1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_395
timestamp 1486834041
transform 1 0 22456 0 1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_427
timestamp 1486834041
transform 1 0 24248 0 1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_443
timestamp 1486834041
transform 1 0 25144 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_451
timestamp 1486834041
transform 1 0 25592 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_457
timestamp 1486834041
transform 1 0 25928 0 1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_489
timestamp 1486834041
transform 1 0 27720 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_497
timestamp 1486834041
transform 1 0 28168 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_501
timestamp 1486834041
transform 1 0 28392 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_513
timestamp 1486834041
transform 1 0 29064 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_527
timestamp 1486834041
transform 1 0 29848 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_531
timestamp 1486834041
transform 1 0 30072 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_2
timestamp 1486834041
transform 1 0 448 0 -1 3528
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_66
timestamp 1486834041
transform 1 0 4032 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_72
timestamp 1486834041
transform 1 0 4368 0 -1 3528
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_136
timestamp 1486834041
transform 1 0 7952 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_142
timestamp 1486834041
transform 1 0 8288 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_146
timestamp 1486834041
transform 1 0 8512 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_148
timestamp 1486834041
transform 1 0 8624 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_159
timestamp 1486834041
transform 1 0 9240 0 -1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_191
timestamp 1486834041
transform 1 0 11032 0 -1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_207
timestamp 1486834041
transform 1 0 11928 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_209
timestamp 1486834041
transform 1 0 12040 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_212
timestamp 1486834041
transform 1 0 12208 0 -1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_244
timestamp 1486834041
transform 1 0 14000 0 -1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_260
timestamp 1486834041
transform 1 0 14896 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_272
timestamp 1486834041
transform 1 0 15568 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_282
timestamp 1486834041
transform 1 0 16128 0 -1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_314
timestamp 1486834041
transform 1 0 17920 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_316
timestamp 1486834041
transform 1 0 18032 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_327
timestamp 1486834041
transform 1 0 18648 0 -1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_343
timestamp 1486834041
transform 1 0 19544 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_347
timestamp 1486834041
transform 1 0 19768 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_349
timestamp 1486834041
transform 1 0 19880 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_352
timestamp 1486834041
transform 1 0 20048 0 -1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_384
timestamp 1486834041
transform 1 0 21840 0 -1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_400
timestamp 1486834041
transform 1 0 22736 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_408
timestamp 1486834041
transform 1 0 23184 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_422
timestamp 1486834041
transform 1 0 23968 0 -1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_438
timestamp 1486834041
transform 1 0 24864 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_440
timestamp 1486834041
transform 1 0 24976 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_451
timestamp 1486834041
transform 1 0 25592 0 -1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_483
timestamp 1486834041
transform 1 0 27384 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_487
timestamp 1486834041
transform 1 0 27608 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_489
timestamp 1486834041
transform 1 0 27720 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_492
timestamp 1486834041
transform 1 0 27888 0 -1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_508
timestamp 1486834041
transform 1 0 28784 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1486834041
transform 1 0 448 0 1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1486834041
transform 1 0 2240 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_37
timestamp 1486834041
transform 1 0 2408 0 1 3528
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_101
timestamp 1486834041
transform 1 0 5992 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_107
timestamp 1486834041
transform 1 0 6328 0 1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_123
timestamp 1486834041
transform 1 0 7224 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_134
timestamp 1486834041
transform 1 0 7840 0 1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_166
timestamp 1486834041
transform 1 0 9632 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_174
timestamp 1486834041
transform 1 0 10080 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_177
timestamp 1486834041
transform 1 0 10248 0 1 3528
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_241
timestamp 1486834041
transform 1 0 13832 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_247
timestamp 1486834041
transform 1 0 14168 0 1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_279
timestamp 1486834041
transform 1 0 15960 0 1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_295
timestamp 1486834041
transform 1 0 16856 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_299
timestamp 1486834041
transform 1 0 17080 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_301
timestamp 1486834041
transform 1 0 17192 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_312
timestamp 1486834041
transform 1 0 17808 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_314
timestamp 1486834041
transform 1 0 17920 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_317
timestamp 1486834041
transform 1 0 18088 0 1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_349
timestamp 1486834041
transform 1 0 19880 0 1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_375
timestamp 1486834041
transform 1 0 21336 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_383
timestamp 1486834041
transform 1 0 21784 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_387
timestamp 1486834041
transform 1 0 22008 0 1 3528
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_451
timestamp 1486834041
transform 1 0 25592 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_457
timestamp 1486834041
transform 1 0 25928 0 1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_489
timestamp 1486834041
transform 1 0 27720 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_497
timestamp 1486834041
transform 1 0 28168 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_501
timestamp 1486834041
transform 1 0 28392 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_527
timestamp 1486834041
transform 1 0 29848 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_531
timestamp 1486834041
transform 1 0 30072 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_2
timestamp 1486834041
transform 1 0 448 0 -1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_18
timestamp 1486834041
transform 1 0 1344 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_26
timestamp 1486834041
transform 1 0 1792 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_30
timestamp 1486834041
transform 1 0 2016 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_32
timestamp 1486834041
transform 1 0 2128 0 -1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_43
timestamp 1486834041
transform 1 0 2744 0 -1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_59
timestamp 1486834041
transform 1 0 3640 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_67
timestamp 1486834041
transform 1 0 4088 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_69
timestamp 1486834041
transform 1 0 4200 0 -1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_72
timestamp 1486834041
transform 1 0 4368 0 -1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_88
timestamp 1486834041
transform 1 0 5264 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_96
timestamp 1486834041
transform 1 0 5712 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_100
timestamp 1486834041
transform 1 0 5936 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_112
timestamp 1486834041
transform 1 0 6608 0 -1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_128
timestamp 1486834041
transform 1 0 7504 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_136
timestamp 1486834041
transform 1 0 7952 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_142
timestamp 1486834041
transform 1 0 8288 0 -1 4312
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_206
timestamp 1486834041
transform 1 0 11872 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_212
timestamp 1486834041
transform 1 0 12208 0 -1 4312
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_276
timestamp 1486834041
transform 1 0 15792 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_282
timestamp 1486834041
transform 1 0 16128 0 -1 4312
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_346
timestamp 1486834041
transform 1 0 19712 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_352
timestamp 1486834041
transform 1 0 20048 0 -1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_368
timestamp 1486834041
transform 1 0 20944 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_376
timestamp 1486834041
transform 1 0 21392 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_390
timestamp 1486834041
transform 1 0 22176 0 -1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_406
timestamp 1486834041
transform 1 0 23072 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_414
timestamp 1486834041
transform 1 0 23520 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_418
timestamp 1486834041
transform 1 0 23744 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_422
timestamp 1486834041
transform 1 0 23968 0 -1 4312
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_486
timestamp 1486834041
transform 1 0 27552 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_500
timestamp 1486834041
transform 1 0 28336 0 -1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_2
timestamp 1486834041
transform 1 0 448 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_10
timestamp 1486834041
transform 1 0 896 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_14
timestamp 1486834041
transform 1 0 1120 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_16
timestamp 1486834041
transform 1 0 1232 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_27
timestamp 1486834041
transform 1 0 1848 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_31
timestamp 1486834041
transform 1 0 2072 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_45
timestamp 1486834041
transform 1 0 2856 0 1 4312
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_77
timestamp 1486834041
transform 1 0 4648 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_93
timestamp 1486834041
transform 1 0 5544 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_101
timestamp 1486834041
transform 1 0 5992 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_107
timestamp 1486834041
transform 1 0 6328 0 1 4312
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_139
timestamp 1486834041
transform 1 0 8120 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_143
timestamp 1486834041
transform 1 0 8344 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_155
timestamp 1486834041
transform 1 0 9016 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_171
timestamp 1486834041
transform 1 0 9912 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_177
timestamp 1486834041
transform 1 0 10248 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_181
timestamp 1486834041
transform 1 0 10472 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_183
timestamp 1486834041
transform 1 0 10584 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_194
timestamp 1486834041
transform 1 0 11200 0 1 4312
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_226
timestamp 1486834041
transform 1 0 12992 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_242
timestamp 1486834041
transform 1 0 13888 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_244
timestamp 1486834041
transform 1 0 14000 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_247
timestamp 1486834041
transform 1 0 14168 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_251
timestamp 1486834041
transform 1 0 14392 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_262
timestamp 1486834041
transform 1 0 15008 0 1 4312
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_294
timestamp 1486834041
transform 1 0 16800 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_310
timestamp 1486834041
transform 1 0 17696 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_314
timestamp 1486834041
transform 1 0 17920 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_317
timestamp 1486834041
transform 1 0 18088 0 1 4312
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_349
timestamp 1486834041
transform 1 0 19880 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_353
timestamp 1486834041
transform 1 0 20104 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_364
timestamp 1486834041
transform 1 0 20720 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_380
timestamp 1486834041
transform 1 0 21616 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_384
timestamp 1486834041
transform 1 0 21840 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_387
timestamp 1486834041
transform 1 0 22008 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_403
timestamp 1486834041
transform 1 0 22904 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_411
timestamp 1486834041
transform 1 0 23352 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_415
timestamp 1486834041
transform 1 0 23576 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_426
timestamp 1486834041
transform 1 0 24192 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_442
timestamp 1486834041
transform 1 0 25088 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_450
timestamp 1486834041
transform 1 0 25536 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_454
timestamp 1486834041
transform 1 0 25760 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_457
timestamp 1486834041
transform 1 0 25928 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_461
timestamp 1486834041
transform 1 0 26152 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_472
timestamp 1486834041
transform 1 0 26768 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_488
timestamp 1486834041
transform 1 0 27664 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_492
timestamp 1486834041
transform 1 0 27888 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_527
timestamp 1486834041
transform 1 0 29848 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_531
timestamp 1486834041
transform 1 0 30072 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_2
timestamp 1486834041
transform 1 0 448 0 -1 5096
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_34
timestamp 1486834041
transform 1 0 2240 0 -1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_50
timestamp 1486834041
transform 1 0 3136 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_58
timestamp 1486834041
transform 1 0 3584 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_72
timestamp 1486834041
transform 1 0 4368 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_80
timestamp 1486834041
transform 1 0 4816 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_84
timestamp 1486834041
transform 1 0 5040 0 -1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_99
timestamp 1486834041
transform 1 0 5880 0 -1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_115
timestamp 1486834041
transform 1 0 6776 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_131
timestamp 1486834041
transform 1 0 7672 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_139
timestamp 1486834041
transform 1 0 8120 0 -1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_142
timestamp 1486834041
transform 1 0 8288 0 -1 5096
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_206
timestamp 1486834041
transform 1 0 11872 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_212
timestamp 1486834041
transform 1 0 12208 0 -1 5096
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_276
timestamp 1486834041
transform 1 0 15792 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_282
timestamp 1486834041
transform 1 0 16128 0 -1 5096
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_346
timestamp 1486834041
transform 1 0 19712 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_352
timestamp 1486834041
transform 1 0 20048 0 -1 5096
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_416
timestamp 1486834041
transform 1 0 23632 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_422
timestamp 1486834041
transform 1 0 23968 0 -1 5096
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_486
timestamp 1486834041
transform 1 0 27552 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_500
timestamp 1486834041
transform 1 0 28336 0 -1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_2
timestamp 1486834041
transform 1 0 448 0 1 5096
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1486834041
transform 1 0 2240 0 1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_37
timestamp 1486834041
transform 1 0 2408 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_45
timestamp 1486834041
transform 1 0 2856 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_117
timestamp 1486834041
transform 1 0 6888 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_177
timestamp 1486834041
transform 1 0 10248 0 1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_188
timestamp 1486834041
transform 1 0 10864 0 1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_203
timestamp 1486834041
transform 1 0 11704 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_219
timestamp 1486834041
transform 1 0 12600 0 1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_235
timestamp 1486834041
transform 1 0 13496 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_243
timestamp 1486834041
transform 1 0 13944 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_247
timestamp 1486834041
transform 1 0 14168 0 1 5096
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_311
timestamp 1486834041
transform 1 0 17752 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_317
timestamp 1486834041
transform 1 0 18088 0 1 5096
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_349
timestamp 1486834041
transform 1 0 19880 0 1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_365
timestamp 1486834041
transform 1 0 20776 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_373
timestamp 1486834041
transform 1 0 21224 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_387
timestamp 1486834041
transform 1 0 22008 0 1 5096
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_451
timestamp 1486834041
transform 1 0 25592 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_457
timestamp 1486834041
transform 1 0 25928 0 1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_473
timestamp 1486834041
transform 1 0 26824 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_481
timestamp 1486834041
transform 1 0 27272 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_527
timestamp 1486834041
transform 1 0 29848 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_531
timestamp 1486834041
transform 1 0 30072 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_2
timestamp 1486834041
transform 1 0 448 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_6
timestamp 1486834041
transform 1 0 672 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_8
timestamp 1486834041
transform 1 0 784 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_19
timestamp 1486834041
transform 1 0 1400 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_27
timestamp 1486834041
transform 1 0 1848 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_72
timestamp 1486834041
transform 1 0 4368 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_80
timestamp 1486834041
transform 1 0 4816 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_142
timestamp 1486834041
transform 1 0 8288 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_150
timestamp 1486834041
transform 1 0 8736 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_212
timestamp 1486834041
transform 1 0 12208 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_220
timestamp 1486834041
transform 1 0 12656 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_224
timestamp 1486834041
transform 1 0 12880 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_239
timestamp 1486834041
transform 1 0 13720 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_251
timestamp 1486834041
transform 1 0 14392 0 -1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_267
timestamp 1486834041
transform 1 0 15288 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_275
timestamp 1486834041
transform 1 0 15736 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_279
timestamp 1486834041
transform 1 0 15960 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_282
timestamp 1486834041
transform 1 0 16128 0 -1 5880
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_346
timestamp 1486834041
transform 1 0 19712 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_352
timestamp 1486834041
transform 1 0 20048 0 -1 5880
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_384
timestamp 1486834041
transform 1 0 21840 0 -1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_400
timestamp 1486834041
transform 1 0 22736 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_404
timestamp 1486834041
transform 1 0 22960 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_415
timestamp 1486834041
transform 1 0 23576 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_419
timestamp 1486834041
transform 1 0 23800 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_422
timestamp 1486834041
transform 1 0 23968 0 -1 5880
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_454
timestamp 1486834041
transform 1 0 25760 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_458
timestamp 1486834041
transform 1 0 25984 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_460
timestamp 1486834041
transform 1 0 26096 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_489
timestamp 1486834041
transform 1 0 27720 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_558
timestamp 1486834041
transform 1 0 31584 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_2
timestamp 1486834041
transform 1 0 448 0 1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_18
timestamp 1486834041
transform 1 0 1344 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_20
timestamp 1486834041
transform 1 0 1456 0 1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_37
timestamp 1486834041
transform 1 0 2408 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_45
timestamp 1486834041
transform 1 0 2856 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_107
timestamp 1486834041
transform 1 0 6328 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_115
timestamp 1486834041
transform 1 0 6776 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_177
timestamp 1486834041
transform 1 0 10248 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_185
timestamp 1486834041
transform 1 0 10696 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_243
timestamp 1486834041
transform 1 0 13944 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_247
timestamp 1486834041
transform 1 0 14168 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_251
timestamp 1486834041
transform 1 0 14392 0 1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_262
timestamp 1486834041
transform 1 0 15008 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_274
timestamp 1486834041
transform 1 0 15680 0 1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_290
timestamp 1486834041
transform 1 0 16576 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_298
timestamp 1486834041
transform 1 0 17024 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_302
timestamp 1486834041
transform 1 0 17248 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_304
timestamp 1486834041
transform 1 0 17360 0 1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_317
timestamp 1486834041
transform 1 0 18088 0 1 5880
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_349
timestamp 1486834041
transform 1 0 19880 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_353
timestamp 1486834041
transform 1 0 20104 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_365
timestamp 1486834041
transform 1 0 20776 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_373
timestamp 1486834041
transform 1 0 21224 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_387
timestamp 1486834041
transform 1 0 22008 0 1 5880
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_451
timestamp 1486834041
transform 1 0 25592 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_513
timestamp 1486834041
transform 1 0 29064 0 1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_524
timestamp 1486834041
transform 1 0 29680 0 1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_555
timestamp 1486834041
transform 1 0 31416 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_559
timestamp 1486834041
transform 1 0 31640 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_2
timestamp 1486834041
transform 1 0 448 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_36
timestamp 1486834041
transform 1 0 2352 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_70
timestamp 1486834041
transform 1 0 4256 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_104
timestamp 1486834041
transform 1 0 6160 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_138
timestamp 1486834041
transform 1 0 8064 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_172
timestamp 1486834041
transform 1 0 9968 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_206
timestamp 1486834041
transform 1 0 11872 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_254
timestamp 1486834041
transform 1 0 14560 0 -1 6664
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_270
timestamp 1486834041
transform 1 0 15456 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_274
timestamp 1486834041
transform 1 0 15680 0 -1 6664
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_308
timestamp 1486834041
transform 1 0 17584 0 -1 6664
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_342
timestamp 1486834041
transform 1 0 19488 0 -1 6664
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_376
timestamp 1486834041
transform 1 0 21392 0 -1 6664
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_410
timestamp 1486834041
transform 1 0 23296 0 -1 6664
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_444
timestamp 1486834041
transform 1 0 25200 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_446
timestamp 1486834041
transform 1 0 25312 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_467
timestamp 1486834041
transform 1 0 26488 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_475
timestamp 1486834041
transform 1 0 26936 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_506
timestamp 1486834041
transform 1 0 28672 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_540
timestamp 1486834041
transform 1 0 30576 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_560
timestamp 1486834041
transform 1 0 31696 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output1
timestamp 1486834041
transform 1 0 30184 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output2
timestamp 1486834041
transform 1 0 30072 0 -1 2744
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output3
timestamp 1486834041
transform 1 0 30968 0 1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output4
timestamp 1486834041
transform 1 0 30856 0 -1 2744
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output5
timestamp 1486834041
transform 1 0 30072 0 -1 3528
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output6
timestamp 1486834041
transform 1 0 30968 0 1 2744
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output7
timestamp 1486834041
transform 1 0 30184 0 1 3528
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output8
timestamp 1486834041
transform 1 0 30856 0 -1 3528
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output9
timestamp 1486834041
transform 1 0 30856 0 -1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output10
timestamp 1486834041
transform 1 0 30968 0 1 3528
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output11
timestamp 1486834041
transform 1 0 30968 0 1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output12
timestamp 1486834041
transform 1 0 29232 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output13
timestamp 1486834041
transform 1 0 30856 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output14
timestamp 1486834041
transform 1 0 30968 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output15
timestamp 1486834041
transform 1 0 30184 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output16
timestamp 1486834041
transform 1 0 30072 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output17
timestamp 1486834041
transform 1 0 30184 0 1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output18
timestamp 1486834041
transform 1 0 29288 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output19
timestamp 1486834041
transform 1 0 30072 0 -1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output20
timestamp 1486834041
transform -1 0 29736 0 1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output21
timestamp 1486834041
transform 1 0 29288 0 -1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output22
timestamp 1486834041
transform 1 0 28504 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output23
timestamp 1486834041
transform 1 0 30016 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output24
timestamp 1486834041
transform 1 0 30184 0 1 2744
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output25
timestamp 1486834041
transform -1 0 28168 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output26
timestamp 1486834041
transform 1 0 30072 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output27
timestamp 1486834041
transform 1 0 30968 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output28
timestamp 1486834041
transform 1 0 30856 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output29
timestamp 1486834041
transform 1 0 30072 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output30
timestamp 1486834041
transform 1 0 30968 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output31
timestamp 1486834041
transform 1 0 30184 0 1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output32
timestamp 1486834041
transform 1 0 30856 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output33
timestamp 1486834041
transform 1 0 25704 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output34
timestamp 1486834041
transform 1 0 29008 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output35
timestamp 1486834041
transform 1 0 28168 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output36
timestamp 1486834041
transform 1 0 28672 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output37
timestamp 1486834041
transform 1 0 29792 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output38
timestamp 1486834041
transform 1 0 28952 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output39
timestamp 1486834041
transform 1 0 29848 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output40
timestamp 1486834041
transform 1 0 29456 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output41
timestamp 1486834041
transform 1 0 30912 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output42
timestamp 1486834041
transform 1 0 30632 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output43
timestamp 1486834041
transform 1 0 30240 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output44
timestamp 1486834041
transform 1 0 25928 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output45
timestamp 1486834041
transform 1 0 26152 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output46
timestamp 1486834041
transform 1 0 26712 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output47
timestamp 1486834041
transform 1 0 27104 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output48
timestamp 1486834041
transform 1 0 26936 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output49
timestamp 1486834041
transform 1 0 27496 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output50
timestamp 1486834041
transform 1 0 27888 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output51
timestamp 1486834041
transform 1 0 28280 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output52
timestamp 1486834041
transform 1 0 27888 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output53
timestamp 1486834041
transform 1 0 672 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output54
timestamp 1486834041
transform -1 0 2296 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output55
timestamp 1486834041
transform -1 0 2688 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output56
timestamp 1486834041
transform -1 0 2240 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output57
timestamp 1486834041
transform -1 0 3472 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output58
timestamp 1486834041
transform -1 0 3864 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output59
timestamp 1486834041
transform -1 0 3360 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output60
timestamp 1486834041
transform -1 0 3864 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output61
timestamp 1486834041
transform -1 0 4648 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output62
timestamp 1486834041
transform -1 0 4256 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output63
timestamp 1486834041
transform -1 0 4144 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output64
timestamp 1486834041
transform -1 0 5432 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output65
timestamp 1486834041
transform -1 0 4648 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output66
timestamp 1486834041
transform -1 0 5880 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output67
timestamp 1486834041
transform -1 0 5432 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output68
timestamp 1486834041
transform -1 0 6216 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output69
timestamp 1486834041
transform -1 0 5824 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output70
timestamp 1486834041
transform -1 0 5264 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output71
timestamp 1486834041
transform -1 0 6608 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output72
timestamp 1486834041
transform -1 0 6216 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output73
timestamp 1486834041
transform -1 0 6048 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output74
timestamp 1486834041
transform 1 0 8568 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output75
timestamp 1486834041
transform 1 0 8960 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output76
timestamp 1486834041
transform -1 0 10136 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output77
timestamp 1486834041
transform -1 0 9352 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output78
timestamp 1486834041
transform -1 0 9072 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output79
timestamp 1486834041
transform 1 0 9352 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output80
timestamp 1486834041
transform -1 0 7672 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output81
timestamp 1486834041
transform -1 0 7784 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output82
timestamp 1486834041
transform 1 0 6608 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output83
timestamp 1486834041
transform 1 0 6384 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output84
timestamp 1486834041
transform 1 0 7784 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output85
timestamp 1486834041
transform 1 0 7000 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output86
timestamp 1486834041
transform 1 0 7392 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output87
timestamp 1486834041
transform -1 0 7952 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output88
timestamp 1486834041
transform -1 0 8568 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output89
timestamp 1486834041
transform -1 0 10528 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output90
timestamp 1486834041
transform -1 0 13160 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output91
timestamp 1486834041
transform -1 0 12880 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output92
timestamp 1486834041
transform -1 0 13720 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output93
timestamp 1486834041
transform -1 0 13944 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output94
timestamp 1486834041
transform -1 0 13664 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output95
timestamp 1486834041
transform -1 0 14560 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output96
timestamp 1486834041
transform -1 0 9856 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output97
timestamp 1486834041
transform -1 0 11312 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output98
timestamp 1486834041
transform -1 0 11704 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output99
timestamp 1486834041
transform -1 0 10976 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output100
timestamp 1486834041
transform -1 0 11592 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output101
timestamp 1486834041
transform -1 0 12096 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output102
timestamp 1486834041
transform -1 0 12600 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output103
timestamp 1486834041
transform -1 0 11760 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output104
timestamp 1486834041
transform -1 0 12376 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output105
timestamp 1486834041
transform -1 0 25704 0 -1 6664
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_16
timestamp 1486834041
transform 1 0 336 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1486834041
transform -1 0 31864 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_17
timestamp 1486834041
transform 1 0 336 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1486834041
transform -1 0 31864 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_18
timestamp 1486834041
transform 1 0 336 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1486834041
transform -1 0 31864 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_19
timestamp 1486834041
transform 1 0 336 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1486834041
transform -1 0 31864 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_20
timestamp 1486834041
transform 1 0 336 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1486834041
transform -1 0 31864 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_21
timestamp 1486834041
transform 1 0 336 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1486834041
transform -1 0 31864 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_22
timestamp 1486834041
transform 1 0 336 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1486834041
transform -1 0 31864 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_23
timestamp 1486834041
transform 1 0 336 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1486834041
transform -1 0 31864 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_24
timestamp 1486834041
transform 1 0 336 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1486834041
transform -1 0 31864 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_25
timestamp 1486834041
transform 1 0 336 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1486834041
transform -1 0 31864 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_26
timestamp 1486834041
transform 1 0 336 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1486834041
transform -1 0 31864 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_27
timestamp 1486834041
transform 1 0 336 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1486834041
transform -1 0 31864 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_28
timestamp 1486834041
transform 1 0 336 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1486834041
transform -1 0 31864 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_29
timestamp 1486834041
transform 1 0 336 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1486834041
transform -1 0 31864 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_30
timestamp 1486834041
transform 1 0 336 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1486834041
transform -1 0 31864 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_31
timestamp 1486834041
transform 1 0 336 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1486834041
transform -1 0 31864 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_32
timestamp 1486834041
transform 1 0 2240 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_33
timestamp 1486834041
transform 1 0 4144 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_34
timestamp 1486834041
transform 1 0 6048 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_35
timestamp 1486834041
transform 1 0 7952 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_36
timestamp 1486834041
transform 1 0 9856 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_37
timestamp 1486834041
transform 1 0 11760 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_38
timestamp 1486834041
transform 1 0 13664 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_39
timestamp 1486834041
transform 1 0 15568 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_40
timestamp 1486834041
transform 1 0 17472 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_41
timestamp 1486834041
transform 1 0 19376 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_42
timestamp 1486834041
transform 1 0 21280 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_43
timestamp 1486834041
transform 1 0 23184 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_44
timestamp 1486834041
transform 1 0 25088 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_45
timestamp 1486834041
transform 1 0 26992 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_46
timestamp 1486834041
transform 1 0 28896 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_47
timestamp 1486834041
transform 1 0 30800 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_48
timestamp 1486834041
transform 1 0 4256 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_49
timestamp 1486834041
transform 1 0 8176 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_50
timestamp 1486834041
transform 1 0 12096 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_51
timestamp 1486834041
transform 1 0 16016 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_52
timestamp 1486834041
transform 1 0 19936 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_53
timestamp 1486834041
transform 1 0 23856 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_54
timestamp 1486834041
transform 1 0 27776 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_55
timestamp 1486834041
transform 1 0 31640 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_56
timestamp 1486834041
transform 1 0 2296 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_57
timestamp 1486834041
transform 1 0 6216 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_58
timestamp 1486834041
transform 1 0 10136 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_59
timestamp 1486834041
transform 1 0 14056 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_60
timestamp 1486834041
transform 1 0 17976 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_61
timestamp 1486834041
transform 1 0 21896 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_62
timestamp 1486834041
transform 1 0 25816 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_63
timestamp 1486834041
transform 1 0 29736 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_64
timestamp 1486834041
transform 1 0 4256 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_65
timestamp 1486834041
transform 1 0 8176 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_66
timestamp 1486834041
transform 1 0 12096 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_67
timestamp 1486834041
transform 1 0 16016 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_68
timestamp 1486834041
transform 1 0 19936 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_69
timestamp 1486834041
transform 1 0 23856 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_70
timestamp 1486834041
transform 1 0 27776 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_71
timestamp 1486834041
transform 1 0 31640 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_72
timestamp 1486834041
transform 1 0 2296 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_73
timestamp 1486834041
transform 1 0 6216 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_74
timestamp 1486834041
transform 1 0 10136 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_75
timestamp 1486834041
transform 1 0 14056 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_76
timestamp 1486834041
transform 1 0 17976 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_77
timestamp 1486834041
transform 1 0 21896 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_78
timestamp 1486834041
transform 1 0 25816 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_79
timestamp 1486834041
transform 1 0 29736 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_80
timestamp 1486834041
transform 1 0 4256 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_81
timestamp 1486834041
transform 1 0 8176 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_82
timestamp 1486834041
transform 1 0 12096 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_83
timestamp 1486834041
transform 1 0 16016 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_84
timestamp 1486834041
transform 1 0 19936 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_85
timestamp 1486834041
transform 1 0 23856 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_86
timestamp 1486834041
transform 1 0 27776 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_87
timestamp 1486834041
transform 1 0 31640 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_88
timestamp 1486834041
transform 1 0 2296 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_89
timestamp 1486834041
transform 1 0 6216 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_90
timestamp 1486834041
transform 1 0 10136 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_91
timestamp 1486834041
transform 1 0 14056 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_92
timestamp 1486834041
transform 1 0 17976 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_93
timestamp 1486834041
transform 1 0 21896 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_94
timestamp 1486834041
transform 1 0 25816 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_95
timestamp 1486834041
transform 1 0 29736 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_96
timestamp 1486834041
transform 1 0 4256 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_97
timestamp 1486834041
transform 1 0 8176 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_98
timestamp 1486834041
transform 1 0 12096 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_99
timestamp 1486834041
transform 1 0 16016 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_100
timestamp 1486834041
transform 1 0 19936 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_101
timestamp 1486834041
transform 1 0 23856 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_102
timestamp 1486834041
transform 1 0 27776 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_103
timestamp 1486834041
transform 1 0 31640 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_104
timestamp 1486834041
transform 1 0 2296 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_105
timestamp 1486834041
transform 1 0 6216 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_106
timestamp 1486834041
transform 1 0 10136 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_107
timestamp 1486834041
transform 1 0 14056 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_108
timestamp 1486834041
transform 1 0 17976 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_109
timestamp 1486834041
transform 1 0 21896 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_110
timestamp 1486834041
transform 1 0 25816 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_111
timestamp 1486834041
transform 1 0 29736 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_112
timestamp 1486834041
transform 1 0 4256 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_113
timestamp 1486834041
transform 1 0 8176 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_114
timestamp 1486834041
transform 1 0 12096 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_115
timestamp 1486834041
transform 1 0 16016 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_116
timestamp 1486834041
transform 1 0 19936 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_117
timestamp 1486834041
transform 1 0 23856 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_118
timestamp 1486834041
transform 1 0 27776 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_119
timestamp 1486834041
transform 1 0 31640 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_120
timestamp 1486834041
transform 1 0 2296 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_121
timestamp 1486834041
transform 1 0 6216 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_122
timestamp 1486834041
transform 1 0 10136 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_123
timestamp 1486834041
transform 1 0 14056 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_124
timestamp 1486834041
transform 1 0 17976 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_125
timestamp 1486834041
transform 1 0 21896 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_126
timestamp 1486834041
transform 1 0 25816 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_127
timestamp 1486834041
transform 1 0 29736 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_128
timestamp 1486834041
transform 1 0 4256 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_129
timestamp 1486834041
transform 1 0 8176 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_130
timestamp 1486834041
transform 1 0 12096 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_131
timestamp 1486834041
transform 1 0 16016 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_132
timestamp 1486834041
transform 1 0 19936 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_133
timestamp 1486834041
transform 1 0 23856 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_134
timestamp 1486834041
transform 1 0 27776 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_135
timestamp 1486834041
transform 1 0 31640 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_136
timestamp 1486834041
transform 1 0 2296 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_137
timestamp 1486834041
transform 1 0 6216 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_138
timestamp 1486834041
transform 1 0 10136 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_139
timestamp 1486834041
transform 1 0 14056 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_140
timestamp 1486834041
transform 1 0 17976 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_141
timestamp 1486834041
transform 1 0 21896 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_142
timestamp 1486834041
transform 1 0 25816 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_143
timestamp 1486834041
transform 1 0 29736 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_144
timestamp 1486834041
transform 1 0 4256 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_145
timestamp 1486834041
transform 1 0 8176 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_146
timestamp 1486834041
transform 1 0 12096 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_147
timestamp 1486834041
transform 1 0 16016 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_148
timestamp 1486834041
transform 1 0 19936 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_149
timestamp 1486834041
transform 1 0 23856 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_150
timestamp 1486834041
transform 1 0 27776 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_151
timestamp 1486834041
transform 1 0 31640 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_152
timestamp 1486834041
transform 1 0 2296 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_153
timestamp 1486834041
transform 1 0 6216 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_154
timestamp 1486834041
transform 1 0 10136 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_155
timestamp 1486834041
transform 1 0 14056 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_156
timestamp 1486834041
transform 1 0 17976 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_157
timestamp 1486834041
transform 1 0 21896 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1486834041
transform 1 0 25816 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1486834041
transform 1 0 29736 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_160
timestamp 1486834041
transform 1 0 2240 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_161
timestamp 1486834041
transform 1 0 4144 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_162
timestamp 1486834041
transform 1 0 6048 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1486834041
transform 1 0 7952 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1486834041
transform 1 0 9856 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1486834041
transform 1 0 11760 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1486834041
transform 1 0 13664 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_167
timestamp 1486834041
transform 1 0 15568 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_168
timestamp 1486834041
transform 1 0 17472 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_169
timestamp 1486834041
transform 1 0 19376 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_170
timestamp 1486834041
transform 1 0 21280 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_171
timestamp 1486834041
transform 1 0 23184 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_172
timestamp 1486834041
transform 1 0 25088 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_173
timestamp 1486834041
transform 1 0 26992 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_174
timestamp 1486834041
transform 1 0 28896 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_175
timestamp 1486834041
transform 1 0 30800 0 -1 6664
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 0 56 56 0 FreeSans 224 0 0 0 FrameData[0]
port 0 nsew signal input
flabel metal3 s 0 2240 56 2296 0 FreeSans 224 0 0 0 FrameData[10]
port 1 nsew signal input
flabel metal3 s 0 2464 56 2520 0 FreeSans 224 0 0 0 FrameData[11]
port 2 nsew signal input
flabel metal3 s 0 2688 56 2744 0 FreeSans 224 0 0 0 FrameData[12]
port 3 nsew signal input
flabel metal3 s 0 2912 56 2968 0 FreeSans 224 0 0 0 FrameData[13]
port 4 nsew signal input
flabel metal3 s 0 3136 56 3192 0 FreeSans 224 0 0 0 FrameData[14]
port 5 nsew signal input
flabel metal3 s 0 3360 56 3416 0 FreeSans 224 0 0 0 FrameData[15]
port 6 nsew signal input
flabel metal3 s 0 3584 56 3640 0 FreeSans 224 0 0 0 FrameData[16]
port 7 nsew signal input
flabel metal3 s 0 3808 56 3864 0 FreeSans 224 0 0 0 FrameData[17]
port 8 nsew signal input
flabel metal3 s 0 4032 56 4088 0 FreeSans 224 0 0 0 FrameData[18]
port 9 nsew signal input
flabel metal3 s 0 4256 56 4312 0 FreeSans 224 0 0 0 FrameData[19]
port 10 nsew signal input
flabel metal3 s 0 224 56 280 0 FreeSans 224 0 0 0 FrameData[1]
port 11 nsew signal input
flabel metal3 s 0 4480 56 4536 0 FreeSans 224 0 0 0 FrameData[20]
port 12 nsew signal input
flabel metal3 s 0 4704 56 4760 0 FreeSans 224 0 0 0 FrameData[21]
port 13 nsew signal input
flabel metal3 s 0 4928 56 4984 0 FreeSans 224 0 0 0 FrameData[22]
port 14 nsew signal input
flabel metal3 s 0 5152 56 5208 0 FreeSans 224 0 0 0 FrameData[23]
port 15 nsew signal input
flabel metal3 s 0 5376 56 5432 0 FreeSans 224 0 0 0 FrameData[24]
port 16 nsew signal input
flabel metal3 s 0 5600 56 5656 0 FreeSans 224 0 0 0 FrameData[25]
port 17 nsew signal input
flabel metal3 s 0 5824 56 5880 0 FreeSans 224 0 0 0 FrameData[26]
port 18 nsew signal input
flabel metal3 s 0 6048 56 6104 0 FreeSans 224 0 0 0 FrameData[27]
port 19 nsew signal input
flabel metal3 s 0 6272 56 6328 0 FreeSans 224 0 0 0 FrameData[28]
port 20 nsew signal input
flabel metal3 s 0 6496 56 6552 0 FreeSans 224 0 0 0 FrameData[29]
port 21 nsew signal input
flabel metal3 s 0 448 56 504 0 FreeSans 224 0 0 0 FrameData[2]
port 22 nsew signal input
flabel metal3 s 0 6720 56 6776 0 FreeSans 224 0 0 0 FrameData[30]
port 23 nsew signal input
flabel metal3 s 0 6944 56 7000 0 FreeSans 224 0 0 0 FrameData[31]
port 24 nsew signal input
flabel metal3 s 0 672 56 728 0 FreeSans 224 0 0 0 FrameData[3]
port 25 nsew signal input
flabel metal3 s 0 896 56 952 0 FreeSans 224 0 0 0 FrameData[4]
port 26 nsew signal input
flabel metal3 s 0 1120 56 1176 0 FreeSans 224 0 0 0 FrameData[5]
port 27 nsew signal input
flabel metal3 s 0 1344 56 1400 0 FreeSans 224 0 0 0 FrameData[6]
port 28 nsew signal input
flabel metal3 s 0 1568 56 1624 0 FreeSans 224 0 0 0 FrameData[7]
port 29 nsew signal input
flabel metal3 s 0 1792 56 1848 0 FreeSans 224 0 0 0 FrameData[8]
port 30 nsew signal input
flabel metal3 s 0 2016 56 2072 0 FreeSans 224 0 0 0 FrameData[9]
port 31 nsew signal input
flabel metal3 s 32144 0 32200 56 0 FreeSans 224 0 0 0 FrameData_O[0]
port 32 nsew signal output
flabel metal3 s 32144 2240 32200 2296 0 FreeSans 224 0 0 0 FrameData_O[10]
port 33 nsew signal output
flabel metal3 s 32144 2464 32200 2520 0 FreeSans 224 0 0 0 FrameData_O[11]
port 34 nsew signal output
flabel metal3 s 32144 2688 32200 2744 0 FreeSans 224 0 0 0 FrameData_O[12]
port 35 nsew signal output
flabel metal3 s 32144 2912 32200 2968 0 FreeSans 224 0 0 0 FrameData_O[13]
port 36 nsew signal output
flabel metal3 s 32144 3136 32200 3192 0 FreeSans 224 0 0 0 FrameData_O[14]
port 37 nsew signal output
flabel metal3 s 32144 3360 32200 3416 0 FreeSans 224 0 0 0 FrameData_O[15]
port 38 nsew signal output
flabel metal3 s 32144 3584 32200 3640 0 FreeSans 224 0 0 0 FrameData_O[16]
port 39 nsew signal output
flabel metal3 s 32144 3808 32200 3864 0 FreeSans 224 0 0 0 FrameData_O[17]
port 40 nsew signal output
flabel metal3 s 32144 4032 32200 4088 0 FreeSans 224 0 0 0 FrameData_O[18]
port 41 nsew signal output
flabel metal3 s 32144 4256 32200 4312 0 FreeSans 224 0 0 0 FrameData_O[19]
port 42 nsew signal output
flabel metal3 s 32144 224 32200 280 0 FreeSans 224 0 0 0 FrameData_O[1]
port 43 nsew signal output
flabel metal3 s 32144 4480 32200 4536 0 FreeSans 224 0 0 0 FrameData_O[20]
port 44 nsew signal output
flabel metal3 s 32144 4704 32200 4760 0 FreeSans 224 0 0 0 FrameData_O[21]
port 45 nsew signal output
flabel metal3 s 32144 4928 32200 4984 0 FreeSans 224 0 0 0 FrameData_O[22]
port 46 nsew signal output
flabel metal3 s 32144 5152 32200 5208 0 FreeSans 224 0 0 0 FrameData_O[23]
port 47 nsew signal output
flabel metal3 s 32144 5376 32200 5432 0 FreeSans 224 0 0 0 FrameData_O[24]
port 48 nsew signal output
flabel metal3 s 32144 5600 32200 5656 0 FreeSans 224 0 0 0 FrameData_O[25]
port 49 nsew signal output
flabel metal3 s 32144 5824 32200 5880 0 FreeSans 224 0 0 0 FrameData_O[26]
port 50 nsew signal output
flabel metal3 s 32144 6048 32200 6104 0 FreeSans 224 0 0 0 FrameData_O[27]
port 51 nsew signal output
flabel metal3 s 32144 6272 32200 6328 0 FreeSans 224 0 0 0 FrameData_O[28]
port 52 nsew signal output
flabel metal3 s 32144 6496 32200 6552 0 FreeSans 224 0 0 0 FrameData_O[29]
port 53 nsew signal output
flabel metal3 s 32144 448 32200 504 0 FreeSans 224 0 0 0 FrameData_O[2]
port 54 nsew signal output
flabel metal3 s 32144 6720 32200 6776 0 FreeSans 224 0 0 0 FrameData_O[30]
port 55 nsew signal output
flabel metal3 s 32144 6944 32200 7000 0 FreeSans 224 0 0 0 FrameData_O[31]
port 56 nsew signal output
flabel metal3 s 32144 672 32200 728 0 FreeSans 224 0 0 0 FrameData_O[3]
port 57 nsew signal output
flabel metal3 s 32144 896 32200 952 0 FreeSans 224 0 0 0 FrameData_O[4]
port 58 nsew signal output
flabel metal3 s 32144 1120 32200 1176 0 FreeSans 224 0 0 0 FrameData_O[5]
port 59 nsew signal output
flabel metal3 s 32144 1344 32200 1400 0 FreeSans 224 0 0 0 FrameData_O[6]
port 60 nsew signal output
flabel metal3 s 32144 1568 32200 1624 0 FreeSans 224 0 0 0 FrameData_O[7]
port 61 nsew signal output
flabel metal3 s 32144 1792 32200 1848 0 FreeSans 224 0 0 0 FrameData_O[8]
port 62 nsew signal output
flabel metal3 s 32144 2016 32200 2072 0 FreeSans 224 0 0 0 FrameData_O[9]
port 63 nsew signal output
flabel metal2 s 2912 0 2968 56 0 FreeSans 224 0 0 0 FrameStrobe[0]
port 64 nsew signal input
flabel metal2 s 17472 0 17528 56 0 FreeSans 224 0 0 0 FrameStrobe[10]
port 65 nsew signal input
flabel metal2 s 18928 0 18984 56 0 FreeSans 224 0 0 0 FrameStrobe[11]
port 66 nsew signal input
flabel metal2 s 20384 0 20440 56 0 FreeSans 224 0 0 0 FrameStrobe[12]
port 67 nsew signal input
flabel metal2 s 21840 0 21896 56 0 FreeSans 224 0 0 0 FrameStrobe[13]
port 68 nsew signal input
flabel metal2 s 23296 0 23352 56 0 FreeSans 224 0 0 0 FrameStrobe[14]
port 69 nsew signal input
flabel metal2 s 24752 0 24808 56 0 FreeSans 224 0 0 0 FrameStrobe[15]
port 70 nsew signal input
flabel metal2 s 26208 0 26264 56 0 FreeSans 224 0 0 0 FrameStrobe[16]
port 71 nsew signal input
flabel metal2 s 27664 0 27720 56 0 FreeSans 224 0 0 0 FrameStrobe[17]
port 72 nsew signal input
flabel metal2 s 29120 0 29176 56 0 FreeSans 224 0 0 0 FrameStrobe[18]
port 73 nsew signal input
flabel metal2 s 30576 0 30632 56 0 FreeSans 224 0 0 0 FrameStrobe[19]
port 74 nsew signal input
flabel metal2 s 4368 0 4424 56 0 FreeSans 224 0 0 0 FrameStrobe[1]
port 75 nsew signal input
flabel metal2 s 5824 0 5880 56 0 FreeSans 224 0 0 0 FrameStrobe[2]
port 76 nsew signal input
flabel metal2 s 7280 0 7336 56 0 FreeSans 224 0 0 0 FrameStrobe[3]
port 77 nsew signal input
flabel metal2 s 8736 0 8792 56 0 FreeSans 224 0 0 0 FrameStrobe[4]
port 78 nsew signal input
flabel metal2 s 10192 0 10248 56 0 FreeSans 224 0 0 0 FrameStrobe[5]
port 79 nsew signal input
flabel metal2 s 11648 0 11704 56 0 FreeSans 224 0 0 0 FrameStrobe[6]
port 80 nsew signal input
flabel metal2 s 13104 0 13160 56 0 FreeSans 224 0 0 0 FrameStrobe[7]
port 81 nsew signal input
flabel metal2 s 14560 0 14616 56 0 FreeSans 224 0 0 0 FrameStrobe[8]
port 82 nsew signal input
flabel metal2 s 16016 0 16072 56 0 FreeSans 224 0 0 0 FrameStrobe[9]
port 83 nsew signal input
flabel metal2 s 25648 7056 25704 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[0]
port 84 nsew signal output
flabel metal2 s 27888 7056 27944 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[10]
port 85 nsew signal output
flabel metal2 s 28112 7056 28168 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[11]
port 86 nsew signal output
flabel metal2 s 28336 7056 28392 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[12]
port 87 nsew signal output
flabel metal2 s 28560 7056 28616 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[13]
port 88 nsew signal output
flabel metal2 s 28784 7056 28840 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[14]
port 89 nsew signal output
flabel metal2 s 29008 7056 29064 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[15]
port 90 nsew signal output
flabel metal2 s 29232 7056 29288 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[16]
port 91 nsew signal output
flabel metal2 s 29456 7056 29512 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[17]
port 92 nsew signal output
flabel metal2 s 29680 7056 29736 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[18]
port 93 nsew signal output
flabel metal2 s 29904 7056 29960 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[19]
port 94 nsew signal output
flabel metal2 s 25872 7056 25928 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[1]
port 95 nsew signal output
flabel metal2 s 26096 7056 26152 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[2]
port 96 nsew signal output
flabel metal2 s 26320 7056 26376 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[3]
port 97 nsew signal output
flabel metal2 s 26544 7056 26600 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[4]
port 98 nsew signal output
flabel metal2 s 26768 7056 26824 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[5]
port 99 nsew signal output
flabel metal2 s 26992 7056 27048 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[6]
port 100 nsew signal output
flabel metal2 s 27216 7056 27272 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[7]
port 101 nsew signal output
flabel metal2 s 27440 7056 27496 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[8]
port 102 nsew signal output
flabel metal2 s 27664 7056 27720 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[9]
port 103 nsew signal output
flabel metal2 s 2128 7056 2184 7112 0 FreeSans 224 0 0 0 N1BEG[0]
port 104 nsew signal output
flabel metal2 s 2352 7056 2408 7112 0 FreeSans 224 0 0 0 N1BEG[1]
port 105 nsew signal output
flabel metal2 s 2576 7056 2632 7112 0 FreeSans 224 0 0 0 N1BEG[2]
port 106 nsew signal output
flabel metal2 s 2800 7056 2856 7112 0 FreeSans 224 0 0 0 N1BEG[3]
port 107 nsew signal output
flabel metal2 s 3024 7056 3080 7112 0 FreeSans 224 0 0 0 N2BEG[0]
port 108 nsew signal output
flabel metal2 s 3248 7056 3304 7112 0 FreeSans 224 0 0 0 N2BEG[1]
port 109 nsew signal output
flabel metal2 s 3472 7056 3528 7112 0 FreeSans 224 0 0 0 N2BEG[2]
port 110 nsew signal output
flabel metal2 s 3696 7056 3752 7112 0 FreeSans 224 0 0 0 N2BEG[3]
port 111 nsew signal output
flabel metal2 s 3920 7056 3976 7112 0 FreeSans 224 0 0 0 N2BEG[4]
port 112 nsew signal output
flabel metal2 s 4144 7056 4200 7112 0 FreeSans 224 0 0 0 N2BEG[5]
port 113 nsew signal output
flabel metal2 s 4368 7056 4424 7112 0 FreeSans 224 0 0 0 N2BEG[6]
port 114 nsew signal output
flabel metal2 s 4592 7056 4648 7112 0 FreeSans 224 0 0 0 N2BEG[7]
port 115 nsew signal output
flabel metal2 s 4816 7056 4872 7112 0 FreeSans 224 0 0 0 N2BEGb[0]
port 116 nsew signal output
flabel metal2 s 5040 7056 5096 7112 0 FreeSans 224 0 0 0 N2BEGb[1]
port 117 nsew signal output
flabel metal2 s 5264 7056 5320 7112 0 FreeSans 224 0 0 0 N2BEGb[2]
port 118 nsew signal output
flabel metal2 s 5488 7056 5544 7112 0 FreeSans 224 0 0 0 N2BEGb[3]
port 119 nsew signal output
flabel metal2 s 5712 7056 5768 7112 0 FreeSans 224 0 0 0 N2BEGb[4]
port 120 nsew signal output
flabel metal2 s 5936 7056 5992 7112 0 FreeSans 224 0 0 0 N2BEGb[5]
port 121 nsew signal output
flabel metal2 s 6160 7056 6216 7112 0 FreeSans 224 0 0 0 N2BEGb[6]
port 122 nsew signal output
flabel metal2 s 6384 7056 6440 7112 0 FreeSans 224 0 0 0 N2BEGb[7]
port 123 nsew signal output
flabel metal2 s 6608 7056 6664 7112 0 FreeSans 224 0 0 0 N4BEG[0]
port 124 nsew signal output
flabel metal2 s 8848 7056 8904 7112 0 FreeSans 224 0 0 0 N4BEG[10]
port 125 nsew signal output
flabel metal2 s 9072 7056 9128 7112 0 FreeSans 224 0 0 0 N4BEG[11]
port 126 nsew signal output
flabel metal2 s 9296 7056 9352 7112 0 FreeSans 224 0 0 0 N4BEG[12]
port 127 nsew signal output
flabel metal2 s 9520 7056 9576 7112 0 FreeSans 224 0 0 0 N4BEG[13]
port 128 nsew signal output
flabel metal2 s 9744 7056 9800 7112 0 FreeSans 224 0 0 0 N4BEG[14]
port 129 nsew signal output
flabel metal2 s 9968 7056 10024 7112 0 FreeSans 224 0 0 0 N4BEG[15]
port 130 nsew signal output
flabel metal2 s 6832 7056 6888 7112 0 FreeSans 224 0 0 0 N4BEG[1]
port 131 nsew signal output
flabel metal2 s 7056 7056 7112 7112 0 FreeSans 224 0 0 0 N4BEG[2]
port 132 nsew signal output
flabel metal2 s 7280 7056 7336 7112 0 FreeSans 224 0 0 0 N4BEG[3]
port 133 nsew signal output
flabel metal2 s 7504 7056 7560 7112 0 FreeSans 224 0 0 0 N4BEG[4]
port 134 nsew signal output
flabel metal2 s 7728 7056 7784 7112 0 FreeSans 224 0 0 0 N4BEG[5]
port 135 nsew signal output
flabel metal2 s 7952 7056 8008 7112 0 FreeSans 224 0 0 0 N4BEG[6]
port 136 nsew signal output
flabel metal2 s 8176 7056 8232 7112 0 FreeSans 224 0 0 0 N4BEG[7]
port 137 nsew signal output
flabel metal2 s 8400 7056 8456 7112 0 FreeSans 224 0 0 0 N4BEG[8]
port 138 nsew signal output
flabel metal2 s 8624 7056 8680 7112 0 FreeSans 224 0 0 0 N4BEG[9]
port 139 nsew signal output
flabel metal2 s 10192 7056 10248 7112 0 FreeSans 224 0 0 0 NN4BEG[0]
port 140 nsew signal output
flabel metal2 s 12432 7056 12488 7112 0 FreeSans 224 0 0 0 NN4BEG[10]
port 141 nsew signal output
flabel metal2 s 12656 7056 12712 7112 0 FreeSans 224 0 0 0 NN4BEG[11]
port 142 nsew signal output
flabel metal2 s 12880 7056 12936 7112 0 FreeSans 224 0 0 0 NN4BEG[12]
port 143 nsew signal output
flabel metal2 s 13104 7056 13160 7112 0 FreeSans 224 0 0 0 NN4BEG[13]
port 144 nsew signal output
flabel metal2 s 13328 7056 13384 7112 0 FreeSans 224 0 0 0 NN4BEG[14]
port 145 nsew signal output
flabel metal2 s 13552 7056 13608 7112 0 FreeSans 224 0 0 0 NN4BEG[15]
port 146 nsew signal output
flabel metal2 s 10416 7056 10472 7112 0 FreeSans 224 0 0 0 NN4BEG[1]
port 147 nsew signal output
flabel metal2 s 10640 7056 10696 7112 0 FreeSans 224 0 0 0 NN4BEG[2]
port 148 nsew signal output
flabel metal2 s 10864 7056 10920 7112 0 FreeSans 224 0 0 0 NN4BEG[3]
port 149 nsew signal output
flabel metal2 s 11088 7056 11144 7112 0 FreeSans 224 0 0 0 NN4BEG[4]
port 150 nsew signal output
flabel metal2 s 11312 7056 11368 7112 0 FreeSans 224 0 0 0 NN4BEG[5]
port 151 nsew signal output
flabel metal2 s 11536 7056 11592 7112 0 FreeSans 224 0 0 0 NN4BEG[6]
port 152 nsew signal output
flabel metal2 s 11760 7056 11816 7112 0 FreeSans 224 0 0 0 NN4BEG[7]
port 153 nsew signal output
flabel metal2 s 11984 7056 12040 7112 0 FreeSans 224 0 0 0 NN4BEG[8]
port 154 nsew signal output
flabel metal2 s 12208 7056 12264 7112 0 FreeSans 224 0 0 0 NN4BEG[9]
port 155 nsew signal output
flabel metal2 s 13776 7056 13832 7112 0 FreeSans 224 0 0 0 S1END[0]
port 156 nsew signal input
flabel metal2 s 14000 7056 14056 7112 0 FreeSans 224 0 0 0 S1END[1]
port 157 nsew signal input
flabel metal2 s 14224 7056 14280 7112 0 FreeSans 224 0 0 0 S1END[2]
port 158 nsew signal input
flabel metal2 s 14448 7056 14504 7112 0 FreeSans 224 0 0 0 S1END[3]
port 159 nsew signal input
flabel metal2 s 16464 7056 16520 7112 0 FreeSans 224 0 0 0 S2END[0]
port 160 nsew signal input
flabel metal2 s 16688 7056 16744 7112 0 FreeSans 224 0 0 0 S2END[1]
port 161 nsew signal input
flabel metal2 s 16912 7056 16968 7112 0 FreeSans 224 0 0 0 S2END[2]
port 162 nsew signal input
flabel metal2 s 17136 7056 17192 7112 0 FreeSans 224 0 0 0 S2END[3]
port 163 nsew signal input
flabel metal2 s 17360 7056 17416 7112 0 FreeSans 224 0 0 0 S2END[4]
port 164 nsew signal input
flabel metal2 s 17584 7056 17640 7112 0 FreeSans 224 0 0 0 S2END[5]
port 165 nsew signal input
flabel metal2 s 17808 7056 17864 7112 0 FreeSans 224 0 0 0 S2END[6]
port 166 nsew signal input
flabel metal2 s 18032 7056 18088 7112 0 FreeSans 224 0 0 0 S2END[7]
port 167 nsew signal input
flabel metal2 s 14672 7056 14728 7112 0 FreeSans 224 0 0 0 S2MID[0]
port 168 nsew signal input
flabel metal2 s 14896 7056 14952 7112 0 FreeSans 224 0 0 0 S2MID[1]
port 169 nsew signal input
flabel metal2 s 15120 7056 15176 7112 0 FreeSans 224 0 0 0 S2MID[2]
port 170 nsew signal input
flabel metal2 s 15344 7056 15400 7112 0 FreeSans 224 0 0 0 S2MID[3]
port 171 nsew signal input
flabel metal2 s 15568 7056 15624 7112 0 FreeSans 224 0 0 0 S2MID[4]
port 172 nsew signal input
flabel metal2 s 15792 7056 15848 7112 0 FreeSans 224 0 0 0 S2MID[5]
port 173 nsew signal input
flabel metal2 s 16016 7056 16072 7112 0 FreeSans 224 0 0 0 S2MID[6]
port 174 nsew signal input
flabel metal2 s 16240 7056 16296 7112 0 FreeSans 224 0 0 0 S2MID[7]
port 175 nsew signal input
flabel metal2 s 18256 7056 18312 7112 0 FreeSans 224 0 0 0 S4END[0]
port 176 nsew signal input
flabel metal2 s 20496 7056 20552 7112 0 FreeSans 224 0 0 0 S4END[10]
port 177 nsew signal input
flabel metal2 s 20720 7056 20776 7112 0 FreeSans 224 0 0 0 S4END[11]
port 178 nsew signal input
flabel metal2 s 20944 7056 21000 7112 0 FreeSans 224 0 0 0 S4END[12]
port 179 nsew signal input
flabel metal2 s 21168 7056 21224 7112 0 FreeSans 224 0 0 0 S4END[13]
port 180 nsew signal input
flabel metal2 s 21392 7056 21448 7112 0 FreeSans 224 0 0 0 S4END[14]
port 181 nsew signal input
flabel metal2 s 21616 7056 21672 7112 0 FreeSans 224 0 0 0 S4END[15]
port 182 nsew signal input
flabel metal2 s 18480 7056 18536 7112 0 FreeSans 224 0 0 0 S4END[1]
port 183 nsew signal input
flabel metal2 s 18704 7056 18760 7112 0 FreeSans 224 0 0 0 S4END[2]
port 184 nsew signal input
flabel metal2 s 18928 7056 18984 7112 0 FreeSans 224 0 0 0 S4END[3]
port 185 nsew signal input
flabel metal2 s 19152 7056 19208 7112 0 FreeSans 224 0 0 0 S4END[4]
port 186 nsew signal input
flabel metal2 s 19376 7056 19432 7112 0 FreeSans 224 0 0 0 S4END[5]
port 187 nsew signal input
flabel metal2 s 19600 7056 19656 7112 0 FreeSans 224 0 0 0 S4END[6]
port 188 nsew signal input
flabel metal2 s 19824 7056 19880 7112 0 FreeSans 224 0 0 0 S4END[7]
port 189 nsew signal input
flabel metal2 s 20048 7056 20104 7112 0 FreeSans 224 0 0 0 S4END[8]
port 190 nsew signal input
flabel metal2 s 20272 7056 20328 7112 0 FreeSans 224 0 0 0 S4END[9]
port 191 nsew signal input
flabel metal2 s 21840 7056 21896 7112 0 FreeSans 224 0 0 0 SS4END[0]
port 192 nsew signal input
flabel metal2 s 24080 7056 24136 7112 0 FreeSans 224 0 0 0 SS4END[10]
port 193 nsew signal input
flabel metal2 s 24304 7056 24360 7112 0 FreeSans 224 0 0 0 SS4END[11]
port 194 nsew signal input
flabel metal2 s 24528 7056 24584 7112 0 FreeSans 224 0 0 0 SS4END[12]
port 195 nsew signal input
flabel metal2 s 24752 7056 24808 7112 0 FreeSans 224 0 0 0 SS4END[13]
port 196 nsew signal input
flabel metal2 s 24976 7056 25032 7112 0 FreeSans 224 0 0 0 SS4END[14]
port 197 nsew signal input
flabel metal2 s 25200 7056 25256 7112 0 FreeSans 224 0 0 0 SS4END[15]
port 198 nsew signal input
flabel metal2 s 22064 7056 22120 7112 0 FreeSans 224 0 0 0 SS4END[1]
port 199 nsew signal input
flabel metal2 s 22288 7056 22344 7112 0 FreeSans 224 0 0 0 SS4END[2]
port 200 nsew signal input
flabel metal2 s 22512 7056 22568 7112 0 FreeSans 224 0 0 0 SS4END[3]
port 201 nsew signal input
flabel metal2 s 22736 7056 22792 7112 0 FreeSans 224 0 0 0 SS4END[4]
port 202 nsew signal input
flabel metal2 s 22960 7056 23016 7112 0 FreeSans 224 0 0 0 SS4END[5]
port 203 nsew signal input
flabel metal2 s 23184 7056 23240 7112 0 FreeSans 224 0 0 0 SS4END[6]
port 204 nsew signal input
flabel metal2 s 23408 7056 23464 7112 0 FreeSans 224 0 0 0 SS4END[7]
port 205 nsew signal input
flabel metal2 s 23632 7056 23688 7112 0 FreeSans 224 0 0 0 SS4END[8]
port 206 nsew signal input
flabel metal2 s 23856 7056 23912 7112 0 FreeSans 224 0 0 0 SS4END[9]
port 207 nsew signal input
flabel metal2 s 1456 0 1512 56 0 FreeSans 224 0 0 0 UserCLK
port 208 nsew signal input
flabel metal2 s 25424 7056 25480 7112 0 FreeSans 224 0 0 0 UserCLKo
port 209 nsew signal output
flabel metal4 s 1888 0 2048 7112 0 FreeSans 736 90 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 1888 0 2048 28 0 FreeSans 184 0 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 1888 7084 2048 7112 0 FreeSans 184 0 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 11888 0 12048 7112 0 FreeSans 736 90 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 11888 0 12048 28 0 FreeSans 184 0 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 11888 7084 12048 7112 0 FreeSans 184 0 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 21888 0 22048 7112 0 FreeSans 736 90 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 21888 0 22048 28 0 FreeSans 184 0 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 21888 7084 22048 7112 0 FreeSans 184 0 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 2218 0 2378 7112 0 FreeSans 736 90 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 2218 0 2378 28 0 FreeSans 184 0 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 2218 7084 2378 7112 0 FreeSans 184 0 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 12218 0 12378 7112 0 FreeSans 736 90 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 12218 0 12378 28 0 FreeSans 184 0 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 12218 7084 12378 7112 0 FreeSans 184 0 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 22218 0 22378 7112 0 FreeSans 736 90 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 22218 0 22378 28 0 FreeSans 184 0 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 22218 7084 22378 7112 0 FreeSans 184 0 0 0 VSS
port 211 nsew ground bidirectional
rlabel metal1 16100 6272 16100 6272 0 VDD
rlabel metal1 16100 6664 16100 6664 0 VSS
rlabel metal2 4788 252 4788 252 0 FrameData[0]
rlabel metal3 12852 2940 12852 2940 0 FrameData[10]
rlabel metal2 10108 2660 10108 2660 0 FrameData[11]
rlabel metal3 11284 4340 11284 4340 0 FrameData[12]
rlabel metal2 6076 3500 6076 3500 0 FrameData[13]
rlabel metal2 8596 4396 8596 4396 0 FrameData[14]
rlabel metal2 10444 5180 10444 5180 0 FrameData[15]
rlabel metal2 10724 4648 10724 4648 0 FrameData[16]
rlabel metal2 10836 3080 10836 3080 0 FrameData[17]
rlabel metal3 259 4060 259 4060 0 FrameData[18]
rlabel metal3 12740 252 12740 252 0 FrameData[19]
rlabel metal2 4844 364 4844 364 0 FrameData[1]
rlabel metal2 12180 2016 12180 2016 0 FrameData[20]
rlabel metal3 861 4732 861 4732 0 FrameData[21]
rlabel metal2 13020 3388 13020 3388 0 FrameData[22]
rlabel metal2 3752 5012 3752 5012 0 FrameData[23]
rlabel metal2 11340 1148 11340 1148 0 FrameData[24]
rlabel metal3 868 5600 868 5600 0 FrameData[25]
rlabel metal2 12600 3724 12600 3724 0 FrameData[26]
rlabel metal3 427 6076 427 6076 0 FrameData[27]
rlabel metal2 12908 1708 12908 1708 0 FrameData[28]
rlabel metal4 10668 5516 10668 5516 0 FrameData[29]
rlabel metal3 259 476 259 476 0 FrameData[2]
rlabel metal3 861 6748 861 6748 0 FrameData[30]
rlabel metal3 91 6972 91 6972 0 FrameData[31]
rlabel metal2 12124 2156 12124 2156 0 FrameData[3]
rlabel metal3 483 924 483 924 0 FrameData[4]
rlabel metal3 1071 1148 1071 1148 0 FrameData[5]
rlabel metal4 13076 2324 13076 2324 0 FrameData[6]
rlabel metal3 931 1596 931 1596 0 FrameData[7]
rlabel metal4 10108 672 10108 672 0 FrameData[8]
rlabel metal3 1092 2072 1092 2072 0 FrameData[9]
rlabel metal3 31773 28 31773 28 0 FrameData_O[0]
rlabel metal3 31717 2268 31717 2268 0 FrameData_O[10]
rlabel metal2 31556 2380 31556 2380 0 FrameData_O[11]
rlabel metal2 31332 2660 31332 2660 0 FrameData_O[12]
rlabel metal3 31409 2940 31409 2940 0 FrameData_O[13]
rlabel metal2 31556 3108 31556 3108 0 FrameData_O[14]
rlabel metal3 31465 3388 31465 3388 0 FrameData_O[15]
rlabel metal2 31444 3444 31444 3444 0 FrameData_O[16]
rlabel metal3 31801 3836 31801 3836 0 FrameData_O[17]
rlabel metal2 31556 3948 31556 3948 0 FrameData_O[18]
rlabel metal3 31801 4284 31801 4284 0 FrameData_O[19]
rlabel metal3 30989 252 30989 252 0 FrameData_O[1]
rlabel metal3 31773 4508 31773 4508 0 FrameData_O[20]
rlabel metal3 31801 4732 31801 4732 0 FrameData_O[21]
rlabel metal3 31745 4956 31745 4956 0 FrameData_O[22]
rlabel metal3 30856 4956 30856 4956 0 FrameData_O[23]
rlabel metal3 31052 4620 31052 4620 0 FrameData_O[24]
rlabel metal3 30744 4844 30744 4844 0 FrameData_O[25]
rlabel metal3 30884 4172 30884 4172 0 FrameData_O[26]
rlabel metal3 31941 6076 31941 6076 0 FrameData_O[27]
rlabel metal2 29876 4088 29876 4088 0 FrameData_O[28]
rlabel metal3 29372 4844 29372 4844 0 FrameData_O[29]
rlabel metal3 31381 476 31381 476 0 FrameData_O[2]
rlabel metal3 31444 3052 31444 3052 0 FrameData_O[30]
rlabel metal2 27692 5432 27692 5432 0 FrameData_O[31]
rlabel metal3 31717 700 31717 700 0 FrameData_O[3]
rlabel metal2 31556 812 31556 812 0 FrameData_O[4]
rlabel metal2 31444 1036 31444 1036 0 FrameData_O[5]
rlabel metal3 31745 1372 31745 1372 0 FrameData_O[6]
rlabel metal2 31556 1540 31556 1540 0 FrameData_O[7]
rlabel metal3 31409 1820 31409 1820 0 FrameData_O[8]
rlabel metal2 31444 1876 31444 1876 0 FrameData_O[9]
rlabel metal2 2940 91 2940 91 0 FrameStrobe[0]
rlabel metal2 25004 588 25004 588 0 FrameStrobe[10]
rlabel metal2 23716 4592 23716 4592 0 FrameStrobe[11]
rlabel metal2 25032 2548 25032 2548 0 FrameStrobe[12]
rlabel metal2 25060 3080 25060 3080 0 FrameStrobe[13]
rlabel metal2 14924 3052 14924 3052 0 FrameStrobe[14]
rlabel metal2 24780 1155 24780 1155 0 FrameStrobe[15]
rlabel metal2 22036 4172 22036 4172 0 FrameStrobe[16]
rlabel metal2 27692 287 27692 287 0 FrameStrobe[17]
rlabel metal3 26376 1260 26376 1260 0 FrameStrobe[18]
rlabel metal3 29400 2044 29400 2044 0 FrameStrobe[19]
rlabel metal3 13356 5964 13356 5964 0 FrameStrobe[1]
rlabel metal2 13524 6244 13524 6244 0 FrameStrobe[2]
rlabel metal2 13636 1512 13636 1512 0 FrameStrobe[3]
rlabel metal2 10892 2128 10892 2128 0 FrameStrobe[4]
rlabel metal2 10220 399 10220 399 0 FrameStrobe[5]
rlabel metal2 11676 343 11676 343 0 FrameStrobe[6]
rlabel metal2 13132 175 13132 175 0 FrameStrobe[7]
rlabel metal2 14588 91 14588 91 0 FrameStrobe[8]
rlabel metal3 23968 924 23968 924 0 FrameStrobe[9]
rlabel metal2 25676 6825 25676 6825 0 FrameStrobe_O[0]
rlabel metal2 27916 6909 27916 6909 0 FrameStrobe_O[10]
rlabel metal2 28140 6601 28140 6601 0 FrameStrobe_O[11]
rlabel metal2 28364 6685 28364 6685 0 FrameStrobe_O[12]
rlabel metal2 28588 6797 28588 6797 0 FrameStrobe_O[13]
rlabel metal2 28812 6601 28812 6601 0 FrameStrobe_O[14]
rlabel metal2 29036 6769 29036 6769 0 FrameStrobe_O[15]
rlabel metal2 29260 6657 29260 6657 0 FrameStrobe_O[16]
rlabel metal2 29484 6825 29484 6825 0 FrameStrobe_O[17]
rlabel metal2 29708 6601 29708 6601 0 FrameStrobe_O[18]
rlabel metal2 29932 6713 29932 6713 0 FrameStrobe_O[19]
rlabel metal2 25900 6629 25900 6629 0 FrameStrobe_O[1]
rlabel metal2 26124 6433 26124 6433 0 FrameStrobe_O[2]
rlabel metal2 26348 6797 26348 6797 0 FrameStrobe_O[3]
rlabel metal2 26572 6909 26572 6909 0 FrameStrobe_O[4]
rlabel metal2 26796 6713 26796 6713 0 FrameStrobe_O[5]
rlabel metal2 27020 6629 27020 6629 0 FrameStrobe_O[6]
rlabel metal2 27244 6825 27244 6825 0 FrameStrobe_O[7]
rlabel metal2 27468 6965 27468 6965 0 FrameStrobe_O[8]
rlabel metal2 27692 6769 27692 6769 0 FrameStrobe_O[9]
rlabel metal2 1260 6496 1260 6496 0 N1BEG[0]
rlabel metal2 2380 6909 2380 6909 0 N1BEG[1]
rlabel metal3 2464 5796 2464 5796 0 N1BEG[2]
rlabel metal2 2828 6937 2828 6937 0 N1BEG[3]
rlabel metal2 3052 6349 3052 6349 0 N2BEG[0]
rlabel metal2 3444 5964 3444 5964 0 N2BEG[1]
rlabel metal2 2996 6608 2996 6608 0 N2BEG[2]
rlabel metal2 3724 6629 3724 6629 0 N2BEG[3]
rlabel metal2 4060 5992 4060 5992 0 N2BEG[4]
rlabel metal3 4032 5796 4032 5796 0 N2BEG[5]
rlabel metal2 3780 6608 3780 6608 0 N2BEG[6]
rlabel metal2 4732 5404 4732 5404 0 N2BEG[7]
rlabel metal2 4844 6629 4844 6629 0 N2BEGb[0]
rlabel metal2 5068 6685 5068 6685 0 N2BEGb[1]
rlabel metal2 5292 6629 5292 6629 0 N2BEGb[2]
rlabel metal2 5628 5768 5628 5768 0 N2BEGb[3]
rlabel metal3 5600 5796 5600 5796 0 N2BEGb[4]
rlabel metal2 4900 6664 4900 6664 0 N2BEGb[5]
rlabel metal2 6188 6349 6188 6349 0 N2BEGb[6]
rlabel metal2 6412 6629 6412 6629 0 N2BEGb[7]
rlabel metal2 5684 6608 5684 6608 0 N4BEG[0]
rlabel metal2 8876 6237 8876 6237 0 N4BEG[10]
rlabel metal2 9100 6797 9100 6797 0 N4BEG[11]
rlabel metal2 9548 5656 9548 5656 0 N4BEG[12]
rlabel metal2 9548 6629 9548 6629 0 N4BEG[13]
rlabel metal2 8708 6608 8708 6608 0 N4BEG[14]
rlabel metal2 9968 6188 9968 6188 0 N4BEG[15]
rlabel metal2 6860 6965 6860 6965 0 N4BEG[1]
rlabel metal2 7168 5404 7168 5404 0 N4BEG[2]
rlabel metal2 7196 5964 7196 5964 0 N4BEG[3]
rlabel metal2 6972 6580 6972 6580 0 N4BEG[4]
rlabel metal2 7756 6237 7756 6237 0 N4BEG[5]
rlabel metal2 7980 6769 7980 6769 0 N4BEG[6]
rlabel metal2 7980 5992 7980 5992 0 N4BEG[7]
rlabel metal2 8428 6797 8428 6797 0 N4BEG[8]
rlabel metal2 8652 6629 8652 6629 0 N4BEG[9]
rlabel metal2 10192 5796 10192 5796 0 NN4BEG[0]
rlabel metal2 12516 6188 12516 6188 0 NN4BEG[10]
rlabel metal2 12516 6636 12516 6636 0 NN4BEG[11]
rlabel metal2 12908 6349 12908 6349 0 NN4BEG[12]
rlabel metal3 13300 6132 13300 6132 0 NN4BEG[13]
rlabel metal2 13328 6580 13328 6580 0 NN4BEG[14]
rlabel metal2 13580 6909 13580 6909 0 NN4BEG[15]
rlabel metal2 10444 6825 10444 6825 0 NN4BEG[1]
rlabel metal2 10668 6349 10668 6349 0 NN4BEG[2]
rlabel metal3 10976 5404 10976 5404 0 NN4BEG[3]
rlabel metal3 10864 6580 10864 6580 0 NN4BEG[4]
rlabel metal2 11340 6629 11340 6629 0 NN4BEG[5]
rlabel metal2 11564 6349 11564 6349 0 NN4BEG[6]
rlabel metal2 11928 5404 11928 5404 0 NN4BEG[7]
rlabel metal3 11704 6580 11704 6580 0 NN4BEG[8]
rlabel metal2 12236 6909 12236 6909 0 NN4BEG[9]
rlabel metal2 11620 2240 11620 2240 0 S1END[0]
rlabel metal2 14028 6685 14028 6685 0 S1END[1]
rlabel metal2 14252 7049 14252 7049 0 S1END[2]
rlabel metal3 1344 2548 1344 2548 0 S1END[3]
rlabel metal2 21364 2744 21364 2744 0 S2END[0]
rlabel metal2 19908 3052 19908 3052 0 S2END[1]
rlabel metal3 24780 4368 24780 4368 0 S2END[2]
rlabel metal2 23492 3304 23492 3304 0 S2END[3]
rlabel metal2 22092 3192 22092 3192 0 S2END[4]
rlabel metal2 23268 6216 23268 6216 0 S2END[5]
rlabel metal3 17892 3780 17892 3780 0 S2END[6]
rlabel metal3 26320 4508 26320 4508 0 S2END[7]
rlabel metal3 13104 2660 13104 2660 0 S2MID[0]
rlabel metal2 14924 6853 14924 6853 0 S2MID[1]
rlabel metal2 14924 4928 14924 4928 0 S2MID[2]
rlabel metal2 12376 1876 12376 1876 0 S2MID[3]
rlabel metal4 11564 1932 11564 1932 0 S2MID[4]
rlabel metal3 11452 3472 11452 3472 0 S2MID[5]
rlabel metal2 8820 3220 8820 3220 0 S2MID[6]
rlabel metal3 9352 1876 9352 1876 0 S2MID[7]
rlabel metal2 9828 5600 9828 5600 0 S4END[0]
rlabel metal2 1428 1204 1428 1204 0 S4END[10]
rlabel metal3 1400 1764 1400 1764 0 S4END[11]
rlabel metal3 1260 2044 1260 2044 0 S4END[12]
rlabel metal2 13468 1428 13468 1428 0 S4END[13]
rlabel metal3 15148 2884 15148 2884 0 S4END[14]
rlabel metal2 16436 1008 16436 1008 0 S4END[15]
rlabel metal2 18508 3332 18508 3332 0 S4END[1]
rlabel metal2 13580 2968 13580 2968 0 S4END[2]
rlabel metal2 15372 3304 15372 3304 0 S4END[3]
rlabel metal3 11508 3388 11508 3388 0 S4END[4]
rlabel metal2 1372 5516 1372 5516 0 S4END[5]
rlabel metal3 11032 2660 11032 2660 0 S4END[6]
rlabel metal3 13076 3080 13076 3080 0 S4END[7]
rlabel metal2 1372 3164 1372 3164 0 S4END[8]
rlabel metal3 1260 476 1260 476 0 S4END[9]
rlabel metal2 15596 6244 15596 6244 0 SS4END[0]
rlabel metal2 22708 1820 22708 1820 0 SS4END[10]
rlabel metal3 23072 980 23072 980 0 SS4END[11]
rlabel metal3 23800 1092 23800 1092 0 SS4END[12]
rlabel metal2 24612 2212 24612 2212 0 SS4END[13]
rlabel metal2 23716 2044 23716 2044 0 SS4END[14]
rlabel metal2 25340 1876 25340 1876 0 SS4END[15]
rlabel metal2 22092 6965 22092 6965 0 SS4END[1]
rlabel metal2 22316 6909 22316 6909 0 SS4END[2]
rlabel metal2 22540 6741 22540 6741 0 SS4END[3]
rlabel metal2 22764 4753 22764 4753 0 SS4END[4]
rlabel metal2 22988 6489 22988 6489 0 SS4END[5]
rlabel metal2 23212 5425 23212 5425 0 SS4END[6]
rlabel metal2 23324 3206 23324 3206 0 SS4END[7]
rlabel metal2 23660 6993 23660 6993 0 SS4END[8]
rlabel metal3 22820 1120 22820 1120 0 SS4END[9]
rlabel metal2 1484 455 1484 455 0 UserCLK
rlabel metal2 25452 6825 25452 6825 0 UserCLKo
rlabel metal3 22092 840 22092 840 0 net1
rlabel metal3 12460 1232 12460 1232 0 net10
rlabel metal3 11928 1652 11928 1652 0 net100
rlabel metal3 13888 1876 13888 1876 0 net101
rlabel metal3 14308 5040 14308 5040 0 net102
rlabel metal2 15204 5460 15204 5460 0 net103
rlabel metal3 13328 3948 13328 3948 0 net104
rlabel metal2 15428 1176 15428 1176 0 net105
rlabel metal2 31108 5068 31108 5068 0 net11
rlabel metal2 13020 1260 13020 1260 0 net12
rlabel metal3 30492 3332 30492 3332 0 net13
rlabel metal4 11844 3220 11844 3220 0 net14
rlabel metal2 28980 3136 28980 3136 0 net15
rlabel metal4 14252 4928 14252 4928 0 net16
rlabel metal3 29260 4172 29260 4172 0 net17
rlabel metal4 14196 4956 14196 4956 0 net18
rlabel metal3 29204 4452 29204 4452 0 net19
rlabel metal3 28980 2548 28980 2548 0 net2
rlabel metal2 29596 5264 29596 5264 0 net20
rlabel metal2 29288 4116 29288 4116 0 net21
rlabel metal2 28812 4732 28812 4732 0 net22
rlabel metal2 30100 952 30100 952 0 net23
rlabel metal3 10836 2632 10836 2632 0 net24
rlabel metal2 29596 3990 29596 3990 0 net25
rlabel metal3 29484 1036 29484 1036 0 net26
rlabel metal2 4900 560 4900 560 0 net27
rlabel metal3 30464 980 30464 980 0 net28
rlabel metal2 30072 1764 30072 1764 0 net29
rlabel metal2 31164 2408 31164 2408 0 net3
rlabel metal3 30380 1372 30380 1372 0 net30
rlabel metal2 29260 1064 29260 1064 0 net31
rlabel metal2 13300 1932 13300 1932 0 net32
rlabel metal2 23324 5628 23324 5628 0 net33
rlabel metal2 25452 1708 25452 1708 0 net34
rlabel metal2 24108 4788 24108 4788 0 net35
rlabel metal3 26292 2604 26292 2604 0 net36
rlabel metal3 25984 3332 25984 3332 0 net37
rlabel metal3 15232 2604 15232 2604 0 net38
rlabel metal3 23380 1988 23380 1988 0 net39
rlabel metal3 30464 2548 30464 2548 0 net4
rlabel metal2 21756 4032 21756 4032 0 net40
rlabel metal3 24836 5740 24836 5740 0 net41
rlabel metal2 26068 1456 26068 1456 0 net42
rlabel metal3 29120 2212 29120 2212 0 net43
rlabel metal2 14924 6328 14924 6328 0 net44
rlabel metal2 17892 5852 17892 5852 0 net45
rlabel metal3 23744 6076 23744 6076 0 net46
rlabel metal2 27188 6244 27188 6244 0 net47
rlabel metal2 27020 5460 27020 5460 0 net48
rlabel metal2 22400 2884 22400 2884 0 net49
rlabel metal3 12572 1932 12572 1932 0 net5
rlabel metal2 22484 1960 22484 1960 0 net50
rlabel metal3 27188 1624 27188 1624 0 net51
rlabel metal3 26460 1036 26460 1036 0 net52
rlabel metal2 1008 2604 1008 2604 0 net53
rlabel metal2 4116 4424 4116 4424 0 net54
rlabel metal2 7812 1876 7812 1876 0 net55
rlabel metal2 10500 2772 10500 2772 0 net56
rlabel metal3 7966 1820 7966 1820 0 net57
rlabel metal2 5012 3192 5012 3192 0 net58
rlabel metal2 3248 2604 3248 2604 0 net59
rlabel metal3 11844 4732 11844 4732 0 net6
rlabel metal2 7364 1064 7364 1064 0 net60
rlabel metal2 11788 1960 11788 1960 0 net61
rlabel metal2 6244 5096 6244 5096 0 net62
rlabel metal2 17668 3724 17668 3724 0 net63
rlabel metal2 12180 2828 12180 2828 0 net64
rlabel metal2 13524 5012 13524 5012 0 net65
rlabel metal2 13412 4200 13412 4200 0 net66
rlabel metal3 12488 4172 12488 4172 0 net67
rlabel metal3 22932 5544 22932 5544 0 net68
rlabel metal3 10080 3192 10080 3192 0 net69
rlabel metal3 18956 3892 18956 3892 0 net7
rlabel metal2 13524 980 13524 980 0 net70
rlabel metal4 16100 5236 16100 5236 0 net71
rlabel metal2 13524 3136 13524 3136 0 net72
rlabel metal2 12180 1092 12180 1092 0 net73
rlabel metal2 8652 5460 8652 5460 0 net74
rlabel metal2 7420 4732 7420 4732 0 net75
rlabel metal3 12180 2688 12180 2688 0 net76
rlabel metal2 13300 3136 13300 3136 0 net77
rlabel metal3 12180 2800 12180 2800 0 net78
rlabel metal2 6916 5320 6916 5320 0 net79
rlabel metal3 13300 4900 13300 4900 0 net8
rlabel metal2 14784 2996 14784 2996 0 net80
rlabel metal3 7980 5236 7980 5236 0 net81
rlabel metal2 924 2408 924 2408 0 net82
rlabel metal2 1092 4060 1092 4060 0 net83
rlabel metal2 7924 1484 7924 1484 0 net84
rlabel metal4 4676 476 4676 476 0 net85
rlabel metal2 7084 3724 7084 3724 0 net86
rlabel metal3 8344 3332 8344 3332 0 net87
rlabel metal3 10136 2604 10136 2604 0 net88
rlabel metal2 24948 1820 24948 1820 0 net89
rlabel metal3 30268 2996 30268 2996 0 net9
rlabel metal2 13188 5292 13188 5292 0 net90
rlabel metal3 13496 1932 13496 1932 0 net91
rlabel metal3 14644 5684 14644 5684 0 net92
rlabel metal3 14364 5124 14364 5124 0 net93
rlabel metal2 13804 2674 13804 2674 0 net94
rlabel metal3 14840 6132 14840 6132 0 net95
rlabel metal2 23268 2156 23268 2156 0 net96
rlabel metal2 22652 1876 22652 1876 0 net97
rlabel metal2 22764 924 22764 924 0 net98
rlabel metal3 14644 4172 14644 4172 0 net99
<< properties >>
string FIXED_BBOX 0 0 32200 7112
<< end >>
