magic
tech gf180mcuD
magscale 1 5
timestamp 1764970367
<< metal1 >>
rect 336 6677 28392 6694
rect 336 6651 2233 6677
rect 2259 6651 2285 6677
rect 2311 6651 2337 6677
rect 2363 6651 12233 6677
rect 12259 6651 12285 6677
rect 12311 6651 12337 6677
rect 12363 6651 22233 6677
rect 22259 6651 22285 6677
rect 22311 6651 22337 6677
rect 22363 6651 28392 6677
rect 336 6634 28392 6651
rect 5335 6593 5361 6599
rect 1017 6567 1023 6593
rect 1049 6567 1055 6593
rect 5335 6561 5361 6567
rect 26559 6593 26585 6599
rect 26559 6561 26585 6567
rect 4041 6511 4047 6537
rect 4073 6511 4079 6537
rect 1191 6481 1217 6487
rect 3033 6455 3039 6481
rect 3065 6455 3071 6481
rect 5161 6455 5167 6481
rect 5193 6455 5199 6481
rect 7009 6455 7015 6481
rect 7041 6455 7047 6481
rect 9697 6455 9703 6481
rect 9729 6455 9735 6481
rect 11041 6455 11047 6481
rect 11073 6455 11079 6481
rect 12553 6455 12559 6481
rect 12585 6455 12591 6481
rect 13561 6455 13567 6481
rect 13593 6455 13599 6481
rect 15073 6455 15079 6481
rect 15105 6455 15111 6481
rect 16417 6455 16423 6481
rect 16449 6455 16455 6481
rect 19105 6455 19111 6481
rect 19137 6455 19143 6481
rect 20449 6455 20455 6481
rect 20481 6455 20487 6481
rect 22073 6455 22079 6481
rect 22105 6455 22111 6481
rect 23081 6455 23087 6481
rect 23113 6455 23119 6481
rect 24481 6455 24487 6481
rect 24513 6455 24519 6481
rect 25881 6455 25887 6481
rect 25913 6455 25919 6481
rect 26273 6455 26279 6481
rect 26305 6455 26311 6481
rect 27673 6455 27679 6481
rect 27705 6455 27711 6481
rect 1191 6449 1217 6455
rect 2535 6425 2561 6431
rect 6511 6425 6537 6431
rect 3593 6399 3599 6425
rect 3625 6399 3631 6425
rect 2535 6393 2561 6399
rect 6511 6393 6537 6399
rect 9199 6425 9225 6431
rect 9199 6393 9225 6399
rect 10543 6425 10569 6431
rect 10543 6393 10569 6399
rect 12055 6425 12081 6431
rect 12055 6393 12081 6399
rect 13063 6425 13089 6431
rect 13063 6393 13089 6399
rect 14575 6425 14601 6431
rect 14575 6393 14601 6399
rect 15919 6425 15945 6431
rect 15919 6393 15945 6399
rect 18607 6425 18633 6431
rect 18607 6393 18633 6399
rect 19951 6425 19977 6431
rect 19951 6393 19977 6399
rect 21575 6425 21601 6431
rect 21575 6393 21601 6399
rect 22583 6425 22609 6431
rect 22583 6393 22609 6399
rect 23983 6425 24009 6431
rect 23983 6393 24009 6399
rect 25383 6425 25409 6431
rect 25383 6393 25409 6399
rect 28071 6369 28097 6375
rect 28071 6337 28097 6343
rect 336 6285 28392 6302
rect 336 6259 1903 6285
rect 1929 6259 1955 6285
rect 1981 6259 2007 6285
rect 2033 6259 11903 6285
rect 11929 6259 11955 6285
rect 11981 6259 12007 6285
rect 12033 6259 21903 6285
rect 21929 6259 21955 6285
rect 21981 6259 22007 6285
rect 22033 6259 28392 6285
rect 336 6242 28392 6259
rect 7855 6201 7881 6207
rect 7855 6169 7881 6175
rect 17263 6201 17289 6207
rect 17263 6169 17289 6175
rect 26503 6201 26529 6207
rect 26503 6169 26529 6175
rect 5223 6145 5249 6151
rect 5223 6113 5249 6119
rect 5671 6145 5697 6151
rect 10319 6145 10345 6151
rect 7513 6119 7519 6145
rect 7545 6119 7551 6145
rect 5671 6113 5697 6119
rect 10319 6113 10345 6119
rect 10767 6145 10793 6151
rect 10767 6113 10793 6119
rect 11159 6145 11185 6151
rect 11159 6113 11185 6119
rect 11551 6145 11577 6151
rect 11551 6113 11577 6119
rect 13063 6145 13089 6151
rect 13063 6113 13089 6119
rect 13231 6145 13257 6151
rect 13231 6113 13257 6119
rect 16087 6145 16113 6151
rect 19951 6145 19977 6151
rect 16417 6119 16423 6145
rect 16449 6119 16455 6145
rect 16087 6113 16113 6119
rect 19951 6113 19977 6119
rect 23255 6145 23281 6151
rect 24985 6119 24991 6145
rect 25017 6119 25023 6145
rect 23255 6113 23281 6119
rect 5503 6089 5529 6095
rect 5503 6057 5529 6063
rect 10599 6089 10625 6095
rect 10599 6057 10625 6063
rect 11719 6089 11745 6095
rect 11719 6057 11745 6063
rect 14015 6089 14041 6095
rect 14015 6057 14041 6063
rect 14239 6089 14265 6095
rect 14239 6057 14265 6063
rect 14519 6089 14545 6095
rect 14519 6057 14545 6063
rect 16199 6089 16225 6095
rect 16199 6057 16225 6063
rect 23423 6089 23449 6095
rect 26105 6063 26111 6089
rect 26137 6063 26143 6089
rect 26777 6063 26783 6089
rect 26809 6063 26815 6089
rect 23423 6057 23449 6063
rect 11999 6033 12025 6039
rect 8353 6007 8359 6033
rect 8385 6007 8391 6033
rect 11999 6001 12025 6007
rect 15359 6033 15385 6039
rect 18551 6033 18577 6039
rect 17761 6007 17767 6033
rect 17793 6007 17799 6033
rect 15359 6001 15385 6007
rect 18551 6001 18577 6007
rect 20231 6033 20257 6039
rect 20231 6001 20257 6007
rect 20399 6033 20425 6039
rect 20399 6001 20425 6007
rect 23703 6033 23729 6039
rect 27169 6007 27175 6033
rect 27201 6007 27207 6033
rect 27561 6007 27567 6033
rect 27593 6007 27599 6033
rect 27953 6007 27959 6033
rect 27985 6007 27991 6033
rect 23703 6001 23729 6007
rect 7183 5977 7209 5983
rect 7183 5945 7209 5951
rect 7295 5977 7321 5983
rect 7295 5945 7321 5951
rect 11439 5977 11465 5983
rect 11439 5945 11465 5951
rect 12671 5977 12697 5983
rect 12671 5945 12697 5951
rect 12783 5977 12809 5983
rect 12783 5945 12809 5951
rect 13511 5977 13537 5983
rect 13511 5945 13537 5951
rect 13679 5977 13705 5983
rect 13679 5945 13705 5951
rect 14967 5977 14993 5983
rect 14967 5945 14993 5951
rect 15079 5977 15105 5983
rect 15079 5945 15105 5951
rect 18831 5977 18857 5983
rect 18831 5945 18857 5951
rect 18999 5977 19025 5983
rect 22471 5977 22497 5983
rect 22297 5951 22303 5977
rect 22329 5951 22335 5977
rect 18999 5945 19025 5951
rect 22471 5945 22497 5951
rect 22639 5977 22665 5983
rect 22639 5945 22665 5951
rect 24655 5977 24681 5983
rect 24655 5945 24681 5951
rect 24767 5977 24793 5983
rect 24767 5945 24793 5951
rect 336 5893 28392 5910
rect 336 5867 2233 5893
rect 2259 5867 2285 5893
rect 2311 5867 2337 5893
rect 2363 5867 12233 5893
rect 12259 5867 12285 5893
rect 12311 5867 12337 5893
rect 12363 5867 22233 5893
rect 22259 5867 22285 5893
rect 22311 5867 22337 5893
rect 22363 5867 28392 5893
rect 336 5850 28392 5867
rect 7407 5809 7433 5815
rect 7407 5777 7433 5783
rect 7519 5809 7545 5815
rect 7519 5777 7545 5783
rect 7127 5753 7153 5759
rect 7127 5721 7153 5727
rect 9087 5753 9113 5759
rect 25489 5727 25495 5753
rect 25521 5727 25527 5753
rect 25881 5727 25887 5753
rect 25913 5727 25919 5753
rect 9087 5721 9113 5727
rect 9367 5697 9393 5703
rect 9367 5665 9393 5671
rect 9479 5697 9505 5703
rect 9479 5665 9505 5671
rect 12279 5697 12305 5703
rect 12279 5665 12305 5671
rect 17543 5697 17569 5703
rect 17543 5665 17569 5671
rect 23759 5697 23785 5703
rect 26385 5671 26391 5697
rect 26417 5671 26423 5697
rect 27057 5671 27063 5697
rect 27089 5671 27095 5697
rect 23759 5665 23785 5671
rect 11551 5641 11577 5647
rect 11551 5609 11577 5615
rect 11999 5641 12025 5647
rect 11999 5609 12025 5615
rect 12559 5641 12585 5647
rect 12559 5609 12585 5615
rect 17375 5641 17401 5647
rect 17375 5609 17401 5615
rect 17823 5641 17849 5647
rect 23983 5641 24009 5647
rect 23529 5615 23535 5641
rect 23561 5615 23567 5641
rect 17823 5609 17849 5615
rect 23983 5609 24009 5615
rect 26783 5585 26809 5591
rect 26783 5553 26809 5559
rect 27567 5585 27593 5591
rect 27567 5553 27593 5559
rect 336 5501 28392 5518
rect 336 5475 1903 5501
rect 1929 5475 1955 5501
rect 1981 5475 2007 5501
rect 2033 5475 11903 5501
rect 11929 5475 11955 5501
rect 11981 5475 12007 5501
rect 12033 5475 21903 5501
rect 21929 5475 21955 5501
rect 21981 5475 22007 5501
rect 22033 5475 28392 5501
rect 336 5458 28392 5475
rect 26503 5417 26529 5423
rect 26503 5385 26529 5391
rect 14351 5361 14377 5367
rect 14351 5329 14377 5335
rect 14799 5361 14825 5367
rect 14799 5329 14825 5335
rect 17095 5361 17121 5367
rect 17095 5329 17121 5335
rect 27287 5361 27313 5367
rect 27287 5329 27313 5335
rect 28071 5361 28097 5367
rect 28071 5329 28097 5335
rect 14631 5305 14657 5311
rect 14631 5273 14657 5279
rect 17263 5305 17289 5311
rect 17263 5273 17289 5279
rect 19279 5305 19305 5311
rect 26049 5279 26055 5305
rect 26081 5279 26087 5305
rect 27617 5279 27623 5305
rect 27649 5279 27655 5305
rect 19279 5273 19305 5279
rect 15695 5249 15721 5255
rect 15695 5217 15721 5223
rect 17543 5249 17569 5255
rect 26777 5223 26783 5249
rect 26809 5223 26815 5249
rect 17543 5217 17569 5223
rect 15247 5193 15273 5199
rect 15247 5161 15273 5167
rect 15415 5193 15441 5199
rect 15415 5161 15441 5167
rect 18831 5193 18857 5199
rect 18831 5161 18857 5167
rect 18999 5193 19025 5199
rect 18999 5161 19025 5167
rect 336 5109 28392 5126
rect 336 5083 2233 5109
rect 2259 5083 2285 5109
rect 2311 5083 2337 5109
rect 2363 5083 12233 5109
rect 12259 5083 12285 5109
rect 12311 5083 12337 5109
rect 12363 5083 22233 5109
rect 22259 5083 22285 5109
rect 22311 5083 22337 5109
rect 22363 5083 28392 5109
rect 336 5066 28392 5083
rect 9535 5025 9561 5031
rect 9535 4993 9561 4999
rect 9703 5025 9729 5031
rect 9703 4993 9729 4999
rect 17207 5025 17233 5031
rect 17207 4993 17233 4999
rect 17319 5025 17345 5031
rect 17319 4993 17345 4999
rect 16311 4969 16337 4975
rect 16311 4937 16337 4943
rect 17599 4969 17625 4975
rect 26273 4943 26279 4969
rect 26305 4943 26311 4969
rect 17599 4937 17625 4943
rect 16591 4913 16617 4919
rect 27057 4887 27063 4913
rect 27089 4887 27095 4913
rect 16591 4881 16617 4887
rect 9983 4857 10009 4863
rect 9983 4825 10009 4831
rect 16703 4857 16729 4863
rect 16703 4825 16729 4831
rect 26783 4857 26809 4863
rect 26783 4825 26809 4831
rect 27567 4801 27593 4807
rect 27567 4769 27593 4775
rect 336 4717 28392 4734
rect 336 4691 1903 4717
rect 1929 4691 1955 4717
rect 1981 4691 2007 4717
rect 2033 4691 11903 4717
rect 11929 4691 11955 4717
rect 11981 4691 12007 4717
rect 12033 4691 21903 4717
rect 21929 4691 21955 4717
rect 21981 4691 22007 4717
rect 22033 4691 28392 4717
rect 336 4674 28392 4691
rect 11159 4577 11185 4583
rect 11159 4545 11185 4551
rect 12615 4577 12641 4583
rect 12615 4545 12641 4551
rect 13063 4577 13089 4583
rect 13063 4545 13089 4551
rect 14015 4577 14041 4583
rect 14457 4551 14463 4577
rect 14489 4551 14495 4577
rect 14015 4545 14041 4551
rect 11327 4521 11353 4527
rect 11327 4489 11353 4495
rect 11607 4521 11633 4527
rect 11607 4489 11633 4495
rect 12783 4521 12809 4527
rect 12783 4489 12809 4495
rect 14239 4521 14265 4527
rect 27617 4495 27623 4521
rect 27649 4495 27655 4521
rect 14239 4489 14265 4495
rect 1471 4465 1497 4471
rect 1471 4433 1497 4439
rect 20455 4465 20481 4471
rect 20455 4433 20481 4439
rect 20567 4465 20593 4471
rect 20567 4433 20593 4439
rect 20847 4465 20873 4471
rect 20847 4433 20873 4439
rect 22359 4465 22385 4471
rect 26777 4439 26783 4465
rect 26809 4439 26815 4465
rect 27169 4439 27175 4465
rect 27201 4439 27207 4465
rect 27953 4439 27959 4465
rect 27985 4439 27991 4465
rect 22359 4433 22385 4439
rect 1079 4409 1105 4415
rect 1079 4377 1105 4383
rect 1191 4409 1217 4415
rect 1191 4377 1217 4383
rect 21855 4409 21881 4415
rect 21855 4377 21881 4383
rect 22079 4409 22105 4415
rect 22079 4377 22105 4383
rect 336 4325 28392 4342
rect 336 4299 2233 4325
rect 2259 4299 2285 4325
rect 2311 4299 2337 4325
rect 2363 4299 12233 4325
rect 12259 4299 12285 4325
rect 12311 4299 12337 4325
rect 12363 4299 22233 4325
rect 22259 4299 22285 4325
rect 22311 4299 22337 4325
rect 22363 4299 28392 4325
rect 336 4282 28392 4299
rect 11103 4185 11129 4191
rect 11103 4153 11129 4159
rect 11215 4185 11241 4191
rect 11215 4153 11241 4159
rect 11495 4185 11521 4191
rect 27449 4159 27455 4185
rect 27481 4159 27487 4185
rect 11495 4153 11521 4159
rect 9143 4129 9169 4135
rect 9143 4097 9169 4103
rect 14631 4129 14657 4135
rect 14631 4097 14657 4103
rect 15359 4129 15385 4135
rect 15359 4097 15385 4103
rect 21799 4129 21825 4135
rect 27057 4103 27063 4129
rect 27089 4103 27095 4129
rect 21799 4097 21825 4103
rect 9255 4073 9281 4079
rect 8913 4047 8919 4073
rect 8945 4047 8951 4073
rect 9255 4041 9281 4047
rect 14519 4073 14545 4079
rect 14519 4041 14545 4047
rect 14911 4073 14937 4079
rect 14911 4041 14937 4047
rect 15191 4073 15217 4079
rect 21631 4073 21657 4079
rect 15577 4047 15583 4073
rect 15609 4047 15615 4073
rect 15191 4041 15217 4047
rect 21631 4041 21657 4047
rect 22079 4073 22105 4079
rect 22079 4041 22105 4047
rect 336 3933 28392 3950
rect 336 3907 1903 3933
rect 1929 3907 1955 3933
rect 1981 3907 2007 3933
rect 2033 3907 11903 3933
rect 11929 3907 11955 3933
rect 11981 3907 12007 3933
rect 12033 3907 21903 3933
rect 21929 3907 21955 3933
rect 21981 3907 22007 3933
rect 22033 3907 28392 3933
rect 336 3890 28392 3907
rect 28071 3849 28097 3855
rect 28071 3817 28097 3823
rect 17375 3793 17401 3799
rect 13169 3767 13175 3793
rect 13201 3767 13207 3793
rect 17375 3761 17401 3767
rect 17823 3793 17849 3799
rect 17823 3761 17849 3767
rect 27287 3793 27313 3799
rect 27287 3761 27313 3767
rect 12839 3737 12865 3743
rect 12839 3705 12865 3711
rect 12951 3737 12977 3743
rect 12951 3705 12977 3711
rect 17543 3737 17569 3743
rect 26777 3711 26783 3737
rect 26809 3711 26815 3737
rect 27561 3711 27567 3737
rect 27593 3711 27599 3737
rect 17543 3705 17569 3711
rect 2703 3681 2729 3687
rect 2703 3649 2729 3655
rect 4551 3681 4577 3687
rect 4551 3649 4577 3655
rect 10711 3681 10737 3687
rect 10711 3649 10737 3655
rect 2983 3625 3009 3631
rect 2983 3593 3009 3599
rect 3151 3625 3177 3631
rect 3151 3593 3177 3599
rect 4831 3625 4857 3631
rect 4831 3593 4857 3599
rect 4999 3625 5025 3631
rect 4999 3593 5025 3599
rect 10263 3625 10289 3631
rect 10263 3593 10289 3599
rect 10431 3625 10457 3631
rect 10431 3593 10457 3599
rect 336 3541 28392 3558
rect 336 3515 2233 3541
rect 2259 3515 2285 3541
rect 2311 3515 2337 3541
rect 2363 3515 12233 3541
rect 12259 3515 12285 3541
rect 12311 3515 12337 3541
rect 12363 3515 22233 3541
rect 22259 3515 22285 3541
rect 22311 3515 22337 3541
rect 22363 3515 28392 3541
rect 336 3498 28392 3515
rect 7799 3345 7825 3351
rect 7799 3313 7825 3319
rect 13231 3345 13257 3351
rect 13231 3313 13257 3319
rect 21631 3345 21657 3351
rect 21631 3313 21657 3319
rect 22415 3345 22441 3351
rect 22415 3313 22441 3319
rect 22695 3345 22721 3351
rect 27057 3319 27063 3345
rect 27089 3319 27095 3345
rect 22695 3313 22721 3319
rect 7631 3289 7657 3295
rect 7631 3257 7657 3263
rect 8079 3289 8105 3295
rect 8079 3257 8105 3263
rect 13063 3289 13089 3295
rect 13063 3257 13089 3263
rect 13511 3289 13537 3295
rect 13511 3257 13537 3263
rect 21463 3289 21489 3295
rect 22247 3289 22273 3295
rect 21849 3263 21855 3289
rect 21881 3263 21887 3289
rect 21463 3257 21489 3263
rect 22247 3257 22273 3263
rect 27567 3233 27593 3239
rect 27567 3201 27593 3207
rect 336 3149 28392 3166
rect 336 3123 1903 3149
rect 1929 3123 1955 3149
rect 1981 3123 2007 3149
rect 2033 3123 11903 3149
rect 11929 3123 11955 3149
rect 11981 3123 12007 3149
rect 12033 3123 21903 3149
rect 21929 3123 21955 3149
rect 21981 3123 22007 3149
rect 22033 3123 28392 3149
rect 336 3106 28392 3123
rect 28071 3065 28097 3071
rect 28071 3033 28097 3039
rect 12671 3009 12697 3015
rect 12671 2977 12697 2983
rect 17487 3009 17513 3015
rect 18551 3009 18577 3015
rect 17817 2983 17823 3009
rect 17849 2983 17855 3009
rect 17487 2977 17513 2983
rect 18551 2977 18577 2983
rect 23199 3009 23225 3015
rect 23199 2977 23225 2983
rect 26503 3009 26529 3015
rect 26503 2977 26529 2983
rect 27287 3009 27313 3015
rect 27287 2977 27313 2983
rect 17599 2953 17625 2959
rect 12441 2927 12447 2953
rect 12473 2927 12479 2953
rect 17599 2921 17625 2927
rect 18663 2953 18689 2959
rect 18663 2921 18689 2927
rect 23311 2953 23337 2959
rect 23311 2921 23337 2927
rect 24599 2953 24625 2959
rect 24599 2921 24625 2927
rect 24711 2953 24737 2959
rect 26777 2927 26783 2953
rect 26809 2927 26815 2953
rect 27561 2927 27567 2953
rect 27593 2927 27599 2953
rect 24711 2921 24737 2927
rect 7127 2897 7153 2903
rect 7127 2865 7153 2871
rect 8191 2897 8217 2903
rect 8191 2865 8217 2871
rect 8303 2897 8329 2903
rect 8303 2865 8329 2871
rect 8583 2897 8609 2903
rect 8583 2865 8609 2871
rect 12223 2897 12249 2903
rect 12223 2865 12249 2871
rect 18943 2897 18969 2903
rect 18943 2865 18969 2871
rect 20287 2897 20313 2903
rect 20287 2865 20313 2871
rect 23591 2897 23617 2903
rect 23591 2865 23617 2871
rect 24991 2897 25017 2903
rect 24991 2865 25017 2871
rect 7407 2841 7433 2847
rect 7407 2809 7433 2815
rect 7575 2841 7601 2847
rect 7575 2809 7601 2815
rect 11831 2841 11857 2847
rect 11831 2809 11857 2815
rect 11943 2841 11969 2847
rect 11943 2809 11969 2815
rect 19895 2841 19921 2847
rect 19895 2809 19921 2815
rect 20007 2841 20033 2847
rect 20007 2809 20033 2815
rect 26615 2841 26641 2847
rect 26615 2809 26641 2815
rect 336 2757 28392 2774
rect 336 2731 2233 2757
rect 2259 2731 2285 2757
rect 2311 2731 2337 2757
rect 2363 2731 12233 2757
rect 12259 2731 12285 2757
rect 12311 2731 12337 2757
rect 12363 2731 22233 2757
rect 22259 2731 22285 2757
rect 22311 2731 22337 2757
rect 22363 2731 28392 2757
rect 336 2714 28392 2731
rect 9143 2673 9169 2679
rect 9143 2641 9169 2647
rect 9311 2673 9337 2679
rect 9311 2641 9337 2647
rect 14295 2673 14321 2679
rect 14295 2641 14321 2647
rect 14463 2673 14489 2679
rect 14463 2641 14489 2647
rect 17151 2673 17177 2679
rect 17151 2641 17177 2647
rect 17319 2673 17345 2679
rect 17319 2641 17345 2647
rect 21127 2673 21153 2679
rect 21127 2641 21153 2647
rect 21295 2673 21321 2679
rect 21295 2641 21321 2647
rect 23311 2673 23337 2679
rect 23311 2641 23337 2647
rect 23479 2673 23505 2679
rect 23479 2641 23505 2647
rect 5167 2617 5193 2623
rect 5167 2585 5193 2591
rect 9759 2617 9785 2623
rect 9759 2585 9785 2591
rect 14911 2617 14937 2623
rect 14911 2585 14937 2591
rect 16479 2617 16505 2623
rect 16479 2585 16505 2591
rect 17599 2617 17625 2623
rect 17599 2585 17625 2591
rect 23759 2617 23785 2623
rect 23759 2585 23785 2591
rect 26167 2617 26193 2623
rect 26167 2585 26193 2591
rect 26447 2617 26473 2623
rect 27057 2591 27063 2617
rect 27089 2591 27095 2617
rect 26447 2585 26473 2591
rect 5447 2561 5473 2567
rect 5447 2529 5473 2535
rect 5559 2561 5585 2567
rect 5559 2529 5585 2535
rect 10039 2561 10065 2567
rect 10039 2529 10065 2535
rect 10151 2561 10177 2567
rect 10151 2529 10177 2535
rect 12223 2561 12249 2567
rect 12223 2529 12249 2535
rect 15191 2561 15217 2567
rect 15191 2529 15217 2535
rect 15975 2561 16001 2567
rect 15975 2529 16001 2535
rect 16199 2561 16225 2567
rect 16199 2529 16225 2535
rect 19111 2561 19137 2567
rect 19111 2529 19137 2535
rect 19279 2561 19305 2567
rect 19279 2529 19305 2535
rect 19559 2561 19585 2567
rect 19559 2529 19585 2535
rect 26615 2561 26641 2567
rect 27449 2535 27455 2561
rect 27481 2535 27487 2561
rect 26615 2529 26641 2535
rect 9591 2505 9617 2511
rect 9591 2473 9617 2479
rect 14743 2505 14769 2511
rect 14743 2473 14769 2479
rect 21575 2505 21601 2511
rect 21575 2473 21601 2479
rect 26895 2505 26921 2511
rect 26895 2473 26921 2479
rect 336 2365 28392 2382
rect 336 2339 1903 2365
rect 1929 2339 1955 2365
rect 1981 2339 2007 2365
rect 2033 2339 11903 2365
rect 11929 2339 11955 2365
rect 11981 2339 12007 2365
rect 12033 2339 21903 2365
rect 21929 2339 21955 2365
rect 21981 2339 22007 2365
rect 22033 2339 28392 2365
rect 336 2322 28392 2339
rect 27287 2281 27313 2287
rect 27287 2249 27313 2255
rect 28071 2281 28097 2287
rect 28071 2249 28097 2255
rect 16143 2225 16169 2231
rect 5105 2199 5111 2225
rect 5137 2199 5143 2225
rect 5889 2199 5895 2225
rect 5921 2199 5927 2225
rect 12161 2199 12167 2225
rect 12193 2199 12199 2225
rect 16143 2193 16169 2199
rect 17487 2225 17513 2231
rect 17487 2193 17513 2199
rect 20623 2225 20649 2231
rect 26335 2225 26361 2231
rect 20953 2199 20959 2225
rect 20985 2199 20991 2225
rect 20623 2193 20649 2199
rect 26335 2193 26361 2199
rect 16255 2169 16281 2175
rect 16255 2137 16281 2143
rect 17599 2169 17625 2175
rect 17599 2137 17625 2143
rect 18159 2169 18185 2175
rect 18159 2137 18185 2143
rect 20735 2169 20761 2175
rect 20735 2137 20761 2143
rect 22359 2169 22385 2175
rect 22359 2137 22385 2143
rect 22471 2169 22497 2175
rect 26777 2143 26783 2169
rect 26809 2143 26815 2169
rect 27561 2143 27567 2169
rect 27593 2143 27599 2169
rect 22471 2137 22497 2143
rect 1303 2113 1329 2119
rect 1303 2081 1329 2087
rect 9031 2113 9057 2119
rect 9031 2081 9057 2087
rect 16535 2113 16561 2119
rect 16535 2081 16561 2087
rect 17879 2113 17905 2119
rect 17879 2081 17905 2087
rect 18439 2113 18465 2119
rect 18439 2081 18465 2087
rect 19895 2113 19921 2119
rect 19895 2081 19921 2087
rect 22751 2113 22777 2119
rect 22751 2081 22777 2087
rect 23143 2113 23169 2119
rect 23305 2087 23311 2113
rect 23337 2087 23343 2113
rect 23143 2081 23169 2087
rect 1583 2057 1609 2063
rect 1583 2025 1609 2031
rect 1751 2057 1777 2063
rect 1751 2025 1777 2031
rect 5335 2057 5361 2063
rect 5335 2025 5361 2031
rect 5503 2057 5529 2063
rect 5503 2025 5529 2031
rect 6119 2057 6145 2063
rect 6119 2025 6145 2031
rect 6399 2057 6425 2063
rect 6399 2025 6425 2031
rect 9311 2057 9337 2063
rect 9311 2025 9337 2031
rect 9479 2057 9505 2063
rect 9479 2025 9505 2031
rect 11831 2057 11857 2063
rect 11831 2025 11857 2031
rect 11943 2057 11969 2063
rect 11943 2025 11969 2031
rect 13679 2057 13705 2063
rect 13679 2025 13705 2031
rect 14743 2057 14769 2063
rect 14743 2025 14769 2031
rect 19503 2057 19529 2063
rect 19503 2025 19529 2031
rect 19615 2057 19641 2063
rect 19615 2025 19641 2031
rect 23591 2057 23617 2063
rect 23591 2025 23617 2031
rect 24599 2057 24625 2063
rect 24599 2025 24625 2031
rect 25775 2057 25801 2063
rect 25775 2025 25801 2031
rect 26111 2057 26137 2063
rect 26111 2025 26137 2031
rect 26223 2057 26249 2063
rect 26223 2025 26249 2031
rect 26615 2057 26641 2063
rect 26615 2025 26641 2031
rect 336 1973 28392 1990
rect 336 1947 2233 1973
rect 2259 1947 2285 1973
rect 2311 1947 2337 1973
rect 2363 1947 12233 1973
rect 12259 1947 12285 1973
rect 12311 1947 12337 1973
rect 12363 1947 22233 1973
rect 22259 1947 22285 1973
rect 22311 1947 22337 1973
rect 22363 1947 28392 1973
rect 336 1930 28392 1947
rect 23255 1889 23281 1895
rect 23255 1857 23281 1863
rect 24879 1889 24905 1895
rect 24879 1857 24905 1863
rect 24991 1889 25017 1895
rect 24991 1857 25017 1863
rect 24151 1833 24177 1839
rect 17873 1807 17879 1833
rect 17905 1807 17911 1833
rect 18769 1807 18775 1833
rect 18801 1807 18807 1833
rect 19553 1807 19559 1833
rect 19585 1807 19591 1833
rect 20729 1807 20735 1833
rect 20761 1807 20767 1833
rect 20897 1807 20903 1833
rect 20929 1807 20935 1833
rect 21681 1807 21687 1833
rect 21713 1807 21719 1833
rect 22465 1807 22471 1833
rect 22497 1807 22503 1833
rect 24151 1801 24177 1807
rect 24599 1833 24625 1839
rect 24599 1801 24625 1807
rect 25383 1833 25409 1839
rect 25383 1801 25409 1807
rect 25831 1833 25857 1839
rect 25831 1801 25857 1807
rect 26111 1833 26137 1839
rect 27449 1807 27455 1833
rect 27481 1807 27487 1833
rect 26111 1801 26137 1807
rect 11719 1777 11745 1783
rect 11719 1745 11745 1751
rect 12279 1777 12305 1783
rect 12279 1745 12305 1751
rect 12559 1777 12585 1783
rect 13791 1777 13817 1783
rect 24431 1777 24457 1783
rect 13057 1751 13063 1777
rect 13089 1751 13095 1777
rect 16697 1751 16703 1777
rect 16729 1751 16735 1777
rect 12559 1745 12585 1751
rect 13791 1745 13817 1751
rect 24431 1745 24457 1751
rect 25663 1777 25689 1783
rect 26273 1751 26279 1777
rect 26305 1751 26311 1777
rect 27113 1751 27119 1777
rect 27145 1751 27151 1777
rect 25663 1745 25689 1751
rect 11551 1721 11577 1727
rect 11551 1689 11577 1695
rect 11999 1721 12025 1727
rect 11999 1689 12025 1695
rect 13287 1721 13313 1727
rect 13287 1689 13313 1695
rect 14071 1721 14097 1727
rect 14071 1689 14097 1695
rect 14687 1721 14713 1727
rect 14687 1689 14713 1695
rect 17151 1721 17177 1727
rect 17151 1689 17177 1695
rect 17991 1721 18017 1727
rect 21183 1721 21209 1727
rect 26783 1721 26809 1727
rect 19105 1695 19111 1721
rect 19137 1695 19143 1721
rect 20281 1695 20287 1721
rect 20313 1695 20319 1721
rect 22129 1695 22135 1721
rect 22161 1695 22167 1721
rect 22801 1695 22807 1721
rect 22833 1695 22839 1721
rect 23473 1695 23479 1721
rect 23505 1695 23511 1721
rect 17991 1689 18017 1695
rect 21183 1689 21209 1695
rect 26783 1689 26809 1695
rect 16311 1665 16337 1671
rect 16311 1633 16337 1639
rect 17375 1665 17401 1671
rect 17375 1633 17401 1639
rect 18271 1665 18297 1671
rect 18271 1633 18297 1639
rect 336 1581 28392 1598
rect 336 1555 1903 1581
rect 1929 1555 1955 1581
rect 1981 1555 2007 1581
rect 2033 1555 11903 1581
rect 11929 1555 11955 1581
rect 11981 1555 12007 1581
rect 12033 1555 21903 1581
rect 21929 1555 21955 1581
rect 21981 1555 22007 1581
rect 22033 1555 28392 1581
rect 336 1538 28392 1555
rect 27287 1497 27313 1503
rect 27287 1465 27313 1471
rect 28071 1497 28097 1503
rect 28071 1465 28097 1471
rect 7183 1441 7209 1447
rect 7183 1409 7209 1415
rect 14239 1441 14265 1447
rect 14239 1409 14265 1415
rect 19055 1441 19081 1447
rect 19055 1409 19081 1415
rect 20623 1441 20649 1447
rect 26503 1441 26529 1447
rect 22409 1415 22415 1441
rect 22441 1415 22447 1441
rect 20623 1409 20649 1415
rect 26503 1409 26529 1415
rect 14351 1385 14377 1391
rect 12609 1359 12615 1385
rect 12641 1359 12647 1385
rect 15241 1359 15247 1385
rect 15273 1359 15279 1385
rect 17425 1359 17431 1385
rect 17457 1359 17463 1385
rect 17649 1359 17655 1385
rect 17681 1359 17687 1385
rect 18153 1359 18159 1385
rect 18185 1359 18191 1385
rect 19441 1359 19447 1385
rect 19473 1359 19479 1385
rect 20337 1359 20343 1385
rect 20369 1359 20375 1385
rect 21065 1359 21071 1385
rect 21097 1359 21103 1385
rect 22073 1359 22079 1385
rect 22105 1359 22111 1385
rect 23641 1359 23647 1385
rect 23673 1359 23679 1385
rect 24481 1359 24487 1385
rect 24513 1359 24519 1385
rect 26777 1359 26783 1385
rect 26809 1359 26815 1385
rect 27561 1359 27567 1385
rect 27593 1359 27599 1385
rect 14351 1353 14377 1359
rect 8527 1329 8553 1335
rect 8527 1297 8553 1303
rect 8639 1329 8665 1335
rect 8639 1297 8665 1303
rect 8919 1329 8945 1335
rect 14631 1329 14657 1335
rect 13337 1303 13343 1329
rect 13369 1303 13375 1329
rect 8919 1297 8945 1303
rect 14631 1297 14657 1303
rect 15079 1329 15105 1335
rect 17879 1329 17905 1335
rect 21799 1329 21825 1335
rect 25719 1329 25745 1335
rect 16025 1303 16031 1329
rect 16057 1303 16063 1329
rect 17033 1303 17039 1329
rect 17065 1303 17071 1329
rect 18545 1303 18551 1329
rect 18577 1303 18583 1329
rect 19945 1303 19951 1329
rect 19977 1303 19983 1329
rect 22857 1303 22863 1329
rect 22889 1303 22895 1329
rect 25993 1303 25999 1329
rect 26025 1303 26031 1329
rect 15079 1297 15105 1303
rect 17879 1297 17905 1303
rect 21799 1297 21825 1303
rect 25719 1297 25745 1303
rect 6791 1273 6817 1279
rect 6791 1241 6817 1247
rect 6903 1273 6929 1279
rect 6903 1241 6929 1247
rect 12111 1273 12137 1279
rect 12111 1241 12137 1247
rect 12839 1273 12865 1279
rect 12839 1241 12865 1247
rect 13623 1273 13649 1279
rect 13623 1241 13649 1247
rect 14799 1273 14825 1279
rect 14799 1241 14825 1247
rect 15527 1273 15553 1279
rect 15527 1241 15553 1247
rect 16311 1273 16337 1279
rect 16311 1241 16337 1247
rect 21351 1273 21377 1279
rect 21351 1241 21377 1247
rect 21519 1273 21545 1279
rect 21519 1241 21545 1247
rect 23143 1273 23169 1279
rect 23143 1241 23169 1247
rect 23927 1273 23953 1279
rect 23927 1241 23953 1247
rect 24711 1273 24737 1279
rect 24711 1241 24737 1247
rect 25327 1273 25353 1279
rect 25327 1241 25353 1247
rect 25439 1273 25465 1279
rect 25439 1241 25465 1247
rect 336 1189 28392 1206
rect 336 1163 2233 1189
rect 2259 1163 2285 1189
rect 2311 1163 2337 1189
rect 2363 1163 12233 1189
rect 12259 1163 12285 1189
rect 12311 1163 12337 1189
rect 12363 1163 22233 1189
rect 22259 1163 22285 1189
rect 22311 1163 22337 1189
rect 22363 1163 28392 1189
rect 336 1146 28392 1163
rect 10263 1105 10289 1111
rect 10263 1073 10289 1079
rect 10431 1105 10457 1111
rect 10431 1073 10457 1079
rect 12391 1105 12417 1111
rect 12391 1073 12417 1079
rect 12559 1105 12585 1111
rect 12559 1073 12585 1079
rect 19335 1105 19361 1111
rect 19335 1073 19361 1079
rect 855 1049 881 1055
rect 855 1017 881 1023
rect 9871 1049 9897 1055
rect 9871 1017 9897 1023
rect 10711 1049 10737 1055
rect 10711 1017 10737 1023
rect 11215 1049 11241 1055
rect 15919 1049 15945 1055
rect 25607 1049 25633 1055
rect 11377 1023 11383 1049
rect 11409 1023 11415 1049
rect 13001 1023 13007 1049
rect 13033 1023 13039 1049
rect 14401 1023 14407 1049
rect 14433 1023 14439 1049
rect 15185 1023 15191 1049
rect 15217 1023 15223 1049
rect 16193 1023 16199 1049
rect 16225 1023 16231 1049
rect 17593 1023 17599 1049
rect 17625 1023 17631 1049
rect 22465 1023 22471 1049
rect 22497 1023 22503 1049
rect 24033 1023 24039 1049
rect 24065 1023 24071 1049
rect 24817 1023 24823 1049
rect 24849 1023 24855 1049
rect 27057 1023 27063 1049
rect 27089 1023 27095 1049
rect 27449 1023 27455 1049
rect 27481 1023 27487 1049
rect 11215 1017 11241 1023
rect 15919 1017 15945 1023
rect 25607 1017 25633 1023
rect 1135 993 1161 999
rect 1135 961 1161 967
rect 4775 993 4801 999
rect 4775 961 4801 967
rect 9591 993 9617 999
rect 9591 961 9617 967
rect 10935 993 10961 999
rect 10935 961 10961 967
rect 15639 993 15665 999
rect 19615 993 19641 999
rect 23535 993 23561 999
rect 18377 967 18383 993
rect 18409 967 18415 993
rect 19049 967 19055 993
rect 19081 967 19087 993
rect 20673 967 20679 993
rect 20705 967 20711 993
rect 21457 967 21463 993
rect 21489 967 21495 993
rect 21681 967 21687 993
rect 21713 967 21719 993
rect 15639 961 15665 967
rect 19615 961 19641 967
rect 23535 961 23561 967
rect 25887 993 25913 999
rect 26329 967 26335 993
rect 26361 967 26367 993
rect 25887 961 25913 967
rect 1247 937 1273 943
rect 1247 905 1273 911
rect 4607 937 4633 943
rect 9423 937 9449 943
rect 4993 911 4999 937
rect 5025 911 5031 937
rect 4607 905 4633 911
rect 9423 905 9449 911
rect 12839 937 12865 943
rect 15471 937 15497 943
rect 14009 911 14015 937
rect 14041 911 14047 937
rect 12839 905 12865 911
rect 15471 905 15497 911
rect 22751 937 22777 943
rect 23647 937 23673 943
rect 25999 937 26025 943
rect 23305 911 23311 937
rect 23337 911 23343 937
rect 24369 911 24375 937
rect 24401 911 24407 937
rect 25265 911 25271 937
rect 25297 911 25303 937
rect 22751 905 22777 911
rect 23647 905 23673 911
rect 25999 905 26025 911
rect 26783 937 26809 943
rect 26783 905 26809 911
rect 11887 881 11913 887
rect 11887 849 11913 855
rect 13511 881 13537 887
rect 13511 849 13537 855
rect 14687 881 14713 887
rect 14687 849 14713 855
rect 16479 881 16505 887
rect 16479 849 16505 855
rect 17095 881 17121 887
rect 17095 849 17121 855
rect 17879 881 17905 887
rect 17879 849 17905 855
rect 18663 881 18689 887
rect 18663 849 18689 855
rect 20231 881 20257 887
rect 20231 849 20257 855
rect 21015 881 21041 887
rect 21015 849 21041 855
rect 21967 881 21993 887
rect 21967 849 21993 855
rect 336 797 28392 814
rect 336 771 1903 797
rect 1929 771 1955 797
rect 1981 771 2007 797
rect 2033 771 11903 797
rect 11929 771 11955 797
rect 11981 771 12007 797
rect 12033 771 21903 797
rect 21929 771 21955 797
rect 21981 771 22007 797
rect 22033 771 28392 797
rect 336 754 28392 771
rect 26783 713 26809 719
rect 26783 681 26809 687
rect 28071 713 28097 719
rect 28071 681 28097 687
rect 10767 657 10793 663
rect 10767 625 10793 631
rect 13455 657 13481 663
rect 13455 625 13481 631
rect 19167 657 19193 663
rect 19167 625 19193 631
rect 20455 657 20481 663
rect 20455 625 20481 631
rect 25999 657 26025 663
rect 25999 625 26025 631
rect 11041 575 11047 601
rect 11073 575 11079 601
rect 12161 575 12167 601
rect 12193 575 12199 601
rect 13057 575 13063 601
rect 13089 575 13095 601
rect 14625 575 14631 601
rect 14657 575 14663 601
rect 14849 575 14855 601
rect 14881 575 14887 601
rect 15745 575 15751 601
rect 15777 575 15783 601
rect 16529 575 16535 601
rect 16561 575 16567 601
rect 17649 575 17655 601
rect 17681 575 17687 601
rect 18545 575 18551 601
rect 18577 575 18583 601
rect 20057 575 20063 601
rect 20089 575 20095 601
rect 20953 575 20959 601
rect 20985 575 20991 601
rect 22073 575 22079 601
rect 22105 575 22111 601
rect 22241 575 22247 601
rect 22273 575 22279 601
rect 24145 575 24151 601
rect 24177 575 24183 601
rect 25489 575 25495 601
rect 25521 575 25527 601
rect 26385 575 26391 601
rect 26417 575 26423 601
rect 11433 519 11439 545
rect 11465 519 11471 545
rect 12553 519 12559 545
rect 12585 519 12591 545
rect 14233 519 14239 545
rect 14265 519 14271 545
rect 19777 519 19783 545
rect 19809 519 19815 545
rect 21681 519 21687 545
rect 21713 519 21719 545
rect 23361 519 23367 545
rect 23393 519 23399 545
rect 27561 519 27567 545
rect 27593 519 27599 545
rect 15079 489 15105 495
rect 15079 457 15105 463
rect 16031 489 16057 495
rect 16031 457 16057 463
rect 16815 489 16841 495
rect 16815 457 16841 463
rect 17935 489 17961 495
rect 17935 457 17961 463
rect 18719 489 18745 495
rect 18719 457 18745 463
rect 22527 489 22553 495
rect 22527 457 22553 463
rect 23647 489 23673 495
rect 23647 457 23673 463
rect 24431 489 24457 495
rect 24431 457 24457 463
rect 336 405 28392 422
rect 336 379 2233 405
rect 2259 379 2285 405
rect 2311 379 2337 405
rect 2363 379 12233 405
rect 12259 379 12285 405
rect 12311 379 12337 405
rect 12363 379 22233 405
rect 22259 379 22285 405
rect 22311 379 22337 405
rect 22363 379 28392 405
rect 336 362 28392 379
<< via1 >>
rect 2233 6651 2259 6677
rect 2285 6651 2311 6677
rect 2337 6651 2363 6677
rect 12233 6651 12259 6677
rect 12285 6651 12311 6677
rect 12337 6651 12363 6677
rect 22233 6651 22259 6677
rect 22285 6651 22311 6677
rect 22337 6651 22363 6677
rect 1023 6567 1049 6593
rect 5335 6567 5361 6593
rect 26559 6567 26585 6593
rect 4047 6511 4073 6537
rect 1191 6455 1217 6481
rect 3039 6455 3065 6481
rect 5167 6455 5193 6481
rect 7015 6455 7041 6481
rect 9703 6455 9729 6481
rect 11047 6455 11073 6481
rect 12559 6455 12585 6481
rect 13567 6455 13593 6481
rect 15079 6455 15105 6481
rect 16423 6455 16449 6481
rect 19111 6455 19137 6481
rect 20455 6455 20481 6481
rect 22079 6455 22105 6481
rect 23087 6455 23113 6481
rect 24487 6455 24513 6481
rect 25887 6455 25913 6481
rect 26279 6455 26305 6481
rect 27679 6455 27705 6481
rect 2535 6399 2561 6425
rect 3599 6399 3625 6425
rect 6511 6399 6537 6425
rect 9199 6399 9225 6425
rect 10543 6399 10569 6425
rect 12055 6399 12081 6425
rect 13063 6399 13089 6425
rect 14575 6399 14601 6425
rect 15919 6399 15945 6425
rect 18607 6399 18633 6425
rect 19951 6399 19977 6425
rect 21575 6399 21601 6425
rect 22583 6399 22609 6425
rect 23983 6399 24009 6425
rect 25383 6399 25409 6425
rect 28071 6343 28097 6369
rect 1903 6259 1929 6285
rect 1955 6259 1981 6285
rect 2007 6259 2033 6285
rect 11903 6259 11929 6285
rect 11955 6259 11981 6285
rect 12007 6259 12033 6285
rect 21903 6259 21929 6285
rect 21955 6259 21981 6285
rect 22007 6259 22033 6285
rect 7855 6175 7881 6201
rect 17263 6175 17289 6201
rect 26503 6175 26529 6201
rect 5223 6119 5249 6145
rect 5671 6119 5697 6145
rect 7519 6119 7545 6145
rect 10319 6119 10345 6145
rect 10767 6119 10793 6145
rect 11159 6119 11185 6145
rect 11551 6119 11577 6145
rect 13063 6119 13089 6145
rect 13231 6119 13257 6145
rect 16087 6119 16113 6145
rect 16423 6119 16449 6145
rect 19951 6119 19977 6145
rect 23255 6119 23281 6145
rect 24991 6119 25017 6145
rect 5503 6063 5529 6089
rect 10599 6063 10625 6089
rect 11719 6063 11745 6089
rect 14015 6063 14041 6089
rect 14239 6063 14265 6089
rect 14519 6063 14545 6089
rect 16199 6063 16225 6089
rect 23423 6063 23449 6089
rect 26111 6063 26137 6089
rect 26783 6063 26809 6089
rect 8359 6007 8385 6033
rect 11999 6007 12025 6033
rect 15359 6007 15385 6033
rect 17767 6007 17793 6033
rect 18551 6007 18577 6033
rect 20231 6007 20257 6033
rect 20399 6007 20425 6033
rect 23703 6007 23729 6033
rect 27175 6007 27201 6033
rect 27567 6007 27593 6033
rect 27959 6007 27985 6033
rect 7183 5951 7209 5977
rect 7295 5951 7321 5977
rect 11439 5951 11465 5977
rect 12671 5951 12697 5977
rect 12783 5951 12809 5977
rect 13511 5951 13537 5977
rect 13679 5951 13705 5977
rect 14967 5951 14993 5977
rect 15079 5951 15105 5977
rect 18831 5951 18857 5977
rect 18999 5951 19025 5977
rect 22303 5951 22329 5977
rect 22471 5951 22497 5977
rect 22639 5951 22665 5977
rect 24655 5951 24681 5977
rect 24767 5951 24793 5977
rect 2233 5867 2259 5893
rect 2285 5867 2311 5893
rect 2337 5867 2363 5893
rect 12233 5867 12259 5893
rect 12285 5867 12311 5893
rect 12337 5867 12363 5893
rect 22233 5867 22259 5893
rect 22285 5867 22311 5893
rect 22337 5867 22363 5893
rect 7407 5783 7433 5809
rect 7519 5783 7545 5809
rect 7127 5727 7153 5753
rect 9087 5727 9113 5753
rect 25495 5727 25521 5753
rect 25887 5727 25913 5753
rect 9367 5671 9393 5697
rect 9479 5671 9505 5697
rect 12279 5671 12305 5697
rect 17543 5671 17569 5697
rect 23759 5671 23785 5697
rect 26391 5671 26417 5697
rect 27063 5671 27089 5697
rect 11551 5615 11577 5641
rect 11999 5615 12025 5641
rect 12559 5615 12585 5641
rect 17375 5615 17401 5641
rect 17823 5615 17849 5641
rect 23535 5615 23561 5641
rect 23983 5615 24009 5641
rect 26783 5559 26809 5585
rect 27567 5559 27593 5585
rect 1903 5475 1929 5501
rect 1955 5475 1981 5501
rect 2007 5475 2033 5501
rect 11903 5475 11929 5501
rect 11955 5475 11981 5501
rect 12007 5475 12033 5501
rect 21903 5475 21929 5501
rect 21955 5475 21981 5501
rect 22007 5475 22033 5501
rect 26503 5391 26529 5417
rect 14351 5335 14377 5361
rect 14799 5335 14825 5361
rect 17095 5335 17121 5361
rect 27287 5335 27313 5361
rect 28071 5335 28097 5361
rect 14631 5279 14657 5305
rect 17263 5279 17289 5305
rect 19279 5279 19305 5305
rect 26055 5279 26081 5305
rect 27623 5279 27649 5305
rect 15695 5223 15721 5249
rect 17543 5223 17569 5249
rect 26783 5223 26809 5249
rect 15247 5167 15273 5193
rect 15415 5167 15441 5193
rect 18831 5167 18857 5193
rect 18999 5167 19025 5193
rect 2233 5083 2259 5109
rect 2285 5083 2311 5109
rect 2337 5083 2363 5109
rect 12233 5083 12259 5109
rect 12285 5083 12311 5109
rect 12337 5083 12363 5109
rect 22233 5083 22259 5109
rect 22285 5083 22311 5109
rect 22337 5083 22363 5109
rect 9535 4999 9561 5025
rect 9703 4999 9729 5025
rect 17207 4999 17233 5025
rect 17319 4999 17345 5025
rect 16311 4943 16337 4969
rect 17599 4943 17625 4969
rect 26279 4943 26305 4969
rect 16591 4887 16617 4913
rect 27063 4887 27089 4913
rect 9983 4831 10009 4857
rect 16703 4831 16729 4857
rect 26783 4831 26809 4857
rect 27567 4775 27593 4801
rect 1903 4691 1929 4717
rect 1955 4691 1981 4717
rect 2007 4691 2033 4717
rect 11903 4691 11929 4717
rect 11955 4691 11981 4717
rect 12007 4691 12033 4717
rect 21903 4691 21929 4717
rect 21955 4691 21981 4717
rect 22007 4691 22033 4717
rect 11159 4551 11185 4577
rect 12615 4551 12641 4577
rect 13063 4551 13089 4577
rect 14015 4551 14041 4577
rect 14463 4551 14489 4577
rect 11327 4495 11353 4521
rect 11607 4495 11633 4521
rect 12783 4495 12809 4521
rect 14239 4495 14265 4521
rect 27623 4495 27649 4521
rect 1471 4439 1497 4465
rect 20455 4439 20481 4465
rect 20567 4439 20593 4465
rect 20847 4439 20873 4465
rect 22359 4439 22385 4465
rect 26783 4439 26809 4465
rect 27175 4439 27201 4465
rect 27959 4439 27985 4465
rect 1079 4383 1105 4409
rect 1191 4383 1217 4409
rect 21855 4383 21881 4409
rect 22079 4383 22105 4409
rect 2233 4299 2259 4325
rect 2285 4299 2311 4325
rect 2337 4299 2363 4325
rect 12233 4299 12259 4325
rect 12285 4299 12311 4325
rect 12337 4299 12363 4325
rect 22233 4299 22259 4325
rect 22285 4299 22311 4325
rect 22337 4299 22363 4325
rect 11103 4159 11129 4185
rect 11215 4159 11241 4185
rect 11495 4159 11521 4185
rect 27455 4159 27481 4185
rect 9143 4103 9169 4129
rect 14631 4103 14657 4129
rect 15359 4103 15385 4129
rect 21799 4103 21825 4129
rect 27063 4103 27089 4129
rect 8919 4047 8945 4073
rect 9255 4047 9281 4073
rect 14519 4047 14545 4073
rect 14911 4047 14937 4073
rect 15191 4047 15217 4073
rect 15583 4047 15609 4073
rect 21631 4047 21657 4073
rect 22079 4047 22105 4073
rect 1903 3907 1929 3933
rect 1955 3907 1981 3933
rect 2007 3907 2033 3933
rect 11903 3907 11929 3933
rect 11955 3907 11981 3933
rect 12007 3907 12033 3933
rect 21903 3907 21929 3933
rect 21955 3907 21981 3933
rect 22007 3907 22033 3933
rect 28071 3823 28097 3849
rect 13175 3767 13201 3793
rect 17375 3767 17401 3793
rect 17823 3767 17849 3793
rect 27287 3767 27313 3793
rect 12839 3711 12865 3737
rect 12951 3711 12977 3737
rect 17543 3711 17569 3737
rect 26783 3711 26809 3737
rect 27567 3711 27593 3737
rect 2703 3655 2729 3681
rect 4551 3655 4577 3681
rect 10711 3655 10737 3681
rect 2983 3599 3009 3625
rect 3151 3599 3177 3625
rect 4831 3599 4857 3625
rect 4999 3599 5025 3625
rect 10263 3599 10289 3625
rect 10431 3599 10457 3625
rect 2233 3515 2259 3541
rect 2285 3515 2311 3541
rect 2337 3515 2363 3541
rect 12233 3515 12259 3541
rect 12285 3515 12311 3541
rect 12337 3515 12363 3541
rect 22233 3515 22259 3541
rect 22285 3515 22311 3541
rect 22337 3515 22363 3541
rect 7799 3319 7825 3345
rect 13231 3319 13257 3345
rect 21631 3319 21657 3345
rect 22415 3319 22441 3345
rect 22695 3319 22721 3345
rect 27063 3319 27089 3345
rect 7631 3263 7657 3289
rect 8079 3263 8105 3289
rect 13063 3263 13089 3289
rect 13511 3263 13537 3289
rect 21463 3263 21489 3289
rect 21855 3263 21881 3289
rect 22247 3263 22273 3289
rect 27567 3207 27593 3233
rect 1903 3123 1929 3149
rect 1955 3123 1981 3149
rect 2007 3123 2033 3149
rect 11903 3123 11929 3149
rect 11955 3123 11981 3149
rect 12007 3123 12033 3149
rect 21903 3123 21929 3149
rect 21955 3123 21981 3149
rect 22007 3123 22033 3149
rect 28071 3039 28097 3065
rect 12671 2983 12697 3009
rect 17487 2983 17513 3009
rect 17823 2983 17849 3009
rect 18551 2983 18577 3009
rect 23199 2983 23225 3009
rect 26503 2983 26529 3009
rect 27287 2983 27313 3009
rect 12447 2927 12473 2953
rect 17599 2927 17625 2953
rect 18663 2927 18689 2953
rect 23311 2927 23337 2953
rect 24599 2927 24625 2953
rect 24711 2927 24737 2953
rect 26783 2927 26809 2953
rect 27567 2927 27593 2953
rect 7127 2871 7153 2897
rect 8191 2871 8217 2897
rect 8303 2871 8329 2897
rect 8583 2871 8609 2897
rect 12223 2871 12249 2897
rect 18943 2871 18969 2897
rect 20287 2871 20313 2897
rect 23591 2871 23617 2897
rect 24991 2871 25017 2897
rect 7407 2815 7433 2841
rect 7575 2815 7601 2841
rect 11831 2815 11857 2841
rect 11943 2815 11969 2841
rect 19895 2815 19921 2841
rect 20007 2815 20033 2841
rect 26615 2815 26641 2841
rect 2233 2731 2259 2757
rect 2285 2731 2311 2757
rect 2337 2731 2363 2757
rect 12233 2731 12259 2757
rect 12285 2731 12311 2757
rect 12337 2731 12363 2757
rect 22233 2731 22259 2757
rect 22285 2731 22311 2757
rect 22337 2731 22363 2757
rect 9143 2647 9169 2673
rect 9311 2647 9337 2673
rect 14295 2647 14321 2673
rect 14463 2647 14489 2673
rect 17151 2647 17177 2673
rect 17319 2647 17345 2673
rect 21127 2647 21153 2673
rect 21295 2647 21321 2673
rect 23311 2647 23337 2673
rect 23479 2647 23505 2673
rect 5167 2591 5193 2617
rect 9759 2591 9785 2617
rect 14911 2591 14937 2617
rect 16479 2591 16505 2617
rect 17599 2591 17625 2617
rect 23759 2591 23785 2617
rect 26167 2591 26193 2617
rect 26447 2591 26473 2617
rect 27063 2591 27089 2617
rect 5447 2535 5473 2561
rect 5559 2535 5585 2561
rect 10039 2535 10065 2561
rect 10151 2535 10177 2561
rect 12223 2535 12249 2561
rect 15191 2535 15217 2561
rect 15975 2535 16001 2561
rect 16199 2535 16225 2561
rect 19111 2535 19137 2561
rect 19279 2535 19305 2561
rect 19559 2535 19585 2561
rect 26615 2535 26641 2561
rect 27455 2535 27481 2561
rect 9591 2479 9617 2505
rect 14743 2479 14769 2505
rect 21575 2479 21601 2505
rect 26895 2479 26921 2505
rect 1903 2339 1929 2365
rect 1955 2339 1981 2365
rect 2007 2339 2033 2365
rect 11903 2339 11929 2365
rect 11955 2339 11981 2365
rect 12007 2339 12033 2365
rect 21903 2339 21929 2365
rect 21955 2339 21981 2365
rect 22007 2339 22033 2365
rect 27287 2255 27313 2281
rect 28071 2255 28097 2281
rect 5111 2199 5137 2225
rect 5895 2199 5921 2225
rect 12167 2199 12193 2225
rect 16143 2199 16169 2225
rect 17487 2199 17513 2225
rect 20623 2199 20649 2225
rect 20959 2199 20985 2225
rect 26335 2199 26361 2225
rect 16255 2143 16281 2169
rect 17599 2143 17625 2169
rect 18159 2143 18185 2169
rect 20735 2143 20761 2169
rect 22359 2143 22385 2169
rect 22471 2143 22497 2169
rect 26783 2143 26809 2169
rect 27567 2143 27593 2169
rect 1303 2087 1329 2113
rect 9031 2087 9057 2113
rect 16535 2087 16561 2113
rect 17879 2087 17905 2113
rect 18439 2087 18465 2113
rect 19895 2087 19921 2113
rect 22751 2087 22777 2113
rect 23143 2087 23169 2113
rect 23311 2087 23337 2113
rect 1583 2031 1609 2057
rect 1751 2031 1777 2057
rect 5335 2031 5361 2057
rect 5503 2031 5529 2057
rect 6119 2031 6145 2057
rect 6399 2031 6425 2057
rect 9311 2031 9337 2057
rect 9479 2031 9505 2057
rect 11831 2031 11857 2057
rect 11943 2031 11969 2057
rect 13679 2031 13705 2057
rect 14743 2031 14769 2057
rect 19503 2031 19529 2057
rect 19615 2031 19641 2057
rect 23591 2031 23617 2057
rect 24599 2031 24625 2057
rect 25775 2031 25801 2057
rect 26111 2031 26137 2057
rect 26223 2031 26249 2057
rect 26615 2031 26641 2057
rect 2233 1947 2259 1973
rect 2285 1947 2311 1973
rect 2337 1947 2363 1973
rect 12233 1947 12259 1973
rect 12285 1947 12311 1973
rect 12337 1947 12363 1973
rect 22233 1947 22259 1973
rect 22285 1947 22311 1973
rect 22337 1947 22363 1973
rect 23255 1863 23281 1889
rect 24879 1863 24905 1889
rect 24991 1863 25017 1889
rect 17879 1807 17905 1833
rect 18775 1807 18801 1833
rect 19559 1807 19585 1833
rect 20735 1807 20761 1833
rect 20903 1807 20929 1833
rect 21687 1807 21713 1833
rect 22471 1807 22497 1833
rect 24151 1807 24177 1833
rect 24599 1807 24625 1833
rect 25383 1807 25409 1833
rect 25831 1807 25857 1833
rect 26111 1807 26137 1833
rect 27455 1807 27481 1833
rect 11719 1751 11745 1777
rect 12279 1751 12305 1777
rect 12559 1751 12585 1777
rect 13063 1751 13089 1777
rect 13791 1751 13817 1777
rect 16703 1751 16729 1777
rect 24431 1751 24457 1777
rect 25663 1751 25689 1777
rect 26279 1751 26305 1777
rect 27119 1751 27145 1777
rect 11551 1695 11577 1721
rect 11999 1695 12025 1721
rect 13287 1695 13313 1721
rect 14071 1695 14097 1721
rect 14687 1695 14713 1721
rect 17151 1695 17177 1721
rect 17991 1695 18017 1721
rect 19111 1695 19137 1721
rect 20287 1695 20313 1721
rect 21183 1695 21209 1721
rect 22135 1695 22161 1721
rect 22807 1695 22833 1721
rect 23479 1695 23505 1721
rect 26783 1695 26809 1721
rect 16311 1639 16337 1665
rect 17375 1639 17401 1665
rect 18271 1639 18297 1665
rect 1903 1555 1929 1581
rect 1955 1555 1981 1581
rect 2007 1555 2033 1581
rect 11903 1555 11929 1581
rect 11955 1555 11981 1581
rect 12007 1555 12033 1581
rect 21903 1555 21929 1581
rect 21955 1555 21981 1581
rect 22007 1555 22033 1581
rect 27287 1471 27313 1497
rect 28071 1471 28097 1497
rect 7183 1415 7209 1441
rect 14239 1415 14265 1441
rect 19055 1415 19081 1441
rect 20623 1415 20649 1441
rect 22415 1415 22441 1441
rect 26503 1415 26529 1441
rect 12615 1359 12641 1385
rect 14351 1359 14377 1385
rect 15247 1359 15273 1385
rect 17431 1359 17457 1385
rect 17655 1359 17681 1385
rect 18159 1359 18185 1385
rect 19447 1359 19473 1385
rect 20343 1359 20369 1385
rect 21071 1359 21097 1385
rect 22079 1359 22105 1385
rect 23647 1359 23673 1385
rect 24487 1359 24513 1385
rect 26783 1359 26809 1385
rect 27567 1359 27593 1385
rect 8527 1303 8553 1329
rect 8639 1303 8665 1329
rect 8919 1303 8945 1329
rect 13343 1303 13369 1329
rect 14631 1303 14657 1329
rect 15079 1303 15105 1329
rect 16031 1303 16057 1329
rect 17039 1303 17065 1329
rect 17879 1303 17905 1329
rect 18551 1303 18577 1329
rect 19951 1303 19977 1329
rect 21799 1303 21825 1329
rect 22863 1303 22889 1329
rect 25719 1303 25745 1329
rect 25999 1303 26025 1329
rect 6791 1247 6817 1273
rect 6903 1247 6929 1273
rect 12111 1247 12137 1273
rect 12839 1247 12865 1273
rect 13623 1247 13649 1273
rect 14799 1247 14825 1273
rect 15527 1247 15553 1273
rect 16311 1247 16337 1273
rect 21351 1247 21377 1273
rect 21519 1247 21545 1273
rect 23143 1247 23169 1273
rect 23927 1247 23953 1273
rect 24711 1247 24737 1273
rect 25327 1247 25353 1273
rect 25439 1247 25465 1273
rect 2233 1163 2259 1189
rect 2285 1163 2311 1189
rect 2337 1163 2363 1189
rect 12233 1163 12259 1189
rect 12285 1163 12311 1189
rect 12337 1163 12363 1189
rect 22233 1163 22259 1189
rect 22285 1163 22311 1189
rect 22337 1163 22363 1189
rect 10263 1079 10289 1105
rect 10431 1079 10457 1105
rect 12391 1079 12417 1105
rect 12559 1079 12585 1105
rect 19335 1079 19361 1105
rect 855 1023 881 1049
rect 9871 1023 9897 1049
rect 10711 1023 10737 1049
rect 11215 1023 11241 1049
rect 11383 1023 11409 1049
rect 13007 1023 13033 1049
rect 14407 1023 14433 1049
rect 15191 1023 15217 1049
rect 15919 1023 15945 1049
rect 16199 1023 16225 1049
rect 17599 1023 17625 1049
rect 22471 1023 22497 1049
rect 24039 1023 24065 1049
rect 24823 1023 24849 1049
rect 25607 1023 25633 1049
rect 27063 1023 27089 1049
rect 27455 1023 27481 1049
rect 1135 967 1161 993
rect 4775 967 4801 993
rect 9591 967 9617 993
rect 10935 967 10961 993
rect 15639 967 15665 993
rect 18383 967 18409 993
rect 19055 967 19081 993
rect 19615 967 19641 993
rect 20679 967 20705 993
rect 21463 967 21489 993
rect 21687 967 21713 993
rect 23535 967 23561 993
rect 25887 967 25913 993
rect 26335 967 26361 993
rect 1247 911 1273 937
rect 4607 911 4633 937
rect 4999 911 5025 937
rect 9423 911 9449 937
rect 12839 911 12865 937
rect 14015 911 14041 937
rect 15471 911 15497 937
rect 22751 911 22777 937
rect 23311 911 23337 937
rect 23647 911 23673 937
rect 24375 911 24401 937
rect 25271 911 25297 937
rect 25999 911 26025 937
rect 26783 911 26809 937
rect 11887 855 11913 881
rect 13511 855 13537 881
rect 14687 855 14713 881
rect 16479 855 16505 881
rect 17095 855 17121 881
rect 17879 855 17905 881
rect 18663 855 18689 881
rect 20231 855 20257 881
rect 21015 855 21041 881
rect 21967 855 21993 881
rect 1903 771 1929 797
rect 1955 771 1981 797
rect 2007 771 2033 797
rect 11903 771 11929 797
rect 11955 771 11981 797
rect 12007 771 12033 797
rect 21903 771 21929 797
rect 21955 771 21981 797
rect 22007 771 22033 797
rect 26783 687 26809 713
rect 28071 687 28097 713
rect 10767 631 10793 657
rect 13455 631 13481 657
rect 19167 631 19193 657
rect 20455 631 20481 657
rect 25999 631 26025 657
rect 11047 575 11073 601
rect 12167 575 12193 601
rect 13063 575 13089 601
rect 14631 575 14657 601
rect 14855 575 14881 601
rect 15751 575 15777 601
rect 16535 575 16561 601
rect 17655 575 17681 601
rect 18551 575 18577 601
rect 20063 575 20089 601
rect 20959 575 20985 601
rect 22079 575 22105 601
rect 22247 575 22273 601
rect 24151 575 24177 601
rect 25495 575 25521 601
rect 26391 575 26417 601
rect 11439 519 11465 545
rect 12559 519 12585 545
rect 14239 519 14265 545
rect 19783 519 19809 545
rect 21687 519 21713 545
rect 23367 519 23393 545
rect 27567 519 27593 545
rect 15079 463 15105 489
rect 16031 463 16057 489
rect 16815 463 16841 489
rect 17935 463 17961 489
rect 18719 463 18745 489
rect 22527 463 22553 489
rect 23647 463 23673 489
rect 24431 463 24457 489
rect 2233 379 2259 405
rect 2285 379 2311 405
rect 2337 379 2363 405
rect 12233 379 12259 405
rect 12285 379 12311 405
rect 12337 379 12363 405
rect 22233 379 22259 405
rect 22285 379 22311 405
rect 22337 379 22363 405
<< metal2 >>
rect 896 7056 952 7112
rect 2240 7056 2296 7112
rect 3584 7056 3640 7112
rect 4928 7056 4984 7112
rect 6272 7056 6328 7112
rect 7616 7056 7672 7112
rect 8960 7056 9016 7112
rect 10304 7056 10360 7112
rect 11648 7056 11704 7112
rect 12992 7056 13048 7112
rect 14336 7056 14392 7112
rect 15680 7056 15736 7112
rect 17024 7056 17080 7112
rect 18368 7056 18424 7112
rect 19712 7056 19768 7112
rect 21056 7056 21112 7112
rect 22400 7056 22456 7112
rect 23744 7056 23800 7112
rect 25088 7056 25144 7112
rect 26432 7056 26488 7112
rect 27776 7056 27832 7112
rect 910 6818 938 7056
rect 2254 7042 2282 7056
rect 2254 7009 2282 7014
rect 2534 7042 2562 7047
rect 910 6790 1050 6818
rect 1022 6593 1050 6790
rect 2232 6678 2364 6683
rect 2260 6650 2284 6678
rect 2312 6650 2336 6678
rect 2232 6645 2364 6650
rect 1022 6567 1023 6593
rect 1049 6567 1050 6593
rect 1022 6561 1050 6567
rect 798 6538 826 6543
rect 406 6090 434 6095
rect 406 5250 434 6062
rect 798 5306 826 6510
rect 1190 6481 1218 6487
rect 1190 6455 1191 6481
rect 1217 6455 1218 6481
rect 1190 5586 1218 6455
rect 2534 6425 2562 7014
rect 3542 6986 3570 6991
rect 2534 6399 2535 6425
rect 2561 6399 2562 6425
rect 2534 6393 2562 6399
rect 3038 6481 3066 6487
rect 3038 6455 3039 6481
rect 3065 6455 3066 6481
rect 1902 6286 2034 6291
rect 1930 6258 1954 6286
rect 1982 6258 2006 6286
rect 1902 6253 2034 6258
rect 2232 5894 2364 5899
rect 2260 5866 2284 5894
rect 2312 5866 2336 5894
rect 2232 5861 2364 5866
rect 3038 5754 3066 6455
rect 3486 6482 3514 6487
rect 3374 6202 3402 6207
rect 3374 5866 3402 6174
rect 3374 5833 3402 5838
rect 3430 6034 3458 6039
rect 3038 5721 3066 5726
rect 1190 5553 1218 5558
rect 3374 5642 3402 5647
rect 2926 5530 2954 5535
rect 1902 5502 2034 5507
rect 1930 5474 1954 5502
rect 1982 5474 2006 5502
rect 1902 5469 2034 5474
rect 798 5273 826 5278
rect 406 5217 434 5222
rect 798 5194 826 5199
rect 574 4970 602 4975
rect 294 4186 322 4191
rect 70 2730 98 2735
rect 98 2702 154 2730
rect 70 2697 98 2702
rect 126 1666 154 2702
rect 126 1633 154 1638
rect 294 490 322 4158
rect 574 3738 602 4942
rect 574 3705 602 3710
rect 742 4634 770 4639
rect 742 3402 770 4606
rect 798 4578 826 5166
rect 2232 5110 2364 5115
rect 2260 5082 2284 5110
rect 2312 5082 2336 5110
rect 2232 5077 2364 5082
rect 2086 4858 2114 4863
rect 1902 4718 2034 4723
rect 1930 4690 1954 4718
rect 1982 4690 2006 4718
rect 1902 4685 2034 4690
rect 798 4545 826 4550
rect 1470 4466 1498 4471
rect 1470 4419 1498 4438
rect 742 3369 770 3374
rect 1078 4410 1106 4415
rect 1190 4410 1218 4415
rect 1078 4409 1218 4410
rect 1078 4383 1079 4409
rect 1105 4383 1191 4409
rect 1217 4383 1218 4409
rect 1078 4382 1218 4383
rect 294 457 322 462
rect 350 2898 378 2903
rect 350 56 378 2870
rect 1022 2842 1050 2847
rect 518 2562 546 2567
rect 518 1386 546 2534
rect 518 1353 546 1358
rect 798 1330 826 1335
rect 574 826 602 831
rect 462 490 490 495
rect 336 0 392 56
rect 462 42 490 462
rect 574 56 602 798
rect 798 56 826 1302
rect 854 1050 882 1055
rect 854 1003 882 1022
rect 1022 56 1050 2814
rect 1078 938 1106 4382
rect 1190 4377 1218 4382
rect 1806 4018 1834 4023
rect 1358 3010 1386 3015
rect 1302 2113 1330 2119
rect 1302 2087 1303 2113
rect 1329 2087 1330 2113
rect 1302 1890 1330 2087
rect 1302 1857 1330 1862
rect 1078 905 1106 910
rect 1134 993 1162 999
rect 1134 967 1135 993
rect 1161 967 1162 993
rect 1134 938 1162 967
rect 1246 938 1274 943
rect 1134 937 1274 938
rect 1134 911 1247 937
rect 1273 911 1274 937
rect 1134 910 1274 911
rect 1134 98 1162 910
rect 1246 905 1274 910
rect 1358 826 1386 2982
rect 1134 65 1162 70
rect 1246 798 1386 826
rect 1470 2170 1498 2175
rect 1246 56 1274 798
rect 1470 56 1498 2142
rect 1582 2058 1610 2063
rect 1750 2058 1778 2063
rect 1582 2057 1778 2058
rect 1582 2031 1583 2057
rect 1609 2031 1751 2057
rect 1777 2031 1778 2057
rect 1582 2030 1778 2031
rect 1582 2025 1610 2030
rect 1750 1778 1778 2030
rect 1750 1745 1778 1750
rect 1806 1666 1834 3990
rect 1902 3934 2034 3939
rect 1930 3906 1954 3934
rect 1982 3906 2006 3934
rect 1902 3901 2034 3906
rect 1902 3150 2034 3155
rect 1930 3122 1954 3150
rect 1982 3122 2006 3150
rect 1902 3117 2034 3122
rect 1902 2366 2034 2371
rect 1930 2338 1954 2366
rect 1982 2338 2006 2366
rect 1902 2333 2034 2338
rect 1694 1638 1834 1666
rect 1694 56 1722 1638
rect 1902 1582 2034 1587
rect 1930 1554 1954 1582
rect 1982 1554 2006 1582
rect 1902 1549 2034 1554
rect 1902 798 2034 803
rect 1930 770 1954 798
rect 1982 770 2006 798
rect 1902 765 2034 770
rect 2086 714 2114 4830
rect 2232 4326 2364 4331
rect 2260 4298 2284 4326
rect 2312 4298 2336 4326
rect 2232 4293 2364 4298
rect 2702 3681 2730 3687
rect 2702 3655 2703 3681
rect 2729 3655 2730 3681
rect 2702 3570 2730 3655
rect 2232 3542 2364 3547
rect 2260 3514 2284 3542
rect 2312 3514 2336 3542
rect 2702 3537 2730 3542
rect 2232 3509 2364 3514
rect 2232 2758 2364 2763
rect 2260 2730 2284 2758
rect 2312 2730 2336 2758
rect 2232 2725 2364 2730
rect 2814 2002 2842 2007
rect 2232 1974 2364 1979
rect 2260 1946 2284 1974
rect 2312 1946 2336 1974
rect 2232 1941 2364 1946
rect 2232 1190 2364 1195
rect 2260 1162 2284 1190
rect 2312 1162 2336 1190
rect 2232 1157 2364 1162
rect 2590 826 2618 831
rect 1918 686 2114 714
rect 2142 770 2170 775
rect 1918 56 1946 686
rect 2142 56 2170 742
rect 2232 406 2364 411
rect 2260 378 2284 406
rect 2312 378 2336 406
rect 2232 373 2364 378
rect 2366 322 2394 327
rect 2366 56 2394 294
rect 2590 56 2618 798
rect 2814 56 2842 1974
rect 2926 714 2954 5502
rect 3374 5026 3402 5614
rect 3430 5418 3458 6006
rect 3430 5385 3458 5390
rect 3374 4993 3402 4998
rect 3430 5082 3458 5087
rect 3430 4410 3458 5054
rect 3430 4377 3458 4382
rect 3430 4242 3458 4247
rect 2982 3626 3010 3631
rect 2982 3579 3010 3598
rect 3150 3626 3178 3631
rect 3150 3579 3178 3598
rect 3374 3626 3402 3631
rect 3374 3122 3402 3598
rect 3374 3089 3402 3094
rect 3430 2954 3458 4214
rect 3430 2921 3458 2926
rect 2926 681 2954 686
rect 3038 2730 3066 2735
rect 3038 56 3066 2702
rect 3430 1778 3458 1783
rect 3374 994 3402 999
rect 3374 490 3402 966
rect 3262 462 3402 490
rect 3262 56 3290 462
rect 3430 154 3458 1750
rect 3430 121 3458 126
rect 3486 56 3514 6454
rect 3542 5474 3570 6958
rect 3598 6425 3626 7056
rect 4942 7042 4970 7056
rect 4942 7009 4970 7014
rect 5334 7042 5362 7047
rect 3598 6399 3599 6425
rect 3625 6399 3626 6425
rect 3598 6393 3626 6399
rect 3654 6930 3682 6935
rect 3542 5441 3570 5446
rect 3542 3794 3570 3799
rect 3542 1834 3570 3766
rect 3542 1801 3570 1806
rect 3598 2618 3626 2623
rect 3542 1554 3570 1559
rect 3542 322 3570 1526
rect 3598 1050 3626 2590
rect 3654 1498 3682 6902
rect 4046 6818 4074 6823
rect 4046 6537 4074 6790
rect 4046 6511 4047 6537
rect 4073 6511 4074 6537
rect 4046 6505 4074 6511
rect 5278 6594 5306 6599
rect 5166 6481 5194 6487
rect 5166 6455 5167 6481
rect 5193 6455 5194 6481
rect 3878 6146 3906 6151
rect 5166 6146 5194 6455
rect 5222 6146 5250 6151
rect 5166 6145 5250 6146
rect 5166 6119 5223 6145
rect 5249 6119 5250 6145
rect 5166 6118 5250 6119
rect 3822 5250 3850 5255
rect 3710 2898 3738 2903
rect 3710 1666 3738 2870
rect 3710 1633 3738 1638
rect 3766 2170 3794 2175
rect 3654 1465 3682 1470
rect 3598 1017 3626 1022
rect 3710 1442 3738 1447
rect 3542 289 3570 294
rect 3710 56 3738 1414
rect 3766 882 3794 2142
rect 3766 849 3794 854
rect 3822 714 3850 5222
rect 3878 2562 3906 6118
rect 5222 6113 5250 6118
rect 5110 5642 5138 5647
rect 4326 4970 4354 4975
rect 4270 4466 4298 4471
rect 4158 3738 4186 3743
rect 3878 2529 3906 2534
rect 3990 3682 4018 3687
rect 3822 681 3850 686
rect 3934 1050 3962 1055
rect 3934 56 3962 1022
rect 3990 770 4018 3654
rect 4158 2338 4186 3710
rect 4270 2450 4298 4438
rect 4270 2417 4298 2422
rect 4158 2305 4186 2310
rect 4326 2058 4354 4942
rect 5054 4242 5082 4247
rect 4942 4074 4970 4079
rect 4550 3681 4578 3687
rect 4550 3655 4551 3681
rect 4577 3655 4578 3681
rect 4550 3458 4578 3655
rect 4830 3626 4858 3631
rect 4830 3579 4858 3598
rect 4550 3425 4578 3430
rect 4942 3290 4970 4046
rect 4998 3626 5026 3631
rect 4998 3579 5026 3598
rect 4942 3257 4970 3262
rect 5054 2394 5082 4214
rect 5110 2730 5138 5614
rect 5166 4690 5194 4695
rect 5166 3010 5194 4662
rect 5166 2977 5194 2982
rect 5222 3514 5250 3519
rect 5110 2697 5138 2702
rect 5166 2786 5194 2791
rect 5166 2617 5194 2758
rect 5166 2591 5167 2617
rect 5193 2591 5194 2617
rect 5166 2585 5194 2591
rect 5054 2361 5082 2366
rect 5110 2226 5138 2231
rect 5110 2179 5138 2198
rect 4326 2025 4354 2030
rect 4550 1722 4578 1727
rect 3990 737 4018 742
rect 4158 1218 4186 1223
rect 4158 56 4186 1190
rect 4382 770 4410 775
rect 4382 56 4410 742
rect 4550 714 4578 1694
rect 4774 993 4802 999
rect 4774 967 4775 993
rect 4801 967 4802 993
rect 4606 938 4634 943
rect 4774 938 4802 967
rect 4606 937 4802 938
rect 4606 911 4607 937
rect 4633 911 4802 937
rect 4606 910 4802 911
rect 4998 938 5026 943
rect 4606 826 4634 910
rect 4998 891 5026 910
rect 4606 793 4634 798
rect 4830 826 4858 831
rect 4550 686 4634 714
rect 4606 56 4634 686
rect 4830 56 4858 798
rect 5222 826 5250 3486
rect 5222 793 5250 798
rect 5054 322 5082 327
rect 5054 56 5082 294
rect 5278 56 5306 6566
rect 5334 6593 5362 7014
rect 6286 7042 6314 7056
rect 6286 7009 6314 7014
rect 6510 7042 6538 7047
rect 5334 6567 5335 6593
rect 5361 6567 5362 6593
rect 5334 6561 5362 6567
rect 6510 6425 6538 7014
rect 7630 6538 7658 7056
rect 8974 7042 9002 7056
rect 8974 7009 9002 7014
rect 9198 7042 9226 7047
rect 8470 6874 8498 6879
rect 8414 6706 8442 6711
rect 7630 6510 7882 6538
rect 7014 6482 7042 6487
rect 7014 6481 7154 6482
rect 7014 6455 7015 6481
rect 7041 6455 7154 6481
rect 7014 6454 7154 6455
rect 7014 6449 7042 6454
rect 6510 6399 6511 6425
rect 6537 6399 6538 6425
rect 6510 6393 6538 6399
rect 5670 6370 5698 6375
rect 5670 6146 5698 6342
rect 5502 6145 5698 6146
rect 5502 6119 5671 6145
rect 5697 6119 5698 6145
rect 5502 6118 5698 6119
rect 5502 6089 5530 6118
rect 5670 6113 5698 6118
rect 6846 6202 6874 6207
rect 5502 6063 5503 6089
rect 5529 6063 5530 6089
rect 5502 6057 5530 6063
rect 6678 6090 6706 6095
rect 6622 6034 6650 6039
rect 6622 5138 6650 6006
rect 6678 5810 6706 6062
rect 6678 5777 6706 5782
rect 6846 5754 6874 6174
rect 6846 5721 6874 5726
rect 7126 5753 7154 6454
rect 7518 6426 7546 6431
rect 7518 6145 7546 6398
rect 7854 6201 7882 6510
rect 7854 6175 7855 6201
rect 7881 6175 7882 6201
rect 7854 6169 7882 6175
rect 8190 6482 8218 6487
rect 7518 6119 7519 6145
rect 7545 6119 7546 6145
rect 7518 6113 7546 6119
rect 7126 5727 7127 5753
rect 7153 5727 7154 5753
rect 7126 5721 7154 5727
rect 7182 5978 7210 5983
rect 7294 5978 7322 5983
rect 7182 5977 7322 5978
rect 7182 5951 7183 5977
rect 7209 5951 7295 5977
rect 7321 5951 7322 5977
rect 7182 5950 7322 5951
rect 6622 5105 6650 5110
rect 7182 4970 7210 5950
rect 7294 5945 7322 5950
rect 7406 5810 7434 5815
rect 7406 5763 7434 5782
rect 7518 5810 7546 5815
rect 7518 5763 7546 5782
rect 7182 4937 7210 4942
rect 7350 5418 7378 5423
rect 7126 4914 7154 4919
rect 6510 4466 6538 4471
rect 5446 2562 5474 2567
rect 5446 2515 5474 2534
rect 5558 2562 5586 2567
rect 5558 2515 5586 2534
rect 6454 2506 6482 2511
rect 5894 2225 5922 2231
rect 5894 2199 5895 2225
rect 5921 2199 5922 2225
rect 5334 2058 5362 2063
rect 5502 2058 5530 2063
rect 5334 2057 5530 2058
rect 5334 2031 5335 2057
rect 5361 2031 5503 2057
rect 5529 2031 5530 2057
rect 5334 2030 5530 2031
rect 5334 2025 5362 2030
rect 5502 434 5530 2030
rect 5502 401 5530 406
rect 5726 1834 5754 1839
rect 5502 210 5530 215
rect 5502 56 5530 182
rect 5726 56 5754 1806
rect 5894 1778 5922 2199
rect 6118 2058 6146 2063
rect 6398 2058 6426 2063
rect 6118 2057 6426 2058
rect 6118 2031 6119 2057
rect 6145 2031 6399 2057
rect 6425 2031 6426 2057
rect 6118 2030 6426 2031
rect 6118 2025 6146 2030
rect 5894 1745 5922 1750
rect 6174 1890 6202 1895
rect 5950 1498 5978 1503
rect 5950 56 5978 1470
rect 6174 56 6202 1862
rect 6398 714 6426 2030
rect 6454 1162 6482 2478
rect 6510 2226 6538 4438
rect 7126 4298 7154 4886
rect 7126 4265 7154 4270
rect 7182 4746 7210 4751
rect 7014 3178 7042 3183
rect 6510 2193 6538 2198
rect 6566 2842 6594 2847
rect 6566 1554 6594 2814
rect 6958 2562 6986 2567
rect 6566 1521 6594 1526
rect 6622 2058 6650 2063
rect 6454 1129 6482 1134
rect 6398 681 6426 686
rect 6398 602 6426 607
rect 6398 56 6426 574
rect 6622 56 6650 2030
rect 6734 1722 6762 1727
rect 6734 1386 6762 1694
rect 6734 1353 6762 1358
rect 6790 1274 6818 1279
rect 6902 1274 6930 1279
rect 6678 1273 6930 1274
rect 6678 1247 6791 1273
rect 6817 1247 6903 1273
rect 6929 1247 6930 1273
rect 6678 1246 6930 1247
rect 6678 770 6706 1246
rect 6790 1241 6818 1246
rect 6902 1241 6930 1246
rect 6678 737 6706 742
rect 6846 546 6874 551
rect 6846 56 6874 518
rect 6958 378 6986 2534
rect 6958 345 6986 350
rect 7014 322 7042 3150
rect 7126 2897 7154 2903
rect 7126 2871 7127 2897
rect 7153 2871 7154 2897
rect 7126 2506 7154 2871
rect 7126 2473 7154 2478
rect 7182 2338 7210 4718
rect 7350 3346 7378 5390
rect 8134 5306 8162 5311
rect 7574 5250 7602 5255
rect 7518 5082 7546 5087
rect 7518 4970 7546 5054
rect 7518 4937 7546 4942
rect 7574 4858 7602 5222
rect 7574 4825 7602 4830
rect 7462 4410 7490 4415
rect 7462 4186 7490 4382
rect 7462 4153 7490 4158
rect 7910 3850 7938 3855
rect 7350 3313 7378 3318
rect 7574 3626 7602 3631
rect 7182 2305 7210 2310
rect 7238 3234 7266 3239
rect 7182 1666 7210 1671
rect 7182 1441 7210 1638
rect 7182 1415 7183 1441
rect 7209 1415 7210 1441
rect 7182 1409 7210 1415
rect 7126 994 7154 999
rect 7014 289 7042 294
rect 7070 826 7098 831
rect 7070 56 7098 798
rect 7126 266 7154 966
rect 7126 233 7154 238
rect 7238 210 7266 3206
rect 7294 3122 7322 3127
rect 7294 322 7322 3094
rect 7350 3066 7378 3071
rect 7350 1890 7378 3038
rect 7574 2954 7602 3598
rect 7854 3458 7882 3463
rect 7798 3345 7826 3351
rect 7798 3319 7799 3345
rect 7825 3319 7826 3345
rect 7574 2921 7602 2926
rect 7630 3290 7658 3295
rect 7798 3290 7826 3319
rect 7630 3289 7826 3290
rect 7630 3263 7631 3289
rect 7657 3263 7826 3289
rect 7630 3262 7826 3263
rect 7406 2842 7434 2847
rect 7574 2842 7602 2847
rect 7406 2841 7602 2842
rect 7406 2815 7407 2841
rect 7433 2815 7575 2841
rect 7601 2815 7602 2841
rect 7406 2814 7602 2815
rect 7406 2809 7434 2814
rect 7350 1857 7378 1862
rect 7462 1610 7490 1615
rect 7462 490 7490 1582
rect 7518 1218 7546 1223
rect 7518 602 7546 1190
rect 7574 770 7602 2814
rect 7630 2674 7658 3262
rect 7630 2641 7658 2646
rect 7686 2730 7714 2735
rect 7686 1218 7714 2702
rect 7854 1890 7882 3430
rect 7910 3122 7938 3822
rect 8078 3289 8106 3295
rect 8078 3263 8079 3289
rect 8105 3263 8106 3289
rect 8078 3178 8106 3263
rect 8078 3145 8106 3150
rect 7910 3089 7938 3094
rect 7854 1857 7882 1862
rect 7686 1185 7714 1190
rect 7966 1610 7994 1615
rect 7574 737 7602 742
rect 7518 569 7546 574
rect 7742 658 7770 663
rect 7462 462 7546 490
rect 7294 289 7322 294
rect 7238 182 7322 210
rect 7294 56 7322 182
rect 7518 56 7546 462
rect 7742 56 7770 630
rect 7966 56 7994 1582
rect 8134 826 8162 5278
rect 8190 3570 8218 6454
rect 8358 6033 8386 6039
rect 8358 6007 8359 6033
rect 8385 6007 8386 6033
rect 8358 5754 8386 6007
rect 8414 5810 8442 6678
rect 8414 5777 8442 5782
rect 8358 5721 8386 5726
rect 8470 5642 8498 6846
rect 9198 6425 9226 7014
rect 9926 7042 9954 7047
rect 9702 6482 9730 6487
rect 9702 6435 9730 6454
rect 9198 6399 9199 6425
rect 9225 6399 9226 6425
rect 9198 6393 9226 6399
rect 9086 5754 9114 5759
rect 9086 5707 9114 5726
rect 9366 5698 9394 5703
rect 9366 5651 9394 5670
rect 9478 5698 9506 5703
rect 9478 5651 9506 5670
rect 8470 5609 8498 5614
rect 8582 5530 8610 5535
rect 8526 5502 8582 5530
rect 8414 5138 8442 5143
rect 8358 5110 8414 5138
rect 8358 4634 8386 5110
rect 8414 5105 8442 5110
rect 8358 4601 8386 4606
rect 8470 4634 8498 4639
rect 8470 4466 8498 4606
rect 8470 4433 8498 4438
rect 8190 3537 8218 3542
rect 8246 4298 8274 4303
rect 8190 2898 8218 2903
rect 8190 2851 8218 2870
rect 8246 1050 8274 4270
rect 8526 4214 8554 5502
rect 8582 5497 8610 5502
rect 9366 5474 9394 5479
rect 9198 4802 9226 4807
rect 8974 4690 9002 4695
rect 8806 4466 8834 4471
rect 8470 4186 8554 4214
rect 8582 4354 8610 4359
rect 8302 2898 8330 2903
rect 8302 2851 8330 2870
rect 8414 2674 8442 2679
rect 8358 2646 8414 2674
rect 8302 2618 8330 2623
rect 8302 2450 8330 2590
rect 8302 2417 8330 2422
rect 8358 2170 8386 2646
rect 8414 2641 8442 2646
rect 8470 2562 8498 4186
rect 8470 2529 8498 2534
rect 8526 3122 8554 3127
rect 8526 2282 8554 3094
rect 8582 3066 8610 4326
rect 8806 3514 8834 4438
rect 8918 4073 8946 4079
rect 8918 4047 8919 4073
rect 8945 4047 8946 4073
rect 8918 3962 8946 4047
rect 8918 3929 8946 3934
rect 8806 3481 8834 3486
rect 8918 3514 8946 3519
rect 8582 3033 8610 3038
rect 8862 2954 8890 2959
rect 8526 2249 8554 2254
rect 8582 2897 8610 2903
rect 8582 2871 8583 2897
rect 8609 2871 8610 2897
rect 8358 2137 8386 2142
rect 8246 1017 8274 1022
rect 8470 1442 8498 1447
rect 8414 882 8442 887
rect 8134 793 8162 798
rect 8358 854 8414 882
rect 8358 490 8386 854
rect 8414 849 8442 854
rect 8358 457 8386 462
rect 8414 154 8442 159
rect 8470 154 8498 1414
rect 8582 1442 8610 2871
rect 8694 2730 8722 2735
rect 8694 2562 8722 2702
rect 8694 2529 8722 2534
rect 8582 1409 8610 1414
rect 8694 2114 8722 2119
rect 8526 1330 8554 1335
rect 8638 1330 8666 1335
rect 8554 1329 8666 1330
rect 8554 1303 8639 1329
rect 8665 1303 8666 1329
rect 8554 1302 8666 1303
rect 8526 1283 8554 1302
rect 8638 1297 8666 1302
rect 8638 322 8666 327
rect 8526 154 8554 159
rect 8470 126 8526 154
rect 8190 98 8218 103
rect 8190 56 8218 70
rect 8414 56 8442 126
rect 8526 121 8554 126
rect 8638 56 8666 294
rect 8694 210 8722 2086
rect 8694 177 8722 182
rect 8862 56 8890 2926
rect 8918 1498 8946 3486
rect 8974 2730 9002 4662
rect 9198 4186 9226 4774
rect 9198 4153 9226 4158
rect 9142 4129 9170 4135
rect 9142 4103 9143 4129
rect 9169 4103 9170 4129
rect 9142 4074 9170 4103
rect 9254 4074 9282 4079
rect 9142 4046 9254 4074
rect 9254 4027 9282 4046
rect 9254 3906 9282 3911
rect 9254 3346 9282 3878
rect 9254 3313 9282 3318
rect 8974 2697 9002 2702
rect 9254 3122 9282 3127
rect 9142 2674 9170 2679
rect 9142 2627 9170 2646
rect 9254 2394 9282 3094
rect 9310 2674 9338 2679
rect 9310 2627 9338 2646
rect 9254 2361 9282 2366
rect 9366 2338 9394 5446
rect 9590 5194 9618 5199
rect 9870 5194 9898 5199
rect 9618 5166 9870 5194
rect 9590 5161 9618 5166
rect 9870 5161 9898 5166
rect 9534 5138 9562 5143
rect 9534 5026 9562 5110
rect 9926 5082 9954 7014
rect 10318 6762 10346 7056
rect 11550 6762 11578 6767
rect 10318 6734 10402 6762
rect 10318 6482 10346 6487
rect 10318 6145 10346 6454
rect 10374 6426 10402 6734
rect 10766 6538 10794 6543
rect 10542 6426 10570 6431
rect 10374 6425 10570 6426
rect 10374 6399 10543 6425
rect 10569 6399 10570 6425
rect 10374 6398 10570 6399
rect 10542 6393 10570 6398
rect 10766 6146 10794 6510
rect 11046 6482 11074 6487
rect 11046 6481 11186 6482
rect 11046 6455 11047 6481
rect 11073 6455 11186 6481
rect 11046 6454 11186 6455
rect 11046 6449 11074 6454
rect 10318 6119 10319 6145
rect 10345 6119 10346 6145
rect 10318 6113 10346 6119
rect 10598 6145 10794 6146
rect 10598 6119 10767 6145
rect 10793 6119 10794 6145
rect 10598 6118 10794 6119
rect 10598 6089 10626 6118
rect 10766 6113 10794 6118
rect 11158 6145 11186 6454
rect 11158 6119 11159 6145
rect 11185 6119 11186 6145
rect 11158 6113 11186 6119
rect 11550 6146 11578 6734
rect 11662 6762 11690 7056
rect 12838 6874 12866 6879
rect 11662 6729 11690 6734
rect 12054 6762 12082 6767
rect 12054 6425 12082 6734
rect 12232 6678 12364 6683
rect 12260 6650 12284 6678
rect 12312 6650 12336 6678
rect 12232 6645 12364 6650
rect 12054 6399 12055 6425
rect 12081 6399 12082 6425
rect 12054 6393 12082 6399
rect 12558 6481 12586 6487
rect 12558 6455 12559 6481
rect 12585 6455 12586 6481
rect 11902 6286 12034 6291
rect 11930 6258 11954 6286
rect 11982 6258 12006 6286
rect 11902 6253 12034 6258
rect 12558 6146 12586 6455
rect 11550 6145 11746 6146
rect 11550 6119 11551 6145
rect 11577 6119 11746 6145
rect 11550 6118 11746 6119
rect 11550 6113 11578 6118
rect 10598 6063 10599 6089
rect 10625 6063 10626 6089
rect 10598 6057 10626 6063
rect 11718 6089 11746 6118
rect 12558 6113 12586 6118
rect 11718 6063 11719 6089
rect 11745 6063 11746 6089
rect 11718 6057 11746 6063
rect 11998 6034 12026 6039
rect 11998 6033 12138 6034
rect 11998 6007 11999 6033
rect 12025 6007 12138 6033
rect 11998 6006 12138 6007
rect 11998 6001 12026 6006
rect 11438 5977 11466 5983
rect 11438 5951 11439 5977
rect 11465 5951 11466 5977
rect 11438 5642 11466 5951
rect 11550 5642 11578 5647
rect 11998 5642 12026 5647
rect 11438 5641 11578 5642
rect 11438 5615 11551 5641
rect 11577 5615 11578 5641
rect 11438 5614 11578 5615
rect 11550 5586 11578 5614
rect 11550 5553 11578 5558
rect 11830 5614 11998 5642
rect 11774 5530 11802 5535
rect 10206 5362 10234 5367
rect 9814 5054 9954 5082
rect 10150 5082 10178 5087
rect 9702 5026 9730 5031
rect 9534 5025 9730 5026
rect 9534 4999 9535 5025
rect 9561 4999 9703 5025
rect 9729 4999 9730 5025
rect 9534 4998 9730 4999
rect 9534 4993 9562 4998
rect 9702 4993 9730 4998
rect 9758 3850 9786 3855
rect 9646 3234 9674 3239
rect 9422 2674 9450 2679
rect 9422 2562 9450 2646
rect 9422 2529 9450 2534
rect 9366 2305 9394 2310
rect 9590 2505 9618 2511
rect 9590 2479 9591 2505
rect 9617 2479 9618 2505
rect 9366 2170 9394 2175
rect 9030 2114 9058 2119
rect 9030 2067 9058 2086
rect 9310 2058 9338 2063
rect 9310 2011 9338 2030
rect 9254 1890 9282 1895
rect 9254 1778 9282 1862
rect 9254 1745 9282 1750
rect 8918 1465 8946 1470
rect 9254 1498 9282 1503
rect 8918 1329 8946 1335
rect 8918 1303 8919 1329
rect 8945 1303 8946 1329
rect 8918 602 8946 1303
rect 9254 826 9282 1470
rect 9366 1106 9394 2142
rect 9478 2058 9506 2063
rect 9478 2011 9506 2030
rect 9590 1330 9618 2479
rect 9590 1297 9618 1302
rect 9366 1073 9394 1078
rect 9590 993 9618 999
rect 9590 967 9591 993
rect 9617 967 9618 993
rect 9422 937 9450 943
rect 9422 911 9423 937
rect 9449 911 9450 937
rect 9422 882 9450 911
rect 9422 849 9450 854
rect 9590 882 9618 967
rect 9590 849 9618 854
rect 9254 793 9282 798
rect 8918 569 8946 574
rect 9534 714 9562 719
rect 9086 434 9114 439
rect 9086 56 9114 406
rect 9310 378 9338 383
rect 9310 56 9338 350
rect 9534 56 9562 686
rect 9646 266 9674 3206
rect 9758 2617 9786 3822
rect 9758 2591 9759 2617
rect 9785 2591 9786 2617
rect 9758 2585 9786 2591
rect 9814 1610 9842 5054
rect 9870 4970 9898 4975
rect 9870 3458 9898 4942
rect 9982 4858 10010 4863
rect 9982 4811 10010 4830
rect 10038 4746 10066 4751
rect 9870 3425 9898 3430
rect 9926 4410 9954 4415
rect 9814 1577 9842 1582
rect 9870 1162 9898 1167
rect 9870 1049 9898 1134
rect 9870 1023 9871 1049
rect 9897 1023 9898 1049
rect 9870 1017 9898 1023
rect 9926 826 9954 4382
rect 9926 793 9954 798
rect 9982 4074 10010 4079
rect 10038 4074 10066 4718
rect 10150 4522 10178 5054
rect 10150 4489 10178 4494
rect 10094 4074 10122 4079
rect 10038 4046 10094 4074
rect 9646 233 9674 238
rect 9758 770 9786 775
rect 9758 56 9786 742
rect 9982 56 10010 4046
rect 10094 4041 10122 4046
rect 10094 3794 10122 3799
rect 10094 3066 10122 3766
rect 10206 3122 10234 5334
rect 11718 5306 11746 5311
rect 11774 5306 11802 5502
rect 11830 5418 11858 5614
rect 11998 5595 12026 5614
rect 11902 5502 12034 5507
rect 11930 5474 11954 5502
rect 11982 5474 12006 5502
rect 11902 5469 12034 5474
rect 11942 5418 11970 5423
rect 11830 5385 11858 5390
rect 11886 5390 11942 5418
rect 11886 5306 11914 5390
rect 11942 5385 11970 5390
rect 11774 5278 11914 5306
rect 11270 5250 11298 5255
rect 11046 4802 11074 4807
rect 11046 3794 11074 4774
rect 11158 4578 11186 4583
rect 11158 4531 11186 4550
rect 11102 4186 11130 4191
rect 11102 4139 11130 4158
rect 11214 4186 11242 4191
rect 11214 4139 11242 4158
rect 11270 3906 11298 5222
rect 11662 5138 11690 5143
rect 11662 4634 11690 5110
rect 11718 5026 11746 5278
rect 11718 4993 11746 4998
rect 12110 4746 12138 6006
rect 12670 5978 12698 5983
rect 12782 5978 12810 5983
rect 12670 5977 12810 5978
rect 12670 5951 12671 5977
rect 12697 5951 12783 5977
rect 12809 5951 12810 5977
rect 12670 5950 12810 5951
rect 12670 5945 12698 5950
rect 12232 5894 12364 5899
rect 12260 5866 12284 5894
rect 12312 5866 12336 5894
rect 12232 5861 12364 5866
rect 12278 5697 12306 5703
rect 12278 5671 12279 5697
rect 12305 5671 12306 5697
rect 12278 5642 12306 5671
rect 12278 5609 12306 5614
rect 12558 5642 12586 5647
rect 12558 5641 12698 5642
rect 12558 5615 12559 5641
rect 12585 5615 12698 5641
rect 12558 5614 12698 5615
rect 12558 5609 12586 5614
rect 12166 5474 12194 5479
rect 12166 5082 12194 5446
rect 12232 5110 12364 5115
rect 12260 5082 12284 5110
rect 12312 5082 12336 5110
rect 12232 5077 12364 5082
rect 12166 5049 12194 5054
rect 11902 4718 12034 4723
rect 11930 4690 11954 4718
rect 11982 4690 12006 4718
rect 12110 4713 12138 4718
rect 12614 4970 12642 4975
rect 11902 4685 12034 4690
rect 12166 4690 12194 4695
rect 11662 4601 11690 4606
rect 11326 4578 11354 4583
rect 11326 4521 11354 4550
rect 11326 4495 11327 4521
rect 11353 4495 11354 4521
rect 11326 4489 11354 4495
rect 11606 4522 11634 4527
rect 11606 4475 11634 4494
rect 11494 4410 11522 4415
rect 11494 4185 11522 4382
rect 12166 4354 12194 4662
rect 12614 4578 12642 4942
rect 12614 4531 12642 4550
rect 12614 4466 12642 4471
rect 12614 4354 12642 4438
rect 12166 4321 12194 4326
rect 12232 4326 12364 4331
rect 12260 4298 12284 4326
rect 12312 4298 12336 4326
rect 12614 4321 12642 4326
rect 12232 4293 12364 4298
rect 11494 4159 11495 4185
rect 11521 4159 11522 4185
rect 11494 4153 11522 4159
rect 11270 3873 11298 3878
rect 11494 3962 11522 3967
rect 12614 3962 12642 3967
rect 11046 3761 11074 3766
rect 10710 3681 10738 3687
rect 10710 3655 10711 3681
rect 10737 3655 10738 3681
rect 10262 3626 10290 3631
rect 10430 3626 10458 3631
rect 10262 3625 10458 3626
rect 10262 3599 10263 3625
rect 10289 3599 10431 3625
rect 10457 3599 10458 3625
rect 10262 3598 10458 3599
rect 10262 3402 10290 3598
rect 10430 3593 10458 3598
rect 10710 3626 10738 3655
rect 10710 3593 10738 3598
rect 10262 3369 10290 3374
rect 10206 3089 10234 3094
rect 11438 3290 11466 3295
rect 10094 3033 10122 3038
rect 10038 2562 10066 2567
rect 10094 2562 10122 2567
rect 10150 2562 10178 2567
rect 10038 2561 10094 2562
rect 10038 2535 10039 2561
rect 10065 2535 10094 2561
rect 10038 2534 10094 2535
rect 10122 2561 10178 2562
rect 10122 2535 10151 2561
rect 10177 2535 10178 2561
rect 10122 2534 10178 2535
rect 10038 2529 10066 2534
rect 10094 2529 10122 2534
rect 10150 2529 10178 2534
rect 10486 2562 10514 2567
rect 10206 2058 10234 2063
rect 10206 56 10234 2030
rect 10262 1554 10290 1559
rect 10262 1106 10290 1526
rect 10430 1106 10458 1111
rect 10262 1105 10458 1106
rect 10262 1079 10263 1105
rect 10289 1079 10431 1105
rect 10457 1079 10458 1105
rect 10262 1078 10458 1079
rect 10262 1073 10290 1078
rect 10430 1073 10458 1078
rect 10486 994 10514 2534
rect 11326 2562 11354 2567
rect 10710 2506 10738 2511
rect 10710 1834 10738 2478
rect 10878 2282 10906 2287
rect 11214 2282 11242 2287
rect 10906 2254 10962 2282
rect 10878 2249 10906 2254
rect 10710 1801 10738 1806
rect 10934 1666 10962 2254
rect 10934 1633 10962 1638
rect 10710 1386 10738 1391
rect 10710 1049 10738 1358
rect 10710 1023 10711 1049
rect 10737 1023 10738 1049
rect 10710 1017 10738 1023
rect 11102 1218 11130 1223
rect 10430 966 10514 994
rect 10598 994 10626 999
rect 10934 994 10962 999
rect 10430 56 10458 966
rect 10598 714 10626 966
rect 10598 681 10626 686
rect 10766 993 10962 994
rect 10766 967 10935 993
rect 10961 967 10962 993
rect 10766 966 10962 967
rect 10766 658 10794 966
rect 10934 961 10962 966
rect 10654 657 10794 658
rect 10654 631 10767 657
rect 10793 631 10794 657
rect 10654 630 10794 631
rect 10654 56 10682 630
rect 10766 625 10794 630
rect 10878 882 10906 887
rect 10878 56 10906 854
rect 11046 602 11074 607
rect 11046 555 11074 574
rect 11102 56 11130 1190
rect 11214 1049 11242 2254
rect 11214 1023 11215 1049
rect 11241 1023 11242 1049
rect 11214 1017 11242 1023
rect 11214 546 11242 551
rect 11214 98 11242 518
rect 11214 65 11242 70
rect 11326 56 11354 2534
rect 11382 1442 11410 1447
rect 11382 1049 11410 1414
rect 11382 1023 11383 1049
rect 11409 1023 11410 1049
rect 11382 1017 11410 1023
rect 11438 770 11466 3262
rect 11494 2898 11522 3934
rect 11902 3934 12034 3939
rect 11930 3906 11954 3934
rect 11982 3906 12006 3934
rect 11902 3901 12034 3906
rect 12166 3906 12194 3911
rect 11886 3682 11914 3687
rect 11886 3458 11914 3654
rect 12166 3570 12194 3878
rect 12558 3794 12586 3799
rect 12614 3794 12642 3934
rect 12586 3766 12642 3794
rect 12670 3794 12698 5614
rect 12726 4914 12754 5950
rect 12782 5945 12810 5950
rect 12726 4881 12754 4886
rect 12782 4578 12810 4583
rect 12782 4521 12810 4550
rect 12782 4495 12783 4521
rect 12809 4495 12810 4521
rect 12782 4489 12810 4495
rect 12838 4242 12866 6846
rect 12838 4209 12866 4214
rect 12894 6706 12922 6711
rect 12894 4214 12922 6678
rect 13006 6426 13034 7056
rect 13118 6650 13146 6655
rect 13062 6426 13090 6431
rect 13006 6425 13090 6426
rect 13006 6399 13063 6425
rect 13089 6399 13090 6425
rect 13006 6398 13090 6399
rect 13062 6393 13090 6398
rect 13062 6146 13090 6151
rect 13118 6146 13146 6622
rect 13286 6594 13314 6599
rect 13062 6145 13146 6146
rect 13062 6119 13063 6145
rect 13089 6119 13146 6145
rect 13062 6118 13146 6119
rect 13230 6146 13258 6151
rect 13062 6113 13090 6118
rect 13230 6099 13258 6118
rect 12950 6034 12978 6039
rect 12950 5082 12978 6006
rect 12950 5049 12978 5054
rect 13006 5586 13034 5591
rect 13006 4690 13034 5558
rect 13006 4657 13034 4662
rect 13118 5250 13146 5255
rect 13062 4578 13090 4583
rect 13062 4531 13090 4550
rect 13118 4298 13146 5222
rect 13286 4410 13314 6566
rect 13566 6481 13594 6487
rect 13566 6455 13567 6481
rect 13593 6455 13594 6481
rect 13510 5977 13538 5983
rect 13510 5951 13511 5977
rect 13537 5951 13538 5977
rect 13510 5866 13538 5951
rect 13510 5833 13538 5838
rect 13454 5754 13482 5759
rect 13454 4690 13482 5726
rect 13510 5418 13538 5423
rect 13510 4746 13538 5390
rect 13566 5362 13594 6455
rect 14350 6426 14378 7056
rect 15190 6762 15218 6767
rect 15694 6762 15722 7056
rect 16086 6930 16114 6935
rect 15694 6734 15946 6762
rect 15078 6481 15106 6487
rect 15078 6455 15079 6481
rect 15105 6455 15106 6481
rect 14574 6426 14602 6431
rect 14350 6425 14602 6426
rect 14350 6399 14575 6425
rect 14601 6399 14602 6425
rect 14350 6398 14602 6399
rect 14574 6393 14602 6398
rect 14014 6090 14042 6095
rect 14014 6043 14042 6062
rect 14238 6090 14266 6095
rect 14238 6043 14266 6062
rect 14518 6090 14546 6095
rect 15078 6090 15106 6455
rect 15078 6062 15162 6090
rect 14518 6043 14546 6062
rect 15134 6034 15162 6062
rect 15134 6001 15162 6006
rect 13678 5977 13706 5983
rect 13678 5951 13679 5977
rect 13705 5951 13706 5977
rect 13678 5866 13706 5951
rect 13678 5418 13706 5838
rect 14966 5978 14994 5983
rect 15078 5978 15106 5983
rect 14966 5977 15106 5978
rect 14966 5951 14967 5977
rect 14993 5951 15079 5977
rect 15105 5951 15106 5977
rect 14966 5950 15106 5951
rect 13678 5385 13706 5390
rect 14294 5474 14322 5479
rect 13566 5329 13594 5334
rect 13510 4713 13538 4718
rect 13902 5250 13930 5255
rect 13454 4657 13482 4662
rect 13454 4466 13482 4471
rect 13286 4382 13370 4410
rect 13118 4270 13314 4298
rect 12558 3761 12586 3766
rect 12670 3761 12698 3766
rect 12782 4186 12810 4191
rect 12894 4186 13034 4214
rect 12166 3537 12194 3542
rect 12232 3542 12364 3547
rect 12260 3514 12284 3542
rect 12312 3514 12336 3542
rect 12232 3509 12364 3514
rect 11886 3425 11914 3430
rect 12726 3346 12754 3351
rect 12558 3178 12586 3183
rect 11902 3150 12034 3155
rect 11494 2865 11522 2870
rect 11774 3122 11802 3127
rect 11930 3122 11954 3150
rect 11982 3122 12006 3150
rect 11902 3117 12034 3122
rect 11774 2170 11802 3094
rect 12054 2954 12082 2959
rect 11830 2842 11858 2847
rect 11830 2795 11858 2814
rect 11942 2842 11970 2847
rect 11942 2795 11970 2814
rect 12054 2674 12082 2926
rect 12446 2953 12474 2959
rect 12446 2927 12447 2953
rect 12473 2927 12474 2953
rect 12054 2641 12082 2646
rect 12110 2898 12138 2903
rect 12110 2394 12138 2870
rect 12222 2898 12250 2903
rect 12222 2851 12250 2870
rect 12232 2758 12364 2763
rect 12260 2730 12284 2758
rect 12312 2730 12336 2758
rect 12232 2725 12364 2730
rect 12222 2562 12250 2567
rect 12222 2515 12250 2534
rect 12446 2562 12474 2927
rect 12446 2529 12474 2534
rect 12558 2506 12586 3150
rect 12670 3066 12698 3071
rect 12670 3009 12698 3038
rect 12670 2983 12671 3009
rect 12697 2983 12698 3009
rect 12670 2977 12698 2983
rect 12558 2473 12586 2478
rect 12614 2954 12642 2959
rect 11902 2366 12034 2371
rect 11930 2338 11954 2366
rect 11982 2338 12006 2366
rect 12110 2361 12138 2366
rect 11902 2333 12034 2338
rect 11774 2137 11802 2142
rect 12166 2225 12194 2231
rect 12166 2199 12167 2225
rect 12193 2199 12194 2225
rect 11830 2058 11858 2063
rect 11942 2058 11970 2063
rect 11830 2057 11970 2058
rect 11830 2031 11831 2057
rect 11857 2031 11943 2057
rect 11969 2031 11970 2057
rect 11830 2030 11970 2031
rect 11830 2002 11858 2030
rect 11942 2025 11970 2030
rect 11830 1969 11858 1974
rect 11718 1777 11746 1783
rect 11718 1751 11719 1777
rect 11745 1751 11746 1777
rect 11494 1722 11522 1727
rect 11494 1442 11522 1694
rect 11494 1409 11522 1414
rect 11550 1722 11578 1727
rect 11718 1722 11746 1751
rect 11550 1721 11746 1722
rect 11550 1695 11551 1721
rect 11577 1695 11746 1721
rect 11550 1694 11746 1695
rect 11998 1722 12026 1727
rect 11550 882 11578 1694
rect 11998 1675 12026 1694
rect 11830 1610 11858 1615
rect 12110 1610 12138 1615
rect 11830 1050 11858 1582
rect 11902 1582 12034 1587
rect 11930 1554 11954 1582
rect 11982 1554 12006 1582
rect 11902 1549 12034 1554
rect 12110 1273 12138 1582
rect 12110 1247 12111 1273
rect 12137 1247 12138 1273
rect 12110 1218 12138 1247
rect 12110 1185 12138 1190
rect 11830 1017 11858 1022
rect 11550 849 11578 854
rect 11886 882 11914 887
rect 11886 881 12138 882
rect 11886 855 11887 881
rect 11913 855 12138 881
rect 11886 854 12138 855
rect 11886 849 11914 854
rect 11902 798 12034 803
rect 11930 770 11954 798
rect 11982 770 12006 798
rect 11438 742 11578 770
rect 11902 765 12034 770
rect 11438 546 11466 551
rect 11438 499 11466 518
rect 11550 56 11578 742
rect 11774 602 11802 607
rect 11774 56 11802 574
rect 12110 322 12138 854
rect 12166 601 12194 2199
rect 12232 1974 12364 1979
rect 12260 1946 12284 1974
rect 12312 1946 12336 1974
rect 12232 1941 12364 1946
rect 12278 1777 12306 1783
rect 12278 1751 12279 1777
rect 12305 1751 12306 1777
rect 12278 1610 12306 1751
rect 12558 1778 12586 1783
rect 12558 1731 12586 1750
rect 12278 1577 12306 1582
rect 12502 1722 12530 1727
rect 12446 1274 12474 1279
rect 12232 1190 12364 1195
rect 12260 1162 12284 1190
rect 12312 1162 12336 1190
rect 12232 1157 12364 1162
rect 12390 1106 12418 1111
rect 12446 1106 12474 1246
rect 12502 1218 12530 1694
rect 12614 1498 12642 2926
rect 12558 1470 12642 1498
rect 12670 2506 12698 2511
rect 12558 1218 12586 1470
rect 12614 1385 12642 1391
rect 12614 1359 12615 1385
rect 12641 1359 12642 1385
rect 12614 1330 12642 1359
rect 12614 1297 12642 1302
rect 12558 1190 12642 1218
rect 12502 1185 12530 1190
rect 12558 1106 12586 1111
rect 12390 1105 12586 1106
rect 12390 1079 12391 1105
rect 12417 1079 12559 1105
rect 12585 1079 12586 1105
rect 12390 1078 12586 1079
rect 12390 1073 12418 1078
rect 12558 1073 12586 1078
rect 12166 575 12167 601
rect 12193 575 12194 601
rect 12166 569 12194 575
rect 12446 546 12474 551
rect 12232 406 12364 411
rect 12260 378 12284 406
rect 12312 378 12336 406
rect 12232 373 12364 378
rect 12110 294 12250 322
rect 12222 56 12250 294
rect 12446 56 12474 518
rect 12558 546 12586 551
rect 12558 499 12586 518
rect 12614 378 12642 1190
rect 12670 658 12698 2478
rect 12670 625 12698 630
rect 12726 602 12754 3318
rect 12782 2954 12810 4158
rect 12838 3738 12866 3743
rect 12838 3691 12866 3710
rect 12950 3738 12978 3743
rect 12950 3691 12978 3710
rect 12782 2921 12810 2926
rect 12894 2898 12922 2903
rect 12838 2618 12866 2623
rect 12838 1890 12866 2590
rect 12838 1857 12866 1862
rect 12838 1273 12866 1279
rect 12838 1247 12839 1273
rect 12865 1247 12866 1273
rect 12838 1050 12866 1247
rect 12726 569 12754 574
rect 12782 1022 12866 1050
rect 12894 1050 12922 2870
rect 13006 2450 13034 4186
rect 13174 3793 13202 3799
rect 13174 3767 13175 3793
rect 13201 3767 13202 3793
rect 13118 3514 13146 3519
rect 13062 3290 13090 3295
rect 13062 3243 13090 3262
rect 13118 2898 13146 3486
rect 13118 2865 13146 2870
rect 13006 2417 13034 2422
rect 13062 1777 13090 1783
rect 13062 1751 13063 1777
rect 13089 1751 13090 1777
rect 13062 1386 13090 1751
rect 13174 1666 13202 3767
rect 13286 3570 13314 4270
rect 13286 3537 13314 3542
rect 13230 3345 13258 3351
rect 13230 3319 13231 3345
rect 13257 3319 13258 3345
rect 13230 3290 13258 3319
rect 13230 3257 13258 3262
rect 13286 2226 13314 2231
rect 13286 1890 13314 2198
rect 13342 2002 13370 4382
rect 13398 4354 13426 4359
rect 13398 4186 13426 4326
rect 13398 4153 13426 4158
rect 13398 3010 13426 3015
rect 13454 3010 13482 4438
rect 13734 4354 13762 4359
rect 13426 2982 13482 3010
rect 13510 3289 13538 3295
rect 13510 3263 13511 3289
rect 13537 3263 13538 3289
rect 13398 2977 13426 2982
rect 13342 1969 13370 1974
rect 13398 2394 13426 2399
rect 13286 1862 13370 1890
rect 13286 1722 13314 1727
rect 13062 1353 13090 1358
rect 13118 1638 13202 1666
rect 13230 1721 13314 1722
rect 13230 1695 13287 1721
rect 13313 1695 13314 1721
rect 13230 1694 13314 1695
rect 13118 1218 13146 1638
rect 13062 1190 13146 1218
rect 13006 1050 13034 1055
rect 12894 1049 13034 1050
rect 12894 1023 13007 1049
rect 13033 1023 13034 1049
rect 12894 1022 13034 1023
rect 12782 490 12810 1022
rect 13006 1017 13034 1022
rect 12838 937 12866 943
rect 12838 911 12839 937
rect 12865 911 12866 937
rect 12838 602 12866 911
rect 12838 569 12866 574
rect 12894 658 12922 663
rect 12614 345 12642 350
rect 12670 462 12810 490
rect 12670 56 12698 462
rect 12894 56 12922 630
rect 13062 601 13090 1190
rect 13230 658 13258 1694
rect 13286 1689 13314 1694
rect 13342 1554 13370 1862
rect 13286 1526 13370 1554
rect 13286 770 13314 1526
rect 13398 1386 13426 2366
rect 13398 1353 13426 1358
rect 13454 2226 13482 2231
rect 13342 1329 13370 1335
rect 13342 1303 13343 1329
rect 13369 1303 13370 1329
rect 13342 938 13370 1303
rect 13398 994 13426 999
rect 13454 994 13482 2198
rect 13426 966 13482 994
rect 13510 994 13538 3263
rect 13734 2506 13762 4326
rect 13902 3682 13930 5222
rect 13958 4802 13986 4807
rect 13958 4214 13986 4774
rect 14014 4634 14042 4639
rect 14014 4577 14042 4606
rect 14014 4551 14015 4577
rect 14041 4551 14042 4577
rect 14014 4545 14042 4551
rect 14238 4634 14266 4639
rect 14238 4521 14266 4606
rect 14238 4495 14239 4521
rect 14265 4495 14266 4521
rect 14238 4489 14266 4495
rect 14182 4298 14210 4303
rect 13958 4186 14042 4214
rect 13902 3649 13930 3654
rect 13734 2473 13762 2478
rect 13678 2057 13706 2063
rect 13678 2031 13679 2057
rect 13705 2031 13706 2057
rect 13678 1778 13706 2031
rect 13790 1778 13818 1783
rect 13678 1777 13818 1778
rect 13678 1751 13791 1777
rect 13817 1751 13818 1777
rect 13678 1750 13818 1751
rect 13398 961 13426 966
rect 13510 961 13538 966
rect 13622 1273 13650 1279
rect 13622 1247 13623 1273
rect 13649 1247 13650 1273
rect 13342 905 13370 910
rect 13510 882 13538 887
rect 13510 881 13594 882
rect 13510 855 13511 881
rect 13537 855 13594 881
rect 13510 854 13594 855
rect 13510 849 13538 854
rect 13286 737 13314 742
rect 13230 625 13258 630
rect 13454 658 13482 663
rect 13454 611 13482 630
rect 13062 575 13063 601
rect 13089 575 13090 601
rect 13062 569 13090 575
rect 13118 546 13146 551
rect 13118 56 13146 518
rect 13342 546 13370 551
rect 13342 56 13370 518
rect 13566 56 13594 854
rect 13622 546 13650 1247
rect 13790 1050 13818 1750
rect 14014 1498 14042 4186
rect 14126 1778 14154 1783
rect 14070 1722 14098 1727
rect 14070 1675 14098 1694
rect 14014 1465 14042 1470
rect 13790 1017 13818 1022
rect 14014 937 14042 943
rect 14014 911 14015 937
rect 14041 911 14042 937
rect 13622 513 13650 518
rect 13790 658 13818 663
rect 13790 56 13818 630
rect 14014 56 14042 911
rect 14126 714 14154 1750
rect 14182 1442 14210 4270
rect 14294 4214 14322 5446
rect 14350 5362 14378 5367
rect 14350 5315 14378 5334
rect 14630 5362 14658 5367
rect 14630 5305 14658 5334
rect 14798 5362 14826 5367
rect 14798 5315 14826 5334
rect 14630 5279 14631 5305
rect 14657 5279 14658 5305
rect 14630 5273 14658 5279
rect 14854 5306 14882 5311
rect 14350 5138 14378 5143
rect 14350 5026 14378 5110
rect 14350 4993 14378 4998
rect 14462 4577 14490 4583
rect 14462 4551 14463 4577
rect 14489 4551 14490 4577
rect 14462 4214 14490 4551
rect 14294 4186 14378 4214
rect 14294 2674 14322 2679
rect 14294 2627 14322 2646
rect 14350 2506 14378 4186
rect 14350 2473 14378 2478
rect 14406 4186 14490 4214
rect 14238 1442 14266 1447
rect 14182 1441 14378 1442
rect 14182 1415 14239 1441
rect 14265 1415 14378 1441
rect 14182 1414 14378 1415
rect 14238 1409 14266 1414
rect 14350 1385 14378 1414
rect 14350 1359 14351 1385
rect 14377 1359 14378 1385
rect 14350 1353 14378 1359
rect 14406 1049 14434 4186
rect 14630 4129 14658 4135
rect 14630 4103 14631 4129
rect 14657 4103 14658 4129
rect 14518 4074 14546 4079
rect 14630 4074 14658 4103
rect 14854 4130 14882 5278
rect 14854 4097 14882 4102
rect 14546 4046 14658 4074
rect 14910 4073 14938 4079
rect 14910 4047 14911 4073
rect 14937 4047 14938 4073
rect 14518 4027 14546 4046
rect 14910 3682 14938 4047
rect 14966 4074 14994 5950
rect 15078 5945 15106 5950
rect 15190 5866 15218 6734
rect 15918 6425 15946 6734
rect 15918 6399 15919 6425
rect 15945 6399 15946 6425
rect 15918 6393 15946 6399
rect 16086 6146 16114 6902
rect 17038 6594 17066 7056
rect 18382 6762 18410 7056
rect 19726 7042 19754 7056
rect 19726 7009 19754 7014
rect 19950 7042 19978 7047
rect 18382 6729 18410 6734
rect 18438 6930 18466 6935
rect 17038 6566 17290 6594
rect 16422 6482 16450 6487
rect 16422 6435 16450 6454
rect 17038 6482 17066 6487
rect 16534 6258 16562 6263
rect 16086 6145 16226 6146
rect 16086 6119 16087 6145
rect 16113 6119 16226 6145
rect 16086 6118 16226 6119
rect 16086 6113 16114 6118
rect 16198 6089 16226 6118
rect 16198 6063 16199 6089
rect 16225 6063 16226 6089
rect 16198 6057 16226 6063
rect 16422 6145 16450 6151
rect 16422 6119 16423 6145
rect 16449 6119 16450 6145
rect 15190 5833 15218 5838
rect 15358 6033 15386 6039
rect 15358 6007 15359 6033
rect 15385 6007 15386 6033
rect 15246 5194 15274 5199
rect 15246 5147 15274 5166
rect 14966 4041 14994 4046
rect 15022 4410 15050 4415
rect 14910 3649 14938 3654
rect 14462 2674 14490 2679
rect 14462 2627 14490 2646
rect 14910 2618 14938 2623
rect 14686 2617 14938 2618
rect 14686 2591 14911 2617
rect 14937 2591 14938 2617
rect 14686 2590 14938 2591
rect 14686 2058 14714 2590
rect 14910 2585 14938 2590
rect 14742 2506 14770 2511
rect 14742 2505 14882 2506
rect 14742 2479 14743 2505
rect 14769 2479 14882 2505
rect 14742 2478 14882 2479
rect 14742 2473 14770 2478
rect 14742 2058 14770 2063
rect 14686 2057 14770 2058
rect 14686 2031 14743 2057
rect 14769 2031 14770 2057
rect 14686 2030 14770 2031
rect 14742 1834 14770 2030
rect 14406 1023 14407 1049
rect 14433 1023 14434 1049
rect 14406 1017 14434 1023
rect 14574 1806 14770 1834
rect 14574 938 14602 1806
rect 14686 1721 14714 1727
rect 14686 1695 14687 1721
rect 14713 1695 14714 1721
rect 14630 1329 14658 1335
rect 14630 1303 14631 1329
rect 14657 1303 14658 1329
rect 14630 1050 14658 1303
rect 14686 1274 14714 1695
rect 14798 1274 14826 1279
rect 14686 1273 14826 1274
rect 14686 1247 14799 1273
rect 14825 1247 14826 1273
rect 14686 1246 14826 1247
rect 14630 1017 14658 1022
rect 14126 681 14154 686
rect 14406 910 14602 938
rect 14742 994 14770 999
rect 14238 545 14266 551
rect 14238 519 14239 545
rect 14265 519 14266 545
rect 14238 56 14266 519
rect 14406 210 14434 910
rect 14686 882 14714 887
rect 14406 177 14434 182
rect 14462 881 14714 882
rect 14462 855 14687 881
rect 14713 855 14714 881
rect 14462 854 14714 855
rect 14462 56 14490 854
rect 14686 849 14714 854
rect 14630 602 14658 607
rect 14742 602 14770 966
rect 14798 882 14826 1246
rect 14798 849 14826 854
rect 14630 601 14770 602
rect 14630 575 14631 601
rect 14657 575 14770 601
rect 14630 574 14770 575
rect 14854 601 14882 2478
rect 15022 2394 15050 4382
rect 15358 4214 15386 6007
rect 16310 6034 16338 6039
rect 15974 5474 16002 5479
rect 15694 5249 15722 5255
rect 15694 5223 15695 5249
rect 15721 5223 15722 5249
rect 15414 5194 15442 5199
rect 15414 5147 15442 5166
rect 15358 4186 15498 4214
rect 15358 4129 15386 4135
rect 15358 4103 15359 4129
rect 15385 4103 15386 4129
rect 15190 4073 15218 4079
rect 15190 4047 15191 4073
rect 15217 4047 15218 4073
rect 15190 4018 15218 4047
rect 15190 3985 15218 3990
rect 15358 4018 15386 4103
rect 15358 3985 15386 3990
rect 15470 4018 15498 4186
rect 15470 3985 15498 3990
rect 15582 4073 15610 4079
rect 15582 4047 15583 4073
rect 15609 4047 15610 4073
rect 15078 3906 15106 3911
rect 15106 3878 15162 3906
rect 15078 3873 15106 3878
rect 15022 2361 15050 2366
rect 15134 2226 15162 3878
rect 15190 3122 15218 3127
rect 15190 3010 15218 3094
rect 15190 2977 15218 2982
rect 15134 2193 15162 2198
rect 15190 2561 15218 2567
rect 15190 2535 15191 2561
rect 15217 2535 15218 2561
rect 15078 2058 15106 2063
rect 15078 1666 15106 2030
rect 15078 1633 15106 1638
rect 15078 1329 15106 1335
rect 15078 1303 15079 1329
rect 15105 1303 15106 1329
rect 15078 1106 15106 1303
rect 15078 1073 15106 1078
rect 15190 1049 15218 2535
rect 15246 1442 15274 1447
rect 15246 1385 15274 1414
rect 15246 1359 15247 1385
rect 15273 1359 15274 1385
rect 15246 1353 15274 1359
rect 15526 1274 15554 1279
rect 15190 1023 15191 1049
rect 15217 1023 15218 1049
rect 15190 1017 15218 1023
rect 15302 1273 15554 1274
rect 15302 1247 15527 1273
rect 15553 1247 15554 1273
rect 15302 1246 15554 1247
rect 15302 658 15330 1246
rect 15526 1241 15554 1246
rect 15582 994 15610 4047
rect 15694 3514 15722 5223
rect 15974 5026 16002 5446
rect 15918 4998 16002 5026
rect 15694 3481 15722 3486
rect 15806 4242 15834 4247
rect 15694 2562 15722 2567
rect 15582 961 15610 966
rect 15638 993 15666 999
rect 15638 967 15639 993
rect 15665 967 15666 993
rect 14854 575 14855 601
rect 14881 575 14882 601
rect 14630 569 14658 574
rect 14854 569 14882 575
rect 15134 630 15330 658
rect 15470 937 15498 943
rect 15470 911 15471 937
rect 15497 911 15498 937
rect 15470 826 15498 911
rect 14686 490 14714 495
rect 14686 56 14714 462
rect 15078 490 15106 495
rect 15078 443 15106 462
rect 14910 434 14938 439
rect 14910 56 14938 406
rect 15134 56 15162 630
rect 15358 210 15386 215
rect 15358 56 15386 182
rect 15470 154 15498 798
rect 15470 121 15498 126
rect 15582 882 15610 887
rect 15582 56 15610 854
rect 15638 826 15666 967
rect 15638 793 15666 798
rect 15694 98 15722 2534
rect 15750 1722 15778 1727
rect 15750 601 15778 1694
rect 15806 1554 15834 4214
rect 15918 3010 15946 4998
rect 16310 4969 16338 6006
rect 16310 4943 16311 4969
rect 16337 4943 16338 4969
rect 16310 4937 16338 4943
rect 15974 4634 16002 4639
rect 15974 3906 16002 4606
rect 16422 4214 16450 6119
rect 15974 3873 16002 3878
rect 16254 4186 16450 4214
rect 16478 5530 16506 5535
rect 15918 2977 15946 2982
rect 15974 2562 16002 2567
rect 16198 2562 16226 2567
rect 15974 2561 16226 2562
rect 15974 2535 15975 2561
rect 16001 2535 16199 2561
rect 16225 2535 16226 2561
rect 15974 2534 16226 2535
rect 15974 2506 16002 2534
rect 16198 2529 16226 2534
rect 15974 2473 16002 2478
rect 16254 2338 16282 4186
rect 16254 2305 16282 2310
rect 16422 3570 16450 3575
rect 16142 2226 16170 2231
rect 16170 2198 16282 2226
rect 16142 2179 16170 2198
rect 16254 2169 16282 2198
rect 16254 2143 16255 2169
rect 16281 2143 16282 2169
rect 16254 2137 16282 2143
rect 16310 1666 16338 1671
rect 15806 1521 15834 1526
rect 16086 1665 16338 1666
rect 16086 1639 16311 1665
rect 16337 1639 16338 1665
rect 16086 1638 16338 1639
rect 16030 1330 16058 1335
rect 15918 1329 16058 1330
rect 15918 1303 16031 1329
rect 16057 1303 16058 1329
rect 15918 1302 16058 1303
rect 15918 1049 15946 1302
rect 16030 1297 16058 1302
rect 15918 1023 15919 1049
rect 15945 1023 15946 1049
rect 15918 1017 15946 1023
rect 15750 575 15751 601
rect 15777 575 15778 601
rect 15750 569 15778 575
rect 15806 658 15834 663
rect 15694 65 15722 70
rect 15806 56 15834 630
rect 16030 489 16058 495
rect 16030 463 16031 489
rect 16057 463 16058 489
rect 16030 434 16058 463
rect 16030 401 16058 406
rect 16086 322 16114 1638
rect 16310 1633 16338 1638
rect 16310 1273 16338 1279
rect 16310 1247 16311 1273
rect 16337 1247 16338 1273
rect 16198 1050 16226 1055
rect 16198 1003 16226 1022
rect 16310 658 16338 1247
rect 16310 625 16338 630
rect 16030 294 16114 322
rect 16254 434 16282 439
rect 16030 56 16058 294
rect 16254 56 16282 406
rect 16422 266 16450 3542
rect 16478 2617 16506 5502
rect 16534 4214 16562 6230
rect 16758 6202 16786 6207
rect 16758 5754 16786 6174
rect 16758 5721 16786 5726
rect 16758 5250 16786 5255
rect 16590 4913 16618 4919
rect 16590 4887 16591 4913
rect 16617 4887 16618 4913
rect 16590 4858 16618 4887
rect 16702 4858 16730 4863
rect 16590 4857 16730 4858
rect 16590 4831 16703 4857
rect 16729 4831 16730 4857
rect 16590 4830 16730 4831
rect 16702 4802 16730 4830
rect 16702 4769 16730 4774
rect 16534 4186 16674 4214
rect 16478 2591 16479 2617
rect 16505 2591 16506 2617
rect 16478 2585 16506 2591
rect 16646 2170 16674 4186
rect 16758 3794 16786 5222
rect 16758 3761 16786 3766
rect 16814 4746 16842 4751
rect 16814 2674 16842 4718
rect 17038 4634 17066 6454
rect 17262 6201 17290 6566
rect 17262 6175 17263 6201
rect 17289 6175 17290 6201
rect 17262 6169 17290 6175
rect 18214 6370 18242 6375
rect 17766 6034 17794 6039
rect 17766 5987 17794 6006
rect 18046 5978 18074 5983
rect 17094 5810 17122 5815
rect 17094 5362 17122 5782
rect 17206 5810 17234 5815
rect 17206 5530 17234 5782
rect 17542 5697 17570 5703
rect 17542 5671 17543 5697
rect 17569 5671 17570 5697
rect 17206 5497 17234 5502
rect 17374 5642 17402 5647
rect 17542 5642 17570 5671
rect 17374 5641 17570 5642
rect 17374 5615 17375 5641
rect 17401 5615 17570 5641
rect 17374 5614 17570 5615
rect 17822 5641 17850 5647
rect 17822 5615 17823 5641
rect 17849 5615 17850 5641
rect 17374 5474 17402 5614
rect 17374 5441 17402 5446
rect 17710 5586 17738 5591
rect 17094 5361 17290 5362
rect 17094 5335 17095 5361
rect 17121 5335 17290 5361
rect 17094 5334 17290 5335
rect 17094 5329 17122 5334
rect 17262 5305 17290 5334
rect 17262 5279 17263 5305
rect 17289 5279 17290 5305
rect 17262 5273 17290 5279
rect 17542 5249 17570 5255
rect 17542 5223 17543 5249
rect 17569 5223 17570 5249
rect 17542 5194 17570 5223
rect 17542 5161 17570 5166
rect 17206 5082 17234 5087
rect 17206 5026 17234 5054
rect 17318 5026 17346 5031
rect 17206 5025 17346 5026
rect 17206 4999 17207 5025
rect 17233 4999 17319 5025
rect 17345 4999 17346 5025
rect 17206 4998 17346 4999
rect 17206 4993 17234 4998
rect 17318 4993 17346 4998
rect 17598 5026 17626 5031
rect 17598 4969 17626 4998
rect 17598 4943 17599 4969
rect 17625 4943 17626 4969
rect 17598 4937 17626 4943
rect 17038 4601 17066 4606
rect 17374 3794 17402 3799
rect 17402 3766 17570 3794
rect 17374 3747 17402 3766
rect 17542 3737 17570 3766
rect 17542 3711 17543 3737
rect 17569 3711 17570 3737
rect 17542 3705 17570 3711
rect 17486 3346 17514 3351
rect 17486 3010 17514 3318
rect 17486 3009 17626 3010
rect 17486 2983 17487 3009
rect 17513 2983 17626 3009
rect 17486 2982 17626 2983
rect 17486 2977 17514 2982
rect 17598 2953 17626 2982
rect 17598 2927 17599 2953
rect 17625 2927 17626 2953
rect 17598 2921 17626 2927
rect 16814 2641 16842 2646
rect 17150 2898 17178 2903
rect 17150 2674 17178 2870
rect 17318 2674 17346 2679
rect 17150 2673 17346 2674
rect 17150 2647 17151 2673
rect 17177 2647 17319 2673
rect 17345 2647 17346 2673
rect 17150 2646 17346 2647
rect 17150 2641 17178 2646
rect 17318 2641 17346 2646
rect 17598 2618 17626 2623
rect 17598 2571 17626 2590
rect 17430 2394 17458 2399
rect 17430 2226 17458 2366
rect 17710 2282 17738 5558
rect 17822 5586 17850 5615
rect 17822 5553 17850 5558
rect 17822 3794 17850 3799
rect 17822 3747 17850 3766
rect 17710 2249 17738 2254
rect 17822 3009 17850 3015
rect 17822 2983 17823 3009
rect 17849 2983 17850 3009
rect 17486 2226 17514 2231
rect 17430 2225 17626 2226
rect 17430 2199 17487 2225
rect 17513 2199 17626 2225
rect 17430 2198 17626 2199
rect 17486 2193 17514 2198
rect 16646 2142 16786 2170
rect 16534 2114 16562 2119
rect 16534 2113 16730 2114
rect 16534 2087 16535 2113
rect 16561 2087 16730 2113
rect 16534 2086 16730 2087
rect 16534 2081 16562 2086
rect 16702 1777 16730 2086
rect 16702 1751 16703 1777
rect 16729 1751 16730 1777
rect 16702 1745 16730 1751
rect 16534 1330 16562 1335
rect 16478 882 16506 887
rect 16478 835 16506 854
rect 16534 714 16562 1302
rect 16422 233 16450 238
rect 16478 686 16562 714
rect 16646 770 16674 775
rect 16478 56 16506 686
rect 16646 658 16674 742
rect 16758 770 16786 2142
rect 17598 2169 17626 2198
rect 17598 2143 17599 2169
rect 17625 2143 17626 2169
rect 17598 2137 17626 2143
rect 17430 2114 17458 2119
rect 17094 2002 17122 2007
rect 17094 1834 17122 1974
rect 17094 1801 17122 1806
rect 17150 1722 17178 1727
rect 17150 1675 17178 1694
rect 17374 1666 17402 1671
rect 17206 1665 17402 1666
rect 17206 1639 17375 1665
rect 17401 1639 17402 1665
rect 17206 1638 17402 1639
rect 17038 1330 17066 1335
rect 17038 1283 17066 1302
rect 16758 737 16786 742
rect 17094 881 17122 887
rect 17094 855 17095 881
rect 17121 855 17122 881
rect 16646 625 16674 630
rect 16534 602 16562 607
rect 16534 555 16562 574
rect 16702 490 16730 495
rect 16702 56 16730 462
rect 16814 489 16842 495
rect 16814 463 16815 489
rect 16841 463 16842 489
rect 16814 210 16842 463
rect 17094 434 17122 855
rect 17206 826 17234 1638
rect 17374 1633 17402 1638
rect 17430 1385 17458 2086
rect 17430 1359 17431 1385
rect 17457 1359 17458 1385
rect 17430 1353 17458 1359
rect 17654 1722 17682 1727
rect 17654 1385 17682 1694
rect 17654 1359 17655 1385
rect 17681 1359 17682 1385
rect 17654 1353 17682 1359
rect 17822 1386 17850 2983
rect 18046 2954 18074 5950
rect 18046 2921 18074 2926
rect 18158 4354 18186 4359
rect 18158 2169 18186 4326
rect 18214 2562 18242 6342
rect 18438 5866 18466 6902
rect 18606 6762 18634 6767
rect 18606 6425 18634 6734
rect 18606 6399 18607 6425
rect 18633 6399 18634 6425
rect 18606 6393 18634 6399
rect 19110 6481 19138 6487
rect 19110 6455 19111 6481
rect 19137 6455 19138 6481
rect 19110 6146 19138 6455
rect 19950 6425 19978 7014
rect 21070 6762 21098 7056
rect 22414 7042 22442 7056
rect 22414 7009 22442 7014
rect 22582 7042 22610 7047
rect 21070 6729 21098 6734
rect 21574 6762 21602 6767
rect 21406 6650 21434 6655
rect 20454 6482 20482 6487
rect 20454 6481 20538 6482
rect 20454 6455 20455 6481
rect 20481 6455 20538 6481
rect 20454 6454 20538 6455
rect 20454 6449 20482 6454
rect 19950 6399 19951 6425
rect 19977 6399 19978 6425
rect 19950 6393 19978 6399
rect 19110 6113 19138 6118
rect 19950 6146 19978 6151
rect 19950 6099 19978 6118
rect 18550 6034 18578 6039
rect 18550 5987 18578 6006
rect 20230 6034 20258 6039
rect 20230 5987 20258 6006
rect 20398 6034 20426 6039
rect 20398 5987 20426 6006
rect 18830 5978 18858 5983
rect 18998 5978 19026 5983
rect 18830 5977 19082 5978
rect 18830 5951 18831 5977
rect 18857 5951 18999 5977
rect 19025 5951 19082 5977
rect 18830 5950 19082 5951
rect 18830 5945 18858 5950
rect 18998 5945 19026 5950
rect 18438 5838 18522 5866
rect 18326 5138 18354 5143
rect 18326 2954 18354 5110
rect 18438 4410 18466 4415
rect 18326 2921 18354 2926
rect 18382 4298 18410 4303
rect 18382 2730 18410 4270
rect 18382 2697 18410 2702
rect 18214 2529 18242 2534
rect 18438 2226 18466 4382
rect 18438 2193 18466 2198
rect 18158 2143 18159 2169
rect 18185 2143 18186 2169
rect 17878 2114 17906 2119
rect 17878 2067 17906 2086
rect 17878 1834 17906 1839
rect 17878 1787 17906 1806
rect 17990 1722 18018 1727
rect 18158 1722 18186 2143
rect 18438 2113 18466 2119
rect 18438 2087 18439 2113
rect 18465 2087 18466 2113
rect 18438 1834 18466 2087
rect 18438 1801 18466 1806
rect 17990 1721 18186 1722
rect 17990 1695 17991 1721
rect 18017 1695 18186 1721
rect 17990 1694 18186 1695
rect 17990 1689 18018 1694
rect 18270 1666 18298 1671
rect 17822 1353 17850 1358
rect 18046 1665 18298 1666
rect 18046 1639 18271 1665
rect 18297 1639 18298 1665
rect 18046 1638 18298 1639
rect 17878 1329 17906 1335
rect 17878 1303 17879 1329
rect 17905 1303 17906 1329
rect 17598 1050 17626 1055
rect 17598 1003 17626 1022
rect 17878 1050 17906 1303
rect 17878 1017 17906 1022
rect 17094 401 17122 406
rect 17150 798 17234 826
rect 17598 882 17626 887
rect 16814 177 16842 182
rect 16926 378 16954 383
rect 16926 56 16954 350
rect 17150 56 17178 798
rect 17486 658 17514 663
rect 17486 546 17514 630
rect 17486 513 17514 518
rect 17374 434 17402 439
rect 17374 56 17402 406
rect 17598 56 17626 854
rect 17878 881 17906 887
rect 17878 855 17879 881
rect 17905 855 17906 881
rect 17654 826 17682 831
rect 17654 601 17682 798
rect 17654 575 17655 601
rect 17681 575 17682 601
rect 17654 569 17682 575
rect 17878 378 17906 855
rect 17934 490 17962 495
rect 17934 443 17962 462
rect 17878 345 17906 350
rect 17822 210 17850 215
rect 17822 56 17850 182
rect 18046 56 18074 1638
rect 18270 1633 18298 1638
rect 18494 1666 18522 5838
rect 18830 5194 18858 5199
rect 18998 5194 19026 5199
rect 18830 5193 19026 5194
rect 18830 5167 18831 5193
rect 18857 5167 18999 5193
rect 19025 5167 19026 5193
rect 18830 5166 19026 5167
rect 18718 4074 18746 4079
rect 18550 3906 18578 3911
rect 18550 3010 18578 3878
rect 18550 3009 18690 3010
rect 18550 2983 18551 3009
rect 18577 2983 18690 3009
rect 18550 2982 18690 2983
rect 18550 2977 18578 2982
rect 18662 2953 18690 2982
rect 18662 2927 18663 2953
rect 18689 2927 18690 2953
rect 18662 2921 18690 2927
rect 18494 1633 18522 1638
rect 18606 2618 18634 2623
rect 18158 1386 18186 1391
rect 18158 1339 18186 1358
rect 18494 1386 18522 1391
rect 18494 1218 18522 1358
rect 18494 1185 18522 1190
rect 18550 1329 18578 1335
rect 18550 1303 18551 1329
rect 18577 1303 18578 1329
rect 18494 1106 18522 1111
rect 18382 994 18410 999
rect 18382 947 18410 966
rect 18270 546 18298 551
rect 18270 56 18298 518
rect 18494 56 18522 1078
rect 18550 882 18578 1303
rect 18550 849 18578 854
rect 18550 602 18578 607
rect 18606 602 18634 2590
rect 18718 2338 18746 4046
rect 18830 3962 18858 5166
rect 18998 5161 19026 5166
rect 18830 3929 18858 3934
rect 18830 3570 18858 3575
rect 18718 2305 18746 2310
rect 18774 2450 18802 2455
rect 18774 1833 18802 2422
rect 18774 1807 18775 1833
rect 18801 1807 18802 1833
rect 18774 1801 18802 1807
rect 18830 1554 18858 3542
rect 18942 2898 18970 2903
rect 18942 2897 19026 2898
rect 18942 2871 18943 2897
rect 18969 2871 19026 2897
rect 18942 2870 19026 2871
rect 18942 2865 18970 2870
rect 18886 2114 18914 2119
rect 18886 1946 18914 2086
rect 18886 1913 18914 1918
rect 18830 1521 18858 1526
rect 18998 994 19026 2870
rect 19054 1610 19082 5950
rect 19670 5362 19698 5367
rect 19278 5306 19306 5311
rect 19278 5259 19306 5278
rect 19446 2898 19474 2903
rect 19110 2561 19138 2567
rect 19110 2535 19111 2561
rect 19137 2535 19138 2561
rect 19110 2506 19138 2535
rect 19110 2473 19138 2478
rect 19278 2561 19306 2567
rect 19278 2535 19279 2561
rect 19305 2535 19306 2561
rect 19278 2506 19306 2535
rect 19278 2473 19306 2478
rect 19054 1577 19082 1582
rect 19110 1721 19138 1727
rect 19110 1695 19111 1721
rect 19137 1695 19138 1721
rect 19054 1441 19082 1447
rect 19054 1415 19055 1441
rect 19081 1415 19082 1441
rect 19054 1106 19082 1415
rect 19054 1073 19082 1078
rect 19054 994 19082 999
rect 18998 993 19082 994
rect 18998 967 19055 993
rect 19081 967 19082 993
rect 18998 966 19082 967
rect 19054 961 19082 966
rect 18550 601 18634 602
rect 18550 575 18551 601
rect 18577 575 18634 601
rect 18550 574 18634 575
rect 18662 881 18690 887
rect 18662 855 18663 881
rect 18689 855 18690 881
rect 18550 569 18578 574
rect 18662 210 18690 855
rect 19110 546 19138 1695
rect 19334 1666 19362 1671
rect 19334 1106 19362 1638
rect 19446 1385 19474 2870
rect 19558 2561 19586 2567
rect 19558 2535 19559 2561
rect 19585 2535 19586 2561
rect 19558 2450 19586 2535
rect 19558 2417 19586 2422
rect 19558 2226 19586 2231
rect 19502 2058 19530 2063
rect 19502 2011 19530 2030
rect 19558 1833 19586 2198
rect 19614 2058 19642 2063
rect 19614 2011 19642 2030
rect 19558 1807 19559 1833
rect 19585 1807 19586 1833
rect 19558 1801 19586 1807
rect 19446 1359 19447 1385
rect 19473 1359 19474 1385
rect 19446 1353 19474 1359
rect 19166 1105 19362 1106
rect 19166 1079 19335 1105
rect 19361 1079 19362 1105
rect 19166 1078 19362 1079
rect 19166 657 19194 1078
rect 19334 1073 19362 1078
rect 19614 994 19642 999
rect 19614 947 19642 966
rect 19166 631 19167 657
rect 19193 631 19194 657
rect 19166 625 19194 631
rect 19614 882 19642 887
rect 18774 518 19138 546
rect 18718 490 18746 495
rect 18718 443 18746 462
rect 18774 378 18802 518
rect 18662 177 18690 182
rect 18718 350 18802 378
rect 19166 378 19194 383
rect 18718 56 18746 350
rect 18942 266 18970 271
rect 18942 56 18970 238
rect 19166 56 19194 350
rect 19390 322 19418 327
rect 19390 56 19418 294
rect 19614 56 19642 854
rect 19670 714 19698 5334
rect 20454 4466 20482 4471
rect 20454 4419 20482 4438
rect 20342 3178 20370 3183
rect 20286 2898 20314 2903
rect 20286 2851 20314 2870
rect 19894 2842 19922 2847
rect 20006 2842 20034 2847
rect 19894 2841 20034 2842
rect 19894 2815 19895 2841
rect 19921 2815 20007 2841
rect 20033 2815 20034 2841
rect 19894 2814 20034 2815
rect 19894 2226 19922 2814
rect 20006 2809 20034 2814
rect 19782 2198 19922 2226
rect 19726 826 19754 831
rect 19782 826 19810 2198
rect 19894 2114 19922 2119
rect 19894 2113 20034 2114
rect 19894 2087 19895 2113
rect 19921 2087 20034 2113
rect 19894 2086 20034 2087
rect 19894 2081 19922 2086
rect 19950 1329 19978 1335
rect 19950 1303 19951 1329
rect 19977 1303 19978 1329
rect 19894 1218 19922 1223
rect 19754 798 19810 826
rect 19838 826 19866 831
rect 19726 793 19754 798
rect 19670 686 19754 714
rect 19726 98 19754 686
rect 19782 546 19810 551
rect 19782 499 19810 518
rect 19726 65 19754 70
rect 19838 56 19866 798
rect 19894 770 19922 1190
rect 19894 737 19922 742
rect 19950 378 19978 1303
rect 20006 602 20034 2086
rect 20286 1721 20314 1727
rect 20286 1695 20287 1721
rect 20313 1695 20314 1721
rect 20230 881 20258 887
rect 20230 855 20231 881
rect 20257 855 20258 881
rect 20062 602 20090 607
rect 20006 601 20090 602
rect 20006 575 20063 601
rect 20089 575 20090 601
rect 20006 574 20090 575
rect 20062 569 20090 574
rect 19950 345 19978 350
rect 20062 490 20090 495
rect 20062 56 20090 462
rect 20230 322 20258 855
rect 20286 826 20314 1695
rect 20342 1385 20370 3150
rect 20510 2450 20538 6454
rect 20566 4466 20594 4471
rect 20566 4419 20594 4438
rect 20846 4466 20874 4471
rect 20846 4419 20874 4438
rect 21182 4466 21210 4471
rect 20510 2417 20538 2422
rect 20790 3346 20818 3351
rect 20622 2282 20650 2287
rect 20622 2226 20650 2254
rect 20622 2225 20762 2226
rect 20622 2199 20623 2225
rect 20649 2199 20762 2225
rect 20622 2198 20762 2199
rect 20622 2193 20650 2198
rect 20734 2169 20762 2198
rect 20734 2143 20735 2169
rect 20761 2143 20762 2169
rect 20734 2137 20762 2143
rect 20734 1834 20762 1839
rect 20790 1834 20818 3318
rect 20734 1833 20818 1834
rect 20734 1807 20735 1833
rect 20761 1807 20818 1833
rect 20734 1806 20818 1807
rect 20902 3066 20930 3071
rect 20902 1833 20930 3038
rect 21070 3010 21098 3015
rect 20958 2226 20986 2231
rect 20958 2179 20986 2198
rect 20902 1807 20903 1833
rect 20929 1807 20930 1833
rect 20734 1801 20762 1806
rect 20902 1801 20930 1807
rect 20678 1778 20706 1783
rect 20342 1359 20343 1385
rect 20369 1359 20370 1385
rect 20342 1353 20370 1359
rect 20622 1441 20650 1447
rect 20622 1415 20623 1441
rect 20649 1415 20650 1441
rect 20286 793 20314 798
rect 20510 826 20538 831
rect 20454 657 20482 663
rect 20454 631 20455 657
rect 20481 631 20482 657
rect 20230 289 20258 294
rect 20286 546 20314 551
rect 20286 56 20314 518
rect 20454 266 20482 631
rect 20454 233 20482 238
rect 20510 56 20538 798
rect 20622 490 20650 1415
rect 20678 993 20706 1750
rect 20678 967 20679 993
rect 20705 967 20706 993
rect 20678 961 20706 967
rect 20790 1722 20818 1727
rect 20790 826 20818 1694
rect 21070 1385 21098 2982
rect 21126 2674 21154 2679
rect 21126 2627 21154 2646
rect 21182 2226 21210 4438
rect 21406 3066 21434 6622
rect 21574 6425 21602 6734
rect 22232 6678 22364 6683
rect 22260 6650 22284 6678
rect 22312 6650 22336 6678
rect 22232 6645 22364 6650
rect 22078 6482 22106 6487
rect 22078 6435 22106 6454
rect 21574 6399 21575 6425
rect 21601 6399 21602 6425
rect 21574 6393 21602 6399
rect 22582 6425 22610 7014
rect 23758 7042 23786 7056
rect 23758 7009 23786 7014
rect 23982 7042 24010 7047
rect 23254 6594 23282 6599
rect 22582 6399 22583 6425
rect 22609 6399 22610 6425
rect 22582 6393 22610 6399
rect 23086 6481 23114 6487
rect 23086 6455 23087 6481
rect 23113 6455 23114 6481
rect 21902 6286 22034 6291
rect 21930 6258 21954 6286
rect 21982 6258 22006 6286
rect 21902 6253 22034 6258
rect 22414 6034 22442 6039
rect 22302 5978 22330 5997
rect 22302 5945 22330 5950
rect 22232 5894 22364 5899
rect 22134 5866 22162 5871
rect 22260 5866 22284 5894
rect 22312 5866 22336 5894
rect 22232 5861 22364 5866
rect 21902 5502 22034 5507
rect 21930 5474 21954 5502
rect 21982 5474 22006 5502
rect 21902 5469 22034 5474
rect 22134 5362 22162 5838
rect 22134 5329 22162 5334
rect 22232 5110 22364 5115
rect 22260 5082 22284 5110
rect 22312 5082 22336 5110
rect 22232 5077 22364 5082
rect 21902 4718 22034 4723
rect 21930 4690 21954 4718
rect 21982 4690 22006 4718
rect 21902 4685 22034 4690
rect 22358 4466 22386 4471
rect 22358 4419 22386 4438
rect 21854 4410 21882 4415
rect 22078 4410 22106 4415
rect 21882 4409 22106 4410
rect 21882 4383 22079 4409
rect 22105 4383 22106 4409
rect 21882 4382 22106 4383
rect 21854 4363 21882 4382
rect 22078 4377 22106 4382
rect 22232 4326 22364 4331
rect 22260 4298 22284 4326
rect 22312 4298 22336 4326
rect 22232 4293 22364 4298
rect 21798 4129 21826 4135
rect 21798 4103 21799 4129
rect 21825 4103 21826 4129
rect 21630 4074 21658 4079
rect 21630 4027 21658 4046
rect 21798 4074 21826 4103
rect 21798 4041 21826 4046
rect 22078 4074 22106 4079
rect 22078 4027 22106 4046
rect 21902 3934 22034 3939
rect 21930 3906 21954 3934
rect 21982 3906 22006 3934
rect 21902 3901 22034 3906
rect 21910 3850 21938 3855
rect 22134 3850 22162 3855
rect 21630 3345 21658 3351
rect 21630 3319 21631 3345
rect 21657 3319 21658 3345
rect 21462 3290 21490 3295
rect 21630 3290 21658 3319
rect 21462 3289 21658 3290
rect 21462 3263 21463 3289
rect 21489 3263 21658 3289
rect 21462 3262 21658 3263
rect 21854 3289 21882 3295
rect 21854 3263 21855 3289
rect 21881 3263 21882 3289
rect 21462 3122 21490 3262
rect 21854 3234 21882 3263
rect 21910 3290 21938 3822
rect 21966 3822 22134 3850
rect 21966 3402 21994 3822
rect 22134 3817 22162 3822
rect 21966 3369 21994 3374
rect 22134 3570 22162 3575
rect 21910 3262 22106 3290
rect 21798 3206 21882 3234
rect 21798 3178 21826 3206
rect 21798 3145 21826 3150
rect 21902 3150 22034 3155
rect 21930 3122 21954 3150
rect 21982 3122 22006 3150
rect 21902 3117 22034 3122
rect 21462 3089 21490 3094
rect 21406 3033 21434 3038
rect 21294 2674 21322 2679
rect 21294 2627 21322 2646
rect 21182 2193 21210 2198
rect 21574 2505 21602 2511
rect 21574 2479 21575 2505
rect 21601 2479 21602 2505
rect 21182 1722 21210 1727
rect 21182 1675 21210 1694
rect 21462 1722 21490 1727
rect 21070 1359 21071 1385
rect 21097 1359 21098 1385
rect 21070 1353 21098 1359
rect 21070 1274 21098 1279
rect 21014 882 21042 887
rect 21014 835 21042 854
rect 20622 457 20650 462
rect 20734 798 20818 826
rect 20734 56 20762 798
rect 20958 770 20986 775
rect 20958 601 20986 742
rect 20958 575 20959 601
rect 20985 575 20986 601
rect 20958 569 20986 575
rect 20958 434 20986 439
rect 20958 56 20986 406
rect 21070 210 21098 1246
rect 21350 1273 21378 1279
rect 21350 1247 21351 1273
rect 21377 1247 21378 1273
rect 21350 1218 21378 1247
rect 21350 1185 21378 1190
rect 21070 177 21098 182
rect 21182 994 21210 999
rect 21182 56 21210 966
rect 21462 993 21490 1694
rect 21518 1273 21546 1279
rect 21518 1247 21519 1273
rect 21545 1247 21546 1273
rect 21518 1218 21546 1247
rect 21518 1185 21546 1190
rect 21462 967 21463 993
rect 21489 967 21490 993
rect 21462 961 21490 967
rect 21574 770 21602 2479
rect 21686 2394 21714 2399
rect 21686 1833 21714 2366
rect 21902 2366 22034 2371
rect 21930 2338 21954 2366
rect 21982 2338 22006 2366
rect 21902 2333 22034 2338
rect 21686 1807 21687 1833
rect 21713 1807 21714 1833
rect 21686 1801 21714 1807
rect 21902 1582 22034 1587
rect 21930 1554 21954 1582
rect 21982 1554 22006 1582
rect 21902 1549 22034 1554
rect 22022 1498 22050 1503
rect 21798 1329 21826 1335
rect 21798 1303 21799 1329
rect 21825 1303 21826 1329
rect 21686 993 21714 999
rect 21686 967 21687 993
rect 21713 967 21714 993
rect 21686 938 21714 967
rect 21686 905 21714 910
rect 21574 737 21602 742
rect 21630 714 21658 719
rect 21798 714 21826 1303
rect 22022 938 22050 1470
rect 22078 1385 22106 3262
rect 22134 3122 22162 3542
rect 22232 3542 22364 3547
rect 22260 3514 22284 3542
rect 22312 3514 22336 3542
rect 22232 3509 22364 3514
rect 22414 3514 22442 6006
rect 22470 5978 22498 5983
rect 22638 5978 22666 5983
rect 22470 5977 22666 5978
rect 22470 5951 22471 5977
rect 22497 5951 22639 5977
rect 22665 5951 22666 5977
rect 22470 5950 22666 5951
rect 22470 5945 22498 5950
rect 22414 3481 22442 3486
rect 22470 5362 22498 5367
rect 22414 3345 22442 3351
rect 22414 3319 22415 3345
rect 22441 3319 22442 3345
rect 22134 3089 22162 3094
rect 22246 3290 22274 3295
rect 22414 3290 22442 3319
rect 22246 3289 22442 3290
rect 22246 3263 22247 3289
rect 22273 3263 22442 3289
rect 22246 3262 22442 3263
rect 22246 2842 22274 3262
rect 22134 2814 22274 2842
rect 22134 1890 22162 2814
rect 22232 2758 22364 2763
rect 22260 2730 22284 2758
rect 22312 2730 22336 2758
rect 22232 2725 22364 2730
rect 22470 2338 22498 5334
rect 22470 2305 22498 2310
rect 22358 2170 22386 2175
rect 22358 2123 22386 2142
rect 22470 2170 22498 2175
rect 22470 2123 22498 2142
rect 22232 1974 22364 1979
rect 22260 1946 22284 1974
rect 22312 1946 22336 1974
rect 22232 1941 22364 1946
rect 22134 1862 22218 1890
rect 22078 1359 22079 1385
rect 22105 1359 22106 1385
rect 22078 1353 22106 1359
rect 22134 1721 22162 1727
rect 22134 1695 22135 1721
rect 22161 1695 22162 1721
rect 22022 905 22050 910
rect 21966 882 21994 901
rect 21966 849 21994 854
rect 21902 798 22034 803
rect 21930 770 21954 798
rect 21982 770 22006 798
rect 21902 765 22034 770
rect 22078 770 22106 775
rect 21798 686 21882 714
rect 21406 434 21434 439
rect 21406 56 21434 406
rect 21630 56 21658 686
rect 21686 546 21714 551
rect 21686 499 21714 518
rect 21854 546 21882 686
rect 22078 601 22106 742
rect 22078 575 22079 601
rect 22105 575 22106 601
rect 22078 569 22106 575
rect 21854 513 21882 518
rect 22134 434 22162 1695
rect 22190 1498 22218 1862
rect 22470 1834 22498 1839
rect 22470 1787 22498 1806
rect 22638 1666 22666 5950
rect 22974 4466 23002 4471
rect 22750 4074 22778 4079
rect 22694 3346 22722 3351
rect 22694 3299 22722 3318
rect 22750 2786 22778 4046
rect 22974 3906 23002 4438
rect 23086 4214 23114 6455
rect 23254 6146 23282 6566
rect 23646 6538 23674 6543
rect 23254 6145 23450 6146
rect 23254 6119 23255 6145
rect 23281 6119 23450 6145
rect 23254 6118 23450 6119
rect 23254 6113 23282 6118
rect 23422 6089 23450 6118
rect 23422 6063 23423 6089
rect 23449 6063 23450 6089
rect 23422 6057 23450 6063
rect 23534 5754 23562 5759
rect 23534 5641 23562 5726
rect 23534 5615 23535 5641
rect 23561 5615 23562 5641
rect 23534 5609 23562 5615
rect 23646 4214 23674 6510
rect 23982 6425 24010 7014
rect 25102 7042 25130 7056
rect 25102 7009 25130 7014
rect 25382 7042 25410 7047
rect 24990 6818 25018 6823
rect 23982 6399 23983 6425
rect 24009 6399 24010 6425
rect 23982 6393 24010 6399
rect 24486 6481 24514 6487
rect 24486 6455 24487 6481
rect 24513 6455 24514 6481
rect 23702 6034 23730 6039
rect 23702 5987 23730 6006
rect 23758 5697 23786 5703
rect 23758 5671 23759 5697
rect 23785 5671 23786 5697
rect 23758 5586 23786 5671
rect 24262 5698 24290 5703
rect 23982 5641 24010 5647
rect 23982 5615 23983 5641
rect 24009 5615 24010 5641
rect 23982 5586 24010 5615
rect 23758 5558 24010 5586
rect 23982 4214 24010 5558
rect 24206 4802 24234 4807
rect 24150 4634 24178 4639
rect 23086 4186 23450 4214
rect 23646 4186 23954 4214
rect 23982 4186 24122 4214
rect 22974 3873 23002 3878
rect 23366 4018 23394 4023
rect 23198 3122 23226 3127
rect 23198 3010 23226 3094
rect 23198 3009 23338 3010
rect 23198 2983 23199 3009
rect 23225 2983 23338 3009
rect 23198 2982 23338 2983
rect 23198 2977 23226 2982
rect 23310 2953 23338 2982
rect 23310 2927 23311 2953
rect 23337 2927 23338 2953
rect 23310 2921 23338 2927
rect 22750 2753 22778 2758
rect 23310 2674 23338 2679
rect 23310 2627 23338 2646
rect 22918 2618 22946 2623
rect 22750 2113 22778 2119
rect 22750 2087 22751 2113
rect 22777 2087 22778 2113
rect 22750 1778 22778 2087
rect 22750 1745 22778 1750
rect 22638 1633 22666 1638
rect 22806 1721 22834 1727
rect 22806 1695 22807 1721
rect 22833 1695 22834 1721
rect 22190 1465 22218 1470
rect 22414 1441 22442 1447
rect 22414 1415 22415 1441
rect 22441 1415 22442 1441
rect 22232 1190 22364 1195
rect 22260 1162 22284 1190
rect 22312 1162 22336 1190
rect 22232 1157 22364 1162
rect 22414 714 22442 1415
rect 22470 1386 22498 1391
rect 22470 1049 22498 1358
rect 22470 1023 22471 1049
rect 22497 1023 22498 1049
rect 22470 1017 22498 1023
rect 22750 994 22778 999
rect 22750 937 22778 966
rect 22750 911 22751 937
rect 22777 911 22778 937
rect 22750 905 22778 911
rect 22414 681 22442 686
rect 22246 602 22274 607
rect 22246 555 22274 574
rect 22526 490 22554 495
rect 22526 443 22554 462
rect 22750 434 22778 439
rect 22134 401 22162 406
rect 22232 406 22364 411
rect 22260 378 22284 406
rect 22312 378 22336 406
rect 22232 373 22364 378
rect 22302 322 22330 327
rect 21854 266 21882 271
rect 21854 56 21882 238
rect 22078 98 22106 103
rect 22078 56 22106 70
rect 22302 56 22330 294
rect 22526 210 22554 215
rect 22526 56 22554 182
rect 22750 56 22778 406
rect 22806 322 22834 1695
rect 22862 1330 22890 1335
rect 22862 1283 22890 1302
rect 22918 490 22946 2590
rect 23030 2506 23058 2511
rect 22918 457 22946 462
rect 22974 882 23002 887
rect 22806 289 22834 294
rect 22974 56 23002 854
rect 23030 770 23058 2478
rect 23366 2170 23394 3990
rect 23366 2137 23394 2142
rect 23142 2114 23170 2119
rect 23170 2086 23282 2114
rect 23142 2067 23170 2086
rect 23254 1889 23282 2086
rect 23310 2113 23338 2119
rect 23310 2087 23311 2113
rect 23337 2087 23338 2113
rect 23310 2058 23338 2087
rect 23310 2025 23338 2030
rect 23254 1863 23255 1889
rect 23281 1863 23282 1889
rect 23254 1857 23282 1863
rect 23198 1778 23226 1783
rect 23142 1274 23170 1279
rect 23030 737 23058 742
rect 23086 1273 23170 1274
rect 23086 1247 23143 1273
rect 23169 1247 23170 1273
rect 23086 1246 23170 1247
rect 23086 98 23114 1246
rect 23142 1241 23170 1246
rect 23086 65 23114 70
rect 23198 56 23226 1750
rect 23310 938 23338 943
rect 23422 938 23450 4186
rect 23758 3010 23786 3015
rect 23590 2897 23618 2903
rect 23590 2871 23591 2897
rect 23617 2871 23618 2897
rect 23478 2674 23506 2679
rect 23478 2627 23506 2646
rect 23590 2562 23618 2871
rect 23758 2617 23786 2982
rect 23758 2591 23759 2617
rect 23785 2591 23786 2617
rect 23758 2585 23786 2591
rect 23926 2618 23954 4186
rect 23926 2585 23954 2590
rect 24038 2842 24066 2847
rect 23590 2529 23618 2534
rect 23590 2057 23618 2063
rect 23590 2031 23591 2057
rect 23617 2031 23618 2057
rect 23590 1778 23618 2031
rect 23590 1745 23618 1750
rect 23478 1722 23506 1727
rect 23478 1675 23506 1694
rect 23870 1666 23898 1671
rect 23646 1442 23674 1447
rect 23646 1385 23674 1414
rect 23646 1359 23647 1385
rect 23673 1359 23674 1385
rect 23646 1353 23674 1359
rect 23310 937 23450 938
rect 23310 911 23311 937
rect 23337 911 23450 937
rect 23310 910 23450 911
rect 23534 993 23562 999
rect 23534 967 23535 993
rect 23561 967 23562 993
rect 23534 938 23562 967
rect 23646 938 23674 943
rect 23534 910 23646 938
rect 23310 905 23338 910
rect 23646 891 23674 910
rect 23422 602 23450 607
rect 23366 545 23394 551
rect 23366 519 23367 545
rect 23393 519 23394 545
rect 23366 154 23394 519
rect 23366 121 23394 126
rect 23422 56 23450 574
rect 23646 489 23674 495
rect 23646 463 23647 489
rect 23673 463 23674 489
rect 23646 266 23674 463
rect 23646 233 23674 238
rect 23646 154 23674 159
rect 23646 56 23674 126
rect 23870 56 23898 1638
rect 23926 1273 23954 1279
rect 23926 1247 23927 1273
rect 23953 1247 23954 1273
rect 23926 882 23954 1247
rect 24038 1049 24066 2814
rect 24038 1023 24039 1049
rect 24065 1023 24066 1049
rect 24038 1017 24066 1023
rect 23926 849 23954 854
rect 24094 56 24122 4186
rect 24150 1833 24178 4606
rect 24150 1807 24151 1833
rect 24177 1807 24178 1833
rect 24150 1801 24178 1807
rect 24206 714 24234 4774
rect 24262 826 24290 5670
rect 24318 5250 24346 5255
rect 24318 3682 24346 5222
rect 24486 4214 24514 6455
rect 24542 6482 24570 6487
rect 24542 5362 24570 6454
rect 24990 6145 25018 6790
rect 25382 6425 25410 7014
rect 26446 6594 26474 7056
rect 26558 6594 26586 6599
rect 26446 6593 26586 6594
rect 26446 6567 26559 6593
rect 26585 6567 26586 6593
rect 26446 6566 26586 6567
rect 26558 6561 26586 6566
rect 25886 6482 25914 6487
rect 26278 6482 26306 6487
rect 25886 6435 25914 6454
rect 26166 6481 26306 6482
rect 26166 6455 26279 6481
rect 26305 6455 26306 6481
rect 26166 6454 26306 6455
rect 25382 6399 25383 6425
rect 25409 6399 25410 6425
rect 25382 6393 25410 6399
rect 24990 6119 24991 6145
rect 25017 6119 25018 6145
rect 24990 6113 25018 6119
rect 26110 6089 26138 6095
rect 26110 6063 26111 6089
rect 26137 6063 26138 6089
rect 25494 6034 25522 6039
rect 24654 5978 24682 5983
rect 24766 5978 24794 5983
rect 24654 5977 24794 5978
rect 24654 5951 24655 5977
rect 24681 5951 24767 5977
rect 24793 5951 24794 5977
rect 24654 5950 24794 5951
rect 24654 5945 24682 5950
rect 24542 5329 24570 5334
rect 24486 4186 24570 4214
rect 24318 3649 24346 3654
rect 24486 3850 24514 3855
rect 24374 2282 24402 2287
rect 24262 793 24290 798
rect 24318 1666 24346 1671
rect 24206 681 24234 686
rect 24150 658 24178 663
rect 24150 601 24178 630
rect 24150 575 24151 601
rect 24177 575 24178 601
rect 24150 569 24178 575
rect 24318 56 24346 1638
rect 24374 1386 24402 2254
rect 24430 1777 24458 1783
rect 24430 1751 24431 1777
rect 24457 1751 24458 1777
rect 24430 1722 24458 1751
rect 24430 1689 24458 1694
rect 24374 1353 24402 1358
rect 24486 1385 24514 3822
rect 24542 1834 24570 4186
rect 24598 2954 24626 2959
rect 24598 2907 24626 2926
rect 24710 2954 24738 2959
rect 24710 2907 24738 2926
rect 24710 2338 24738 2343
rect 24598 2058 24626 2063
rect 24598 2057 24682 2058
rect 24598 2031 24599 2057
rect 24625 2031 24682 2057
rect 24598 2030 24682 2031
rect 24598 2025 24626 2030
rect 24598 1834 24626 1839
rect 24542 1833 24626 1834
rect 24542 1807 24599 1833
rect 24625 1807 24626 1833
rect 24542 1806 24626 1807
rect 24598 1801 24626 1806
rect 24654 1722 24682 2030
rect 24654 1689 24682 1694
rect 24710 1554 24738 2310
rect 24766 1666 24794 5950
rect 25270 5922 25298 5927
rect 25046 5642 25074 5647
rect 24990 2898 25018 2903
rect 24990 2851 25018 2870
rect 24990 1946 25018 1951
rect 24766 1633 24794 1638
rect 24822 1890 24850 1895
rect 24710 1526 24794 1554
rect 24486 1359 24487 1385
rect 24513 1359 24514 1385
rect 24486 1353 24514 1359
rect 24710 1273 24738 1279
rect 24710 1247 24711 1273
rect 24737 1247 24738 1273
rect 24374 937 24402 943
rect 24374 911 24375 937
rect 24401 911 24402 937
rect 24374 434 24402 911
rect 24710 602 24738 1247
rect 24710 569 24738 574
rect 24374 401 24402 406
rect 24430 489 24458 495
rect 24430 463 24431 489
rect 24457 463 24458 489
rect 24430 210 24458 463
rect 24430 177 24458 182
rect 24542 490 24570 495
rect 24542 56 24570 462
rect 24766 56 24794 1526
rect 24822 1049 24850 1862
rect 24878 1890 24906 1895
rect 24990 1890 25018 1918
rect 24878 1889 25018 1890
rect 24878 1863 24879 1889
rect 24905 1863 24991 1889
rect 25017 1863 25018 1889
rect 24878 1862 25018 1863
rect 24878 1857 24906 1862
rect 24990 1857 25018 1862
rect 24822 1023 24823 1049
rect 24849 1023 24850 1049
rect 24822 1017 24850 1023
rect 24990 826 25018 831
rect 24990 56 25018 798
rect 25046 770 25074 5614
rect 25158 4858 25186 4863
rect 25158 3010 25186 4830
rect 25270 4522 25298 5894
rect 25494 5753 25522 6006
rect 25494 5727 25495 5753
rect 25521 5727 25522 5753
rect 25494 5721 25522 5727
rect 25886 5754 25914 5759
rect 25886 5707 25914 5726
rect 25270 4489 25298 4494
rect 25718 5418 25746 5423
rect 25214 4466 25242 4471
rect 25214 3794 25242 4438
rect 25214 3761 25242 3766
rect 25158 2977 25186 2982
rect 25046 737 25074 742
rect 25102 2618 25130 2623
rect 25102 98 25130 2590
rect 25494 2562 25522 2567
rect 25382 1890 25410 1895
rect 25382 1833 25410 1862
rect 25382 1807 25383 1833
rect 25409 1807 25410 1833
rect 25382 1801 25410 1807
rect 25326 1274 25354 1279
rect 25326 1227 25354 1246
rect 25438 1274 25466 1279
rect 25438 1227 25466 1246
rect 25270 937 25298 943
rect 25270 911 25271 937
rect 25297 911 25298 937
rect 25270 154 25298 911
rect 25270 121 25298 126
rect 25438 770 25466 775
rect 25102 65 25130 70
rect 25214 98 25242 103
rect 25214 56 25242 70
rect 25438 56 25466 742
rect 25494 601 25522 2534
rect 25606 2450 25634 2455
rect 25606 1049 25634 2422
rect 25662 1778 25690 1783
rect 25662 1731 25690 1750
rect 25718 1666 25746 5390
rect 25830 5362 25858 5367
rect 25774 2057 25802 2063
rect 25774 2031 25775 2057
rect 25801 2031 25802 2057
rect 25774 1778 25802 2031
rect 25830 1833 25858 5334
rect 26054 5305 26082 5311
rect 26054 5279 26055 5305
rect 26081 5279 26082 5305
rect 26054 5194 26082 5279
rect 26054 5161 26082 5166
rect 26110 5138 26138 6063
rect 26110 5105 26138 5110
rect 26166 2617 26194 6454
rect 26278 6449 26306 6454
rect 26334 6482 26362 6487
rect 26222 5586 26250 5591
rect 26222 4802 26250 5558
rect 26278 4970 26306 4975
rect 26278 4923 26306 4942
rect 26222 4769 26250 4774
rect 26166 2591 26167 2617
rect 26193 2591 26194 2617
rect 26166 2585 26194 2591
rect 26278 4242 26306 4247
rect 26278 2114 26306 4214
rect 26334 2225 26362 6454
rect 27678 6481 27706 6487
rect 27678 6455 27679 6481
rect 27705 6455 27706 6481
rect 27510 6426 27538 6431
rect 26502 6202 26530 6207
rect 26502 6155 26530 6174
rect 26782 6090 26810 6095
rect 26782 6043 26810 6062
rect 27174 6034 27202 6039
rect 27174 5987 27202 6006
rect 26390 5697 26418 5703
rect 26390 5671 26391 5697
rect 26417 5671 26418 5697
rect 26390 5026 26418 5671
rect 27062 5697 27090 5703
rect 27062 5671 27063 5697
rect 27089 5671 27090 5697
rect 26782 5585 26810 5591
rect 26782 5559 26783 5585
rect 26809 5559 26810 5585
rect 26782 5530 26810 5559
rect 26782 5497 26810 5502
rect 26502 5474 26530 5479
rect 26502 5417 26530 5446
rect 26502 5391 26503 5417
rect 26529 5391 26530 5417
rect 26502 5385 26530 5391
rect 27062 5306 27090 5671
rect 27062 5273 27090 5278
rect 27286 5361 27314 5367
rect 27286 5335 27287 5361
rect 27313 5335 27314 5361
rect 26782 5250 26810 5255
rect 26782 5203 26810 5222
rect 26390 4993 26418 4998
rect 26838 5138 26866 5143
rect 26782 4858 26810 4863
rect 26782 4811 26810 4830
rect 26782 4466 26810 4471
rect 26782 4419 26810 4438
rect 26782 3738 26810 3743
rect 26782 3691 26810 3710
rect 26726 3514 26754 3519
rect 26502 3290 26530 3295
rect 26502 3009 26530 3262
rect 26502 2983 26503 3009
rect 26529 2983 26530 3009
rect 26334 2199 26335 2225
rect 26361 2199 26362 2225
rect 26334 2193 26362 2199
rect 26390 2898 26418 2903
rect 26278 2086 26362 2114
rect 26110 2058 26138 2063
rect 26110 2011 26138 2030
rect 26222 2057 26250 2063
rect 26222 2031 26223 2057
rect 26249 2031 26250 2057
rect 25830 1807 25831 1833
rect 25857 1807 25858 1833
rect 25830 1801 25858 1807
rect 26110 1834 26138 1839
rect 26110 1787 26138 1806
rect 26222 1834 26250 2031
rect 26222 1801 26250 1806
rect 25774 1745 25802 1750
rect 26278 1777 26306 1783
rect 26278 1751 26279 1777
rect 26305 1751 26306 1777
rect 25606 1023 25607 1049
rect 25633 1023 25634 1049
rect 25606 1017 25634 1023
rect 25662 1638 25746 1666
rect 26222 1722 26250 1727
rect 25494 575 25495 601
rect 25521 575 25522 601
rect 25494 569 25522 575
rect 25662 56 25690 1638
rect 25718 1329 25746 1335
rect 25718 1303 25719 1329
rect 25745 1303 25746 1329
rect 25718 1050 25746 1303
rect 25998 1329 26026 1335
rect 25998 1303 25999 1329
rect 26025 1303 26026 1329
rect 25998 1106 26026 1303
rect 25998 1073 26026 1078
rect 25718 1017 25746 1022
rect 25886 993 25914 999
rect 25886 967 25887 993
rect 25913 967 25914 993
rect 25886 938 25914 967
rect 25998 938 26026 943
rect 25886 937 26026 938
rect 25886 911 25999 937
rect 26025 911 26026 937
rect 25886 910 26026 911
rect 25998 882 26026 910
rect 26222 882 26250 1694
rect 26278 994 26306 1751
rect 26278 961 26306 966
rect 26334 993 26362 2086
rect 26334 967 26335 993
rect 26361 967 26362 993
rect 26334 961 26362 967
rect 26222 854 26362 882
rect 25998 849 26026 854
rect 26110 714 26138 719
rect 25998 657 26026 663
rect 25998 631 25999 657
rect 26025 631 26026 657
rect 25998 490 26026 631
rect 25998 457 26026 462
rect 25886 98 25914 103
rect 25886 56 25914 70
rect 26110 56 26138 686
rect 26334 56 26362 854
rect 26390 601 26418 2870
rect 26446 2618 26474 2623
rect 26446 2571 26474 2590
rect 26502 2562 26530 2983
rect 26614 2841 26642 2847
rect 26614 2815 26615 2841
rect 26641 2815 26642 2841
rect 26614 2674 26642 2815
rect 26614 2641 26642 2646
rect 26614 2562 26642 2567
rect 26502 2561 26642 2562
rect 26502 2535 26615 2561
rect 26641 2535 26642 2561
rect 26502 2534 26642 2535
rect 26614 2529 26642 2534
rect 26614 2058 26642 2063
rect 26614 2011 26642 2030
rect 26558 1610 26586 1615
rect 26502 1442 26530 1447
rect 26502 1395 26530 1414
rect 26390 575 26391 601
rect 26417 575 26418 601
rect 26390 569 26418 575
rect 26558 56 26586 1582
rect 26726 602 26754 3486
rect 26782 3066 26810 3071
rect 26782 2953 26810 3038
rect 26782 2927 26783 2953
rect 26809 2927 26810 2953
rect 26782 2921 26810 2927
rect 26782 2170 26810 2175
rect 26782 2123 26810 2142
rect 26838 1890 26866 5110
rect 27286 5082 27314 5335
rect 27286 5049 27314 5054
rect 27062 4914 27090 4919
rect 27062 4867 27090 4886
rect 27118 4802 27146 4807
rect 27062 4129 27090 4135
rect 27062 4103 27063 4129
rect 27089 4103 27090 4129
rect 27062 3458 27090 4103
rect 27062 3425 27090 3430
rect 27062 3345 27090 3351
rect 27062 3319 27063 3345
rect 27089 3319 27090 3345
rect 27062 3234 27090 3319
rect 27062 3201 27090 3206
rect 27062 2786 27090 2791
rect 27062 2617 27090 2758
rect 27062 2591 27063 2617
rect 27089 2591 27090 2617
rect 27062 2585 27090 2591
rect 26894 2506 26922 2511
rect 26894 2459 26922 2478
rect 26838 1857 26866 1862
rect 27118 1777 27146 4774
rect 27174 4465 27202 4471
rect 27174 4439 27175 4465
rect 27201 4439 27202 4465
rect 27174 4298 27202 4439
rect 27174 4265 27202 4270
rect 27454 4186 27482 4191
rect 27454 4139 27482 4158
rect 27286 3793 27314 3799
rect 27286 3767 27287 3793
rect 27313 3767 27314 3793
rect 27286 3626 27314 3767
rect 27286 3593 27314 3598
rect 27286 3009 27314 3015
rect 27286 2983 27287 3009
rect 27313 2983 27314 3009
rect 27286 2954 27314 2983
rect 27286 2921 27314 2926
rect 27454 2562 27482 2567
rect 27454 2515 27482 2534
rect 27286 2282 27314 2287
rect 27286 2235 27314 2254
rect 27118 1751 27119 1777
rect 27145 1751 27146 1777
rect 27118 1745 27146 1751
rect 27230 1834 27258 1839
rect 26782 1722 26810 1727
rect 26782 1675 26810 1694
rect 26782 1386 26810 1391
rect 26782 1339 26810 1358
rect 27062 1050 27090 1055
rect 27062 1003 27090 1022
rect 26782 938 26810 943
rect 26782 891 26810 910
rect 27006 882 27034 887
rect 26782 714 26810 719
rect 26782 667 26810 686
rect 26726 574 26810 602
rect 26782 56 26810 574
rect 27006 56 27034 854
rect 27230 56 27258 1806
rect 27454 1834 27482 1839
rect 27454 1787 27482 1806
rect 27286 1610 27314 1615
rect 27286 1497 27314 1582
rect 27286 1471 27287 1497
rect 27313 1471 27314 1497
rect 27286 1465 27314 1471
rect 27510 1386 27538 6398
rect 27566 6033 27594 6039
rect 27566 6007 27567 6033
rect 27593 6007 27594 6033
rect 27566 5922 27594 6007
rect 27566 5889 27594 5894
rect 27622 5810 27650 5815
rect 27566 5585 27594 5591
rect 27566 5559 27567 5585
rect 27593 5559 27594 5585
rect 27566 5418 27594 5559
rect 27566 5385 27594 5390
rect 27622 5305 27650 5782
rect 27622 5279 27623 5305
rect 27649 5279 27650 5305
rect 27622 5273 27650 5279
rect 27566 4801 27594 4807
rect 27566 4775 27567 4801
rect 27593 4775 27594 4801
rect 27566 4746 27594 4775
rect 27566 4713 27594 4718
rect 27678 4578 27706 6455
rect 27790 6202 27818 7056
rect 28182 6986 28210 6991
rect 27790 6169 27818 6174
rect 28070 6369 28098 6375
rect 28070 6343 28071 6369
rect 28097 6343 28098 6369
rect 27958 6033 27986 6039
rect 27958 6007 27959 6033
rect 27985 6007 27986 6033
rect 27958 5194 27986 6007
rect 28070 5642 28098 6343
rect 28182 5754 28210 6958
rect 28406 6762 28434 6767
rect 28182 5721 28210 5726
rect 28238 6090 28266 6095
rect 28070 5609 28098 5614
rect 28238 5530 28266 6062
rect 28238 5497 28266 5502
rect 27958 5161 27986 5166
rect 28070 5361 28098 5367
rect 28070 5335 28071 5361
rect 28097 5335 28098 5361
rect 27678 4545 27706 4550
rect 27622 4521 27650 4527
rect 27622 4495 27623 4521
rect 27649 4495 27650 4521
rect 27566 3906 27594 3911
rect 27566 3737 27594 3878
rect 27566 3711 27567 3737
rect 27593 3711 27594 3737
rect 27566 3705 27594 3711
rect 27622 3682 27650 4495
rect 28070 4522 28098 5335
rect 28406 4858 28434 6734
rect 28518 6538 28546 6543
rect 28462 6314 28490 6319
rect 28462 5474 28490 6286
rect 28462 5441 28490 5446
rect 28406 4825 28434 4830
rect 28070 4489 28098 4494
rect 27958 4465 27986 4471
rect 27958 4439 27959 4465
rect 27985 4439 27986 4465
rect 27958 4074 27986 4439
rect 28518 4186 28546 6510
rect 28518 4153 28546 4158
rect 27958 4041 27986 4046
rect 28070 3850 28098 3855
rect 28070 3803 28098 3822
rect 27622 3649 27650 3654
rect 28070 3402 28098 3407
rect 27566 3233 27594 3239
rect 27566 3207 27567 3233
rect 27593 3207 27594 3233
rect 27566 3178 27594 3207
rect 27566 3145 27594 3150
rect 28070 3065 28098 3374
rect 28070 3039 28071 3065
rect 28097 3039 28098 3065
rect 28070 3033 28098 3039
rect 27566 3010 27594 3015
rect 27566 2953 27594 2982
rect 27566 2927 27567 2953
rect 27593 2927 27594 2953
rect 27566 2921 27594 2927
rect 28070 2730 28098 2735
rect 28070 2281 28098 2702
rect 28070 2255 28071 2281
rect 28097 2255 28098 2281
rect 28070 2249 28098 2255
rect 28126 2618 28154 2623
rect 27566 2226 27594 2231
rect 27566 2169 27594 2198
rect 27566 2143 27567 2169
rect 27593 2143 27594 2169
rect 27566 2137 27594 2143
rect 27902 2058 27930 2063
rect 27678 1946 27706 1951
rect 27566 1386 27594 1391
rect 27510 1385 27594 1386
rect 27510 1359 27567 1385
rect 27593 1359 27594 1385
rect 27510 1358 27594 1359
rect 27566 1353 27594 1358
rect 27454 1162 27482 1167
rect 27454 1049 27482 1134
rect 27454 1023 27455 1049
rect 27481 1023 27482 1049
rect 27454 1017 27482 1023
rect 27398 994 27426 999
rect 27398 938 27426 966
rect 27398 910 27482 938
rect 27454 56 27482 910
rect 27566 546 27594 551
rect 27566 499 27594 518
rect 27678 56 27706 1918
rect 27902 56 27930 2030
rect 28070 2058 28098 2063
rect 28070 1497 28098 2030
rect 28070 1471 28071 1497
rect 28097 1471 28098 1497
rect 28070 1465 28098 1471
rect 28070 1386 28098 1391
rect 28070 713 28098 1358
rect 28070 687 28071 713
rect 28097 687 28098 713
rect 28070 681 28098 687
rect 28126 56 28154 2590
rect 28350 1778 28378 1783
rect 28350 56 28378 1750
rect 28462 1722 28490 1727
rect 28462 266 28490 1694
rect 28462 233 28490 238
rect 28518 1442 28546 1447
rect 462 9 490 14
rect 560 0 616 56
rect 784 0 840 56
rect 1008 0 1064 56
rect 1232 0 1288 56
rect 1456 0 1512 56
rect 1680 0 1736 56
rect 1904 0 1960 56
rect 2128 0 2184 56
rect 2352 0 2408 56
rect 2576 0 2632 56
rect 2800 0 2856 56
rect 3024 0 3080 56
rect 3248 0 3304 56
rect 3472 0 3528 56
rect 3696 0 3752 56
rect 3920 0 3976 56
rect 4144 0 4200 56
rect 4368 0 4424 56
rect 4592 0 4648 56
rect 4816 0 4872 56
rect 5040 0 5096 56
rect 5264 0 5320 56
rect 5488 0 5544 56
rect 5712 0 5768 56
rect 5936 0 5992 56
rect 6160 0 6216 56
rect 6384 0 6440 56
rect 6608 0 6664 56
rect 6832 0 6888 56
rect 7056 0 7112 56
rect 7280 0 7336 56
rect 7504 0 7560 56
rect 7728 0 7784 56
rect 7952 0 8008 56
rect 8176 0 8232 56
rect 8400 0 8456 56
rect 8624 0 8680 56
rect 8848 0 8904 56
rect 9072 0 9128 56
rect 9296 0 9352 56
rect 9520 0 9576 56
rect 9744 0 9800 56
rect 9968 0 10024 56
rect 10192 0 10248 56
rect 10416 0 10472 56
rect 10640 0 10696 56
rect 10864 0 10920 56
rect 11088 0 11144 56
rect 11312 0 11368 56
rect 11536 0 11592 56
rect 11760 0 11816 56
rect 11984 0 12040 56
rect 12208 0 12264 56
rect 12432 0 12488 56
rect 12656 0 12712 56
rect 12880 0 12936 56
rect 13104 0 13160 56
rect 13328 0 13384 56
rect 13552 0 13608 56
rect 13776 0 13832 56
rect 14000 0 14056 56
rect 14224 0 14280 56
rect 14448 0 14504 56
rect 14672 0 14728 56
rect 14896 0 14952 56
rect 15120 0 15176 56
rect 15344 0 15400 56
rect 15568 0 15624 56
rect 15792 0 15848 56
rect 16016 0 16072 56
rect 16240 0 16296 56
rect 16464 0 16520 56
rect 16688 0 16744 56
rect 16912 0 16968 56
rect 17136 0 17192 56
rect 17360 0 17416 56
rect 17584 0 17640 56
rect 17808 0 17864 56
rect 18032 0 18088 56
rect 18256 0 18312 56
rect 18480 0 18536 56
rect 18704 0 18760 56
rect 18928 0 18984 56
rect 19152 0 19208 56
rect 19376 0 19432 56
rect 19600 0 19656 56
rect 19824 0 19880 56
rect 20048 0 20104 56
rect 20272 0 20328 56
rect 20496 0 20552 56
rect 20720 0 20776 56
rect 20944 0 21000 56
rect 21168 0 21224 56
rect 21392 0 21448 56
rect 21616 0 21672 56
rect 21840 0 21896 56
rect 22064 0 22120 56
rect 22288 0 22344 56
rect 22512 0 22568 56
rect 22736 0 22792 56
rect 22960 0 23016 56
rect 23184 0 23240 56
rect 23408 0 23464 56
rect 23632 0 23688 56
rect 23856 0 23912 56
rect 24080 0 24136 56
rect 24304 0 24360 56
rect 24528 0 24584 56
rect 24752 0 24808 56
rect 24976 0 25032 56
rect 25200 0 25256 56
rect 25424 0 25480 56
rect 25648 0 25704 56
rect 25872 0 25928 56
rect 26096 0 26152 56
rect 26320 0 26376 56
rect 26544 0 26600 56
rect 26768 0 26824 56
rect 26992 0 27048 56
rect 27216 0 27272 56
rect 27440 0 27496 56
rect 27664 0 27720 56
rect 27888 0 27944 56
rect 28112 0 28168 56
rect 28336 0 28392 56
rect 28518 42 28546 1414
rect 28518 9 28546 14
<< via2 >>
rect 2254 7014 2282 7042
rect 2534 7014 2562 7042
rect 2232 6677 2260 6678
rect 2232 6651 2233 6677
rect 2233 6651 2259 6677
rect 2259 6651 2260 6677
rect 2232 6650 2260 6651
rect 2284 6677 2312 6678
rect 2284 6651 2285 6677
rect 2285 6651 2311 6677
rect 2311 6651 2312 6677
rect 2284 6650 2312 6651
rect 2336 6677 2364 6678
rect 2336 6651 2337 6677
rect 2337 6651 2363 6677
rect 2363 6651 2364 6677
rect 2336 6650 2364 6651
rect 798 6510 826 6538
rect 406 6062 434 6090
rect 3542 6958 3570 6986
rect 1902 6285 1930 6286
rect 1902 6259 1903 6285
rect 1903 6259 1929 6285
rect 1929 6259 1930 6285
rect 1902 6258 1930 6259
rect 1954 6285 1982 6286
rect 1954 6259 1955 6285
rect 1955 6259 1981 6285
rect 1981 6259 1982 6285
rect 1954 6258 1982 6259
rect 2006 6285 2034 6286
rect 2006 6259 2007 6285
rect 2007 6259 2033 6285
rect 2033 6259 2034 6285
rect 2006 6258 2034 6259
rect 2232 5893 2260 5894
rect 2232 5867 2233 5893
rect 2233 5867 2259 5893
rect 2259 5867 2260 5893
rect 2232 5866 2260 5867
rect 2284 5893 2312 5894
rect 2284 5867 2285 5893
rect 2285 5867 2311 5893
rect 2311 5867 2312 5893
rect 2284 5866 2312 5867
rect 2336 5893 2364 5894
rect 2336 5867 2337 5893
rect 2337 5867 2363 5893
rect 2363 5867 2364 5893
rect 2336 5866 2364 5867
rect 3486 6454 3514 6482
rect 3374 6174 3402 6202
rect 3374 5838 3402 5866
rect 3430 6006 3458 6034
rect 3038 5726 3066 5754
rect 1190 5558 1218 5586
rect 3374 5614 3402 5642
rect 1902 5501 1930 5502
rect 1902 5475 1903 5501
rect 1903 5475 1929 5501
rect 1929 5475 1930 5501
rect 1902 5474 1930 5475
rect 1954 5501 1982 5502
rect 1954 5475 1955 5501
rect 1955 5475 1981 5501
rect 1981 5475 1982 5501
rect 1954 5474 1982 5475
rect 2006 5501 2034 5502
rect 2006 5475 2007 5501
rect 2007 5475 2033 5501
rect 2033 5475 2034 5501
rect 2006 5474 2034 5475
rect 2926 5502 2954 5530
rect 798 5278 826 5306
rect 406 5222 434 5250
rect 798 5166 826 5194
rect 574 4942 602 4970
rect 294 4158 322 4186
rect 70 2702 98 2730
rect 126 1638 154 1666
rect 574 3710 602 3738
rect 742 4606 770 4634
rect 2232 5109 2260 5110
rect 2232 5083 2233 5109
rect 2233 5083 2259 5109
rect 2259 5083 2260 5109
rect 2232 5082 2260 5083
rect 2284 5109 2312 5110
rect 2284 5083 2285 5109
rect 2285 5083 2311 5109
rect 2311 5083 2312 5109
rect 2284 5082 2312 5083
rect 2336 5109 2364 5110
rect 2336 5083 2337 5109
rect 2337 5083 2363 5109
rect 2363 5083 2364 5109
rect 2336 5082 2364 5083
rect 2086 4830 2114 4858
rect 1902 4717 1930 4718
rect 1902 4691 1903 4717
rect 1903 4691 1929 4717
rect 1929 4691 1930 4717
rect 1902 4690 1930 4691
rect 1954 4717 1982 4718
rect 1954 4691 1955 4717
rect 1955 4691 1981 4717
rect 1981 4691 1982 4717
rect 1954 4690 1982 4691
rect 2006 4717 2034 4718
rect 2006 4691 2007 4717
rect 2007 4691 2033 4717
rect 2033 4691 2034 4717
rect 2006 4690 2034 4691
rect 798 4550 826 4578
rect 1470 4465 1498 4466
rect 1470 4439 1471 4465
rect 1471 4439 1497 4465
rect 1497 4439 1498 4465
rect 1470 4438 1498 4439
rect 742 3374 770 3402
rect 294 462 322 490
rect 350 2870 378 2898
rect 1022 2814 1050 2842
rect 518 2534 546 2562
rect 518 1358 546 1386
rect 798 1302 826 1330
rect 574 798 602 826
rect 462 462 490 490
rect 854 1049 882 1050
rect 854 1023 855 1049
rect 855 1023 881 1049
rect 881 1023 882 1049
rect 854 1022 882 1023
rect 1806 3990 1834 4018
rect 1358 2982 1386 3010
rect 1302 1862 1330 1890
rect 1078 910 1106 938
rect 1134 70 1162 98
rect 1470 2142 1498 2170
rect 1750 1750 1778 1778
rect 1902 3933 1930 3934
rect 1902 3907 1903 3933
rect 1903 3907 1929 3933
rect 1929 3907 1930 3933
rect 1902 3906 1930 3907
rect 1954 3933 1982 3934
rect 1954 3907 1955 3933
rect 1955 3907 1981 3933
rect 1981 3907 1982 3933
rect 1954 3906 1982 3907
rect 2006 3933 2034 3934
rect 2006 3907 2007 3933
rect 2007 3907 2033 3933
rect 2033 3907 2034 3933
rect 2006 3906 2034 3907
rect 1902 3149 1930 3150
rect 1902 3123 1903 3149
rect 1903 3123 1929 3149
rect 1929 3123 1930 3149
rect 1902 3122 1930 3123
rect 1954 3149 1982 3150
rect 1954 3123 1955 3149
rect 1955 3123 1981 3149
rect 1981 3123 1982 3149
rect 1954 3122 1982 3123
rect 2006 3149 2034 3150
rect 2006 3123 2007 3149
rect 2007 3123 2033 3149
rect 2033 3123 2034 3149
rect 2006 3122 2034 3123
rect 1902 2365 1930 2366
rect 1902 2339 1903 2365
rect 1903 2339 1929 2365
rect 1929 2339 1930 2365
rect 1902 2338 1930 2339
rect 1954 2365 1982 2366
rect 1954 2339 1955 2365
rect 1955 2339 1981 2365
rect 1981 2339 1982 2365
rect 1954 2338 1982 2339
rect 2006 2365 2034 2366
rect 2006 2339 2007 2365
rect 2007 2339 2033 2365
rect 2033 2339 2034 2365
rect 2006 2338 2034 2339
rect 1902 1581 1930 1582
rect 1902 1555 1903 1581
rect 1903 1555 1929 1581
rect 1929 1555 1930 1581
rect 1902 1554 1930 1555
rect 1954 1581 1982 1582
rect 1954 1555 1955 1581
rect 1955 1555 1981 1581
rect 1981 1555 1982 1581
rect 1954 1554 1982 1555
rect 2006 1581 2034 1582
rect 2006 1555 2007 1581
rect 2007 1555 2033 1581
rect 2033 1555 2034 1581
rect 2006 1554 2034 1555
rect 1902 797 1930 798
rect 1902 771 1903 797
rect 1903 771 1929 797
rect 1929 771 1930 797
rect 1902 770 1930 771
rect 1954 797 1982 798
rect 1954 771 1955 797
rect 1955 771 1981 797
rect 1981 771 1982 797
rect 1954 770 1982 771
rect 2006 797 2034 798
rect 2006 771 2007 797
rect 2007 771 2033 797
rect 2033 771 2034 797
rect 2006 770 2034 771
rect 2232 4325 2260 4326
rect 2232 4299 2233 4325
rect 2233 4299 2259 4325
rect 2259 4299 2260 4325
rect 2232 4298 2260 4299
rect 2284 4325 2312 4326
rect 2284 4299 2285 4325
rect 2285 4299 2311 4325
rect 2311 4299 2312 4325
rect 2284 4298 2312 4299
rect 2336 4325 2364 4326
rect 2336 4299 2337 4325
rect 2337 4299 2363 4325
rect 2363 4299 2364 4325
rect 2336 4298 2364 4299
rect 2232 3541 2260 3542
rect 2232 3515 2233 3541
rect 2233 3515 2259 3541
rect 2259 3515 2260 3541
rect 2232 3514 2260 3515
rect 2284 3541 2312 3542
rect 2284 3515 2285 3541
rect 2285 3515 2311 3541
rect 2311 3515 2312 3541
rect 2284 3514 2312 3515
rect 2336 3541 2364 3542
rect 2336 3515 2337 3541
rect 2337 3515 2363 3541
rect 2363 3515 2364 3541
rect 2702 3542 2730 3570
rect 2336 3514 2364 3515
rect 2232 2757 2260 2758
rect 2232 2731 2233 2757
rect 2233 2731 2259 2757
rect 2259 2731 2260 2757
rect 2232 2730 2260 2731
rect 2284 2757 2312 2758
rect 2284 2731 2285 2757
rect 2285 2731 2311 2757
rect 2311 2731 2312 2757
rect 2284 2730 2312 2731
rect 2336 2757 2364 2758
rect 2336 2731 2337 2757
rect 2337 2731 2363 2757
rect 2363 2731 2364 2757
rect 2336 2730 2364 2731
rect 2232 1973 2260 1974
rect 2232 1947 2233 1973
rect 2233 1947 2259 1973
rect 2259 1947 2260 1973
rect 2232 1946 2260 1947
rect 2284 1973 2312 1974
rect 2284 1947 2285 1973
rect 2285 1947 2311 1973
rect 2311 1947 2312 1973
rect 2284 1946 2312 1947
rect 2336 1973 2364 1974
rect 2336 1947 2337 1973
rect 2337 1947 2363 1973
rect 2363 1947 2364 1973
rect 2336 1946 2364 1947
rect 2814 1974 2842 2002
rect 2232 1189 2260 1190
rect 2232 1163 2233 1189
rect 2233 1163 2259 1189
rect 2259 1163 2260 1189
rect 2232 1162 2260 1163
rect 2284 1189 2312 1190
rect 2284 1163 2285 1189
rect 2285 1163 2311 1189
rect 2311 1163 2312 1189
rect 2284 1162 2312 1163
rect 2336 1189 2364 1190
rect 2336 1163 2337 1189
rect 2337 1163 2363 1189
rect 2363 1163 2364 1189
rect 2336 1162 2364 1163
rect 2590 798 2618 826
rect 2142 742 2170 770
rect 2232 405 2260 406
rect 2232 379 2233 405
rect 2233 379 2259 405
rect 2259 379 2260 405
rect 2232 378 2260 379
rect 2284 405 2312 406
rect 2284 379 2285 405
rect 2285 379 2311 405
rect 2311 379 2312 405
rect 2284 378 2312 379
rect 2336 405 2364 406
rect 2336 379 2337 405
rect 2337 379 2363 405
rect 2363 379 2364 405
rect 2336 378 2364 379
rect 2366 294 2394 322
rect 3430 5390 3458 5418
rect 3374 4998 3402 5026
rect 3430 5054 3458 5082
rect 3430 4382 3458 4410
rect 3430 4214 3458 4242
rect 2982 3625 3010 3626
rect 2982 3599 2983 3625
rect 2983 3599 3009 3625
rect 3009 3599 3010 3625
rect 2982 3598 3010 3599
rect 3150 3625 3178 3626
rect 3150 3599 3151 3625
rect 3151 3599 3177 3625
rect 3177 3599 3178 3625
rect 3150 3598 3178 3599
rect 3374 3598 3402 3626
rect 3374 3094 3402 3122
rect 3430 2926 3458 2954
rect 2926 686 2954 714
rect 3038 2702 3066 2730
rect 3430 1750 3458 1778
rect 3374 966 3402 994
rect 3430 126 3458 154
rect 4942 7014 4970 7042
rect 5334 7014 5362 7042
rect 3654 6902 3682 6930
rect 3542 5446 3570 5474
rect 3542 3766 3570 3794
rect 3542 1806 3570 1834
rect 3598 2590 3626 2618
rect 3542 1526 3570 1554
rect 4046 6790 4074 6818
rect 5278 6566 5306 6594
rect 3878 6118 3906 6146
rect 3822 5222 3850 5250
rect 3710 2870 3738 2898
rect 3710 1638 3738 1666
rect 3766 2142 3794 2170
rect 3654 1470 3682 1498
rect 3598 1022 3626 1050
rect 3710 1414 3738 1442
rect 3542 294 3570 322
rect 3766 854 3794 882
rect 5110 5614 5138 5642
rect 4326 4942 4354 4970
rect 4270 4438 4298 4466
rect 4158 3710 4186 3738
rect 3878 2534 3906 2562
rect 3990 3654 4018 3682
rect 3822 686 3850 714
rect 3934 1022 3962 1050
rect 4270 2422 4298 2450
rect 4158 2310 4186 2338
rect 5054 4214 5082 4242
rect 4942 4046 4970 4074
rect 4830 3625 4858 3626
rect 4830 3599 4831 3625
rect 4831 3599 4857 3625
rect 4857 3599 4858 3625
rect 4830 3598 4858 3599
rect 4550 3430 4578 3458
rect 4998 3625 5026 3626
rect 4998 3599 4999 3625
rect 4999 3599 5025 3625
rect 5025 3599 5026 3625
rect 4998 3598 5026 3599
rect 4942 3262 4970 3290
rect 5166 4662 5194 4690
rect 5166 2982 5194 3010
rect 5222 3486 5250 3514
rect 5110 2702 5138 2730
rect 5166 2758 5194 2786
rect 5054 2366 5082 2394
rect 5110 2225 5138 2226
rect 5110 2199 5111 2225
rect 5111 2199 5137 2225
rect 5137 2199 5138 2225
rect 5110 2198 5138 2199
rect 4326 2030 4354 2058
rect 4550 1694 4578 1722
rect 3990 742 4018 770
rect 4158 1190 4186 1218
rect 4382 742 4410 770
rect 4998 937 5026 938
rect 4998 911 4999 937
rect 4999 911 5025 937
rect 5025 911 5026 937
rect 4998 910 5026 911
rect 4606 798 4634 826
rect 4830 798 4858 826
rect 5222 798 5250 826
rect 5054 294 5082 322
rect 6286 7014 6314 7042
rect 6510 7014 6538 7042
rect 8974 7014 9002 7042
rect 9198 7014 9226 7042
rect 8470 6846 8498 6874
rect 8414 6678 8442 6706
rect 5670 6342 5698 6370
rect 6846 6174 6874 6202
rect 6678 6062 6706 6090
rect 6622 6006 6650 6034
rect 6678 5782 6706 5810
rect 6846 5726 6874 5754
rect 7518 6398 7546 6426
rect 8190 6454 8218 6482
rect 6622 5110 6650 5138
rect 7406 5809 7434 5810
rect 7406 5783 7407 5809
rect 7407 5783 7433 5809
rect 7433 5783 7434 5809
rect 7406 5782 7434 5783
rect 7518 5809 7546 5810
rect 7518 5783 7519 5809
rect 7519 5783 7545 5809
rect 7545 5783 7546 5809
rect 7518 5782 7546 5783
rect 7182 4942 7210 4970
rect 7350 5390 7378 5418
rect 7126 4886 7154 4914
rect 6510 4438 6538 4466
rect 5446 2561 5474 2562
rect 5446 2535 5447 2561
rect 5447 2535 5473 2561
rect 5473 2535 5474 2561
rect 5446 2534 5474 2535
rect 5558 2561 5586 2562
rect 5558 2535 5559 2561
rect 5559 2535 5585 2561
rect 5585 2535 5586 2561
rect 5558 2534 5586 2535
rect 6454 2478 6482 2506
rect 5502 406 5530 434
rect 5726 1806 5754 1834
rect 5502 182 5530 210
rect 5894 1750 5922 1778
rect 6174 1862 6202 1890
rect 5950 1470 5978 1498
rect 7126 4270 7154 4298
rect 7182 4718 7210 4746
rect 7014 3150 7042 3178
rect 6510 2198 6538 2226
rect 6566 2814 6594 2842
rect 6958 2534 6986 2562
rect 6566 1526 6594 1554
rect 6622 2030 6650 2058
rect 6454 1134 6482 1162
rect 6398 686 6426 714
rect 6398 574 6426 602
rect 6734 1694 6762 1722
rect 6734 1358 6762 1386
rect 6678 742 6706 770
rect 6846 518 6874 546
rect 6958 350 6986 378
rect 7126 2478 7154 2506
rect 8134 5278 8162 5306
rect 7574 5222 7602 5250
rect 7518 5054 7546 5082
rect 7518 4942 7546 4970
rect 7574 4830 7602 4858
rect 7462 4382 7490 4410
rect 7462 4158 7490 4186
rect 7910 3822 7938 3850
rect 7350 3318 7378 3346
rect 7574 3598 7602 3626
rect 7182 2310 7210 2338
rect 7238 3206 7266 3234
rect 7182 1638 7210 1666
rect 7126 966 7154 994
rect 7014 294 7042 322
rect 7070 798 7098 826
rect 7126 238 7154 266
rect 7294 3094 7322 3122
rect 7350 3038 7378 3066
rect 7854 3430 7882 3458
rect 7574 2926 7602 2954
rect 7350 1862 7378 1890
rect 7462 1582 7490 1610
rect 7518 1190 7546 1218
rect 7630 2646 7658 2674
rect 7686 2702 7714 2730
rect 8078 3150 8106 3178
rect 7910 3094 7938 3122
rect 7854 1862 7882 1890
rect 7686 1190 7714 1218
rect 7966 1582 7994 1610
rect 7574 742 7602 770
rect 7518 574 7546 602
rect 7742 630 7770 658
rect 7294 294 7322 322
rect 8414 5782 8442 5810
rect 8358 5726 8386 5754
rect 9926 7014 9954 7042
rect 9702 6481 9730 6482
rect 9702 6455 9703 6481
rect 9703 6455 9729 6481
rect 9729 6455 9730 6481
rect 9702 6454 9730 6455
rect 9086 5753 9114 5754
rect 9086 5727 9087 5753
rect 9087 5727 9113 5753
rect 9113 5727 9114 5753
rect 9086 5726 9114 5727
rect 9366 5697 9394 5698
rect 9366 5671 9367 5697
rect 9367 5671 9393 5697
rect 9393 5671 9394 5697
rect 9366 5670 9394 5671
rect 9478 5697 9506 5698
rect 9478 5671 9479 5697
rect 9479 5671 9505 5697
rect 9505 5671 9506 5697
rect 9478 5670 9506 5671
rect 8470 5614 8498 5642
rect 8582 5502 8610 5530
rect 8414 5110 8442 5138
rect 8358 4606 8386 4634
rect 8470 4606 8498 4634
rect 8470 4438 8498 4466
rect 8190 3542 8218 3570
rect 8246 4270 8274 4298
rect 8190 2897 8218 2898
rect 8190 2871 8191 2897
rect 8191 2871 8217 2897
rect 8217 2871 8218 2897
rect 8190 2870 8218 2871
rect 9366 5446 9394 5474
rect 9198 4774 9226 4802
rect 8974 4662 9002 4690
rect 8806 4438 8834 4466
rect 8582 4326 8610 4354
rect 8302 2897 8330 2898
rect 8302 2871 8303 2897
rect 8303 2871 8329 2897
rect 8329 2871 8330 2897
rect 8302 2870 8330 2871
rect 8414 2646 8442 2674
rect 8302 2590 8330 2618
rect 8302 2422 8330 2450
rect 8470 2534 8498 2562
rect 8526 3094 8554 3122
rect 8918 3934 8946 3962
rect 8806 3486 8834 3514
rect 8918 3486 8946 3514
rect 8582 3038 8610 3066
rect 8862 2926 8890 2954
rect 8526 2254 8554 2282
rect 8358 2142 8386 2170
rect 8246 1022 8274 1050
rect 8470 1414 8498 1442
rect 8134 798 8162 826
rect 8414 854 8442 882
rect 8358 462 8386 490
rect 8414 126 8442 154
rect 8694 2702 8722 2730
rect 8694 2534 8722 2562
rect 8582 1414 8610 1442
rect 8694 2086 8722 2114
rect 8526 1329 8554 1330
rect 8526 1303 8527 1329
rect 8527 1303 8553 1329
rect 8553 1303 8554 1329
rect 8526 1302 8554 1303
rect 8638 294 8666 322
rect 8526 126 8554 154
rect 8190 70 8218 98
rect 8694 182 8722 210
rect 9198 4158 9226 4186
rect 9254 4073 9282 4074
rect 9254 4047 9255 4073
rect 9255 4047 9281 4073
rect 9281 4047 9282 4073
rect 9254 4046 9282 4047
rect 9254 3878 9282 3906
rect 9254 3318 9282 3346
rect 8974 2702 9002 2730
rect 9254 3094 9282 3122
rect 9142 2673 9170 2674
rect 9142 2647 9143 2673
rect 9143 2647 9169 2673
rect 9169 2647 9170 2673
rect 9142 2646 9170 2647
rect 9310 2673 9338 2674
rect 9310 2647 9311 2673
rect 9311 2647 9337 2673
rect 9337 2647 9338 2673
rect 9310 2646 9338 2647
rect 9254 2366 9282 2394
rect 9590 5166 9618 5194
rect 9870 5166 9898 5194
rect 9534 5110 9562 5138
rect 10318 6454 10346 6482
rect 11550 6734 11578 6762
rect 10766 6510 10794 6538
rect 12838 6846 12866 6874
rect 11662 6734 11690 6762
rect 12054 6734 12082 6762
rect 12232 6677 12260 6678
rect 12232 6651 12233 6677
rect 12233 6651 12259 6677
rect 12259 6651 12260 6677
rect 12232 6650 12260 6651
rect 12284 6677 12312 6678
rect 12284 6651 12285 6677
rect 12285 6651 12311 6677
rect 12311 6651 12312 6677
rect 12284 6650 12312 6651
rect 12336 6677 12364 6678
rect 12336 6651 12337 6677
rect 12337 6651 12363 6677
rect 12363 6651 12364 6677
rect 12336 6650 12364 6651
rect 11902 6285 11930 6286
rect 11902 6259 11903 6285
rect 11903 6259 11929 6285
rect 11929 6259 11930 6285
rect 11902 6258 11930 6259
rect 11954 6285 11982 6286
rect 11954 6259 11955 6285
rect 11955 6259 11981 6285
rect 11981 6259 11982 6285
rect 11954 6258 11982 6259
rect 12006 6285 12034 6286
rect 12006 6259 12007 6285
rect 12007 6259 12033 6285
rect 12033 6259 12034 6285
rect 12006 6258 12034 6259
rect 12558 6118 12586 6146
rect 11550 5558 11578 5586
rect 11998 5641 12026 5642
rect 11998 5615 11999 5641
rect 11999 5615 12025 5641
rect 12025 5615 12026 5641
rect 11998 5614 12026 5615
rect 11774 5502 11802 5530
rect 10206 5334 10234 5362
rect 10150 5054 10178 5082
rect 9758 3822 9786 3850
rect 9646 3206 9674 3234
rect 9422 2646 9450 2674
rect 9422 2534 9450 2562
rect 9366 2310 9394 2338
rect 9366 2142 9394 2170
rect 9030 2113 9058 2114
rect 9030 2087 9031 2113
rect 9031 2087 9057 2113
rect 9057 2087 9058 2113
rect 9030 2086 9058 2087
rect 9310 2057 9338 2058
rect 9310 2031 9311 2057
rect 9311 2031 9337 2057
rect 9337 2031 9338 2057
rect 9310 2030 9338 2031
rect 9254 1862 9282 1890
rect 9254 1750 9282 1778
rect 8918 1470 8946 1498
rect 9254 1470 9282 1498
rect 9478 2057 9506 2058
rect 9478 2031 9479 2057
rect 9479 2031 9505 2057
rect 9505 2031 9506 2057
rect 9478 2030 9506 2031
rect 9590 1302 9618 1330
rect 9366 1078 9394 1106
rect 9422 854 9450 882
rect 9590 854 9618 882
rect 9254 798 9282 826
rect 8918 574 8946 602
rect 9534 686 9562 714
rect 9086 406 9114 434
rect 9310 350 9338 378
rect 9870 4942 9898 4970
rect 9982 4857 10010 4858
rect 9982 4831 9983 4857
rect 9983 4831 10009 4857
rect 10009 4831 10010 4857
rect 9982 4830 10010 4831
rect 10038 4718 10066 4746
rect 9870 3430 9898 3458
rect 9926 4382 9954 4410
rect 9814 1582 9842 1610
rect 9870 1134 9898 1162
rect 9926 798 9954 826
rect 9982 4046 10010 4074
rect 10150 4494 10178 4522
rect 10094 4046 10122 4074
rect 9646 238 9674 266
rect 9758 742 9786 770
rect 10094 3766 10122 3794
rect 11718 5278 11746 5306
rect 11902 5501 11930 5502
rect 11902 5475 11903 5501
rect 11903 5475 11929 5501
rect 11929 5475 11930 5501
rect 11902 5474 11930 5475
rect 11954 5501 11982 5502
rect 11954 5475 11955 5501
rect 11955 5475 11981 5501
rect 11981 5475 11982 5501
rect 11954 5474 11982 5475
rect 12006 5501 12034 5502
rect 12006 5475 12007 5501
rect 12007 5475 12033 5501
rect 12033 5475 12034 5501
rect 12006 5474 12034 5475
rect 11830 5390 11858 5418
rect 11942 5390 11970 5418
rect 11270 5222 11298 5250
rect 11046 4774 11074 4802
rect 11158 4577 11186 4578
rect 11158 4551 11159 4577
rect 11159 4551 11185 4577
rect 11185 4551 11186 4577
rect 11158 4550 11186 4551
rect 11102 4185 11130 4186
rect 11102 4159 11103 4185
rect 11103 4159 11129 4185
rect 11129 4159 11130 4185
rect 11102 4158 11130 4159
rect 11214 4185 11242 4186
rect 11214 4159 11215 4185
rect 11215 4159 11241 4185
rect 11241 4159 11242 4185
rect 11214 4158 11242 4159
rect 11662 5110 11690 5138
rect 11718 4998 11746 5026
rect 12232 5893 12260 5894
rect 12232 5867 12233 5893
rect 12233 5867 12259 5893
rect 12259 5867 12260 5893
rect 12232 5866 12260 5867
rect 12284 5893 12312 5894
rect 12284 5867 12285 5893
rect 12285 5867 12311 5893
rect 12311 5867 12312 5893
rect 12284 5866 12312 5867
rect 12336 5893 12364 5894
rect 12336 5867 12337 5893
rect 12337 5867 12363 5893
rect 12363 5867 12364 5893
rect 12336 5866 12364 5867
rect 12278 5614 12306 5642
rect 12166 5446 12194 5474
rect 12166 5054 12194 5082
rect 12232 5109 12260 5110
rect 12232 5083 12233 5109
rect 12233 5083 12259 5109
rect 12259 5083 12260 5109
rect 12232 5082 12260 5083
rect 12284 5109 12312 5110
rect 12284 5083 12285 5109
rect 12285 5083 12311 5109
rect 12311 5083 12312 5109
rect 12284 5082 12312 5083
rect 12336 5109 12364 5110
rect 12336 5083 12337 5109
rect 12337 5083 12363 5109
rect 12363 5083 12364 5109
rect 12336 5082 12364 5083
rect 11902 4717 11930 4718
rect 11902 4691 11903 4717
rect 11903 4691 11929 4717
rect 11929 4691 11930 4717
rect 11902 4690 11930 4691
rect 11954 4717 11982 4718
rect 11954 4691 11955 4717
rect 11955 4691 11981 4717
rect 11981 4691 11982 4717
rect 11954 4690 11982 4691
rect 12006 4717 12034 4718
rect 12006 4691 12007 4717
rect 12007 4691 12033 4717
rect 12033 4691 12034 4717
rect 12110 4718 12138 4746
rect 12614 4942 12642 4970
rect 12006 4690 12034 4691
rect 11662 4606 11690 4634
rect 12166 4662 12194 4690
rect 11326 4550 11354 4578
rect 11606 4521 11634 4522
rect 11606 4495 11607 4521
rect 11607 4495 11633 4521
rect 11633 4495 11634 4521
rect 11606 4494 11634 4495
rect 11494 4382 11522 4410
rect 12614 4577 12642 4578
rect 12614 4551 12615 4577
rect 12615 4551 12641 4577
rect 12641 4551 12642 4577
rect 12614 4550 12642 4551
rect 12166 4326 12194 4354
rect 12614 4438 12642 4466
rect 12232 4325 12260 4326
rect 12232 4299 12233 4325
rect 12233 4299 12259 4325
rect 12259 4299 12260 4325
rect 12232 4298 12260 4299
rect 12284 4325 12312 4326
rect 12284 4299 12285 4325
rect 12285 4299 12311 4325
rect 12311 4299 12312 4325
rect 12284 4298 12312 4299
rect 12336 4325 12364 4326
rect 12336 4299 12337 4325
rect 12337 4299 12363 4325
rect 12363 4299 12364 4325
rect 12614 4326 12642 4354
rect 12336 4298 12364 4299
rect 11270 3878 11298 3906
rect 11494 3934 11522 3962
rect 11046 3766 11074 3794
rect 10710 3598 10738 3626
rect 10262 3374 10290 3402
rect 10206 3094 10234 3122
rect 11438 3262 11466 3290
rect 10094 3038 10122 3066
rect 10094 2534 10122 2562
rect 10486 2534 10514 2562
rect 10206 2030 10234 2058
rect 10262 1526 10290 1554
rect 11326 2534 11354 2562
rect 10710 2478 10738 2506
rect 10878 2254 10906 2282
rect 10710 1806 10738 1834
rect 10934 1638 10962 1666
rect 11214 2254 11242 2282
rect 10710 1358 10738 1386
rect 11102 1190 11130 1218
rect 10598 966 10626 994
rect 10598 686 10626 714
rect 10878 854 10906 882
rect 11046 601 11074 602
rect 11046 575 11047 601
rect 11047 575 11073 601
rect 11073 575 11074 601
rect 11046 574 11074 575
rect 11214 518 11242 546
rect 11214 70 11242 98
rect 11382 1414 11410 1442
rect 11902 3933 11930 3934
rect 11902 3907 11903 3933
rect 11903 3907 11929 3933
rect 11929 3907 11930 3933
rect 11902 3906 11930 3907
rect 11954 3933 11982 3934
rect 11954 3907 11955 3933
rect 11955 3907 11981 3933
rect 11981 3907 11982 3933
rect 11954 3906 11982 3907
rect 12006 3933 12034 3934
rect 12006 3907 12007 3933
rect 12007 3907 12033 3933
rect 12033 3907 12034 3933
rect 12614 3934 12642 3962
rect 12006 3906 12034 3907
rect 12166 3878 12194 3906
rect 11886 3654 11914 3682
rect 12558 3766 12586 3794
rect 12726 4886 12754 4914
rect 12782 4550 12810 4578
rect 12838 4214 12866 4242
rect 12894 6678 12922 6706
rect 13118 6622 13146 6650
rect 13286 6566 13314 6594
rect 13230 6145 13258 6146
rect 13230 6119 13231 6145
rect 13231 6119 13257 6145
rect 13257 6119 13258 6145
rect 13230 6118 13258 6119
rect 12950 6006 12978 6034
rect 12950 5054 12978 5082
rect 13006 5558 13034 5586
rect 13006 4662 13034 4690
rect 13118 5222 13146 5250
rect 13062 4577 13090 4578
rect 13062 4551 13063 4577
rect 13063 4551 13089 4577
rect 13089 4551 13090 4577
rect 13062 4550 13090 4551
rect 13510 5838 13538 5866
rect 13454 5726 13482 5754
rect 13510 5390 13538 5418
rect 15190 6734 15218 6762
rect 16086 6902 16114 6930
rect 14014 6089 14042 6090
rect 14014 6063 14015 6089
rect 14015 6063 14041 6089
rect 14041 6063 14042 6089
rect 14014 6062 14042 6063
rect 14238 6089 14266 6090
rect 14238 6063 14239 6089
rect 14239 6063 14265 6089
rect 14265 6063 14266 6089
rect 14238 6062 14266 6063
rect 14518 6089 14546 6090
rect 14518 6063 14519 6089
rect 14519 6063 14545 6089
rect 14545 6063 14546 6089
rect 14518 6062 14546 6063
rect 15134 6006 15162 6034
rect 13678 5838 13706 5866
rect 13678 5390 13706 5418
rect 14294 5446 14322 5474
rect 13566 5334 13594 5362
rect 13510 4718 13538 4746
rect 13902 5222 13930 5250
rect 13454 4662 13482 4690
rect 13454 4438 13482 4466
rect 12670 3766 12698 3794
rect 12782 4158 12810 4186
rect 12166 3542 12194 3570
rect 12232 3541 12260 3542
rect 12232 3515 12233 3541
rect 12233 3515 12259 3541
rect 12259 3515 12260 3541
rect 12232 3514 12260 3515
rect 12284 3541 12312 3542
rect 12284 3515 12285 3541
rect 12285 3515 12311 3541
rect 12311 3515 12312 3541
rect 12284 3514 12312 3515
rect 12336 3541 12364 3542
rect 12336 3515 12337 3541
rect 12337 3515 12363 3541
rect 12363 3515 12364 3541
rect 12336 3514 12364 3515
rect 11886 3430 11914 3458
rect 12726 3318 12754 3346
rect 11902 3149 11930 3150
rect 11494 2870 11522 2898
rect 11774 3094 11802 3122
rect 11902 3123 11903 3149
rect 11903 3123 11929 3149
rect 11929 3123 11930 3149
rect 11902 3122 11930 3123
rect 11954 3149 11982 3150
rect 11954 3123 11955 3149
rect 11955 3123 11981 3149
rect 11981 3123 11982 3149
rect 11954 3122 11982 3123
rect 12006 3149 12034 3150
rect 12006 3123 12007 3149
rect 12007 3123 12033 3149
rect 12033 3123 12034 3149
rect 12006 3122 12034 3123
rect 12558 3150 12586 3178
rect 12054 2926 12082 2954
rect 11830 2841 11858 2842
rect 11830 2815 11831 2841
rect 11831 2815 11857 2841
rect 11857 2815 11858 2841
rect 11830 2814 11858 2815
rect 11942 2841 11970 2842
rect 11942 2815 11943 2841
rect 11943 2815 11969 2841
rect 11969 2815 11970 2841
rect 11942 2814 11970 2815
rect 12054 2646 12082 2674
rect 12110 2870 12138 2898
rect 12222 2897 12250 2898
rect 12222 2871 12223 2897
rect 12223 2871 12249 2897
rect 12249 2871 12250 2897
rect 12222 2870 12250 2871
rect 12232 2757 12260 2758
rect 12232 2731 12233 2757
rect 12233 2731 12259 2757
rect 12259 2731 12260 2757
rect 12232 2730 12260 2731
rect 12284 2757 12312 2758
rect 12284 2731 12285 2757
rect 12285 2731 12311 2757
rect 12311 2731 12312 2757
rect 12284 2730 12312 2731
rect 12336 2757 12364 2758
rect 12336 2731 12337 2757
rect 12337 2731 12363 2757
rect 12363 2731 12364 2757
rect 12336 2730 12364 2731
rect 12222 2561 12250 2562
rect 12222 2535 12223 2561
rect 12223 2535 12249 2561
rect 12249 2535 12250 2561
rect 12222 2534 12250 2535
rect 12446 2534 12474 2562
rect 12670 3038 12698 3066
rect 12558 2478 12586 2506
rect 12614 2926 12642 2954
rect 11902 2365 11930 2366
rect 11902 2339 11903 2365
rect 11903 2339 11929 2365
rect 11929 2339 11930 2365
rect 11902 2338 11930 2339
rect 11954 2365 11982 2366
rect 11954 2339 11955 2365
rect 11955 2339 11981 2365
rect 11981 2339 11982 2365
rect 11954 2338 11982 2339
rect 12006 2365 12034 2366
rect 12006 2339 12007 2365
rect 12007 2339 12033 2365
rect 12033 2339 12034 2365
rect 12110 2366 12138 2394
rect 12006 2338 12034 2339
rect 11774 2142 11802 2170
rect 11830 1974 11858 2002
rect 11494 1694 11522 1722
rect 11494 1414 11522 1442
rect 11998 1721 12026 1722
rect 11998 1695 11999 1721
rect 11999 1695 12025 1721
rect 12025 1695 12026 1721
rect 11998 1694 12026 1695
rect 11830 1582 11858 1610
rect 11902 1581 11930 1582
rect 11902 1555 11903 1581
rect 11903 1555 11929 1581
rect 11929 1555 11930 1581
rect 11902 1554 11930 1555
rect 11954 1581 11982 1582
rect 11954 1555 11955 1581
rect 11955 1555 11981 1581
rect 11981 1555 11982 1581
rect 11954 1554 11982 1555
rect 12006 1581 12034 1582
rect 12006 1555 12007 1581
rect 12007 1555 12033 1581
rect 12033 1555 12034 1581
rect 12006 1554 12034 1555
rect 12110 1582 12138 1610
rect 12110 1190 12138 1218
rect 11830 1022 11858 1050
rect 11550 854 11578 882
rect 11902 797 11930 798
rect 11902 771 11903 797
rect 11903 771 11929 797
rect 11929 771 11930 797
rect 11902 770 11930 771
rect 11954 797 11982 798
rect 11954 771 11955 797
rect 11955 771 11981 797
rect 11981 771 11982 797
rect 11954 770 11982 771
rect 12006 797 12034 798
rect 12006 771 12007 797
rect 12007 771 12033 797
rect 12033 771 12034 797
rect 12006 770 12034 771
rect 11438 545 11466 546
rect 11438 519 11439 545
rect 11439 519 11465 545
rect 11465 519 11466 545
rect 11438 518 11466 519
rect 11774 574 11802 602
rect 12232 1973 12260 1974
rect 12232 1947 12233 1973
rect 12233 1947 12259 1973
rect 12259 1947 12260 1973
rect 12232 1946 12260 1947
rect 12284 1973 12312 1974
rect 12284 1947 12285 1973
rect 12285 1947 12311 1973
rect 12311 1947 12312 1973
rect 12284 1946 12312 1947
rect 12336 1973 12364 1974
rect 12336 1947 12337 1973
rect 12337 1947 12363 1973
rect 12363 1947 12364 1973
rect 12336 1946 12364 1947
rect 12558 1777 12586 1778
rect 12558 1751 12559 1777
rect 12559 1751 12585 1777
rect 12585 1751 12586 1777
rect 12558 1750 12586 1751
rect 12278 1582 12306 1610
rect 12502 1694 12530 1722
rect 12446 1246 12474 1274
rect 12232 1189 12260 1190
rect 12232 1163 12233 1189
rect 12233 1163 12259 1189
rect 12259 1163 12260 1189
rect 12232 1162 12260 1163
rect 12284 1189 12312 1190
rect 12284 1163 12285 1189
rect 12285 1163 12311 1189
rect 12311 1163 12312 1189
rect 12284 1162 12312 1163
rect 12336 1189 12364 1190
rect 12336 1163 12337 1189
rect 12337 1163 12363 1189
rect 12363 1163 12364 1189
rect 12336 1162 12364 1163
rect 12502 1190 12530 1218
rect 12670 2478 12698 2506
rect 12614 1302 12642 1330
rect 12446 518 12474 546
rect 12232 405 12260 406
rect 12232 379 12233 405
rect 12233 379 12259 405
rect 12259 379 12260 405
rect 12232 378 12260 379
rect 12284 405 12312 406
rect 12284 379 12285 405
rect 12285 379 12311 405
rect 12311 379 12312 405
rect 12284 378 12312 379
rect 12336 405 12364 406
rect 12336 379 12337 405
rect 12337 379 12363 405
rect 12363 379 12364 405
rect 12336 378 12364 379
rect 12558 545 12586 546
rect 12558 519 12559 545
rect 12559 519 12585 545
rect 12585 519 12586 545
rect 12558 518 12586 519
rect 12670 630 12698 658
rect 12838 3737 12866 3738
rect 12838 3711 12839 3737
rect 12839 3711 12865 3737
rect 12865 3711 12866 3737
rect 12838 3710 12866 3711
rect 12950 3737 12978 3738
rect 12950 3711 12951 3737
rect 12951 3711 12977 3737
rect 12977 3711 12978 3737
rect 12950 3710 12978 3711
rect 12782 2926 12810 2954
rect 12894 2870 12922 2898
rect 12838 2590 12866 2618
rect 12838 1862 12866 1890
rect 12726 574 12754 602
rect 13118 3486 13146 3514
rect 13062 3289 13090 3290
rect 13062 3263 13063 3289
rect 13063 3263 13089 3289
rect 13089 3263 13090 3289
rect 13062 3262 13090 3263
rect 13118 2870 13146 2898
rect 13006 2422 13034 2450
rect 13286 3542 13314 3570
rect 13230 3262 13258 3290
rect 13286 2198 13314 2226
rect 13398 4326 13426 4354
rect 13398 4158 13426 4186
rect 13734 4326 13762 4354
rect 13398 2982 13426 3010
rect 13342 1974 13370 2002
rect 13398 2366 13426 2394
rect 13062 1358 13090 1386
rect 12838 574 12866 602
rect 12894 630 12922 658
rect 12614 350 12642 378
rect 13398 1358 13426 1386
rect 13454 2198 13482 2226
rect 13398 966 13426 994
rect 13958 4774 13986 4802
rect 14014 4606 14042 4634
rect 14238 4606 14266 4634
rect 14182 4270 14210 4298
rect 13902 3654 13930 3682
rect 13734 2478 13762 2506
rect 13510 966 13538 994
rect 13342 910 13370 938
rect 13286 742 13314 770
rect 13230 630 13258 658
rect 13454 657 13482 658
rect 13454 631 13455 657
rect 13455 631 13481 657
rect 13481 631 13482 657
rect 13454 630 13482 631
rect 13118 518 13146 546
rect 13342 518 13370 546
rect 14126 1750 14154 1778
rect 14070 1721 14098 1722
rect 14070 1695 14071 1721
rect 14071 1695 14097 1721
rect 14097 1695 14098 1721
rect 14070 1694 14098 1695
rect 14014 1470 14042 1498
rect 13790 1022 13818 1050
rect 13622 518 13650 546
rect 13790 630 13818 658
rect 14350 5361 14378 5362
rect 14350 5335 14351 5361
rect 14351 5335 14377 5361
rect 14377 5335 14378 5361
rect 14350 5334 14378 5335
rect 14630 5334 14658 5362
rect 14798 5361 14826 5362
rect 14798 5335 14799 5361
rect 14799 5335 14825 5361
rect 14825 5335 14826 5361
rect 14798 5334 14826 5335
rect 14854 5278 14882 5306
rect 14350 5110 14378 5138
rect 14350 4998 14378 5026
rect 14294 2673 14322 2674
rect 14294 2647 14295 2673
rect 14295 2647 14321 2673
rect 14321 2647 14322 2673
rect 14294 2646 14322 2647
rect 14350 2478 14378 2506
rect 14854 4102 14882 4130
rect 14518 4073 14546 4074
rect 14518 4047 14519 4073
rect 14519 4047 14545 4073
rect 14545 4047 14546 4073
rect 14518 4046 14546 4047
rect 19726 7014 19754 7042
rect 19950 7014 19978 7042
rect 18382 6734 18410 6762
rect 18438 6902 18466 6930
rect 16422 6481 16450 6482
rect 16422 6455 16423 6481
rect 16423 6455 16449 6481
rect 16449 6455 16450 6481
rect 16422 6454 16450 6455
rect 17038 6454 17066 6482
rect 16534 6230 16562 6258
rect 15190 5838 15218 5866
rect 15246 5193 15274 5194
rect 15246 5167 15247 5193
rect 15247 5167 15273 5193
rect 15273 5167 15274 5193
rect 15246 5166 15274 5167
rect 14966 4046 14994 4074
rect 15022 4382 15050 4410
rect 14910 3654 14938 3682
rect 14462 2673 14490 2674
rect 14462 2647 14463 2673
rect 14463 2647 14489 2673
rect 14489 2647 14490 2673
rect 14462 2646 14490 2647
rect 14630 1022 14658 1050
rect 14126 686 14154 714
rect 14742 966 14770 994
rect 14406 182 14434 210
rect 14798 854 14826 882
rect 16310 6006 16338 6034
rect 15974 5446 16002 5474
rect 15414 5193 15442 5194
rect 15414 5167 15415 5193
rect 15415 5167 15441 5193
rect 15441 5167 15442 5193
rect 15414 5166 15442 5167
rect 15190 3990 15218 4018
rect 15358 3990 15386 4018
rect 15470 3990 15498 4018
rect 15078 3878 15106 3906
rect 15022 2366 15050 2394
rect 15190 3094 15218 3122
rect 15190 2982 15218 3010
rect 15134 2198 15162 2226
rect 15078 2030 15106 2058
rect 15078 1638 15106 1666
rect 15078 1078 15106 1106
rect 15246 1414 15274 1442
rect 15694 3486 15722 3514
rect 15806 4214 15834 4242
rect 15694 2534 15722 2562
rect 15582 966 15610 994
rect 15470 798 15498 826
rect 14686 462 14714 490
rect 15078 489 15106 490
rect 15078 463 15079 489
rect 15079 463 15105 489
rect 15105 463 15106 489
rect 15078 462 15106 463
rect 14910 406 14938 434
rect 15358 182 15386 210
rect 15470 126 15498 154
rect 15582 854 15610 882
rect 15638 798 15666 826
rect 15750 1694 15778 1722
rect 15974 4606 16002 4634
rect 15974 3878 16002 3906
rect 16478 5502 16506 5530
rect 15918 2982 15946 3010
rect 15974 2478 16002 2506
rect 16254 2310 16282 2338
rect 16422 3542 16450 3570
rect 16142 2225 16170 2226
rect 16142 2199 16143 2225
rect 16143 2199 16169 2225
rect 16169 2199 16170 2225
rect 16142 2198 16170 2199
rect 15806 1526 15834 1554
rect 15806 630 15834 658
rect 15694 70 15722 98
rect 16030 406 16058 434
rect 16198 1049 16226 1050
rect 16198 1023 16199 1049
rect 16199 1023 16225 1049
rect 16225 1023 16226 1049
rect 16198 1022 16226 1023
rect 16310 630 16338 658
rect 16254 406 16282 434
rect 16758 6174 16786 6202
rect 16758 5726 16786 5754
rect 16758 5222 16786 5250
rect 16702 4774 16730 4802
rect 16758 3766 16786 3794
rect 16814 4718 16842 4746
rect 18214 6342 18242 6370
rect 17766 6033 17794 6034
rect 17766 6007 17767 6033
rect 17767 6007 17793 6033
rect 17793 6007 17794 6033
rect 17766 6006 17794 6007
rect 18046 5950 18074 5978
rect 17094 5782 17122 5810
rect 17206 5782 17234 5810
rect 17206 5502 17234 5530
rect 17374 5446 17402 5474
rect 17710 5558 17738 5586
rect 17542 5166 17570 5194
rect 17206 5054 17234 5082
rect 17598 4998 17626 5026
rect 17038 4606 17066 4634
rect 17374 3793 17402 3794
rect 17374 3767 17375 3793
rect 17375 3767 17401 3793
rect 17401 3767 17402 3793
rect 17374 3766 17402 3767
rect 17486 3318 17514 3346
rect 16814 2646 16842 2674
rect 17150 2870 17178 2898
rect 17598 2617 17626 2618
rect 17598 2591 17599 2617
rect 17599 2591 17625 2617
rect 17625 2591 17626 2617
rect 17598 2590 17626 2591
rect 17430 2366 17458 2394
rect 17822 5558 17850 5586
rect 17822 3793 17850 3794
rect 17822 3767 17823 3793
rect 17823 3767 17849 3793
rect 17849 3767 17850 3793
rect 17822 3766 17850 3767
rect 17710 2254 17738 2282
rect 16534 1302 16562 1330
rect 16478 881 16506 882
rect 16478 855 16479 881
rect 16479 855 16505 881
rect 16505 855 16506 881
rect 16478 854 16506 855
rect 16422 238 16450 266
rect 16646 742 16674 770
rect 17430 2086 17458 2114
rect 17094 1974 17122 2002
rect 17094 1806 17122 1834
rect 17150 1721 17178 1722
rect 17150 1695 17151 1721
rect 17151 1695 17177 1721
rect 17177 1695 17178 1721
rect 17150 1694 17178 1695
rect 17038 1329 17066 1330
rect 17038 1303 17039 1329
rect 17039 1303 17065 1329
rect 17065 1303 17066 1329
rect 17038 1302 17066 1303
rect 16758 742 16786 770
rect 16646 630 16674 658
rect 16534 601 16562 602
rect 16534 575 16535 601
rect 16535 575 16561 601
rect 16561 575 16562 601
rect 16534 574 16562 575
rect 16702 462 16730 490
rect 17654 1694 17682 1722
rect 18046 2926 18074 2954
rect 18158 4326 18186 4354
rect 18606 6734 18634 6762
rect 22414 7014 22442 7042
rect 22582 7014 22610 7042
rect 21070 6734 21098 6762
rect 21574 6734 21602 6762
rect 21406 6622 21434 6650
rect 19110 6118 19138 6146
rect 19950 6145 19978 6146
rect 19950 6119 19951 6145
rect 19951 6119 19977 6145
rect 19977 6119 19978 6145
rect 19950 6118 19978 6119
rect 18550 6033 18578 6034
rect 18550 6007 18551 6033
rect 18551 6007 18577 6033
rect 18577 6007 18578 6033
rect 18550 6006 18578 6007
rect 20230 6033 20258 6034
rect 20230 6007 20231 6033
rect 20231 6007 20257 6033
rect 20257 6007 20258 6033
rect 20230 6006 20258 6007
rect 20398 6033 20426 6034
rect 20398 6007 20399 6033
rect 20399 6007 20425 6033
rect 20425 6007 20426 6033
rect 20398 6006 20426 6007
rect 18326 5110 18354 5138
rect 18438 4382 18466 4410
rect 18326 2926 18354 2954
rect 18382 4270 18410 4298
rect 18382 2702 18410 2730
rect 18214 2534 18242 2562
rect 18438 2198 18466 2226
rect 17878 2113 17906 2114
rect 17878 2087 17879 2113
rect 17879 2087 17905 2113
rect 17905 2087 17906 2113
rect 17878 2086 17906 2087
rect 17878 1833 17906 1834
rect 17878 1807 17879 1833
rect 17879 1807 17905 1833
rect 17905 1807 17906 1833
rect 17878 1806 17906 1807
rect 18438 1806 18466 1834
rect 17822 1358 17850 1386
rect 17598 1049 17626 1050
rect 17598 1023 17599 1049
rect 17599 1023 17625 1049
rect 17625 1023 17626 1049
rect 17598 1022 17626 1023
rect 17878 1022 17906 1050
rect 17094 406 17122 434
rect 17598 854 17626 882
rect 16814 182 16842 210
rect 16926 350 16954 378
rect 17486 630 17514 658
rect 17486 518 17514 546
rect 17374 406 17402 434
rect 17654 798 17682 826
rect 17934 489 17962 490
rect 17934 463 17935 489
rect 17935 463 17961 489
rect 17961 463 17962 489
rect 17934 462 17962 463
rect 17878 350 17906 378
rect 17822 182 17850 210
rect 18718 4046 18746 4074
rect 18550 3878 18578 3906
rect 18494 1638 18522 1666
rect 18606 2590 18634 2618
rect 18158 1385 18186 1386
rect 18158 1359 18159 1385
rect 18159 1359 18185 1385
rect 18185 1359 18186 1385
rect 18158 1358 18186 1359
rect 18494 1358 18522 1386
rect 18494 1190 18522 1218
rect 18494 1078 18522 1106
rect 18382 993 18410 994
rect 18382 967 18383 993
rect 18383 967 18409 993
rect 18409 967 18410 993
rect 18382 966 18410 967
rect 18270 518 18298 546
rect 18550 854 18578 882
rect 18830 3934 18858 3962
rect 18830 3542 18858 3570
rect 18718 2310 18746 2338
rect 18774 2422 18802 2450
rect 18886 2086 18914 2114
rect 18886 1918 18914 1946
rect 18830 1526 18858 1554
rect 19670 5334 19698 5362
rect 19278 5305 19306 5306
rect 19278 5279 19279 5305
rect 19279 5279 19305 5305
rect 19305 5279 19306 5305
rect 19278 5278 19306 5279
rect 19446 2870 19474 2898
rect 19110 2478 19138 2506
rect 19278 2478 19306 2506
rect 19054 1582 19082 1610
rect 19054 1078 19082 1106
rect 19334 1638 19362 1666
rect 19558 2422 19586 2450
rect 19558 2198 19586 2226
rect 19502 2057 19530 2058
rect 19502 2031 19503 2057
rect 19503 2031 19529 2057
rect 19529 2031 19530 2057
rect 19502 2030 19530 2031
rect 19614 2057 19642 2058
rect 19614 2031 19615 2057
rect 19615 2031 19641 2057
rect 19641 2031 19642 2057
rect 19614 2030 19642 2031
rect 19614 993 19642 994
rect 19614 967 19615 993
rect 19615 967 19641 993
rect 19641 967 19642 993
rect 19614 966 19642 967
rect 19614 854 19642 882
rect 18718 489 18746 490
rect 18718 463 18719 489
rect 18719 463 18745 489
rect 18745 463 18746 489
rect 18718 462 18746 463
rect 18662 182 18690 210
rect 19166 350 19194 378
rect 18942 238 18970 266
rect 19390 294 19418 322
rect 20454 4465 20482 4466
rect 20454 4439 20455 4465
rect 20455 4439 20481 4465
rect 20481 4439 20482 4465
rect 20454 4438 20482 4439
rect 20342 3150 20370 3178
rect 20286 2897 20314 2898
rect 20286 2871 20287 2897
rect 20287 2871 20313 2897
rect 20313 2871 20314 2897
rect 20286 2870 20314 2871
rect 19894 1190 19922 1218
rect 19726 798 19754 826
rect 19838 798 19866 826
rect 19782 545 19810 546
rect 19782 519 19783 545
rect 19783 519 19809 545
rect 19809 519 19810 545
rect 19782 518 19810 519
rect 19726 70 19754 98
rect 19894 742 19922 770
rect 19950 350 19978 378
rect 20062 462 20090 490
rect 20566 4465 20594 4466
rect 20566 4439 20567 4465
rect 20567 4439 20593 4465
rect 20593 4439 20594 4465
rect 20566 4438 20594 4439
rect 20846 4465 20874 4466
rect 20846 4439 20847 4465
rect 20847 4439 20873 4465
rect 20873 4439 20874 4465
rect 20846 4438 20874 4439
rect 21182 4438 21210 4466
rect 20510 2422 20538 2450
rect 20790 3318 20818 3346
rect 20622 2254 20650 2282
rect 20902 3038 20930 3066
rect 21070 2982 21098 3010
rect 20958 2225 20986 2226
rect 20958 2199 20959 2225
rect 20959 2199 20985 2225
rect 20985 2199 20986 2225
rect 20958 2198 20986 2199
rect 20678 1750 20706 1778
rect 20286 798 20314 826
rect 20510 798 20538 826
rect 20230 294 20258 322
rect 20286 518 20314 546
rect 20454 238 20482 266
rect 20790 1694 20818 1722
rect 21126 2673 21154 2674
rect 21126 2647 21127 2673
rect 21127 2647 21153 2673
rect 21153 2647 21154 2673
rect 21126 2646 21154 2647
rect 22232 6677 22260 6678
rect 22232 6651 22233 6677
rect 22233 6651 22259 6677
rect 22259 6651 22260 6677
rect 22232 6650 22260 6651
rect 22284 6677 22312 6678
rect 22284 6651 22285 6677
rect 22285 6651 22311 6677
rect 22311 6651 22312 6677
rect 22284 6650 22312 6651
rect 22336 6677 22364 6678
rect 22336 6651 22337 6677
rect 22337 6651 22363 6677
rect 22363 6651 22364 6677
rect 22336 6650 22364 6651
rect 22078 6481 22106 6482
rect 22078 6455 22079 6481
rect 22079 6455 22105 6481
rect 22105 6455 22106 6481
rect 22078 6454 22106 6455
rect 23758 7014 23786 7042
rect 23982 7014 24010 7042
rect 23254 6566 23282 6594
rect 21902 6285 21930 6286
rect 21902 6259 21903 6285
rect 21903 6259 21929 6285
rect 21929 6259 21930 6285
rect 21902 6258 21930 6259
rect 21954 6285 21982 6286
rect 21954 6259 21955 6285
rect 21955 6259 21981 6285
rect 21981 6259 21982 6285
rect 21954 6258 21982 6259
rect 22006 6285 22034 6286
rect 22006 6259 22007 6285
rect 22007 6259 22033 6285
rect 22033 6259 22034 6285
rect 22006 6258 22034 6259
rect 22414 6006 22442 6034
rect 22302 5977 22330 5978
rect 22302 5951 22303 5977
rect 22303 5951 22329 5977
rect 22329 5951 22330 5977
rect 22302 5950 22330 5951
rect 22232 5893 22260 5894
rect 22134 5838 22162 5866
rect 22232 5867 22233 5893
rect 22233 5867 22259 5893
rect 22259 5867 22260 5893
rect 22232 5866 22260 5867
rect 22284 5893 22312 5894
rect 22284 5867 22285 5893
rect 22285 5867 22311 5893
rect 22311 5867 22312 5893
rect 22284 5866 22312 5867
rect 22336 5893 22364 5894
rect 22336 5867 22337 5893
rect 22337 5867 22363 5893
rect 22363 5867 22364 5893
rect 22336 5866 22364 5867
rect 21902 5501 21930 5502
rect 21902 5475 21903 5501
rect 21903 5475 21929 5501
rect 21929 5475 21930 5501
rect 21902 5474 21930 5475
rect 21954 5501 21982 5502
rect 21954 5475 21955 5501
rect 21955 5475 21981 5501
rect 21981 5475 21982 5501
rect 21954 5474 21982 5475
rect 22006 5501 22034 5502
rect 22006 5475 22007 5501
rect 22007 5475 22033 5501
rect 22033 5475 22034 5501
rect 22006 5474 22034 5475
rect 22134 5334 22162 5362
rect 22232 5109 22260 5110
rect 22232 5083 22233 5109
rect 22233 5083 22259 5109
rect 22259 5083 22260 5109
rect 22232 5082 22260 5083
rect 22284 5109 22312 5110
rect 22284 5083 22285 5109
rect 22285 5083 22311 5109
rect 22311 5083 22312 5109
rect 22284 5082 22312 5083
rect 22336 5109 22364 5110
rect 22336 5083 22337 5109
rect 22337 5083 22363 5109
rect 22363 5083 22364 5109
rect 22336 5082 22364 5083
rect 21902 4717 21930 4718
rect 21902 4691 21903 4717
rect 21903 4691 21929 4717
rect 21929 4691 21930 4717
rect 21902 4690 21930 4691
rect 21954 4717 21982 4718
rect 21954 4691 21955 4717
rect 21955 4691 21981 4717
rect 21981 4691 21982 4717
rect 21954 4690 21982 4691
rect 22006 4717 22034 4718
rect 22006 4691 22007 4717
rect 22007 4691 22033 4717
rect 22033 4691 22034 4717
rect 22006 4690 22034 4691
rect 22358 4465 22386 4466
rect 22358 4439 22359 4465
rect 22359 4439 22385 4465
rect 22385 4439 22386 4465
rect 22358 4438 22386 4439
rect 21854 4409 21882 4410
rect 21854 4383 21855 4409
rect 21855 4383 21881 4409
rect 21881 4383 21882 4409
rect 21854 4382 21882 4383
rect 22232 4325 22260 4326
rect 22232 4299 22233 4325
rect 22233 4299 22259 4325
rect 22259 4299 22260 4325
rect 22232 4298 22260 4299
rect 22284 4325 22312 4326
rect 22284 4299 22285 4325
rect 22285 4299 22311 4325
rect 22311 4299 22312 4325
rect 22284 4298 22312 4299
rect 22336 4325 22364 4326
rect 22336 4299 22337 4325
rect 22337 4299 22363 4325
rect 22363 4299 22364 4325
rect 22336 4298 22364 4299
rect 21630 4073 21658 4074
rect 21630 4047 21631 4073
rect 21631 4047 21657 4073
rect 21657 4047 21658 4073
rect 21630 4046 21658 4047
rect 21798 4046 21826 4074
rect 22078 4073 22106 4074
rect 22078 4047 22079 4073
rect 22079 4047 22105 4073
rect 22105 4047 22106 4073
rect 22078 4046 22106 4047
rect 21902 3933 21930 3934
rect 21902 3907 21903 3933
rect 21903 3907 21929 3933
rect 21929 3907 21930 3933
rect 21902 3906 21930 3907
rect 21954 3933 21982 3934
rect 21954 3907 21955 3933
rect 21955 3907 21981 3933
rect 21981 3907 21982 3933
rect 21954 3906 21982 3907
rect 22006 3933 22034 3934
rect 22006 3907 22007 3933
rect 22007 3907 22033 3933
rect 22033 3907 22034 3933
rect 22006 3906 22034 3907
rect 21910 3822 21938 3850
rect 22134 3822 22162 3850
rect 21966 3374 21994 3402
rect 22134 3542 22162 3570
rect 21798 3150 21826 3178
rect 21902 3149 21930 3150
rect 21462 3094 21490 3122
rect 21902 3123 21903 3149
rect 21903 3123 21929 3149
rect 21929 3123 21930 3149
rect 21902 3122 21930 3123
rect 21954 3149 21982 3150
rect 21954 3123 21955 3149
rect 21955 3123 21981 3149
rect 21981 3123 21982 3149
rect 21954 3122 21982 3123
rect 22006 3149 22034 3150
rect 22006 3123 22007 3149
rect 22007 3123 22033 3149
rect 22033 3123 22034 3149
rect 22006 3122 22034 3123
rect 21406 3038 21434 3066
rect 21294 2673 21322 2674
rect 21294 2647 21295 2673
rect 21295 2647 21321 2673
rect 21321 2647 21322 2673
rect 21294 2646 21322 2647
rect 21182 2198 21210 2226
rect 21182 1721 21210 1722
rect 21182 1695 21183 1721
rect 21183 1695 21209 1721
rect 21209 1695 21210 1721
rect 21182 1694 21210 1695
rect 21462 1694 21490 1722
rect 21070 1246 21098 1274
rect 21014 881 21042 882
rect 21014 855 21015 881
rect 21015 855 21041 881
rect 21041 855 21042 881
rect 21014 854 21042 855
rect 20622 462 20650 490
rect 20958 742 20986 770
rect 20958 406 20986 434
rect 21350 1190 21378 1218
rect 21070 182 21098 210
rect 21182 966 21210 994
rect 21518 1190 21546 1218
rect 21686 2366 21714 2394
rect 21902 2365 21930 2366
rect 21902 2339 21903 2365
rect 21903 2339 21929 2365
rect 21929 2339 21930 2365
rect 21902 2338 21930 2339
rect 21954 2365 21982 2366
rect 21954 2339 21955 2365
rect 21955 2339 21981 2365
rect 21981 2339 21982 2365
rect 21954 2338 21982 2339
rect 22006 2365 22034 2366
rect 22006 2339 22007 2365
rect 22007 2339 22033 2365
rect 22033 2339 22034 2365
rect 22006 2338 22034 2339
rect 21902 1581 21930 1582
rect 21902 1555 21903 1581
rect 21903 1555 21929 1581
rect 21929 1555 21930 1581
rect 21902 1554 21930 1555
rect 21954 1581 21982 1582
rect 21954 1555 21955 1581
rect 21955 1555 21981 1581
rect 21981 1555 21982 1581
rect 21954 1554 21982 1555
rect 22006 1581 22034 1582
rect 22006 1555 22007 1581
rect 22007 1555 22033 1581
rect 22033 1555 22034 1581
rect 22006 1554 22034 1555
rect 22022 1470 22050 1498
rect 21686 910 21714 938
rect 21574 742 21602 770
rect 21630 686 21658 714
rect 22232 3541 22260 3542
rect 22232 3515 22233 3541
rect 22233 3515 22259 3541
rect 22259 3515 22260 3541
rect 22232 3514 22260 3515
rect 22284 3541 22312 3542
rect 22284 3515 22285 3541
rect 22285 3515 22311 3541
rect 22311 3515 22312 3541
rect 22284 3514 22312 3515
rect 22336 3541 22364 3542
rect 22336 3515 22337 3541
rect 22337 3515 22363 3541
rect 22363 3515 22364 3541
rect 22336 3514 22364 3515
rect 22414 3486 22442 3514
rect 22470 5334 22498 5362
rect 22134 3094 22162 3122
rect 22232 2757 22260 2758
rect 22232 2731 22233 2757
rect 22233 2731 22259 2757
rect 22259 2731 22260 2757
rect 22232 2730 22260 2731
rect 22284 2757 22312 2758
rect 22284 2731 22285 2757
rect 22285 2731 22311 2757
rect 22311 2731 22312 2757
rect 22284 2730 22312 2731
rect 22336 2757 22364 2758
rect 22336 2731 22337 2757
rect 22337 2731 22363 2757
rect 22363 2731 22364 2757
rect 22336 2730 22364 2731
rect 22470 2310 22498 2338
rect 22358 2169 22386 2170
rect 22358 2143 22359 2169
rect 22359 2143 22385 2169
rect 22385 2143 22386 2169
rect 22358 2142 22386 2143
rect 22470 2169 22498 2170
rect 22470 2143 22471 2169
rect 22471 2143 22497 2169
rect 22497 2143 22498 2169
rect 22470 2142 22498 2143
rect 22232 1973 22260 1974
rect 22232 1947 22233 1973
rect 22233 1947 22259 1973
rect 22259 1947 22260 1973
rect 22232 1946 22260 1947
rect 22284 1973 22312 1974
rect 22284 1947 22285 1973
rect 22285 1947 22311 1973
rect 22311 1947 22312 1973
rect 22284 1946 22312 1947
rect 22336 1973 22364 1974
rect 22336 1947 22337 1973
rect 22337 1947 22363 1973
rect 22363 1947 22364 1973
rect 22336 1946 22364 1947
rect 22022 910 22050 938
rect 21966 881 21994 882
rect 21966 855 21967 881
rect 21967 855 21993 881
rect 21993 855 21994 881
rect 21966 854 21994 855
rect 21902 797 21930 798
rect 21902 771 21903 797
rect 21903 771 21929 797
rect 21929 771 21930 797
rect 21902 770 21930 771
rect 21954 797 21982 798
rect 21954 771 21955 797
rect 21955 771 21981 797
rect 21981 771 21982 797
rect 21954 770 21982 771
rect 22006 797 22034 798
rect 22006 771 22007 797
rect 22007 771 22033 797
rect 22033 771 22034 797
rect 22006 770 22034 771
rect 22078 742 22106 770
rect 21406 406 21434 434
rect 21686 545 21714 546
rect 21686 519 21687 545
rect 21687 519 21713 545
rect 21713 519 21714 545
rect 21686 518 21714 519
rect 21854 518 21882 546
rect 22470 1833 22498 1834
rect 22470 1807 22471 1833
rect 22471 1807 22497 1833
rect 22497 1807 22498 1833
rect 22470 1806 22498 1807
rect 22974 4438 23002 4466
rect 22750 4046 22778 4074
rect 22694 3345 22722 3346
rect 22694 3319 22695 3345
rect 22695 3319 22721 3345
rect 22721 3319 22722 3345
rect 22694 3318 22722 3319
rect 23646 6510 23674 6538
rect 23534 5726 23562 5754
rect 25102 7014 25130 7042
rect 25382 7014 25410 7042
rect 24990 6790 25018 6818
rect 23702 6033 23730 6034
rect 23702 6007 23703 6033
rect 23703 6007 23729 6033
rect 23729 6007 23730 6033
rect 23702 6006 23730 6007
rect 24262 5670 24290 5698
rect 24206 4774 24234 4802
rect 24150 4606 24178 4634
rect 22974 3878 23002 3906
rect 23366 3990 23394 4018
rect 23198 3094 23226 3122
rect 22750 2758 22778 2786
rect 23310 2673 23338 2674
rect 23310 2647 23311 2673
rect 23311 2647 23337 2673
rect 23337 2647 23338 2673
rect 23310 2646 23338 2647
rect 22918 2590 22946 2618
rect 22750 1750 22778 1778
rect 22638 1638 22666 1666
rect 22190 1470 22218 1498
rect 22232 1189 22260 1190
rect 22232 1163 22233 1189
rect 22233 1163 22259 1189
rect 22259 1163 22260 1189
rect 22232 1162 22260 1163
rect 22284 1189 22312 1190
rect 22284 1163 22285 1189
rect 22285 1163 22311 1189
rect 22311 1163 22312 1189
rect 22284 1162 22312 1163
rect 22336 1189 22364 1190
rect 22336 1163 22337 1189
rect 22337 1163 22363 1189
rect 22363 1163 22364 1189
rect 22336 1162 22364 1163
rect 22470 1358 22498 1386
rect 22750 966 22778 994
rect 22414 686 22442 714
rect 22246 601 22274 602
rect 22246 575 22247 601
rect 22247 575 22273 601
rect 22273 575 22274 601
rect 22246 574 22274 575
rect 22526 489 22554 490
rect 22526 463 22527 489
rect 22527 463 22553 489
rect 22553 463 22554 489
rect 22526 462 22554 463
rect 22134 406 22162 434
rect 22232 405 22260 406
rect 22232 379 22233 405
rect 22233 379 22259 405
rect 22259 379 22260 405
rect 22232 378 22260 379
rect 22284 405 22312 406
rect 22284 379 22285 405
rect 22285 379 22311 405
rect 22311 379 22312 405
rect 22284 378 22312 379
rect 22336 405 22364 406
rect 22336 379 22337 405
rect 22337 379 22363 405
rect 22363 379 22364 405
rect 22336 378 22364 379
rect 22750 406 22778 434
rect 22302 294 22330 322
rect 21854 238 21882 266
rect 22078 70 22106 98
rect 22526 182 22554 210
rect 22862 1329 22890 1330
rect 22862 1303 22863 1329
rect 22863 1303 22889 1329
rect 22889 1303 22890 1329
rect 22862 1302 22890 1303
rect 23030 2478 23058 2506
rect 22918 462 22946 490
rect 22974 854 23002 882
rect 22806 294 22834 322
rect 23366 2142 23394 2170
rect 23142 2113 23170 2114
rect 23142 2087 23143 2113
rect 23143 2087 23169 2113
rect 23169 2087 23170 2113
rect 23142 2086 23170 2087
rect 23310 2030 23338 2058
rect 23198 1750 23226 1778
rect 23030 742 23058 770
rect 23086 70 23114 98
rect 23758 2982 23786 3010
rect 23478 2673 23506 2674
rect 23478 2647 23479 2673
rect 23479 2647 23505 2673
rect 23505 2647 23506 2673
rect 23478 2646 23506 2647
rect 23926 2590 23954 2618
rect 24038 2814 24066 2842
rect 23590 2534 23618 2562
rect 23590 1750 23618 1778
rect 23478 1721 23506 1722
rect 23478 1695 23479 1721
rect 23479 1695 23505 1721
rect 23505 1695 23506 1721
rect 23478 1694 23506 1695
rect 23870 1638 23898 1666
rect 23646 1414 23674 1442
rect 23646 937 23674 938
rect 23646 911 23647 937
rect 23647 911 23673 937
rect 23673 911 23674 937
rect 23646 910 23674 911
rect 23422 574 23450 602
rect 23366 126 23394 154
rect 23646 238 23674 266
rect 23646 126 23674 154
rect 23926 854 23954 882
rect 24318 5222 24346 5250
rect 24542 6454 24570 6482
rect 25886 6481 25914 6482
rect 25886 6455 25887 6481
rect 25887 6455 25913 6481
rect 25913 6455 25914 6481
rect 25886 6454 25914 6455
rect 25494 6006 25522 6034
rect 24542 5334 24570 5362
rect 24318 3654 24346 3682
rect 24486 3822 24514 3850
rect 24374 2254 24402 2282
rect 24262 798 24290 826
rect 24318 1638 24346 1666
rect 24206 686 24234 714
rect 24150 630 24178 658
rect 24430 1694 24458 1722
rect 24374 1358 24402 1386
rect 24598 2953 24626 2954
rect 24598 2927 24599 2953
rect 24599 2927 24625 2953
rect 24625 2927 24626 2953
rect 24598 2926 24626 2927
rect 24710 2953 24738 2954
rect 24710 2927 24711 2953
rect 24711 2927 24737 2953
rect 24737 2927 24738 2953
rect 24710 2926 24738 2927
rect 24710 2310 24738 2338
rect 24654 1694 24682 1722
rect 25270 5894 25298 5922
rect 25046 5614 25074 5642
rect 24990 2897 25018 2898
rect 24990 2871 24991 2897
rect 24991 2871 25017 2897
rect 25017 2871 25018 2897
rect 24990 2870 25018 2871
rect 24990 1918 25018 1946
rect 24766 1638 24794 1666
rect 24822 1862 24850 1890
rect 24710 574 24738 602
rect 24374 406 24402 434
rect 24430 182 24458 210
rect 24542 462 24570 490
rect 24990 798 25018 826
rect 25158 4830 25186 4858
rect 25886 5753 25914 5754
rect 25886 5727 25887 5753
rect 25887 5727 25913 5753
rect 25913 5727 25914 5753
rect 25886 5726 25914 5727
rect 25270 4494 25298 4522
rect 25718 5390 25746 5418
rect 25214 4438 25242 4466
rect 25214 3766 25242 3794
rect 25158 2982 25186 3010
rect 25046 742 25074 770
rect 25102 2590 25130 2618
rect 25494 2534 25522 2562
rect 25382 1862 25410 1890
rect 25326 1273 25354 1274
rect 25326 1247 25327 1273
rect 25327 1247 25353 1273
rect 25353 1247 25354 1273
rect 25326 1246 25354 1247
rect 25438 1273 25466 1274
rect 25438 1247 25439 1273
rect 25439 1247 25465 1273
rect 25465 1247 25466 1273
rect 25438 1246 25466 1247
rect 25270 126 25298 154
rect 25438 742 25466 770
rect 25102 70 25130 98
rect 25214 70 25242 98
rect 25606 2422 25634 2450
rect 25662 1777 25690 1778
rect 25662 1751 25663 1777
rect 25663 1751 25689 1777
rect 25689 1751 25690 1777
rect 25662 1750 25690 1751
rect 25830 5334 25858 5362
rect 26054 5166 26082 5194
rect 26110 5110 26138 5138
rect 26334 6454 26362 6482
rect 26222 5558 26250 5586
rect 26278 4969 26306 4970
rect 26278 4943 26279 4969
rect 26279 4943 26305 4969
rect 26305 4943 26306 4969
rect 26278 4942 26306 4943
rect 26222 4774 26250 4802
rect 26278 4214 26306 4242
rect 27510 6398 27538 6426
rect 26502 6201 26530 6202
rect 26502 6175 26503 6201
rect 26503 6175 26529 6201
rect 26529 6175 26530 6201
rect 26502 6174 26530 6175
rect 26782 6089 26810 6090
rect 26782 6063 26783 6089
rect 26783 6063 26809 6089
rect 26809 6063 26810 6089
rect 26782 6062 26810 6063
rect 27174 6033 27202 6034
rect 27174 6007 27175 6033
rect 27175 6007 27201 6033
rect 27201 6007 27202 6033
rect 27174 6006 27202 6007
rect 26782 5502 26810 5530
rect 26502 5446 26530 5474
rect 27062 5278 27090 5306
rect 26782 5249 26810 5250
rect 26782 5223 26783 5249
rect 26783 5223 26809 5249
rect 26809 5223 26810 5249
rect 26782 5222 26810 5223
rect 26390 4998 26418 5026
rect 26838 5110 26866 5138
rect 26782 4857 26810 4858
rect 26782 4831 26783 4857
rect 26783 4831 26809 4857
rect 26809 4831 26810 4857
rect 26782 4830 26810 4831
rect 26782 4465 26810 4466
rect 26782 4439 26783 4465
rect 26783 4439 26809 4465
rect 26809 4439 26810 4465
rect 26782 4438 26810 4439
rect 26782 3737 26810 3738
rect 26782 3711 26783 3737
rect 26783 3711 26809 3737
rect 26809 3711 26810 3737
rect 26782 3710 26810 3711
rect 26726 3486 26754 3514
rect 26502 3262 26530 3290
rect 26390 2870 26418 2898
rect 26110 2057 26138 2058
rect 26110 2031 26111 2057
rect 26111 2031 26137 2057
rect 26137 2031 26138 2057
rect 26110 2030 26138 2031
rect 26110 1833 26138 1834
rect 26110 1807 26111 1833
rect 26111 1807 26137 1833
rect 26137 1807 26138 1833
rect 26110 1806 26138 1807
rect 26222 1806 26250 1834
rect 25774 1750 25802 1778
rect 26222 1694 26250 1722
rect 25998 1078 26026 1106
rect 25718 1022 25746 1050
rect 25998 854 26026 882
rect 26278 966 26306 994
rect 26110 686 26138 714
rect 25998 462 26026 490
rect 25886 70 25914 98
rect 26446 2617 26474 2618
rect 26446 2591 26447 2617
rect 26447 2591 26473 2617
rect 26473 2591 26474 2617
rect 26446 2590 26474 2591
rect 26614 2646 26642 2674
rect 26614 2057 26642 2058
rect 26614 2031 26615 2057
rect 26615 2031 26641 2057
rect 26641 2031 26642 2057
rect 26614 2030 26642 2031
rect 26558 1582 26586 1610
rect 26502 1441 26530 1442
rect 26502 1415 26503 1441
rect 26503 1415 26529 1441
rect 26529 1415 26530 1441
rect 26502 1414 26530 1415
rect 26782 3038 26810 3066
rect 26782 2169 26810 2170
rect 26782 2143 26783 2169
rect 26783 2143 26809 2169
rect 26809 2143 26810 2169
rect 26782 2142 26810 2143
rect 27286 5054 27314 5082
rect 27062 4913 27090 4914
rect 27062 4887 27063 4913
rect 27063 4887 27089 4913
rect 27089 4887 27090 4913
rect 27062 4886 27090 4887
rect 27118 4774 27146 4802
rect 27062 3430 27090 3458
rect 27062 3206 27090 3234
rect 27062 2758 27090 2786
rect 26894 2505 26922 2506
rect 26894 2479 26895 2505
rect 26895 2479 26921 2505
rect 26921 2479 26922 2505
rect 26894 2478 26922 2479
rect 26838 1862 26866 1890
rect 27174 4270 27202 4298
rect 27454 4185 27482 4186
rect 27454 4159 27455 4185
rect 27455 4159 27481 4185
rect 27481 4159 27482 4185
rect 27454 4158 27482 4159
rect 27286 3598 27314 3626
rect 27286 2926 27314 2954
rect 27454 2561 27482 2562
rect 27454 2535 27455 2561
rect 27455 2535 27481 2561
rect 27481 2535 27482 2561
rect 27454 2534 27482 2535
rect 27286 2281 27314 2282
rect 27286 2255 27287 2281
rect 27287 2255 27313 2281
rect 27313 2255 27314 2281
rect 27286 2254 27314 2255
rect 27230 1806 27258 1834
rect 26782 1721 26810 1722
rect 26782 1695 26783 1721
rect 26783 1695 26809 1721
rect 26809 1695 26810 1721
rect 26782 1694 26810 1695
rect 26782 1385 26810 1386
rect 26782 1359 26783 1385
rect 26783 1359 26809 1385
rect 26809 1359 26810 1385
rect 26782 1358 26810 1359
rect 27062 1049 27090 1050
rect 27062 1023 27063 1049
rect 27063 1023 27089 1049
rect 27089 1023 27090 1049
rect 27062 1022 27090 1023
rect 26782 937 26810 938
rect 26782 911 26783 937
rect 26783 911 26809 937
rect 26809 911 26810 937
rect 26782 910 26810 911
rect 27006 854 27034 882
rect 26782 713 26810 714
rect 26782 687 26783 713
rect 26783 687 26809 713
rect 26809 687 26810 713
rect 26782 686 26810 687
rect 27454 1833 27482 1834
rect 27454 1807 27455 1833
rect 27455 1807 27481 1833
rect 27481 1807 27482 1833
rect 27454 1806 27482 1807
rect 27286 1582 27314 1610
rect 27566 5894 27594 5922
rect 27622 5782 27650 5810
rect 27566 5390 27594 5418
rect 27566 4718 27594 4746
rect 28182 6958 28210 6986
rect 27790 6174 27818 6202
rect 28406 6734 28434 6762
rect 28182 5726 28210 5754
rect 28238 6062 28266 6090
rect 28070 5614 28098 5642
rect 28238 5502 28266 5530
rect 27958 5166 27986 5194
rect 27678 4550 27706 4578
rect 27566 3878 27594 3906
rect 28518 6510 28546 6538
rect 28462 6286 28490 6314
rect 28462 5446 28490 5474
rect 28406 4830 28434 4858
rect 28070 4494 28098 4522
rect 28518 4158 28546 4186
rect 27958 4046 27986 4074
rect 28070 3849 28098 3850
rect 28070 3823 28071 3849
rect 28071 3823 28097 3849
rect 28097 3823 28098 3849
rect 28070 3822 28098 3823
rect 27622 3654 27650 3682
rect 28070 3374 28098 3402
rect 27566 3150 27594 3178
rect 27566 2982 27594 3010
rect 28070 2702 28098 2730
rect 28126 2590 28154 2618
rect 27566 2198 27594 2226
rect 27902 2030 27930 2058
rect 27678 1918 27706 1946
rect 27454 1134 27482 1162
rect 27398 966 27426 994
rect 27566 545 27594 546
rect 27566 519 27567 545
rect 27567 519 27593 545
rect 27593 519 27594 545
rect 27566 518 27594 519
rect 28070 2030 28098 2058
rect 28070 1358 28098 1386
rect 28350 1750 28378 1778
rect 28462 1694 28490 1722
rect 28462 238 28490 266
rect 28518 1414 28546 1442
rect 462 14 490 42
rect 28518 14 28546 42
<< metal3 >>
rect 2249 7014 2254 7042
rect 2282 7014 2534 7042
rect 2562 7014 2567 7042
rect 4937 7014 4942 7042
rect 4970 7014 5334 7042
rect 5362 7014 5367 7042
rect 6281 7014 6286 7042
rect 6314 7014 6510 7042
rect 6538 7014 6543 7042
rect 8969 7014 8974 7042
rect 9002 7014 9198 7042
rect 9226 7014 9231 7042
rect 9921 7014 9926 7042
rect 9954 7014 18466 7042
rect 19721 7014 19726 7042
rect 19754 7014 19950 7042
rect 19978 7014 19983 7042
rect 22409 7014 22414 7042
rect 22442 7014 22582 7042
rect 22610 7014 22615 7042
rect 23753 7014 23758 7042
rect 23786 7014 23982 7042
rect 24010 7014 24015 7042
rect 25097 7014 25102 7042
rect 25130 7014 25382 7042
rect 25410 7014 25415 7042
rect 0 6986 56 7000
rect 0 6958 3542 6986
rect 3570 6958 3575 6986
rect 0 6944 56 6958
rect 18438 6930 18466 7014
rect 28672 6986 28728 7000
rect 28177 6958 28182 6986
rect 28210 6958 28728 6986
rect 28672 6944 28728 6958
rect 3649 6902 3654 6930
rect 3682 6902 16086 6930
rect 16114 6902 16119 6930
rect 18433 6902 18438 6930
rect 18466 6902 18471 6930
rect 8465 6846 8470 6874
rect 8498 6846 12838 6874
rect 12866 6846 12871 6874
rect 4041 6790 4046 6818
rect 4074 6790 24990 6818
rect 25018 6790 25023 6818
rect 0 6762 56 6776
rect 28672 6762 28728 6776
rect 0 6734 11550 6762
rect 11578 6734 11583 6762
rect 11657 6734 11662 6762
rect 11690 6734 12054 6762
rect 12082 6734 12087 6762
rect 12166 6734 15190 6762
rect 15218 6734 15223 6762
rect 18377 6734 18382 6762
rect 18410 6734 18606 6762
rect 18634 6734 18639 6762
rect 21065 6734 21070 6762
rect 21098 6734 21574 6762
rect 21602 6734 21607 6762
rect 28401 6734 28406 6762
rect 28434 6734 28728 6762
rect 0 6720 56 6734
rect 12166 6706 12194 6734
rect 28672 6720 28728 6734
rect 8409 6678 8414 6706
rect 8442 6678 12194 6706
rect 12889 6678 12894 6706
rect 12922 6678 21854 6706
rect 2227 6650 2232 6678
rect 2260 6650 2284 6678
rect 2312 6650 2336 6678
rect 2364 6650 2369 6678
rect 12227 6650 12232 6678
rect 12260 6650 12284 6678
rect 12312 6650 12336 6678
rect 12364 6650 12369 6678
rect 13113 6622 13118 6650
rect 13146 6622 21406 6650
rect 21434 6622 21439 6650
rect 21826 6594 21854 6678
rect 22227 6650 22232 6678
rect 22260 6650 22284 6678
rect 22312 6650 22336 6678
rect 22364 6650 22369 6678
rect 5273 6566 5278 6594
rect 5306 6566 13286 6594
rect 13314 6566 13319 6594
rect 21826 6566 23254 6594
rect 23282 6566 23287 6594
rect 0 6538 56 6552
rect 28672 6538 28728 6552
rect 0 6510 798 6538
rect 826 6510 831 6538
rect 10761 6510 10766 6538
rect 10794 6510 23646 6538
rect 23674 6510 23679 6538
rect 28513 6510 28518 6538
rect 28546 6510 28728 6538
rect 0 6496 56 6510
rect 28672 6496 28728 6510
rect 3481 6454 3486 6482
rect 3514 6454 8190 6482
rect 8218 6454 8223 6482
rect 9697 6454 9702 6482
rect 9730 6454 10318 6482
rect 10346 6454 10351 6482
rect 16417 6454 16422 6482
rect 16450 6454 17038 6482
rect 17066 6454 17071 6482
rect 22073 6454 22078 6482
rect 22106 6454 24542 6482
rect 24570 6454 24575 6482
rect 25881 6454 25886 6482
rect 25914 6454 26334 6482
rect 26362 6454 26367 6482
rect 7513 6398 7518 6426
rect 7546 6398 27510 6426
rect 27538 6398 27543 6426
rect 5665 6342 5670 6370
rect 5698 6342 18214 6370
rect 18242 6342 18247 6370
rect 0 6314 56 6328
rect 28672 6314 28728 6328
rect 0 6286 1834 6314
rect 28457 6286 28462 6314
rect 28490 6286 28728 6314
rect 0 6272 56 6286
rect 1806 6202 1834 6286
rect 1897 6258 1902 6286
rect 1930 6258 1954 6286
rect 1982 6258 2006 6286
rect 2034 6258 2039 6286
rect 11897 6258 11902 6286
rect 11930 6258 11954 6286
rect 11982 6258 12006 6286
rect 12034 6258 12039 6286
rect 21897 6258 21902 6286
rect 21930 6258 21954 6286
rect 21982 6258 22006 6286
rect 22034 6258 22039 6286
rect 28672 6272 28728 6286
rect 12441 6230 12446 6258
rect 12474 6230 16534 6258
rect 16562 6230 16567 6258
rect 1806 6174 3374 6202
rect 3402 6174 3407 6202
rect 6841 6174 6846 6202
rect 6874 6174 16758 6202
rect 16786 6174 16791 6202
rect 26497 6174 26502 6202
rect 26530 6174 27790 6202
rect 27818 6174 27823 6202
rect 3873 6118 3878 6146
rect 3906 6118 12446 6146
rect 12474 6118 12479 6146
rect 12553 6118 12558 6146
rect 12586 6118 13230 6146
rect 13258 6118 13263 6146
rect 19105 6118 19110 6146
rect 19138 6118 19950 6146
rect 19978 6118 19983 6146
rect 0 6090 56 6104
rect 28672 6090 28728 6104
rect 0 6062 406 6090
rect 434 6062 439 6090
rect 6673 6062 6678 6090
rect 6706 6062 14014 6090
rect 14042 6062 14238 6090
rect 14266 6062 14271 6090
rect 14513 6062 14518 6090
rect 14546 6062 26782 6090
rect 26810 6062 26815 6090
rect 28233 6062 28238 6090
rect 28266 6062 28728 6090
rect 0 6048 56 6062
rect 28672 6048 28728 6062
rect 3425 6006 3430 6034
rect 3458 6006 6622 6034
rect 6650 6006 6655 6034
rect 8017 6006 8022 6034
rect 8050 6006 12950 6034
rect 12978 6006 12983 6034
rect 15129 6006 15134 6034
rect 15162 6006 16310 6034
rect 16338 6006 16343 6034
rect 17761 6006 17766 6034
rect 17794 6006 18550 6034
rect 18578 6006 18583 6034
rect 20225 6006 20230 6034
rect 20258 6006 20398 6034
rect 20426 6006 22414 6034
rect 22442 6006 22447 6034
rect 23697 6006 23702 6034
rect 23730 6006 25494 6034
rect 25522 6006 25527 6034
rect 27169 6006 27174 6034
rect 27202 6006 27734 6034
rect 18041 5950 18046 5978
rect 18074 5950 22302 5978
rect 22330 5950 22335 5978
rect 25265 5894 25270 5922
rect 25298 5894 27566 5922
rect 27594 5894 27599 5922
rect 0 5866 56 5880
rect 2227 5866 2232 5894
rect 2260 5866 2284 5894
rect 2312 5866 2336 5894
rect 2364 5866 2369 5894
rect 12227 5866 12232 5894
rect 12260 5866 12284 5894
rect 12312 5866 12336 5894
rect 12364 5866 12369 5894
rect 22227 5866 22232 5894
rect 22260 5866 22284 5894
rect 22312 5866 22336 5894
rect 22364 5866 22369 5894
rect 27706 5866 27734 6006
rect 28672 5866 28728 5880
rect 0 5838 2114 5866
rect 3369 5838 3374 5866
rect 3402 5838 10094 5866
rect 13505 5838 13510 5866
rect 13538 5838 13678 5866
rect 13706 5838 13711 5866
rect 15185 5838 15190 5866
rect 15218 5838 22134 5866
rect 22162 5838 22167 5866
rect 27706 5838 28728 5866
rect 0 5824 56 5838
rect 2086 5810 2114 5838
rect 10066 5810 10094 5838
rect 28672 5824 28728 5838
rect 2086 5782 6678 5810
rect 6706 5782 6711 5810
rect 7401 5782 7406 5810
rect 7434 5782 7518 5810
rect 7546 5782 8414 5810
rect 8442 5782 8447 5810
rect 10066 5782 17094 5810
rect 17122 5782 17127 5810
rect 17201 5782 17206 5810
rect 17234 5782 27622 5810
rect 27650 5782 27655 5810
rect 3033 5726 3038 5754
rect 3066 5726 6846 5754
rect 6874 5726 6879 5754
rect 8353 5726 8358 5754
rect 8386 5726 9086 5754
rect 9114 5726 9119 5754
rect 11153 5726 11158 5754
rect 11186 5726 13454 5754
rect 13482 5726 13487 5754
rect 16753 5726 16758 5754
rect 16786 5726 23534 5754
rect 23562 5726 23567 5754
rect 25881 5726 25886 5754
rect 25914 5726 28182 5754
rect 28210 5726 28215 5754
rect 9361 5670 9366 5698
rect 9394 5670 9478 5698
rect 9506 5670 24262 5698
rect 24290 5670 24295 5698
rect 0 5642 56 5656
rect 28672 5642 28728 5656
rect 0 5614 3374 5642
rect 3402 5614 3407 5642
rect 5105 5614 5110 5642
rect 5138 5614 8470 5642
rect 8498 5614 8503 5642
rect 11993 5614 11998 5642
rect 12026 5614 12278 5642
rect 12306 5614 12311 5642
rect 12838 5614 25046 5642
rect 25074 5614 25079 5642
rect 28065 5614 28070 5642
rect 28098 5614 28728 5642
rect 0 5600 56 5614
rect 12838 5586 12866 5614
rect 28672 5600 28728 5614
rect 1185 5558 1190 5586
rect 1218 5558 8358 5586
rect 8386 5558 8391 5586
rect 8470 5558 9926 5586
rect 9954 5558 9959 5586
rect 11545 5558 11550 5586
rect 11578 5558 12866 5586
rect 13001 5558 13006 5586
rect 13034 5558 17710 5586
rect 17738 5558 17743 5586
rect 17817 5558 17822 5586
rect 17850 5558 26222 5586
rect 26250 5558 26255 5586
rect 8470 5530 8498 5558
rect 2921 5502 2926 5530
rect 2954 5502 8498 5530
rect 8577 5502 8582 5530
rect 8610 5502 11774 5530
rect 11802 5502 11807 5530
rect 16473 5502 16478 5530
rect 16506 5502 17206 5530
rect 17234 5502 17239 5530
rect 26777 5502 26782 5530
rect 26810 5502 28238 5530
rect 28266 5502 28271 5530
rect 1897 5474 1902 5502
rect 1930 5474 1954 5502
rect 1982 5474 2006 5502
rect 2034 5474 2039 5502
rect 11897 5474 11902 5502
rect 11930 5474 11954 5502
rect 11982 5474 12006 5502
rect 12034 5474 12039 5502
rect 21897 5474 21902 5502
rect 21930 5474 21954 5502
rect 21982 5474 22006 5502
rect 22034 5474 22039 5502
rect 3537 5446 3542 5474
rect 3570 5446 9366 5474
rect 9394 5446 9399 5474
rect 12161 5446 12166 5474
rect 12194 5446 14294 5474
rect 14322 5446 14327 5474
rect 15969 5446 15974 5474
rect 16002 5446 17374 5474
rect 17402 5446 17407 5474
rect 26497 5446 26502 5474
rect 26530 5446 28462 5474
rect 28490 5446 28495 5474
rect 0 5418 56 5432
rect 28672 5418 28728 5432
rect 0 5390 3430 5418
rect 3458 5390 3463 5418
rect 7345 5390 7350 5418
rect 7378 5390 11830 5418
rect 11858 5390 11863 5418
rect 11937 5390 11942 5418
rect 11970 5390 13510 5418
rect 13538 5390 13543 5418
rect 13673 5390 13678 5418
rect 13706 5390 25718 5418
rect 25746 5390 25751 5418
rect 27561 5390 27566 5418
rect 27594 5390 28728 5418
rect 0 5376 56 5390
rect 28672 5376 28728 5390
rect 9921 5334 9926 5362
rect 9954 5334 10094 5362
rect 10201 5334 10206 5362
rect 10234 5334 12586 5362
rect 13561 5334 13566 5362
rect 13594 5334 14350 5362
rect 14378 5334 14383 5362
rect 14625 5334 14630 5362
rect 14658 5334 14798 5362
rect 14826 5334 19670 5362
rect 19698 5334 19703 5362
rect 22129 5334 22134 5362
rect 22162 5334 22470 5362
rect 22498 5334 22503 5362
rect 24537 5334 24542 5362
rect 24570 5334 25830 5362
rect 25858 5334 25863 5362
rect 10066 5306 10094 5334
rect 12558 5306 12586 5334
rect 793 5278 798 5306
rect 826 5278 4214 5306
rect 8129 5278 8134 5306
rect 8162 5278 9786 5306
rect 10066 5278 11718 5306
rect 11746 5278 11751 5306
rect 12558 5278 14854 5306
rect 14882 5278 14887 5306
rect 19273 5278 19278 5306
rect 19306 5278 27062 5306
rect 27090 5278 27095 5306
rect 401 5222 406 5250
rect 434 5222 3822 5250
rect 3850 5222 3855 5250
rect 0 5194 56 5208
rect 4186 5194 4214 5278
rect 9758 5250 9786 5278
rect 7569 5222 7574 5250
rect 7602 5222 9730 5250
rect 9758 5222 11158 5250
rect 11186 5222 11191 5250
rect 11265 5222 11270 5250
rect 11298 5222 13118 5250
rect 13146 5222 13151 5250
rect 13897 5222 13902 5250
rect 13930 5222 16758 5250
rect 16786 5222 16791 5250
rect 24313 5222 24318 5250
rect 24346 5222 26782 5250
rect 26810 5222 26815 5250
rect 0 5166 798 5194
rect 826 5166 831 5194
rect 4186 5166 9590 5194
rect 9618 5166 9623 5194
rect 0 5152 56 5166
rect 9702 5138 9730 5222
rect 28672 5194 28728 5208
rect 9865 5166 9870 5194
rect 9898 5166 15246 5194
rect 15274 5166 15414 5194
rect 15442 5166 15447 5194
rect 17537 5166 17542 5194
rect 17570 5166 26054 5194
rect 26082 5166 26087 5194
rect 27953 5166 27958 5194
rect 27986 5166 28728 5194
rect 28672 5152 28728 5166
rect 6617 5110 6622 5138
rect 6650 5110 7686 5138
rect 7714 5110 7719 5138
rect 8409 5110 8414 5138
rect 8442 5110 9534 5138
rect 9562 5110 9567 5138
rect 9702 5110 11662 5138
rect 11690 5110 11695 5138
rect 14345 5110 14350 5138
rect 14378 5110 18326 5138
rect 18354 5110 18359 5138
rect 26105 5110 26110 5138
rect 26138 5110 26838 5138
rect 26866 5110 26871 5138
rect 2227 5082 2232 5110
rect 2260 5082 2284 5110
rect 2312 5082 2336 5110
rect 2364 5082 2369 5110
rect 12227 5082 12232 5110
rect 12260 5082 12284 5110
rect 12312 5082 12336 5110
rect 12364 5082 12369 5110
rect 22227 5082 22232 5110
rect 22260 5082 22284 5110
rect 22312 5082 22336 5110
rect 22364 5082 22369 5110
rect 3425 5054 3430 5082
rect 3458 5054 7518 5082
rect 7546 5054 7551 5082
rect 8414 5054 10094 5082
rect 10145 5054 10150 5082
rect 10178 5054 12166 5082
rect 12194 5054 12199 5082
rect 12945 5054 12950 5082
rect 12978 5054 17206 5082
rect 17234 5054 17239 5082
rect 27281 5054 27286 5082
rect 27314 5054 27734 5082
rect 8414 5026 8442 5054
rect 3369 4998 3374 5026
rect 3402 4998 8442 5026
rect 10066 5026 10094 5054
rect 10066 4998 11634 5026
rect 11713 4998 11718 5026
rect 11746 4998 14350 5026
rect 14378 4998 14383 5026
rect 17593 4998 17598 5026
rect 17626 4998 26390 5026
rect 26418 4998 26423 5026
rect 0 4970 56 4984
rect 11606 4970 11634 4998
rect 27706 4970 27734 5054
rect 28672 4970 28728 4984
rect 0 4942 574 4970
rect 602 4942 607 4970
rect 4321 4942 4326 4970
rect 4354 4942 7182 4970
rect 7210 4942 7215 4970
rect 7513 4942 7518 4970
rect 7546 4942 9870 4970
rect 9898 4942 9903 4970
rect 11606 4942 12614 4970
rect 12642 4942 12647 4970
rect 13393 4942 13398 4970
rect 13426 4942 26278 4970
rect 26306 4942 26311 4970
rect 27706 4942 28728 4970
rect 0 4928 56 4942
rect 28672 4928 28728 4942
rect 7121 4886 7126 4914
rect 7154 4886 12726 4914
rect 12754 4886 12759 4914
rect 13729 4886 13734 4914
rect 13762 4886 27062 4914
rect 27090 4886 27095 4914
rect 2081 4830 2086 4858
rect 2114 4830 7574 4858
rect 7602 4830 7607 4858
rect 7681 4830 7686 4858
rect 7714 4830 9338 4858
rect 9977 4830 9982 4858
rect 10010 4830 25158 4858
rect 25186 4830 25191 4858
rect 26777 4830 26782 4858
rect 26810 4830 28406 4858
rect 28434 4830 28439 4858
rect 9310 4802 9338 4830
rect 1806 4774 9198 4802
rect 9226 4774 9231 4802
rect 9310 4774 11046 4802
rect 11074 4774 11079 4802
rect 11550 4774 13958 4802
rect 13986 4774 13991 4802
rect 16697 4774 16702 4802
rect 16730 4774 24206 4802
rect 24234 4774 24239 4802
rect 26217 4774 26222 4802
rect 26250 4774 27118 4802
rect 27146 4774 27151 4802
rect 0 4746 56 4760
rect 1806 4746 1834 4774
rect 0 4718 1834 4746
rect 7177 4718 7182 4746
rect 7210 4718 10038 4746
rect 10066 4718 10071 4746
rect 0 4704 56 4718
rect 1897 4690 1902 4718
rect 1930 4690 1954 4718
rect 1982 4690 2006 4718
rect 2034 4690 2039 4718
rect 5161 4662 5166 4690
rect 5194 4662 8974 4690
rect 9002 4662 9007 4690
rect 11550 4634 11578 4774
rect 28672 4746 28728 4760
rect 12105 4718 12110 4746
rect 12138 4718 13398 4746
rect 13426 4718 13431 4746
rect 13505 4718 13510 4746
rect 13538 4718 16814 4746
rect 16842 4718 16847 4746
rect 27561 4718 27566 4746
rect 27594 4718 28728 4746
rect 11897 4690 11902 4718
rect 11930 4690 11954 4718
rect 11982 4690 12006 4718
rect 12034 4690 12039 4718
rect 21897 4690 21902 4718
rect 21930 4690 21954 4718
rect 21982 4690 22006 4718
rect 22034 4690 22039 4718
rect 28672 4704 28728 4718
rect 12161 4662 12166 4690
rect 12194 4662 13006 4690
rect 13034 4662 13039 4690
rect 13449 4662 13454 4690
rect 13482 4662 14378 4690
rect 14350 4634 14378 4662
rect 737 4606 742 4634
rect 770 4606 8358 4634
rect 8386 4606 8391 4634
rect 8465 4606 8470 4634
rect 8498 4606 11578 4634
rect 11657 4606 11662 4634
rect 11690 4606 14014 4634
rect 14042 4606 14238 4634
rect 14266 4606 14271 4634
rect 14350 4606 15974 4634
rect 16002 4606 16007 4634
rect 17033 4606 17038 4634
rect 17066 4606 24150 4634
rect 24178 4606 24183 4634
rect 793 4550 798 4578
rect 826 4550 11158 4578
rect 11186 4550 11326 4578
rect 11354 4550 11359 4578
rect 12609 4550 12614 4578
rect 12642 4550 12782 4578
rect 12810 4550 12815 4578
rect 13057 4550 13062 4578
rect 13090 4550 27678 4578
rect 27706 4550 27711 4578
rect 0 4522 56 4536
rect 28672 4522 28728 4536
rect 0 4494 10150 4522
rect 10178 4494 10183 4522
rect 11601 4494 11606 4522
rect 11634 4494 25270 4522
rect 25298 4494 25303 4522
rect 28065 4494 28070 4522
rect 28098 4494 28728 4522
rect 0 4480 56 4494
rect 28672 4480 28728 4494
rect 1465 4438 1470 4466
rect 1498 4438 4270 4466
rect 4298 4438 4303 4466
rect 6505 4438 6510 4466
rect 6538 4438 8470 4466
rect 8498 4438 8503 4466
rect 8801 4438 8806 4466
rect 8834 4438 12614 4466
rect 12642 4438 12647 4466
rect 13449 4438 13454 4466
rect 13482 4438 20454 4466
rect 20482 4438 20566 4466
rect 20594 4438 20599 4466
rect 20841 4438 20846 4466
rect 20874 4438 21182 4466
rect 21210 4438 21215 4466
rect 22353 4438 22358 4466
rect 22386 4438 22974 4466
rect 23002 4438 23007 4466
rect 25209 4438 25214 4466
rect 25242 4438 26782 4466
rect 26810 4438 26815 4466
rect 2086 4382 3430 4410
rect 3458 4382 3463 4410
rect 7457 4382 7462 4410
rect 7490 4382 9926 4410
rect 9954 4382 9959 4410
rect 11489 4382 11494 4410
rect 11522 4382 13734 4410
rect 13762 4382 13767 4410
rect 13841 4382 13846 4410
rect 13874 4382 15022 4410
rect 15050 4382 15055 4410
rect 18433 4382 18438 4410
rect 18466 4382 21854 4410
rect 21882 4382 21887 4410
rect 0 4298 56 4312
rect 2086 4298 2114 4382
rect 8577 4326 8582 4354
rect 8610 4326 12166 4354
rect 12194 4326 12199 4354
rect 12609 4326 12614 4354
rect 12642 4326 13398 4354
rect 13426 4326 13431 4354
rect 13729 4326 13734 4354
rect 13762 4326 18158 4354
rect 18186 4326 18191 4354
rect 2227 4298 2232 4326
rect 2260 4298 2284 4326
rect 2312 4298 2336 4326
rect 2364 4298 2369 4326
rect 12227 4298 12232 4326
rect 12260 4298 12284 4326
rect 12312 4298 12336 4326
rect 12364 4298 12369 4326
rect 22227 4298 22232 4326
rect 22260 4298 22284 4326
rect 22312 4298 22336 4326
rect 22364 4298 22369 4326
rect 28672 4298 28728 4312
rect 0 4270 2114 4298
rect 4186 4270 7126 4298
rect 7154 4270 7159 4298
rect 8241 4270 8246 4298
rect 8274 4270 12138 4298
rect 0 4256 56 4270
rect 4186 4242 4214 4270
rect 12110 4242 12138 4270
rect 12446 4270 14182 4298
rect 14210 4270 14215 4298
rect 15974 4270 18382 4298
rect 18410 4270 18415 4298
rect 27169 4270 27174 4298
rect 27202 4270 28728 4298
rect 12446 4242 12474 4270
rect 3425 4214 3430 4242
rect 3458 4214 4214 4242
rect 5049 4214 5054 4242
rect 5082 4214 7658 4242
rect 8353 4214 8358 4242
rect 8386 4214 11774 4242
rect 12110 4214 12474 4242
rect 12833 4214 12838 4242
rect 12866 4214 13846 4242
rect 13874 4214 13879 4242
rect 14009 4214 14014 4242
rect 14042 4214 15806 4242
rect 15834 4214 15839 4242
rect 289 4158 294 4186
rect 322 4158 7462 4186
rect 7490 4158 7495 4186
rect 7630 4130 7658 4214
rect 11746 4186 11774 4214
rect 15974 4186 16002 4270
rect 28672 4256 28728 4270
rect 9193 4158 9198 4186
rect 9226 4158 11102 4186
rect 11130 4158 11214 4186
rect 11242 4158 11247 4186
rect 11746 4158 12782 4186
rect 12810 4158 12815 4186
rect 13393 4158 13398 4186
rect 13426 4158 16002 4186
rect 16030 4214 26278 4242
rect 26306 4214 26311 4242
rect 16030 4130 16058 4214
rect 27449 4158 27454 4186
rect 27482 4158 28518 4186
rect 28546 4158 28551 4186
rect 7630 4102 14770 4130
rect 14849 4102 14854 4130
rect 14882 4102 16058 4130
rect 0 4074 56 4088
rect 14742 4074 14770 4102
rect 28672 4074 28728 4088
rect 0 4046 4942 4074
rect 4970 4046 4975 4074
rect 9249 4046 9254 4074
rect 9282 4046 9982 4074
rect 10010 4046 10015 4074
rect 10089 4046 10094 4074
rect 10122 4046 14518 4074
rect 14546 4046 14551 4074
rect 14742 4046 14966 4074
rect 14994 4046 14999 4074
rect 18713 4046 18718 4074
rect 18746 4046 21630 4074
rect 21658 4046 21798 4074
rect 21826 4046 21831 4074
rect 22073 4046 22078 4074
rect 22106 4046 22750 4074
rect 22778 4046 22783 4074
rect 27953 4046 27958 4074
rect 27986 4046 28728 4074
rect 0 4032 56 4046
rect 28672 4032 28728 4046
rect 1801 3990 1806 4018
rect 1834 3990 15190 4018
rect 15218 3990 15358 4018
rect 15386 3990 15391 4018
rect 15465 3990 15470 4018
rect 15498 3990 23366 4018
rect 23394 3990 23399 4018
rect 8913 3934 8918 3962
rect 8946 3934 11494 3962
rect 11522 3934 11527 3962
rect 12609 3934 12614 3962
rect 12642 3934 18830 3962
rect 18858 3934 18863 3962
rect 1897 3906 1902 3934
rect 1930 3906 1954 3934
rect 1982 3906 2006 3934
rect 2034 3906 2039 3934
rect 11897 3906 11902 3934
rect 11930 3906 11954 3934
rect 11982 3906 12006 3934
rect 12034 3906 12039 3934
rect 21897 3906 21902 3934
rect 21930 3906 21954 3934
rect 21982 3906 22006 3934
rect 22034 3906 22039 3934
rect 9249 3878 9254 3906
rect 9282 3878 11270 3906
rect 11298 3878 11303 3906
rect 12161 3878 12166 3906
rect 12194 3878 15078 3906
rect 15106 3878 15111 3906
rect 15969 3878 15974 3906
rect 16002 3878 18550 3906
rect 18578 3878 18583 3906
rect 22969 3878 22974 3906
rect 23002 3878 27566 3906
rect 27594 3878 27599 3906
rect 0 3850 56 3864
rect 28672 3850 28728 3864
rect 0 3822 7910 3850
rect 7938 3822 7943 3850
rect 9753 3822 9758 3850
rect 9786 3822 21910 3850
rect 21938 3822 21943 3850
rect 22129 3822 22134 3850
rect 22162 3822 24486 3850
rect 24514 3822 24519 3850
rect 28065 3822 28070 3850
rect 28098 3822 28728 3850
rect 0 3808 56 3822
rect 28672 3808 28728 3822
rect 3537 3766 3542 3794
rect 3570 3766 10094 3794
rect 10122 3766 10127 3794
rect 11041 3766 11046 3794
rect 11074 3766 12558 3794
rect 12586 3766 12591 3794
rect 12665 3766 12670 3794
rect 12698 3766 15974 3794
rect 16753 3766 16758 3794
rect 16786 3766 17374 3794
rect 17402 3766 17407 3794
rect 17817 3766 17822 3794
rect 17850 3766 25214 3794
rect 25242 3766 25247 3794
rect 15946 3738 15974 3766
rect 569 3710 574 3738
rect 602 3710 4158 3738
rect 4186 3710 4191 3738
rect 10066 3710 12838 3738
rect 12866 3710 12950 3738
rect 12978 3710 12983 3738
rect 15946 3710 26782 3738
rect 26810 3710 26815 3738
rect 10066 3682 10094 3710
rect 3985 3654 3990 3682
rect 4018 3654 10094 3682
rect 11881 3654 11886 3682
rect 11914 3654 13902 3682
rect 13930 3654 13935 3682
rect 14905 3654 14910 3682
rect 14938 3654 24318 3682
rect 24346 3654 24351 3682
rect 24710 3654 27622 3682
rect 27650 3654 27655 3682
rect 0 3626 56 3640
rect 24710 3626 24738 3654
rect 28672 3626 28728 3640
rect 0 3598 2114 3626
rect 2977 3598 2982 3626
rect 3010 3598 3150 3626
rect 3178 3598 3374 3626
rect 3402 3598 3407 3626
rect 4825 3598 4830 3626
rect 4858 3598 4998 3626
rect 5026 3598 7574 3626
rect 7602 3598 7607 3626
rect 10705 3598 10710 3626
rect 10738 3598 24738 3626
rect 27281 3598 27286 3626
rect 27314 3598 28728 3626
rect 0 3584 56 3598
rect 2086 3458 2114 3598
rect 28672 3584 28728 3598
rect 2697 3542 2702 3570
rect 2730 3542 7630 3570
rect 7658 3542 7663 3570
rect 8185 3542 8190 3570
rect 8218 3542 12166 3570
rect 12194 3542 12199 3570
rect 12553 3542 12558 3570
rect 12586 3542 13174 3570
rect 13202 3542 13207 3570
rect 13281 3542 13286 3570
rect 13314 3542 16422 3570
rect 16450 3542 16455 3570
rect 18825 3542 18830 3570
rect 18858 3542 22134 3570
rect 22162 3542 22167 3570
rect 2227 3514 2232 3542
rect 2260 3514 2284 3542
rect 2312 3514 2336 3542
rect 2364 3514 2369 3542
rect 12227 3514 12232 3542
rect 12260 3514 12284 3542
rect 12312 3514 12336 3542
rect 12364 3514 12369 3542
rect 22227 3514 22232 3542
rect 22260 3514 22284 3542
rect 22312 3514 22336 3542
rect 22364 3514 22369 3542
rect 5217 3486 5222 3514
rect 5250 3486 8806 3514
rect 8834 3486 8839 3514
rect 8913 3486 8918 3514
rect 8946 3486 12194 3514
rect 2086 3430 3346 3458
rect 4545 3430 4550 3458
rect 4578 3430 7854 3458
rect 7882 3430 7887 3458
rect 9865 3430 9870 3458
rect 9898 3430 11886 3458
rect 11914 3430 11919 3458
rect 0 3402 56 3416
rect 0 3374 742 3402
rect 770 3374 775 3402
rect 0 3360 56 3374
rect 3318 3346 3346 3430
rect 12166 3402 12194 3486
rect 12502 3486 13118 3514
rect 13146 3486 13151 3514
rect 15689 3486 15694 3514
rect 15722 3486 22106 3514
rect 22409 3486 22414 3514
rect 22442 3486 26726 3514
rect 26754 3486 26759 3514
rect 12502 3402 12530 3486
rect 13225 3430 13230 3458
rect 13258 3430 15974 3458
rect 21826 3430 21882 3486
rect 22078 3458 22106 3486
rect 22078 3430 27062 3458
rect 27090 3430 27095 3458
rect 15946 3402 15974 3430
rect 28672 3402 28728 3416
rect 7462 3374 10262 3402
rect 10290 3374 10295 3402
rect 12166 3374 12530 3402
rect 12558 3374 13482 3402
rect 15946 3374 21966 3402
rect 21994 3374 21999 3402
rect 28065 3374 28070 3402
rect 28098 3374 28728 3402
rect 3318 3318 7350 3346
rect 7378 3318 7383 3346
rect 7462 3290 7490 3374
rect 12558 3346 12586 3374
rect 13454 3346 13482 3374
rect 28672 3360 28728 3374
rect 7569 3318 7574 3346
rect 7602 3318 9254 3346
rect 9282 3318 9287 3346
rect 10066 3318 12586 3346
rect 12721 3318 12726 3346
rect 12754 3318 13370 3346
rect 13454 3318 17486 3346
rect 17514 3318 17519 3346
rect 20785 3318 20790 3346
rect 20818 3318 22694 3346
rect 22722 3318 22727 3346
rect 10066 3290 10094 3318
rect 13342 3290 13370 3318
rect 4937 3262 4942 3290
rect 4970 3262 7490 3290
rect 8414 3262 10094 3290
rect 11433 3262 11438 3290
rect 11466 3262 13062 3290
rect 13090 3262 13230 3290
rect 13258 3262 13263 3290
rect 13342 3262 26502 3290
rect 26530 3262 26535 3290
rect 8414 3234 8442 3262
rect 7233 3206 7238 3234
rect 7266 3206 8442 3234
rect 9641 3206 9646 3234
rect 9674 3206 10934 3234
rect 10962 3206 10967 3234
rect 11830 3206 27062 3234
rect 27090 3206 27095 3234
rect 0 3178 56 3192
rect 11830 3178 11858 3206
rect 28672 3178 28728 3192
rect 0 3150 182 3178
rect 210 3150 215 3178
rect 7009 3150 7014 3178
rect 7042 3150 7574 3178
rect 7602 3150 7607 3178
rect 8073 3150 8078 3178
rect 8106 3150 11858 3178
rect 12553 3150 12558 3178
rect 12586 3150 15890 3178
rect 20337 3150 20342 3178
rect 20370 3150 21798 3178
rect 21826 3150 21831 3178
rect 27561 3150 27566 3178
rect 27594 3150 28728 3178
rect 0 3136 56 3150
rect 1897 3122 1902 3150
rect 1930 3122 1954 3150
rect 1982 3122 2006 3150
rect 2034 3122 2039 3150
rect 11897 3122 11902 3150
rect 11930 3122 11954 3150
rect 11982 3122 12006 3150
rect 12034 3122 12039 3150
rect 15862 3122 15890 3150
rect 21897 3122 21902 3150
rect 21930 3122 21954 3150
rect 21982 3122 22006 3150
rect 22034 3122 22039 3150
rect 28672 3136 28728 3150
rect 3369 3094 3374 3122
rect 3402 3094 7294 3122
rect 7322 3094 7327 3122
rect 7905 3094 7910 3122
rect 7938 3094 8526 3122
rect 8554 3094 8559 3122
rect 9249 3094 9254 3122
rect 9282 3094 10206 3122
rect 10234 3094 10239 3122
rect 10929 3094 10934 3122
rect 10962 3094 11774 3122
rect 11802 3094 11807 3122
rect 12110 3094 15190 3122
rect 15218 3094 15223 3122
rect 15862 3094 21462 3122
rect 21490 3094 21495 3122
rect 22129 3094 22134 3122
rect 22162 3094 23198 3122
rect 23226 3094 23231 3122
rect 12110 3066 12138 3094
rect 7345 3038 7350 3066
rect 7378 3038 8582 3066
rect 8610 3038 8615 3066
rect 10089 3038 10094 3066
rect 10122 3038 12138 3066
rect 12665 3038 12670 3066
rect 12698 3038 20902 3066
rect 20930 3038 20935 3066
rect 21401 3038 21406 3066
rect 21434 3038 26782 3066
rect 26810 3038 26815 3066
rect 1353 2982 1358 3010
rect 1386 2982 5166 3010
rect 5194 2982 5199 3010
rect 8353 2982 8358 3010
rect 8386 2982 13398 3010
rect 13426 2982 13431 3010
rect 15185 2982 15190 3010
rect 15218 2982 15918 3010
rect 15946 2982 15951 3010
rect 21065 2982 21070 3010
rect 21098 2982 23758 3010
rect 23786 2982 23791 3010
rect 25153 2982 25158 3010
rect 25186 2982 27566 3010
rect 27594 2982 27599 3010
rect 0 2954 56 2968
rect 28672 2954 28728 2968
rect 0 2926 3430 2954
rect 3458 2926 3463 2954
rect 7569 2926 7574 2954
rect 7602 2926 8862 2954
rect 8890 2926 8895 2954
rect 12049 2926 12054 2954
rect 12082 2926 12614 2954
rect 12642 2926 12647 2954
rect 12777 2926 12782 2954
rect 12810 2926 18046 2954
rect 18074 2926 18079 2954
rect 18321 2926 18326 2954
rect 18354 2926 24598 2954
rect 24626 2926 24710 2954
rect 24738 2926 24743 2954
rect 27281 2926 27286 2954
rect 27314 2926 28728 2954
rect 0 2912 56 2926
rect 28672 2912 28728 2926
rect 345 2870 350 2898
rect 378 2870 3710 2898
rect 3738 2870 3743 2898
rect 3934 2870 8190 2898
rect 8218 2870 8302 2898
rect 8330 2870 8335 2898
rect 11489 2870 11494 2898
rect 11522 2870 12110 2898
rect 12138 2870 12143 2898
rect 12217 2870 12222 2898
rect 12250 2870 12894 2898
rect 12922 2870 12927 2898
rect 13113 2870 13118 2898
rect 13146 2870 17150 2898
rect 17178 2870 17183 2898
rect 19441 2870 19446 2898
rect 19474 2870 20286 2898
rect 20314 2870 20319 2898
rect 24985 2870 24990 2898
rect 25018 2870 26390 2898
rect 26418 2870 26423 2898
rect 1017 2814 1022 2842
rect 1050 2814 2450 2842
rect 2422 2786 2450 2814
rect 3934 2786 3962 2870
rect 6561 2814 6566 2842
rect 6594 2814 11830 2842
rect 11858 2814 11942 2842
rect 11970 2814 11975 2842
rect 12166 2814 24038 2842
rect 24066 2814 24071 2842
rect 12166 2786 12194 2814
rect 2422 2758 3962 2786
rect 5161 2758 5166 2786
rect 5194 2758 12194 2786
rect 22745 2758 22750 2786
rect 22778 2758 27062 2786
rect 27090 2758 27095 2786
rect 0 2730 56 2744
rect 2227 2730 2232 2758
rect 2260 2730 2284 2758
rect 2312 2730 2336 2758
rect 2364 2730 2369 2758
rect 12227 2730 12232 2758
rect 12260 2730 12284 2758
rect 12312 2730 12336 2758
rect 12364 2730 12369 2758
rect 22227 2730 22232 2758
rect 22260 2730 22284 2758
rect 22312 2730 22336 2758
rect 22364 2730 22369 2758
rect 28672 2730 28728 2744
rect 0 2702 70 2730
rect 98 2702 103 2730
rect 3033 2702 3038 2730
rect 3066 2702 5110 2730
rect 5138 2702 5143 2730
rect 7681 2702 7686 2730
rect 7714 2702 8694 2730
rect 8722 2702 8727 2730
rect 8969 2702 8974 2730
rect 9002 2702 12194 2730
rect 18377 2702 18382 2730
rect 18410 2702 21854 2730
rect 28065 2702 28070 2730
rect 28098 2702 28728 2730
rect 0 2688 56 2702
rect 12166 2674 12194 2702
rect 21826 2674 21854 2702
rect 28672 2688 28728 2702
rect 177 2646 182 2674
rect 210 2646 7630 2674
rect 7658 2646 7663 2674
rect 8409 2646 8414 2674
rect 8442 2646 9142 2674
rect 9170 2646 9310 2674
rect 9338 2646 9343 2674
rect 9417 2646 9422 2674
rect 9450 2646 12054 2674
rect 12082 2646 12087 2674
rect 12166 2646 14294 2674
rect 14322 2646 14462 2674
rect 14490 2646 14495 2674
rect 16809 2646 16814 2674
rect 16842 2646 21126 2674
rect 21154 2646 21294 2674
rect 21322 2646 21327 2674
rect 21826 2646 23310 2674
rect 23338 2646 23478 2674
rect 23506 2646 23511 2674
rect 26609 2646 26614 2674
rect 26642 2646 26647 2674
rect 26614 2618 26642 2646
rect 3593 2590 3598 2618
rect 3626 2590 8302 2618
rect 8330 2590 8335 2618
rect 8582 2590 12838 2618
rect 12866 2590 12871 2618
rect 17593 2590 17598 2618
rect 17626 2590 18606 2618
rect 18634 2590 18639 2618
rect 21826 2590 22918 2618
rect 22946 2590 22951 2618
rect 23921 2590 23926 2618
rect 23954 2590 25102 2618
rect 25130 2590 25135 2618
rect 26441 2590 26446 2618
rect 26474 2590 28126 2618
rect 28154 2590 28159 2618
rect 513 2534 518 2562
rect 546 2534 3878 2562
rect 3906 2534 3911 2562
rect 5441 2534 5446 2562
rect 5474 2534 5558 2562
rect 5586 2534 6958 2562
rect 6986 2534 6991 2562
rect 7569 2534 7574 2562
rect 7602 2534 8470 2562
rect 8498 2534 8503 2562
rect 0 2506 56 2520
rect 8582 2506 8610 2590
rect 21826 2562 21854 2590
rect 8689 2534 8694 2562
rect 8722 2534 9422 2562
rect 9450 2534 9455 2562
rect 10089 2534 10094 2562
rect 10122 2534 10486 2562
rect 10514 2534 10519 2562
rect 11321 2534 11326 2562
rect 11354 2534 12222 2562
rect 12250 2534 12446 2562
rect 12474 2534 12479 2562
rect 15689 2534 15694 2562
rect 15722 2534 17626 2562
rect 18209 2534 18214 2562
rect 18242 2534 21854 2562
rect 23585 2534 23590 2562
rect 23618 2534 25494 2562
rect 25522 2534 25527 2562
rect 27449 2534 27454 2562
rect 27482 2534 27734 2562
rect 17598 2506 17626 2534
rect 27706 2506 27734 2534
rect 28672 2506 28728 2520
rect 0 2478 6454 2506
rect 6482 2478 6487 2506
rect 7121 2478 7126 2506
rect 7154 2478 8610 2506
rect 10705 2478 10710 2506
rect 10738 2478 12558 2506
rect 12586 2478 12591 2506
rect 12665 2478 12670 2506
rect 12698 2478 13734 2506
rect 13762 2478 13767 2506
rect 14345 2478 14350 2506
rect 14378 2478 15974 2506
rect 16002 2478 16007 2506
rect 17598 2478 19110 2506
rect 19138 2478 19278 2506
rect 19306 2478 19311 2506
rect 23025 2478 23030 2506
rect 23058 2478 26894 2506
rect 26922 2478 26927 2506
rect 27706 2478 28728 2506
rect 0 2464 56 2478
rect 28672 2464 28728 2478
rect 4265 2422 4270 2450
rect 4298 2422 5194 2450
rect 8297 2422 8302 2450
rect 8330 2422 11102 2450
rect 11130 2422 11135 2450
rect 11606 2422 13006 2450
rect 13034 2422 13039 2450
rect 13566 2422 18690 2450
rect 18769 2422 18774 2450
rect 18802 2422 19558 2450
rect 19586 2422 19591 2450
rect 20505 2422 20510 2450
rect 20538 2422 25606 2450
rect 25634 2422 25639 2450
rect 5166 2394 5194 2422
rect 3430 2366 5054 2394
rect 5082 2366 5087 2394
rect 5166 2366 9254 2394
rect 9282 2366 9287 2394
rect 1897 2338 1902 2366
rect 1930 2338 1954 2366
rect 1982 2338 2006 2366
rect 2034 2338 2039 2366
rect 0 2282 56 2296
rect 3430 2282 3458 2366
rect 11606 2338 11634 2422
rect 12105 2366 12110 2394
rect 12138 2366 13398 2394
rect 13426 2366 13431 2394
rect 11897 2338 11902 2366
rect 11930 2338 11954 2366
rect 11982 2338 12006 2366
rect 12034 2338 12039 2366
rect 4153 2310 4158 2338
rect 4186 2310 7182 2338
rect 7210 2310 7215 2338
rect 9361 2310 9366 2338
rect 9394 2310 11634 2338
rect 13566 2282 13594 2422
rect 18662 2394 18690 2422
rect 15017 2366 15022 2394
rect 15050 2366 17430 2394
rect 17458 2366 17463 2394
rect 17542 2366 18550 2394
rect 18578 2366 18583 2394
rect 18662 2366 21686 2394
rect 21714 2366 21719 2394
rect 17542 2338 17570 2366
rect 21897 2338 21902 2366
rect 21930 2338 21954 2366
rect 21982 2338 22006 2366
rect 22034 2338 22039 2366
rect 16249 2310 16254 2338
rect 16282 2310 17570 2338
rect 17598 2310 18718 2338
rect 18746 2310 18751 2338
rect 18825 2310 18830 2338
rect 18858 2310 21854 2338
rect 22465 2310 22470 2338
rect 22498 2310 24710 2338
rect 24738 2310 24743 2338
rect 17598 2282 17626 2310
rect 21826 2282 21854 2310
rect 28672 2282 28728 2296
rect 0 2254 3458 2282
rect 3486 2254 4886 2282
rect 4914 2254 4919 2282
rect 4998 2254 8358 2282
rect 8386 2254 8391 2282
rect 8521 2254 8526 2282
rect 8554 2254 10878 2282
rect 10906 2254 10911 2282
rect 11209 2254 11214 2282
rect 11242 2254 13594 2282
rect 13622 2254 17626 2282
rect 17705 2254 17710 2282
rect 17738 2254 20622 2282
rect 20650 2254 20655 2282
rect 21826 2254 24374 2282
rect 24402 2254 24407 2282
rect 27281 2254 27286 2282
rect 27314 2254 28728 2282
rect 0 2240 56 2254
rect 3486 2170 3514 2254
rect 4998 2226 5026 2254
rect 13622 2226 13650 2254
rect 28672 2240 28728 2254
rect 3593 2198 3598 2226
rect 3626 2198 5026 2226
rect 5105 2198 5110 2226
rect 5138 2198 6510 2226
rect 6538 2198 6543 2226
rect 7625 2198 7630 2226
rect 7658 2198 9366 2226
rect 9394 2198 9399 2226
rect 11097 2198 11102 2226
rect 11130 2198 13286 2226
rect 13314 2198 13319 2226
rect 13449 2198 13454 2226
rect 13482 2198 13650 2226
rect 15129 2198 15134 2226
rect 15162 2198 16142 2226
rect 16170 2198 16175 2226
rect 17201 2198 17206 2226
rect 17234 2198 18438 2226
rect 18466 2198 18471 2226
rect 19553 2198 19558 2226
rect 19586 2198 20958 2226
rect 20986 2198 20991 2226
rect 21177 2198 21182 2226
rect 21210 2198 27566 2226
rect 27594 2198 27599 2226
rect 1465 2142 1470 2170
rect 1498 2142 3514 2170
rect 3761 2142 3766 2170
rect 3794 2142 8358 2170
rect 8386 2142 8391 2170
rect 9361 2142 9366 2170
rect 9394 2142 11662 2170
rect 11690 2142 11695 2170
rect 11769 2142 11774 2170
rect 11802 2142 22358 2170
rect 22386 2142 22470 2170
rect 22498 2142 22503 2170
rect 23361 2142 23366 2170
rect 23394 2142 26782 2170
rect 26810 2142 26815 2170
rect 4881 2086 4886 2114
rect 4914 2086 8694 2114
rect 8722 2086 8727 2114
rect 9011 2086 9030 2114
rect 9058 2086 9063 2114
rect 9142 2086 17346 2114
rect 17425 2086 17430 2114
rect 17458 2086 17878 2114
rect 17906 2086 17911 2114
rect 18881 2086 18886 2114
rect 18914 2086 23142 2114
rect 23170 2086 23175 2114
rect 0 2058 56 2072
rect 9142 2058 9170 2086
rect 17318 2058 17346 2086
rect 28672 2058 28728 2072
rect 0 2030 4326 2058
rect 4354 2030 4359 2058
rect 6617 2030 6622 2058
rect 6650 2030 9170 2058
rect 9305 2030 9310 2058
rect 9338 2030 9478 2058
rect 9506 2030 10206 2058
rect 10234 2030 10239 2058
rect 11825 2030 11830 2058
rect 11858 2030 12558 2058
rect 12586 2030 12591 2058
rect 15073 2030 15078 2058
rect 15106 2030 17206 2058
rect 17234 2030 17239 2058
rect 17318 2030 19502 2058
rect 19530 2030 19614 2058
rect 19642 2030 19647 2058
rect 21826 2030 23310 2058
rect 23338 2030 23343 2058
rect 26105 2030 26110 2058
rect 26138 2030 26614 2058
rect 26642 2030 27902 2058
rect 27930 2030 27935 2058
rect 28065 2030 28070 2058
rect 28098 2030 28728 2058
rect 0 2016 56 2030
rect 21826 2002 21854 2030
rect 28672 2016 28728 2030
rect 2809 1974 2814 2002
rect 2842 1974 11830 2002
rect 11858 1974 11863 2002
rect 13337 1974 13342 2002
rect 13370 1974 17010 2002
rect 17089 1974 17094 2002
rect 17122 1974 21854 2002
rect 2227 1946 2232 1974
rect 2260 1946 2284 1974
rect 2312 1946 2336 1974
rect 2364 1946 2369 1974
rect 12227 1946 12232 1974
rect 12260 1946 12284 1974
rect 12312 1946 12336 1974
rect 12364 1946 12369 1974
rect 16982 1946 17010 1974
rect 22227 1946 22232 1974
rect 22260 1946 22284 1974
rect 22312 1946 22336 1974
rect 22364 1946 22369 1974
rect 4186 1918 12194 1946
rect 4186 1890 4214 1918
rect 12166 1890 12194 1918
rect 12446 1918 15974 1946
rect 16982 1918 18886 1946
rect 18914 1918 18919 1946
rect 24985 1918 24990 1946
rect 25018 1918 27678 1946
rect 27706 1918 27711 1946
rect 12446 1890 12474 1918
rect 15946 1890 15974 1918
rect 1297 1862 1302 1890
rect 1330 1862 4214 1890
rect 6169 1862 6174 1890
rect 6202 1862 7350 1890
rect 7378 1862 7383 1890
rect 7849 1862 7854 1890
rect 7882 1862 9254 1890
rect 9282 1862 9287 1890
rect 9361 1862 9366 1890
rect 9394 1862 11830 1890
rect 11858 1862 11863 1890
rect 12166 1862 12474 1890
rect 12833 1862 12838 1890
rect 12866 1862 14238 1890
rect 14266 1862 14271 1890
rect 15946 1862 24822 1890
rect 24850 1862 24855 1890
rect 25377 1862 25382 1890
rect 25410 1862 26838 1890
rect 26866 1862 26871 1890
rect 0 1834 56 1848
rect 28672 1834 28728 1848
rect 0 1806 3542 1834
rect 3570 1806 3575 1834
rect 5721 1806 5726 1834
rect 5754 1806 10710 1834
rect 10738 1806 10743 1834
rect 10934 1806 17094 1834
rect 17122 1806 17127 1834
rect 17873 1806 17878 1834
rect 17906 1806 18438 1834
rect 18466 1806 18471 1834
rect 18886 1806 22470 1834
rect 22498 1806 22503 1834
rect 26105 1806 26110 1834
rect 26138 1806 26222 1834
rect 26250 1806 27230 1834
rect 27258 1806 27263 1834
rect 27449 1806 27454 1834
rect 27482 1806 28728 1834
rect 0 1792 56 1806
rect 10934 1778 10962 1806
rect 18886 1778 18914 1806
rect 28672 1792 28728 1806
rect 1745 1750 1750 1778
rect 1778 1750 3430 1778
rect 3458 1750 3463 1778
rect 5889 1750 5894 1778
rect 5922 1750 8358 1778
rect 8386 1750 8391 1778
rect 9249 1750 9254 1778
rect 9282 1750 10962 1778
rect 11769 1750 11774 1778
rect 11802 1750 12446 1778
rect 12474 1750 12479 1778
rect 12553 1750 12558 1778
rect 12586 1750 14126 1778
rect 14154 1750 14159 1778
rect 14233 1750 14238 1778
rect 14266 1750 18914 1778
rect 20673 1750 20678 1778
rect 20706 1750 22750 1778
rect 22778 1750 22783 1778
rect 23193 1750 23198 1778
rect 23226 1750 23590 1778
rect 23618 1750 23623 1778
rect 25657 1750 25662 1778
rect 25690 1750 25774 1778
rect 25802 1750 28350 1778
rect 28378 1750 28383 1778
rect 4545 1694 4550 1722
rect 4578 1694 6734 1722
rect 6762 1694 6767 1722
rect 8414 1694 11494 1722
rect 11522 1694 11527 1722
rect 11993 1694 11998 1722
rect 12026 1694 12502 1722
rect 12530 1694 12535 1722
rect 12609 1694 12614 1722
rect 12642 1694 13454 1722
rect 13482 1694 13487 1722
rect 14065 1694 14070 1722
rect 14098 1694 15750 1722
rect 15778 1694 15783 1722
rect 15946 1694 17150 1722
rect 17178 1694 17654 1722
rect 17682 1694 17687 1722
rect 20785 1694 20790 1722
rect 20818 1694 21182 1722
rect 21210 1694 21215 1722
rect 21457 1694 21462 1722
rect 21490 1694 23478 1722
rect 23506 1694 23511 1722
rect 24425 1694 24430 1722
rect 24458 1694 24654 1722
rect 24682 1694 26222 1722
rect 26250 1694 26255 1722
rect 26777 1694 26782 1722
rect 26810 1694 28462 1722
rect 28490 1694 28495 1722
rect 8414 1666 8442 1694
rect 121 1638 126 1666
rect 154 1638 3598 1666
rect 3626 1638 3631 1666
rect 3705 1638 3710 1666
rect 3738 1638 6706 1666
rect 7177 1638 7182 1666
rect 7210 1638 8442 1666
rect 10929 1638 10934 1666
rect 10962 1638 15078 1666
rect 15106 1638 15111 1666
rect 0 1610 56 1624
rect 0 1582 378 1610
rect 0 1568 56 1582
rect 350 1498 378 1582
rect 1897 1554 1902 1582
rect 1930 1554 1954 1582
rect 1982 1554 2006 1582
rect 2034 1554 2039 1582
rect 6678 1554 6706 1638
rect 15946 1610 15974 1694
rect 18489 1638 18494 1666
rect 18522 1638 19334 1666
rect 19362 1638 19367 1666
rect 21826 1638 22554 1666
rect 22633 1638 22638 1666
rect 22666 1638 23870 1666
rect 23898 1638 23903 1666
rect 24313 1638 24318 1666
rect 24346 1638 24766 1666
rect 24794 1638 24799 1666
rect 21826 1610 21854 1638
rect 7457 1582 7462 1610
rect 7490 1582 7686 1610
rect 7714 1582 7719 1610
rect 7961 1582 7966 1610
rect 7994 1582 9814 1610
rect 9842 1582 9847 1610
rect 9921 1582 9926 1610
rect 9954 1582 11830 1610
rect 11858 1582 11863 1610
rect 12105 1582 12110 1610
rect 12138 1582 12278 1610
rect 12306 1582 12311 1610
rect 13006 1582 15974 1610
rect 19049 1582 19054 1610
rect 19082 1582 21854 1610
rect 22526 1610 22554 1638
rect 28672 1610 28728 1624
rect 22526 1582 26558 1610
rect 26586 1582 26591 1610
rect 27281 1582 27286 1610
rect 27314 1582 28728 1610
rect 11897 1554 11902 1582
rect 11930 1554 11954 1582
rect 11982 1554 12006 1582
rect 12034 1554 12039 1582
rect 3537 1526 3542 1554
rect 3570 1526 6566 1554
rect 6594 1526 6599 1554
rect 6678 1526 10262 1554
rect 10290 1526 10295 1554
rect 13006 1498 13034 1582
rect 21897 1554 21902 1582
rect 21930 1554 21954 1582
rect 21982 1554 22006 1582
rect 22034 1554 22039 1582
rect 28672 1568 28728 1582
rect 15801 1526 15806 1554
rect 15834 1526 18830 1554
rect 18858 1526 18863 1554
rect 350 1470 3654 1498
rect 3682 1470 3687 1498
rect 5945 1470 5950 1498
rect 5978 1470 7574 1498
rect 7602 1470 7607 1498
rect 7681 1470 7686 1498
rect 7714 1470 8918 1498
rect 8946 1470 8951 1498
rect 9249 1470 9254 1498
rect 9282 1470 13034 1498
rect 14009 1470 14014 1498
rect 14042 1470 15974 1498
rect 22017 1470 22022 1498
rect 22050 1470 22190 1498
rect 22218 1470 22223 1498
rect 15946 1442 15974 1470
rect 3705 1414 3710 1442
rect 3738 1414 8470 1442
rect 8498 1414 8503 1442
rect 8577 1414 8582 1442
rect 8610 1414 11382 1442
rect 11410 1414 11415 1442
rect 11489 1414 11494 1442
rect 11522 1414 15246 1442
rect 15274 1414 15279 1442
rect 15946 1414 23646 1442
rect 23674 1414 23679 1442
rect 26497 1414 26502 1442
rect 26530 1414 28518 1442
rect 28546 1414 28551 1442
rect 0 1386 56 1400
rect 28672 1386 28728 1400
rect 0 1358 518 1386
rect 546 1358 551 1386
rect 6729 1358 6734 1386
rect 6762 1358 9926 1386
rect 9954 1358 9959 1386
rect 10705 1358 10710 1386
rect 10738 1358 13062 1386
rect 13090 1358 13095 1386
rect 13393 1358 13398 1386
rect 13426 1358 17738 1386
rect 17817 1358 17822 1386
rect 17850 1358 18158 1386
rect 18186 1358 18191 1386
rect 18489 1358 18494 1386
rect 18522 1358 22470 1386
rect 22498 1358 22503 1386
rect 24369 1358 24374 1386
rect 24402 1358 26782 1386
rect 26810 1358 26815 1386
rect 28065 1358 28070 1386
rect 28098 1358 28728 1386
rect 0 1344 56 1358
rect 17710 1330 17738 1358
rect 28672 1344 28728 1358
rect 793 1302 798 1330
rect 826 1302 8526 1330
rect 8554 1302 8559 1330
rect 9585 1302 9590 1330
rect 9618 1302 12614 1330
rect 12642 1302 12647 1330
rect 16529 1302 16534 1330
rect 16562 1302 17038 1330
rect 17066 1302 17071 1330
rect 17710 1302 22862 1330
rect 22890 1302 22895 1330
rect 4186 1246 12446 1274
rect 12474 1246 12479 1274
rect 21065 1246 21070 1274
rect 21098 1246 25326 1274
rect 25354 1246 25438 1274
rect 25466 1246 25471 1274
rect 4153 1190 4158 1218
rect 4186 1190 4214 1246
rect 7513 1190 7518 1218
rect 7546 1190 7686 1218
rect 7714 1190 7719 1218
rect 11097 1190 11102 1218
rect 11130 1190 12110 1218
rect 12138 1190 12143 1218
rect 12497 1190 12502 1218
rect 12530 1190 18494 1218
rect 18522 1190 18527 1218
rect 19889 1190 19894 1218
rect 19922 1190 21350 1218
rect 21378 1190 21518 1218
rect 21546 1190 21551 1218
rect 0 1162 56 1176
rect 2227 1162 2232 1190
rect 2260 1162 2284 1190
rect 2312 1162 2336 1190
rect 2364 1162 2369 1190
rect 12227 1162 12232 1190
rect 12260 1162 12284 1190
rect 12312 1162 12336 1190
rect 12364 1162 12369 1190
rect 22227 1162 22232 1190
rect 22260 1162 22284 1190
rect 22312 1162 22336 1190
rect 22364 1162 22369 1190
rect 28672 1162 28728 1176
rect 0 1134 2114 1162
rect 6449 1134 6454 1162
rect 6482 1134 9506 1162
rect 9865 1134 9870 1162
rect 9898 1134 12194 1162
rect 0 1120 56 1134
rect 2086 1106 2114 1134
rect 9478 1106 9506 1134
rect 12166 1106 12194 1134
rect 12446 1134 21854 1162
rect 27449 1134 27454 1162
rect 27482 1134 28728 1162
rect 12446 1106 12474 1134
rect 21826 1106 21854 1134
rect 28672 1120 28728 1134
rect 2086 1078 9366 1106
rect 9394 1078 9399 1106
rect 9478 1078 11774 1106
rect 12166 1078 12474 1106
rect 12553 1078 12558 1106
rect 12586 1078 14014 1106
rect 14042 1078 14047 1106
rect 15073 1078 15078 1106
rect 15106 1078 18298 1106
rect 18489 1078 18494 1106
rect 18522 1078 19054 1106
rect 19082 1078 19087 1106
rect 21826 1078 25998 1106
rect 26026 1078 26031 1106
rect 849 1022 854 1050
rect 882 1022 3598 1050
rect 3626 1022 3631 1050
rect 3929 1022 3934 1050
rect 3962 1022 8246 1050
rect 8274 1022 8279 1050
rect 11746 994 11774 1078
rect 18270 1050 18298 1078
rect 11825 1022 11830 1050
rect 11858 1022 13790 1050
rect 13818 1022 13823 1050
rect 14625 1022 14630 1050
rect 14658 1022 16198 1050
rect 16226 1022 16231 1050
rect 17593 1022 17598 1050
rect 17626 1022 17878 1050
rect 17906 1022 17911 1050
rect 18270 1022 24066 1050
rect 25713 1022 25718 1050
rect 25746 1022 27062 1050
rect 27090 1022 27095 1050
rect 24038 994 24066 1022
rect 3369 966 3374 994
rect 3402 966 4214 994
rect 7121 966 7126 994
rect 7154 966 10598 994
rect 10626 966 10631 994
rect 11746 966 13398 994
rect 13426 966 13431 994
rect 13505 966 13510 994
rect 13538 966 13543 994
rect 14737 966 14742 994
rect 14770 966 15582 994
rect 15610 966 15615 994
rect 18377 966 18382 994
rect 18410 966 19614 994
rect 19642 966 19647 994
rect 21177 966 21182 994
rect 21210 966 22750 994
rect 22778 966 22783 994
rect 24038 966 26278 994
rect 26306 966 26311 994
rect 26390 966 27398 994
rect 27426 966 27431 994
rect 0 938 56 952
rect 0 910 1078 938
rect 1106 910 1111 938
rect 0 896 56 910
rect 4186 882 4214 966
rect 13510 938 13538 966
rect 26390 938 26418 966
rect 28672 938 28728 952
rect 4993 910 4998 938
rect 5026 910 13342 938
rect 13370 910 13375 938
rect 13510 910 21686 938
rect 21714 910 21719 938
rect 21793 910 21798 938
rect 21826 910 22022 938
rect 22050 910 22055 938
rect 23641 910 23646 938
rect 23674 910 26418 938
rect 26777 910 26782 938
rect 26810 910 28728 938
rect 28672 896 28728 910
rect 1694 854 3766 882
rect 3794 854 3799 882
rect 4186 854 8274 882
rect 8409 854 8414 882
rect 8442 854 9422 882
rect 9450 854 9590 882
rect 9618 854 9623 882
rect 10873 854 10878 882
rect 10906 854 11550 882
rect 11578 854 11583 882
rect 11830 854 12558 882
rect 12586 854 12591 882
rect 13174 854 14798 882
rect 14826 854 14831 882
rect 15577 854 15582 882
rect 15610 854 16478 882
rect 16506 854 16511 882
rect 17593 854 17598 882
rect 17626 854 18550 882
rect 18578 854 18583 882
rect 19609 854 19614 882
rect 19642 854 21014 882
rect 21042 854 21047 882
rect 21826 854 21966 882
rect 21994 854 21999 882
rect 22969 854 22974 882
rect 23002 854 23926 882
rect 23954 854 23959 882
rect 25993 854 25998 882
rect 26026 854 27006 882
rect 27034 854 27039 882
rect 1694 826 1722 854
rect 8246 826 8274 854
rect 11830 826 11858 854
rect 569 798 574 826
rect 602 798 1722 826
rect 2585 798 2590 826
rect 2618 798 4606 826
rect 4634 798 4639 826
rect 4825 798 4830 826
rect 4858 798 5222 826
rect 5250 798 5255 826
rect 7065 798 7070 826
rect 7098 798 8134 826
rect 8162 798 8167 826
rect 8246 798 9254 826
rect 9282 798 9287 826
rect 9921 798 9926 826
rect 9954 798 11858 826
rect 1897 770 1902 798
rect 1930 770 1954 798
rect 1982 770 2006 798
rect 2034 770 2039 798
rect 11897 770 11902 798
rect 11930 770 11954 798
rect 11982 770 12006 798
rect 12034 770 12039 798
rect 2137 742 2142 770
rect 2170 742 3990 770
rect 4018 742 4023 770
rect 4377 742 4382 770
rect 4410 742 6678 770
rect 6706 742 6711 770
rect 7569 742 7574 770
rect 7602 742 9758 770
rect 9786 742 9791 770
rect 0 714 56 728
rect 13174 714 13202 854
rect 21826 826 21854 854
rect 15465 798 15470 826
rect 15498 798 15638 826
rect 15666 798 15671 826
rect 15750 798 17654 826
rect 17682 798 17687 826
rect 18769 798 18774 826
rect 18802 798 19726 826
rect 19754 798 19759 826
rect 19833 798 19838 826
rect 19866 798 20286 826
rect 20314 798 20319 826
rect 20505 798 20510 826
rect 20538 798 21854 826
rect 24257 798 24262 826
rect 24290 798 24990 826
rect 25018 798 25023 826
rect 15750 770 15778 798
rect 21897 770 21902 798
rect 21930 770 21954 798
rect 21982 770 22006 798
rect 22034 770 22039 798
rect 13281 742 13286 770
rect 13314 742 15778 770
rect 15857 742 15862 770
rect 15890 742 16646 770
rect 16674 742 16679 770
rect 16753 742 16758 770
rect 16786 742 19894 770
rect 19922 742 19927 770
rect 20953 742 20958 770
rect 20986 742 21574 770
rect 21602 742 21607 770
rect 22073 742 22078 770
rect 22106 742 23030 770
rect 23058 742 23063 770
rect 25041 742 25046 770
rect 25074 742 25438 770
rect 25466 742 25471 770
rect 28672 714 28728 728
rect 0 686 2926 714
rect 2954 686 2959 714
rect 3817 686 3822 714
rect 3850 686 4214 714
rect 6393 686 6398 714
rect 6426 686 9534 714
rect 9562 686 9567 714
rect 10593 686 10598 714
rect 10626 686 13202 714
rect 14121 686 14126 714
rect 14154 686 18886 714
rect 18914 686 18919 714
rect 21625 686 21630 714
rect 21658 686 22414 714
rect 22442 686 22447 714
rect 24201 686 24206 714
rect 24234 686 26110 714
rect 26138 686 26143 714
rect 26777 686 26782 714
rect 26810 686 28728 714
rect 0 672 56 686
rect 4186 658 4214 686
rect 28672 672 28728 686
rect 4186 630 7658 658
rect 7737 630 7742 658
rect 7770 630 12670 658
rect 12698 630 12703 658
rect 12889 630 12894 658
rect 12922 630 13230 658
rect 13258 630 13263 658
rect 13449 630 13454 658
rect 13482 630 13790 658
rect 13818 630 13823 658
rect 15801 630 15806 658
rect 15834 630 16310 658
rect 16338 630 16343 658
rect 16641 630 16646 658
rect 16674 630 17402 658
rect 17481 630 17486 658
rect 17514 630 24150 658
rect 24178 630 24183 658
rect 7630 602 7658 630
rect 17374 602 17402 630
rect 6393 574 6398 602
rect 6426 574 7518 602
rect 7546 574 7551 602
rect 7630 574 8022 602
rect 8050 574 8055 602
rect 8913 574 8918 602
rect 8946 574 11046 602
rect 11074 574 11079 602
rect 11769 574 11774 602
rect 11802 574 12726 602
rect 12754 574 12759 602
rect 12833 574 12838 602
rect 12866 574 16534 602
rect 16562 574 16567 602
rect 17374 574 18774 602
rect 18802 574 18807 602
rect 18881 574 18886 602
rect 18914 574 22246 602
rect 22274 574 22279 602
rect 23417 574 23422 602
rect 23450 574 24710 602
rect 24738 574 24743 602
rect 6841 518 6846 546
rect 6874 518 11214 546
rect 11242 518 11247 546
rect 11433 518 11438 546
rect 11466 518 12446 546
rect 12474 518 12479 546
rect 12553 518 12558 546
rect 12586 518 13118 546
rect 13146 518 13151 546
rect 13337 518 13342 546
rect 13370 518 13622 546
rect 13650 518 13655 546
rect 13734 518 17486 546
rect 17514 518 17519 546
rect 18265 518 18270 546
rect 18298 518 19782 546
rect 19810 518 19815 546
rect 20281 518 20286 546
rect 20314 518 21686 546
rect 21714 518 21719 546
rect 21849 518 21854 546
rect 21882 518 27566 546
rect 27594 518 27599 546
rect 0 490 56 504
rect 13734 490 13762 518
rect 28672 490 28728 504
rect 0 462 294 490
rect 322 462 327 490
rect 457 462 462 490
rect 490 462 8358 490
rect 8386 462 8391 490
rect 8465 462 8470 490
rect 8498 462 13762 490
rect 14681 462 14686 490
rect 14714 462 15078 490
rect 15106 462 15111 490
rect 16697 462 16702 490
rect 16730 462 17934 490
rect 17962 462 17967 490
rect 18713 462 18718 490
rect 18746 462 18751 490
rect 20057 462 20062 490
rect 20090 462 20622 490
rect 20650 462 20655 490
rect 20958 462 22526 490
rect 22554 462 22559 490
rect 22913 462 22918 490
rect 22946 462 24542 490
rect 24570 462 24575 490
rect 25993 462 25998 490
rect 26026 462 28728 490
rect 0 448 56 462
rect 18718 434 18746 462
rect 20958 434 20986 462
rect 28672 448 28728 462
rect 5497 406 5502 434
rect 5530 406 9086 434
rect 9114 406 9119 434
rect 14905 406 14910 434
rect 14938 406 16030 434
rect 16058 406 16063 434
rect 16249 406 16254 434
rect 16282 406 17094 434
rect 17122 406 17127 434
rect 17369 406 17374 434
rect 17402 406 18746 434
rect 18830 406 20090 434
rect 20953 406 20958 434
rect 20986 406 20991 434
rect 21401 406 21406 434
rect 21434 406 22134 434
rect 22162 406 22167 434
rect 22745 406 22750 434
rect 22778 406 24374 434
rect 24402 406 24407 434
rect 2227 378 2232 406
rect 2260 378 2284 406
rect 2312 378 2336 406
rect 2364 378 2369 406
rect 12227 378 12232 406
rect 12260 378 12284 406
rect 12312 378 12336 406
rect 12364 378 12369 406
rect 6953 350 6958 378
rect 6986 350 9310 378
rect 9338 350 9343 378
rect 12609 350 12614 378
rect 12642 350 15806 378
rect 15834 350 15839 378
rect 15913 350 15918 378
rect 15946 350 16842 378
rect 16921 350 16926 378
rect 16954 350 17878 378
rect 17906 350 17911 378
rect 16814 322 16842 350
rect 2361 294 2366 322
rect 2394 294 3542 322
rect 3570 294 3575 322
rect 5049 294 5054 322
rect 5082 294 7014 322
rect 7042 294 7047 322
rect 7289 294 7294 322
rect 7322 294 8638 322
rect 8666 294 8671 322
rect 9025 294 9030 322
rect 9058 294 16702 322
rect 16730 294 16735 322
rect 16814 294 18718 322
rect 18746 294 18751 322
rect 0 266 56 280
rect 18830 266 18858 406
rect 20062 378 20090 406
rect 22227 378 22232 406
rect 22260 378 22284 406
rect 22312 378 22336 406
rect 22364 378 22369 406
rect 19161 350 19166 378
rect 19194 350 19950 378
rect 19978 350 19983 378
rect 20062 350 21798 378
rect 21826 350 21831 378
rect 19385 294 19390 322
rect 19418 294 20230 322
rect 20258 294 20263 322
rect 22297 294 22302 322
rect 22330 294 22806 322
rect 22834 294 22839 322
rect 28672 266 28728 280
rect 0 238 7126 266
rect 7154 238 7159 266
rect 7238 238 9646 266
rect 9674 238 9679 266
rect 13449 238 13454 266
rect 13482 238 15918 266
rect 15946 238 15951 266
rect 16417 238 16422 266
rect 16450 238 18858 266
rect 18937 238 18942 266
rect 18970 238 20454 266
rect 20482 238 20487 266
rect 21849 238 21854 266
rect 21882 238 23646 266
rect 23674 238 23679 266
rect 28457 238 28462 266
rect 28490 238 28728 266
rect 0 224 56 238
rect 7238 210 7266 238
rect 28672 224 28728 238
rect 5497 182 5502 210
rect 5530 182 7266 210
rect 8689 182 8694 210
rect 8722 182 14406 210
rect 14434 182 14439 210
rect 15353 182 15358 210
rect 15386 182 16814 210
rect 16842 182 16847 210
rect 17817 182 17822 210
rect 17850 182 18662 210
rect 18690 182 18695 210
rect 18769 182 18774 210
rect 18802 182 21070 210
rect 21098 182 21103 210
rect 22521 182 22526 210
rect 22554 182 24430 210
rect 24458 182 24463 210
rect 3425 126 3430 154
rect 3458 126 8414 154
rect 8442 126 8447 154
rect 8521 126 8526 154
rect 8554 126 15470 154
rect 15498 126 15503 154
rect 16697 126 16702 154
rect 16730 126 23366 154
rect 23394 126 23399 154
rect 23641 126 23646 154
rect 23674 126 25270 154
rect 25298 126 25303 154
rect 1129 70 1134 98
rect 1162 70 8190 98
rect 8218 70 8223 98
rect 11209 70 11214 98
rect 11242 70 15694 98
rect 15722 70 15727 98
rect 19721 70 19726 98
rect 19754 70 21854 98
rect 22073 70 22078 98
rect 22106 70 23086 98
rect 23114 70 23119 98
rect 25097 70 25102 98
rect 25130 70 25214 98
rect 25242 70 25247 98
rect 25881 70 25886 98
rect 25914 70 25919 98
rect 0 42 56 56
rect 21826 42 21854 70
rect 25886 42 25914 70
rect 28672 42 28728 56
rect 0 14 462 42
rect 490 14 495 42
rect 21826 14 25914 42
rect 28513 14 28518 42
rect 28546 14 28728 42
rect 0 0 56 14
rect 28672 0 28728 14
<< via3 >>
rect 2232 6650 2260 6678
rect 2284 6650 2312 6678
rect 2336 6650 2364 6678
rect 12232 6650 12260 6678
rect 12284 6650 12312 6678
rect 12336 6650 12364 6678
rect 22232 6650 22260 6678
rect 22284 6650 22312 6678
rect 22336 6650 22364 6678
rect 1902 6258 1930 6286
rect 1954 6258 1982 6286
rect 2006 6258 2034 6286
rect 11902 6258 11930 6286
rect 11954 6258 11982 6286
rect 12006 6258 12034 6286
rect 21902 6258 21930 6286
rect 21954 6258 21982 6286
rect 22006 6258 22034 6286
rect 12446 6230 12474 6258
rect 12446 6118 12474 6146
rect 8022 6006 8050 6034
rect 2232 5866 2260 5894
rect 2284 5866 2312 5894
rect 2336 5866 2364 5894
rect 12232 5866 12260 5894
rect 12284 5866 12312 5894
rect 12336 5866 12364 5894
rect 22232 5866 22260 5894
rect 22284 5866 22312 5894
rect 22336 5866 22364 5894
rect 11158 5726 11186 5754
rect 8358 5558 8386 5586
rect 9926 5558 9954 5586
rect 1902 5474 1930 5502
rect 1954 5474 1982 5502
rect 2006 5474 2034 5502
rect 11902 5474 11930 5502
rect 11954 5474 11982 5502
rect 12006 5474 12034 5502
rect 21902 5474 21930 5502
rect 21954 5474 21982 5502
rect 22006 5474 22034 5502
rect 9926 5334 9954 5362
rect 11158 5222 11186 5250
rect 7686 5110 7714 5138
rect 2232 5082 2260 5110
rect 2284 5082 2312 5110
rect 2336 5082 2364 5110
rect 12232 5082 12260 5110
rect 12284 5082 12312 5110
rect 12336 5082 12364 5110
rect 22232 5082 22260 5110
rect 22284 5082 22312 5110
rect 22336 5082 22364 5110
rect 13398 4942 13426 4970
rect 13734 4886 13762 4914
rect 7686 4830 7714 4858
rect 1902 4690 1930 4718
rect 1954 4690 1982 4718
rect 2006 4690 2034 4718
rect 13398 4718 13426 4746
rect 11902 4690 11930 4718
rect 11954 4690 11982 4718
rect 12006 4690 12034 4718
rect 21902 4690 21930 4718
rect 21954 4690 21982 4718
rect 22006 4690 22034 4718
rect 13734 4382 13762 4410
rect 13846 4382 13874 4410
rect 2232 4298 2260 4326
rect 2284 4298 2312 4326
rect 2336 4298 2364 4326
rect 12232 4298 12260 4326
rect 12284 4298 12312 4326
rect 12336 4298 12364 4326
rect 22232 4298 22260 4326
rect 22284 4298 22312 4326
rect 22336 4298 22364 4326
rect 8358 4214 8386 4242
rect 13846 4214 13874 4242
rect 14014 4214 14042 4242
rect 1902 3906 1930 3934
rect 1954 3906 1982 3934
rect 2006 3906 2034 3934
rect 11902 3906 11930 3934
rect 11954 3906 11982 3934
rect 12006 3906 12034 3934
rect 21902 3906 21930 3934
rect 21954 3906 21982 3934
rect 22006 3906 22034 3934
rect 7630 3542 7658 3570
rect 12558 3542 12586 3570
rect 13174 3542 13202 3570
rect 2232 3514 2260 3542
rect 2284 3514 2312 3542
rect 2336 3514 2364 3542
rect 12232 3514 12260 3542
rect 12284 3514 12312 3542
rect 12336 3514 12364 3542
rect 22232 3514 22260 3542
rect 22284 3514 22312 3542
rect 22336 3514 22364 3542
rect 13230 3430 13258 3458
rect 7574 3318 7602 3346
rect 10934 3206 10962 3234
rect 182 3150 210 3178
rect 7574 3150 7602 3178
rect 1902 3122 1930 3150
rect 1954 3122 1982 3150
rect 2006 3122 2034 3150
rect 11902 3122 11930 3150
rect 11954 3122 11982 3150
rect 12006 3122 12034 3150
rect 21902 3122 21930 3150
rect 21954 3122 21982 3150
rect 22006 3122 22034 3150
rect 10934 3094 10962 3122
rect 8358 2982 8386 3010
rect 2232 2730 2260 2758
rect 2284 2730 2312 2758
rect 2336 2730 2364 2758
rect 12232 2730 12260 2758
rect 12284 2730 12312 2758
rect 12336 2730 12364 2758
rect 22232 2730 22260 2758
rect 22284 2730 22312 2758
rect 22336 2730 22364 2758
rect 182 2646 210 2674
rect 7574 2534 7602 2562
rect 11102 2422 11130 2450
rect 1902 2338 1930 2366
rect 1954 2338 1982 2366
rect 2006 2338 2034 2366
rect 11902 2338 11930 2366
rect 11954 2338 11982 2366
rect 12006 2338 12034 2366
rect 18550 2366 18578 2394
rect 21902 2338 21930 2366
rect 21954 2338 21982 2366
rect 22006 2338 22034 2366
rect 18830 2310 18858 2338
rect 4886 2254 4914 2282
rect 8358 2254 8386 2282
rect 3598 2198 3626 2226
rect 7630 2198 7658 2226
rect 9366 2198 9394 2226
rect 11102 2198 11130 2226
rect 17206 2198 17234 2226
rect 11662 2142 11690 2170
rect 4886 2086 4914 2114
rect 9030 2086 9058 2114
rect 11830 2030 11858 2058
rect 12558 2030 12586 2058
rect 17206 2030 17234 2058
rect 2232 1946 2260 1974
rect 2284 1946 2312 1974
rect 2336 1946 2364 1974
rect 12232 1946 12260 1974
rect 12284 1946 12312 1974
rect 12336 1946 12364 1974
rect 22232 1946 22260 1974
rect 22284 1946 22312 1974
rect 22336 1946 22364 1974
rect 9366 1862 9394 1890
rect 11830 1862 11858 1890
rect 14238 1862 14266 1890
rect 8358 1750 8386 1778
rect 11774 1750 11802 1778
rect 12446 1750 12474 1778
rect 14238 1750 14266 1778
rect 12614 1694 12642 1722
rect 13454 1694 13482 1722
rect 3598 1638 3626 1666
rect 1902 1554 1930 1582
rect 1954 1554 1982 1582
rect 2006 1554 2034 1582
rect 7686 1582 7714 1610
rect 9926 1582 9954 1610
rect 11902 1554 11930 1582
rect 11954 1554 11982 1582
rect 12006 1554 12034 1582
rect 21902 1554 21930 1582
rect 21954 1554 21982 1582
rect 22006 1554 22034 1582
rect 7574 1470 7602 1498
rect 7686 1470 7714 1498
rect 9926 1358 9954 1386
rect 2232 1162 2260 1190
rect 2284 1162 2312 1190
rect 2336 1162 2364 1190
rect 12232 1162 12260 1190
rect 12284 1162 12312 1190
rect 12336 1162 12364 1190
rect 22232 1162 22260 1190
rect 22284 1162 22312 1190
rect 22336 1162 22364 1190
rect 12558 1078 12586 1106
rect 14014 1078 14042 1106
rect 21798 910 21826 938
rect 12558 854 12586 882
rect 1902 770 1930 798
rect 1954 770 1982 798
rect 2006 770 2034 798
rect 11902 770 11930 798
rect 11954 770 11982 798
rect 12006 770 12034 798
rect 18774 798 18802 826
rect 21902 770 21930 798
rect 21954 770 21982 798
rect 22006 770 22034 798
rect 15862 742 15890 770
rect 18886 686 18914 714
rect 8022 574 8050 602
rect 18774 574 18802 602
rect 18886 574 18914 602
rect 8470 462 8498 490
rect 2232 378 2260 406
rect 2284 378 2312 406
rect 2336 378 2364 406
rect 12232 378 12260 406
rect 12284 378 12312 406
rect 12336 378 12364 406
rect 15806 350 15834 378
rect 15918 350 15946 378
rect 9030 294 9058 322
rect 16702 294 16730 322
rect 18718 294 18746 322
rect 22232 378 22260 406
rect 22284 378 22312 406
rect 22336 378 22364 406
rect 21798 350 21826 378
rect 13454 238 13482 266
rect 15918 238 15946 266
rect 18774 182 18802 210
rect 16702 126 16730 154
<< metal4 >>
rect 1888 6286 2048 7112
rect 1888 6258 1902 6286
rect 1930 6258 1954 6286
rect 1982 6258 2006 6286
rect 2034 6258 2048 6286
rect 1888 5502 2048 6258
rect 1888 5474 1902 5502
rect 1930 5474 1954 5502
rect 1982 5474 2006 5502
rect 2034 5474 2048 5502
rect 1888 4718 2048 5474
rect 1888 4690 1902 4718
rect 1930 4690 1954 4718
rect 1982 4690 2006 4718
rect 2034 4690 2048 4718
rect 1888 3934 2048 4690
rect 1888 3906 1902 3934
rect 1930 3906 1954 3934
rect 1982 3906 2006 3934
rect 2034 3906 2048 3934
rect 182 3178 210 3183
rect 182 2674 210 3150
rect 182 2641 210 2646
rect 1888 3150 2048 3906
rect 1888 3122 1902 3150
rect 1930 3122 1954 3150
rect 1982 3122 2006 3150
rect 2034 3122 2048 3150
rect 1888 2366 2048 3122
rect 1888 2338 1902 2366
rect 1930 2338 1954 2366
rect 1982 2338 2006 2366
rect 2034 2338 2048 2366
rect 1888 1582 2048 2338
rect 1888 1554 1902 1582
rect 1930 1554 1954 1582
rect 1982 1554 2006 1582
rect 2034 1554 2048 1582
rect 1888 798 2048 1554
rect 1888 770 1902 798
rect 1930 770 1954 798
rect 1982 770 2006 798
rect 2034 770 2048 798
rect 1888 0 2048 770
rect 2218 6678 2378 7112
rect 2218 6650 2232 6678
rect 2260 6650 2284 6678
rect 2312 6650 2336 6678
rect 2364 6650 2378 6678
rect 2218 5894 2378 6650
rect 11888 6286 12048 7112
rect 11888 6258 11902 6286
rect 11930 6258 11954 6286
rect 11982 6258 12006 6286
rect 12034 6258 12048 6286
rect 2218 5866 2232 5894
rect 2260 5866 2284 5894
rect 2312 5866 2336 5894
rect 2364 5866 2378 5894
rect 2218 5110 2378 5866
rect 8022 6034 8050 6039
rect 2218 5082 2232 5110
rect 2260 5082 2284 5110
rect 2312 5082 2336 5110
rect 2364 5082 2378 5110
rect 2218 4326 2378 5082
rect 7686 5138 7714 5143
rect 7686 4858 7714 5110
rect 7686 4825 7714 4830
rect 2218 4298 2232 4326
rect 2260 4298 2284 4326
rect 2312 4298 2336 4326
rect 2364 4298 2378 4326
rect 2218 3542 2378 4298
rect 2218 3514 2232 3542
rect 2260 3514 2284 3542
rect 2312 3514 2336 3542
rect 2364 3514 2378 3542
rect 2218 2758 2378 3514
rect 7630 3570 7658 3575
rect 7574 3346 7602 3351
rect 7574 3178 7602 3318
rect 7574 3145 7602 3150
rect 2218 2730 2232 2758
rect 2260 2730 2284 2758
rect 2312 2730 2336 2758
rect 2364 2730 2378 2758
rect 2218 1974 2378 2730
rect 7574 2562 7602 2567
rect 4886 2282 4914 2287
rect 2218 1946 2232 1974
rect 2260 1946 2284 1974
rect 2312 1946 2336 1974
rect 2364 1946 2378 1974
rect 2218 1190 2378 1946
rect 3598 2226 3626 2231
rect 3598 1666 3626 2198
rect 4886 2114 4914 2254
rect 4886 2081 4914 2086
rect 3598 1633 3626 1638
rect 7574 1498 7602 2534
rect 7630 2226 7658 3542
rect 7630 2193 7658 2198
rect 7574 1465 7602 1470
rect 7686 1610 7714 1615
rect 7686 1498 7714 1582
rect 7686 1465 7714 1470
rect 2218 1162 2232 1190
rect 2260 1162 2284 1190
rect 2312 1162 2336 1190
rect 2364 1162 2378 1190
rect 2218 406 2378 1162
rect 8022 602 8050 6006
rect 11158 5754 11186 5759
rect 8358 5586 8386 5591
rect 8358 4242 8386 5558
rect 9926 5586 9954 5591
rect 9926 5362 9954 5558
rect 9926 5329 9954 5334
rect 11158 5250 11186 5726
rect 11158 5217 11186 5222
rect 11888 5502 12048 6258
rect 11888 5474 11902 5502
rect 11930 5474 11954 5502
rect 11982 5474 12006 5502
rect 12034 5474 12048 5502
rect 8358 4209 8386 4214
rect 11888 4718 12048 5474
rect 11888 4690 11902 4718
rect 11930 4690 11954 4718
rect 11982 4690 12006 4718
rect 12034 4690 12048 4718
rect 11888 3934 12048 4690
rect 11888 3906 11902 3934
rect 11930 3906 11954 3934
rect 11982 3906 12006 3934
rect 12034 3906 12048 3934
rect 10934 3234 10962 3239
rect 10934 3122 10962 3206
rect 10934 3089 10962 3094
rect 11888 3150 12048 3906
rect 11888 3122 11902 3150
rect 11930 3122 11954 3150
rect 11982 3122 12006 3150
rect 12034 3122 12048 3150
rect 8358 3010 8386 3015
rect 8358 2282 8386 2982
rect 8358 2249 8386 2254
rect 11102 2450 11130 2455
rect 9366 2226 9394 2231
rect 9030 2114 9058 2119
rect 8022 569 8050 574
rect 8358 1778 8386 1783
rect 8358 509 8386 1750
rect 8358 490 8498 509
rect 8358 481 8470 490
rect 8470 457 8498 462
rect 2218 378 2232 406
rect 2260 378 2284 406
rect 2312 378 2336 406
rect 2364 378 2378 406
rect 2218 0 2378 378
rect 9030 322 9058 2086
rect 9366 1890 9394 2198
rect 11102 2226 11130 2422
rect 11102 2193 11130 2198
rect 11888 2366 12048 3122
rect 11888 2338 11902 2366
rect 11930 2338 11954 2366
rect 11982 2338 12006 2366
rect 12034 2338 12048 2366
rect 11662 2170 11690 2175
rect 11662 2129 11690 2142
rect 11662 2101 11802 2129
rect 9366 1857 9394 1862
rect 11774 1778 11802 2101
rect 11830 2058 11858 2063
rect 11830 1890 11858 2030
rect 11830 1857 11858 1862
rect 11774 1745 11802 1750
rect 9926 1610 9954 1615
rect 9926 1386 9954 1582
rect 9926 1353 9954 1358
rect 11888 1582 12048 2338
rect 11888 1554 11902 1582
rect 11930 1554 11954 1582
rect 11982 1554 12006 1582
rect 12034 1554 12048 1582
rect 9030 289 9058 294
rect 11888 798 12048 1554
rect 11888 770 11902 798
rect 11930 770 11954 798
rect 11982 770 12006 798
rect 12034 770 12048 798
rect 11888 0 12048 770
rect 12218 6678 12378 7112
rect 12218 6650 12232 6678
rect 12260 6650 12284 6678
rect 12312 6650 12336 6678
rect 12364 6650 12378 6678
rect 12218 5894 12378 6650
rect 21888 6286 22048 7112
rect 12446 6258 12474 6263
rect 12446 6146 12474 6230
rect 12446 6113 12474 6118
rect 21888 6258 21902 6286
rect 21930 6258 21954 6286
rect 21982 6258 22006 6286
rect 22034 6258 22048 6286
rect 12218 5866 12232 5894
rect 12260 5866 12284 5894
rect 12312 5866 12336 5894
rect 12364 5866 12378 5894
rect 12218 5110 12378 5866
rect 12218 5082 12232 5110
rect 12260 5082 12284 5110
rect 12312 5082 12336 5110
rect 12364 5082 12378 5110
rect 12218 4326 12378 5082
rect 21888 5502 22048 6258
rect 21888 5474 21902 5502
rect 21930 5474 21954 5502
rect 21982 5474 22006 5502
rect 22034 5474 22048 5502
rect 13398 4970 13426 4975
rect 13398 4746 13426 4942
rect 13398 4713 13426 4718
rect 13734 4914 13762 4919
rect 13734 4410 13762 4886
rect 21888 4718 22048 5474
rect 21888 4690 21902 4718
rect 21930 4690 21954 4718
rect 21982 4690 22006 4718
rect 22034 4690 22048 4718
rect 13734 4377 13762 4382
rect 13846 4410 13874 4415
rect 12218 4298 12232 4326
rect 12260 4298 12284 4326
rect 12312 4298 12336 4326
rect 12364 4298 12378 4326
rect 12218 3542 12378 4298
rect 13846 4242 13874 4382
rect 13846 4209 13874 4214
rect 14014 4242 14042 4247
rect 12218 3514 12232 3542
rect 12260 3514 12284 3542
rect 12312 3514 12336 3542
rect 12364 3514 12378 3542
rect 12218 2758 12378 3514
rect 12218 2730 12232 2758
rect 12260 2730 12284 2758
rect 12312 2730 12336 2758
rect 12364 2730 12378 2758
rect 12218 1974 12378 2730
rect 12558 3570 12586 3575
rect 12558 2058 12586 3542
rect 13174 3570 13202 3575
rect 13202 3542 13258 3569
rect 13174 3541 13258 3542
rect 13174 3537 13202 3541
rect 13230 3458 13258 3541
rect 13230 3425 13258 3430
rect 12558 2025 12586 2030
rect 12218 1946 12232 1974
rect 12260 1946 12284 1974
rect 12312 1946 12336 1974
rect 12364 1946 12378 1974
rect 12218 1190 12378 1946
rect 12446 1778 12474 1783
rect 12474 1750 12642 1769
rect 12446 1741 12642 1750
rect 12614 1722 12642 1741
rect 12614 1689 12642 1694
rect 13454 1722 13482 1727
rect 12218 1162 12232 1190
rect 12260 1162 12284 1190
rect 12312 1162 12336 1190
rect 12364 1162 12378 1190
rect 12218 406 12378 1162
rect 12558 1106 12586 1111
rect 12558 882 12586 1078
rect 12558 849 12586 854
rect 12218 378 12232 406
rect 12260 378 12284 406
rect 12312 378 12336 406
rect 12364 378 12378 406
rect 12218 0 12378 378
rect 13454 266 13482 1694
rect 14014 1106 14042 4214
rect 21888 3934 22048 4690
rect 21888 3906 21902 3934
rect 21930 3906 21954 3934
rect 21982 3906 22006 3934
rect 22034 3906 22048 3934
rect 21888 3150 22048 3906
rect 21888 3122 21902 3150
rect 21930 3122 21954 3150
rect 21982 3122 22006 3150
rect 22034 3122 22048 3150
rect 18550 2394 18858 2399
rect 18578 2371 18858 2394
rect 18550 2361 18578 2366
rect 18830 2338 18858 2371
rect 18830 2305 18858 2310
rect 21888 2366 22048 3122
rect 21888 2338 21902 2366
rect 21930 2338 21954 2366
rect 21982 2338 22006 2366
rect 22034 2338 22048 2366
rect 17206 2226 17234 2231
rect 17206 2058 17234 2198
rect 17206 2025 17234 2030
rect 14238 1890 14266 1895
rect 14238 1778 14266 1862
rect 14238 1745 14266 1750
rect 14014 1073 14042 1078
rect 21888 1582 22048 2338
rect 21888 1554 21902 1582
rect 21930 1554 21954 1582
rect 21982 1554 22006 1582
rect 22034 1554 22048 1582
rect 21798 938 21826 943
rect 18774 826 18802 831
rect 15862 770 15890 775
rect 15862 509 15890 742
rect 18774 602 18802 798
rect 18774 569 18802 574
rect 18886 714 18914 719
rect 18886 602 18914 686
rect 18886 569 18914 574
rect 15806 481 15890 509
rect 15806 378 15834 481
rect 15806 345 15834 350
rect 15918 378 15946 383
rect 13454 233 13482 238
rect 15918 266 15946 350
rect 21798 378 21826 910
rect 21798 345 21826 350
rect 21888 798 22048 1554
rect 21888 770 21902 798
rect 21930 770 21954 798
rect 21982 770 22006 798
rect 22034 770 22048 798
rect 15918 233 15946 238
rect 16702 322 16730 327
rect 16702 154 16730 294
rect 18718 322 18746 327
rect 18718 239 18746 294
rect 18718 211 18802 239
rect 18774 210 18802 211
rect 18774 177 18802 182
rect 16702 121 16730 126
rect 21888 0 22048 770
rect 22218 6678 22378 7112
rect 22218 6650 22232 6678
rect 22260 6650 22284 6678
rect 22312 6650 22336 6678
rect 22364 6650 22378 6678
rect 22218 5894 22378 6650
rect 22218 5866 22232 5894
rect 22260 5866 22284 5894
rect 22312 5866 22336 5894
rect 22364 5866 22378 5894
rect 22218 5110 22378 5866
rect 22218 5082 22232 5110
rect 22260 5082 22284 5110
rect 22312 5082 22336 5110
rect 22364 5082 22378 5110
rect 22218 4326 22378 5082
rect 22218 4298 22232 4326
rect 22260 4298 22284 4326
rect 22312 4298 22336 4326
rect 22364 4298 22378 4326
rect 22218 3542 22378 4298
rect 22218 3514 22232 3542
rect 22260 3514 22284 3542
rect 22312 3514 22336 3542
rect 22364 3514 22378 3542
rect 22218 2758 22378 3514
rect 22218 2730 22232 2758
rect 22260 2730 22284 2758
rect 22312 2730 22336 2758
rect 22364 2730 22378 2758
rect 22218 1974 22378 2730
rect 22218 1946 22232 1974
rect 22260 1946 22284 1974
rect 22312 1946 22336 1974
rect 22364 1946 22378 1974
rect 22218 1190 22378 1946
rect 22218 1162 22232 1190
rect 22260 1162 22284 1190
rect 22312 1162 22336 1190
rect 22364 1162 22378 1190
rect 22218 406 22378 1162
rect 22218 378 22232 406
rect 22260 378 22284 406
rect 22312 378 22336 406
rect 22364 378 22378 406
rect 22218 0 22378 378
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _000_
timestamp 1486834041
transform 1 0 9520 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _001_
timestamp 1486834041
transform 1 0 14728 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _002_
timestamp 1486834041
transform 1 0 23240 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _003_
timestamp 1486834041
transform 1 0 24640 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _004_
timestamp 1486834041
transform 1 0 1120 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _005_
timestamp 1486834041
transform 1 0 25368 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _006_
timestamp 1486834041
transform 1 0 21448 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _007_
timestamp 1486834041
transform 1 0 16128 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _008_
timestamp 1486834041
transform 1 0 17472 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _009_
timestamp 1486834041
transform 1 0 7224 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _010_
timestamp 1486834041
transform 1 0 15008 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _011_
timestamp 1486834041
transform 1 0 21728 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _012_
timestamp 1486834041
transform 1 0 20496 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _013_
timestamp 1486834041
transform 1 0 12712 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _014_
timestamp 1486834041
transform 1 0 7728 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _015_
timestamp 1486834041
transform 1 0 9632 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _016_
timestamp 1486834041
transform 1 0 12208 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _017_
timestamp 1486834041
transform 1 0 22008 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _018_
timestamp 1486834041
transform 1 0 10360 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _019_
timestamp 1486834041
transform 1 0 17472 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _020_
timestamp 1486834041
transform 1 0 16128 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _021_
timestamp 1486834041
transform 1 0 11144 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _022_
timestamp 1486834041
transform 1 0 14560 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _023_
timestamp 1486834041
transform 1 0 11256 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _024_
timestamp 1486834041
transform 1 0 18928 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _025_
timestamp 1486834041
transform 1 0 12712 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _026_
timestamp 1486834041
transform 1 0 14168 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _027_
timestamp 1486834041
transform 1 0 17248 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _028_
timestamp 1486834041
transform 1 0 17192 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _029_
timestamp 1486834041
transform 1 0 15344 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _030_
timestamp 1486834041
transform 1 0 11648 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _031_
timestamp 1486834041
transform 1 0 23352 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _032_
timestamp 1486834041
transform -1 0 23856 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _033_
timestamp 1486834041
transform 1 0 24696 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _034_
timestamp 1486834041
transform -1 0 5600 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _035_
timestamp 1486834041
transform -1 0 7504 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _036_
timestamp 1486834041
transform -1 0 9464 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _037_
timestamp 1486834041
transform -1 0 10696 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _038_
timestamp 1486834041
transform -1 0 11536 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _039_
timestamp 1486834041
transform -1 0 13608 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _040_
timestamp 1486834041
transform -1 0 14728 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _041_
timestamp 1486834041
transform -1 0 16688 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _042_
timestamp 1486834041
transform -1 0 24528 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _043_
timestamp 1486834041
transform -1 0 18928 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _044_
timestamp 1486834041
transform -1 0 20328 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _045_
timestamp 1486834041
transform -1 0 25984 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _046_
timestamp 1486834041
transform -1 0 26208 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _047_
timestamp 1486834041
transform -1 0 23632 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _048_
timestamp 1486834041
transform -1 0 24976 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _049_
timestamp 1486834041
transform -1 0 26712 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _050_
timestamp 1486834041
transform -1 0 26544 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _051_
timestamp 1486834041
transform -1 0 25760 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _052_
timestamp 1486834041
transform 1 0 8232 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _053_
timestamp 1486834041
transform 1 0 8568 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _054_
timestamp 1486834041
transform 1 0 9240 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _055_
timestamp 1486834041
transform 1 0 10360 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _056_
timestamp 1486834041
transform 1 0 11872 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _057_
timestamp 1486834041
transform 1 0 4704 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _058_
timestamp 1486834041
transform 1 0 11872 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _059_
timestamp 1486834041
transform 1 0 12880 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _060_
timestamp 1486834041
transform 1 0 14168 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _061_
timestamp 1486834041
transform 1 0 15288 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _062_
timestamp 1486834041
transform 1 0 14840 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _063_
timestamp 1486834041
transform 1 0 14392 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _064_
timestamp 1486834041
transform 1 0 13720 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _065_
timestamp 1486834041
transform 1 0 6832 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _066_
timestamp 1486834041
transform 1 0 12488 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _067_
timestamp 1486834041
transform 1 0 14280 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _068_
timestamp 1486834041
transform 1 0 15568 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _069_
timestamp 1486834041
transform 1 0 16184 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _070_
timestamp 1486834041
transform 1 0 17528 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _071_
timestamp 1486834041
transform 1 0 17528 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _072_
timestamp 1486834041
transform -1 0 1232 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _073_
timestamp 1486834041
transform 1 0 19264 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _074_
timestamp 1486834041
transform 1 0 18088 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _075_
timestamp 1486834041
transform 1 0 17248 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _076_
timestamp 1486834041
transform 1 0 17528 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _077_
timestamp 1486834041
transform 1 0 18592 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _078_
timestamp 1486834041
transform 1 0 19208 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _079_
timestamp 1486834041
transform 1 0 19544 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _080_
timestamp 1486834041
transform 1 0 19936 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _081_
timestamp 1486834041
transform 1 0 20664 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _082_
timestamp 1486834041
transform 1 0 21224 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _083_
timestamp 1486834041
transform 1 0 21560 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _084_
timestamp 1486834041
transform 1 0 22400 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _085_
timestamp 1486834041
transform 1 0 23184 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _086_
timestamp 1486834041
transform 1 0 22344 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _087_
timestamp 1486834041
transform 1 0 23408 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _088_
timestamp 1486834041
transform 1 0 26544 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _089_
timestamp 1486834041
transform 1 0 13160 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _090_
timestamp 1486834041
transform 1 0 12320 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _091_
timestamp 1486834041
transform 1 0 12208 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _092_
timestamp 1486834041
transform 1 0 11648 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _093_
timestamp 1486834041
transform 1 0 10864 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _094_
timestamp 1486834041
transform -1 0 10136 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _095_
timestamp 1486834041
transform -1 0 9408 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _096_
timestamp 1486834041
transform -1 0 9240 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _097_
timestamp 1486834041
transform -1 0 7504 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _098_
timestamp 1486834041
transform -1 0 6216 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _099_
timestamp 1486834041
transform -1 0 5544 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _100_
timestamp 1486834041
transform -1 0 5432 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _101_
timestamp 1486834041
transform -1 0 4928 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _102_
timestamp 1486834041
transform -1 0 3080 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _103_
timestamp 1486834041
transform -1 0 1680 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _104_
timestamp 1486834041
transform -1 0 22568 0 1 5880
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__000__I
timestamp 1486834041
transform 1 0 9408 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__001__I
timestamp 1486834041
transform -1 0 14728 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__002__I
timestamp 1486834041
transform -1 0 23240 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__003__I
timestamp 1486834041
transform -1 0 24640 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__004__I
timestamp 1486834041
transform -1 0 1120 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__005__I
timestamp 1486834041
transform -1 0 25368 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__006__I
timestamp 1486834041
transform 1 0 21336 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__007__I
timestamp 1486834041
transform -1 0 16128 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__008__I
timestamp 1486834041
transform 1 0 17360 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__009__I
timestamp 1486834041
transform -1 0 7224 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__010__I
timestamp 1486834041
transform -1 0 15008 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__011__I
timestamp 1486834041
transform 1 0 21616 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__012__I
timestamp 1486834041
transform -1 0 20496 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__013__I
timestamp 1486834041
transform -1 0 12712 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__014__I
timestamp 1486834041
transform 1 0 7616 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__015__I
timestamp 1486834041
transform 1 0 9520 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__016__I
timestamp 1486834041
transform 1 0 11984 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__017__I
timestamp 1486834041
transform -1 0 21896 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__018__I
timestamp 1486834041
transform 1 0 10248 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__019__I
timestamp 1486834041
transform 1 0 17360 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__020__I
timestamp 1486834041
transform -1 0 16016 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__021__I
timestamp 1486834041
transform -1 0 11144 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__022__I
timestamp 1486834041
transform -1 0 14560 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__023__I
timestamp 1486834041
transform 1 0 11144 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__024__I
timestamp 1486834041
transform 1 0 18816 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__025__I
timestamp 1486834041
transform 1 0 12600 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__026__I
timestamp 1486834041
transform -1 0 14056 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__027__I
timestamp 1486834041
transform -1 0 17248 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__028__I
timestamp 1486834041
transform 1 0 17080 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__029__I
timestamp 1486834041
transform 1 0 15232 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__030__I
timestamp 1486834041
transform 1 0 11536 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__031__I
timestamp 1486834041
transform 1 0 23240 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__032__I
timestamp 1486834041
transform 1 0 23968 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__033__I
timestamp 1486834041
transform -1 0 24696 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__034__I
timestamp 1486834041
transform -1 0 5712 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__035__I
timestamp 1486834041
transform 1 0 7504 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__036__I
timestamp 1486834041
transform 1 0 9464 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__037__I
timestamp 1486834041
transform -1 0 10808 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__038__I
timestamp 1486834041
transform 1 0 11536 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__039__I
timestamp 1486834041
transform -1 0 13720 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__040__I
timestamp 1486834041
transform -1 0 14840 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__041__I
timestamp 1486834041
transform 1 0 16688 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__042__I
timestamp 1486834041
transform -1 0 24640 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__043__I
timestamp 1486834041
transform -1 0 19040 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__044__I
timestamp 1486834041
transform -1 0 20440 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__045__I
timestamp 1486834041
transform 1 0 25984 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__046__I
timestamp 1486834041
transform -1 0 26264 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__047__I
timestamp 1486834041
transform 1 0 23632 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__048__I
timestamp 1486834041
transform 1 0 24976 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__049__I
timestamp 1486834041
transform -1 0 26152 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__050__I
timestamp 1486834041
transform -1 0 26656 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__051__I
timestamp 1486834041
transform -1 0 25816 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__052__I
timestamp 1486834041
transform -1 0 8232 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__053__I
timestamp 1486834041
transform -1 0 8568 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__054__I
timestamp 1486834041
transform 1 0 9128 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__055__I
timestamp 1486834041
transform 1 0 10248 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__056__I
timestamp 1486834041
transform -1 0 11872 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__057__I
timestamp 1486834041
transform 1 0 4592 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__058__I
timestamp 1486834041
transform -1 0 11872 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__059__I
timestamp 1486834041
transform -1 0 12880 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__060__I
timestamp 1486834041
transform -1 0 14056 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__061__I
timestamp 1486834041
transform 1 0 15176 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__062__I
timestamp 1486834041
transform 1 0 14728 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__063__I
timestamp 1486834041
transform 1 0 14280 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__064__I
timestamp 1486834041
transform -1 0 13720 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__065__I
timestamp 1486834041
transform -1 0 6832 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__066__I
timestamp 1486834041
transform 1 0 12376 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__067__I
timestamp 1486834041
transform -1 0 14280 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__068__I
timestamp 1486834041
transform 1 0 15456 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__069__I
timestamp 1486834041
transform -1 0 16184 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__070__I
timestamp 1486834041
transform -1 0 17192 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__071__I
timestamp 1486834041
transform -1 0 17528 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__072__I
timestamp 1486834041
transform 1 0 1232 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__073__I
timestamp 1486834041
transform 1 0 19152 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__074__I
timestamp 1486834041
transform 1 0 17976 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__075__I
timestamp 1486834041
transform 1 0 17136 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__076__I
timestamp 1486834041
transform -1 0 17528 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__077__I
timestamp 1486834041
transform -1 0 18592 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__078__I
timestamp 1486834041
transform 1 0 19096 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__079__I
timestamp 1486834041
transform -1 0 19544 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__080__I
timestamp 1486834041
transform -1 0 19936 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__081__I
timestamp 1486834041
transform -1 0 20664 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__082__I
timestamp 1486834041
transform 1 0 21112 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__083__I
timestamp 1486834041
transform 1 0 21448 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__084__I
timestamp 1486834041
transform -1 0 22400 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__085__I
timestamp 1486834041
transform -1 0 23184 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__086__I
timestamp 1486834041
transform 1 0 22232 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__087__I
timestamp 1486834041
transform 1 0 23296 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__088__I
timestamp 1486834041
transform -1 0 26544 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__089__I
timestamp 1486834041
transform 1 0 13048 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__090__I
timestamp 1486834041
transform 1 0 12208 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__091__I
timestamp 1486834041
transform 1 0 12096 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__092__I
timestamp 1486834041
transform 1 0 11536 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__093__I
timestamp 1486834041
transform 1 0 10752 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__094__I
timestamp 1486834041
transform 1 0 10136 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__095__I
timestamp 1486834041
transform -1 0 9520 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__096__I
timestamp 1486834041
transform 1 0 9240 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__097__I
timestamp 1486834041
transform -1 0 7616 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__098__I
timestamp 1486834041
transform -1 0 6440 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__099__I
timestamp 1486834041
transform 1 0 5544 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__100__I
timestamp 1486834041
transform -1 0 5544 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__101__I
timestamp 1486834041
transform -1 0 5040 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__102__I
timestamp 1486834041
transform -1 0 3192 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__103__I
timestamp 1486834041
transform -1 0 1792 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__104__I
timestamp 1486834041
transform -1 0 22680 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2
timestamp 1486834041
transform 1 0 448 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36
timestamp 1486834041
transform 1 0 2352 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_70
timestamp 1486834041
transform 1 0 4256 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_104
timestamp 1486834041
transform 1 0 6160 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_138
timestamp 1486834041
transform 1 0 8064 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_172
timestamp 1486834041
transform 1 0 9968 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_180
timestamp 1486834041
transform 1 0 10416 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_184
timestamp 1486834041
transform 1 0 10640 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_188
timestamp 1486834041
transform 1 0 10864 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_206
timestamp 1486834041
transform 1 0 11872 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_240
timestamp 1486834041
transform 1 0 13776 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_242
timestamp 1486834041
transform 1 0 13888 0 1 392
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_271
timestamp 1486834041
transform 1 0 15512 0 1 392
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_302
timestamp 1486834041
transform 1 0 17248 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_338
timestamp 1486834041
transform 1 0 19264 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_370
timestamp 1486834041
transform 1 0 21056 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_404
timestamp 1486834041
transform 1 0 22960 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_438
timestamp 1486834041
transform 1 0 24864 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_444
timestamp 1486834041
transform 1 0 25200 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_478
timestamp 1486834041
transform 1 0 27104 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_482
timestamp 1486834041
transform 1 0 27328 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_484
timestamp 1486834041
transform 1 0 27440 0 1 392
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_2
timestamp 1486834041
transform 1 0 448 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_6
timestamp 1486834041
transform 1 0 672 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_18
timestamp 1486834041
transform 1 0 1344 0 -1 1176
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_50
timestamp 1486834041
transform 1 0 3136 0 -1 1176
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_66
timestamp 1486834041
transform 1 0 4032 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_72
timestamp 1486834041
transform 1 0 4368 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_86
timestamp 1486834041
transform 1 0 5152 0 -1 1176
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_118
timestamp 1486834041
transform 1 0 6944 0 -1 1176
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_134
timestamp 1486834041
transform 1 0 7840 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_138
timestamp 1486834041
transform 1 0 8064 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_142
timestamp 1486834041
transform 1 0 8288 0 -1 1176
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_158
timestamp 1486834041
transform 1 0 9184 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_172
timestamp 1486834041
transform 1 0 9968 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_176
timestamp 1486834041
transform 1 0 10192 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_187
timestamp 1486834041
transform 1 0 10808 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_212
timestamp 1486834041
transform 1 0 12208 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_214
timestamp 1486834041
transform 1 0 12320 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_267
timestamp 1486834041
transform 1 0 15288 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_269
timestamp 1486834041
transform 1 0 15400 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_346
timestamp 1486834041
transform 1 0 19712 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_418
timestamp 1486834041
transform 1 0 23744 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_460
timestamp 1486834041
transform 1 0 26096 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_492
timestamp 1486834041
transform 1 0 27888 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_496
timestamp 1486834041
transform 1 0 28112 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_498
timestamp 1486834041
transform 1 0 28224 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_2
timestamp 1486834041
transform 1 0 448 0 1 1176
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1486834041
transform 1 0 2240 0 1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_37
timestamp 1486834041
transform 1 0 2408 0 1 1176
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_101
timestamp 1486834041
transform 1 0 5992 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_107
timestamp 1486834041
transform 1 0 6328 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_111
timestamp 1486834041
transform 1 0 6552 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_113
timestamp 1486834041
transform 1 0 6664 0 1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_124
timestamp 1486834041
transform 1 0 7280 0 1 1176
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_140
timestamp 1486834041
transform 1 0 8176 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_144
timestamp 1486834041
transform 1 0 8400 0 1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_155
timestamp 1486834041
transform 1 0 9016 0 1 1176
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_171
timestamp 1486834041
transform 1 0 9912 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_177
timestamp 1486834041
transform 1 0 10248 0 1 1176
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_209
timestamp 1486834041
transform 1 0 12040 0 1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_212
timestamp 1486834041
transform 1 0 12208 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_216
timestamp 1486834041
transform 1 0 12432 0 1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_373
timestamp 1486834041
transform 1 0 21224 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_443
timestamp 1486834041
transform 1 0 25144 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_2
timestamp 1486834041
transform 1 0 448 0 -1 1960
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_66
timestamp 1486834041
transform 1 0 4032 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_72
timestamp 1486834041
transform 1 0 4368 0 -1 1960
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_136
timestamp 1486834041
transform 1 0 7952 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_142
timestamp 1486834041
transform 1 0 8288 0 -1 1960
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_174
timestamp 1486834041
transform 1 0 10080 0 -1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_190
timestamp 1486834041
transform 1 0 10976 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_198
timestamp 1486834041
transform 1 0 11424 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_220
timestamp 1486834041
transform 1 0 12656 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_224
timestamp 1486834041
transform 1 0 12880 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_247
timestamp 1486834041
transform 1 0 14168 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_257
timestamp 1486834041
transform 1 0 14728 0 -1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_273
timestamp 1486834041
transform 1 0 15624 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_277
timestamp 1486834041
transform 1 0 15848 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_279
timestamp 1486834041
transform 1 0 15960 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_296
timestamp 1486834041
transform 1 0 16912 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_298
timestamp 1486834041
transform 1 0 17024 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_345
timestamp 1486834041
transform 1 0 19656 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_349
timestamp 1486834041
transform 1 0 19880 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_416
timestamp 1486834041
transform 1 0 23632 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_422
timestamp 1486834041
transform 1 0 23968 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_442
timestamp 1486834041
transform 1 0 25088 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_492
timestamp 1486834041
transform 1 0 27888 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_496
timestamp 1486834041
transform 1 0 28112 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_498
timestamp 1486834041
transform 1 0 28224 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_2
timestamp 1486834041
transform 1 0 448 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_10
timestamp 1486834041
transform 1 0 896 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_14
timestamp 1486834041
transform 1 0 1120 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_26
timestamp 1486834041
transform 1 0 1792 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1486834041
transform 1 0 2240 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_37
timestamp 1486834041
transform 1 0 2408 0 1 1960
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_69
timestamp 1486834041
transform 1 0 4200 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_77
timestamp 1486834041
transform 1 0 4648 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_81
timestamp 1486834041
transform 1 0 4872 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_93
timestamp 1486834041
transform 1 0 5544 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_109
timestamp 1486834041
transform 1 0 6440 0 1 1960
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_141
timestamp 1486834041
transform 1 0 8232 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_149
timestamp 1486834041
transform 1 0 8680 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_153
timestamp 1486834041
transform 1 0 8904 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_164
timestamp 1486834041
transform 1 0 9520 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_172
timestamp 1486834041
transform 1 0 9968 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_174
timestamp 1486834041
transform 1 0 10080 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_177
timestamp 1486834041
transform 1 0 10248 0 1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_193
timestamp 1486834041
transform 1 0 11144 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_201
timestamp 1486834041
transform 1 0 11592 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_203
timestamp 1486834041
transform 1 0 11704 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_214
timestamp 1486834041
transform 1 0 12320 0 1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_230
timestamp 1486834041
transform 1 0 13216 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_234
timestamp 1486834041
transform 1 0 13440 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_236
timestamp 1486834041
transform 1 0 13552 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_239
timestamp 1486834041
transform 1 0 13720 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_243
timestamp 1486834041
transform 1 0 13944 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_247
timestamp 1486834041
transform 1 0 14168 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_255
timestamp 1486834041
transform 1 0 14616 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_259
timestamp 1486834041
transform 1 0 14840 0 1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_275
timestamp 1486834041
transform 1 0 15736 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_279
timestamp 1486834041
transform 1 0 15960 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_291
timestamp 1486834041
transform 1 0 16632 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_299
timestamp 1486834041
transform 1 0 17080 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_303
timestamp 1486834041
transform 1 0 17304 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_325
timestamp 1486834041
transform 1 0 18536 0 1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_351
timestamp 1486834041
transform 1 0 19992 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_359
timestamp 1486834041
transform 1 0 20440 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_371
timestamp 1486834041
transform 1 0 21112 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_379
timestamp 1486834041
transform 1 0 21560 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_383
timestamp 1486834041
transform 1 0 21784 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_387
timestamp 1486834041
transform 1 0 22008 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_391
timestamp 1486834041
transform 1 0 22232 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_402
timestamp 1486834041
transform 1 0 22848 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_408
timestamp 1486834041
transform 1 0 23184 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_423
timestamp 1486834041
transform 1 0 24024 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_431
timestamp 1486834041
transform 1 0 24472 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_434
timestamp 1486834041
transform 1 0 24640 0 1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_450
timestamp 1486834041
transform 1 0 25536 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_452
timestamp 1486834041
transform 1 0 25648 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_457
timestamp 1486834041
transform 1 0 25928 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_2
timestamp 1486834041
transform 1 0 448 0 -1 2744
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_66
timestamp 1486834041
transform 1 0 4032 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_72
timestamp 1486834041
transform 1 0 4368 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_80
timestamp 1486834041
transform 1 0 4816 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_84
timestamp 1486834041
transform 1 0 5040 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_95
timestamp 1486834041
transform 1 0 5656 0 -1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_127
timestamp 1486834041
transform 1 0 7448 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_135
timestamp 1486834041
transform 1 0 7896 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_139
timestamp 1486834041
transform 1 0 8120 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_142
timestamp 1486834041
transform 1 0 8288 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_150
timestamp 1486834041
transform 1 0 8736 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_154
timestamp 1486834041
transform 1 0 8960 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_156
timestamp 1486834041
transform 1 0 9072 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_177
timestamp 1486834041
transform 1 0 10248 0 -1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_209
timestamp 1486834041
transform 1 0 12040 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_214
timestamp 1486834041
transform 1 0 12320 0 -1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_246
timestamp 1486834041
transform 1 0 14112 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_248
timestamp 1486834041
transform 1 0 14224 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_267
timestamp 1486834041
transform 1 0 15288 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_275
timestamp 1486834041
transform 1 0 15736 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_277
timestamp 1486834041
transform 1 0 15848 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_290
timestamp 1486834041
transform 1 0 16576 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_298
timestamp 1486834041
transform 1 0 17024 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_310
timestamp 1486834041
transform 1 0 17696 0 -1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_326
timestamp 1486834041
transform 1 0 18592 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_334
timestamp 1486834041
transform 1 0 19040 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_345
timestamp 1486834041
transform 1 0 19656 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_349
timestamp 1486834041
transform 1 0 19880 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_352
timestamp 1486834041
transform 1 0 20048 0 -1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_368
timestamp 1486834041
transform 1 0 20944 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_370
timestamp 1486834041
transform 1 0 21056 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_381
timestamp 1486834041
transform 1 0 21672 0 -1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_397
timestamp 1486834041
transform 1 0 22568 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_405
timestamp 1486834041
transform 1 0 23016 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_409
timestamp 1486834041
transform 1 0 23240 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_422
timestamp 1486834041
transform 1 0 23968 0 -1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_454
timestamp 1486834041
transform 1 0 25760 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_458
timestamp 1486834041
transform 1 0 25984 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_492
timestamp 1486834041
transform 1 0 27888 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_496
timestamp 1486834041
transform 1 0 28112 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_498
timestamp 1486834041
transform 1 0 28224 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1486834041
transform 1 0 448 0 1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1486834041
transform 1 0 2240 0 1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_37
timestamp 1486834041
transform 1 0 2408 0 1 2744
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_101
timestamp 1486834041
transform 1 0 5992 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_107
timestamp 1486834041
transform 1 0 6328 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_115
timestamp 1486834041
transform 1 0 6776 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_119
timestamp 1486834041
transform 1 0 7000 0 1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_130
timestamp 1486834041
transform 1 0 7616 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_138
timestamp 1486834041
transform 1 0 8064 0 1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_149
timestamp 1486834041
transform 1 0 8680 0 1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_165
timestamp 1486834041
transform 1 0 9576 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_173
timestamp 1486834041
transform 1 0 10024 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_177
timestamp 1486834041
transform 1 0 10248 0 1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_193
timestamp 1486834041
transform 1 0 11144 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_201
timestamp 1486834041
transform 1 0 11592 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_203
timestamp 1486834041
transform 1 0 11704 0 1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_222
timestamp 1486834041
transform 1 0 12768 0 1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_238
timestamp 1486834041
transform 1 0 13664 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_242
timestamp 1486834041
transform 1 0 13888 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_244
timestamp 1486834041
transform 1 0 14000 0 1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_247
timestamp 1486834041
transform 1 0 14168 0 1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_279
timestamp 1486834041
transform 1 0 15960 0 1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_295
timestamp 1486834041
transform 1 0 16856 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_303
timestamp 1486834041
transform 1 0 17304 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_317
timestamp 1486834041
transform 1 0 18088 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_321
timestamp 1486834041
transform 1 0 18312 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_323
timestamp 1486834041
transform 1 0 18424 0 1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_334
timestamp 1486834041
transform 1 0 19040 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_342
timestamp 1486834041
transform 1 0 19488 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_346
timestamp 1486834041
transform 1 0 19712 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_358
timestamp 1486834041
transform 1 0 20384 0 1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_374
timestamp 1486834041
transform 1 0 21280 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_382
timestamp 1486834041
transform 1 0 21728 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_384
timestamp 1486834041
transform 1 0 21840 0 1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_387
timestamp 1486834041
transform 1 0 22008 0 1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_403
timestamp 1486834041
transform 1 0 22904 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_417
timestamp 1486834041
transform 1 0 23688 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_425
timestamp 1486834041
transform 1 0 24136 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_429
timestamp 1486834041
transform 1 0 24360 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_431
timestamp 1486834041
transform 1 0 24472 0 1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_442
timestamp 1486834041
transform 1 0 25088 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_450
timestamp 1486834041
transform 1 0 25536 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_454
timestamp 1486834041
transform 1 0 25760 0 1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_457
timestamp 1486834041
transform 1 0 25928 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_465
timestamp 1486834041
transform 1 0 26376 0 1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_470
timestamp 1486834041
transform 1 0 26656 0 1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_2
timestamp 1486834041
transform 1 0 448 0 -1 3528
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_66
timestamp 1486834041
transform 1 0 4032 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_72
timestamp 1486834041
transform 1 0 4368 0 -1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_104
timestamp 1486834041
transform 1 0 6160 0 -1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_120
timestamp 1486834041
transform 1 0 7056 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_128
timestamp 1486834041
transform 1 0 7504 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_142
timestamp 1486834041
transform 1 0 8288 0 -1 3528
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_206
timestamp 1486834041
transform 1 0 11872 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_212
timestamp 1486834041
transform 1 0 12208 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_220
timestamp 1486834041
transform 1 0 12656 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_224
timestamp 1486834041
transform 1 0 12880 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_226
timestamp 1486834041
transform 1 0 12992 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_237
timestamp 1486834041
transform 1 0 13608 0 -1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_269
timestamp 1486834041
transform 1 0 15400 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_277
timestamp 1486834041
transform 1 0 15848 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_279
timestamp 1486834041
transform 1 0 15960 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_282
timestamp 1486834041
transform 1 0 16128 0 -1 3528
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_346
timestamp 1486834041
transform 1 0 19712 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_352
timestamp 1486834041
transform 1 0 20048 0 -1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_368
timestamp 1486834041
transform 1 0 20944 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_376
timestamp 1486834041
transform 1 0 21392 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_387
timestamp 1486834041
transform 1 0 22008 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_401
timestamp 1486834041
transform 1 0 22792 0 -1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_417
timestamp 1486834041
transform 1 0 23688 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_419
timestamp 1486834041
transform 1 0 23800 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_422
timestamp 1486834041
transform 1 0 23968 0 -1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_454
timestamp 1486834041
transform 1 0 25760 0 -1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_470
timestamp 1486834041
transform 1 0 26656 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_474
timestamp 1486834041
transform 1 0 26880 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_492
timestamp 1486834041
transform 1 0 27888 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_496
timestamp 1486834041
transform 1 0 28112 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_498
timestamp 1486834041
transform 1 0 28224 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1486834041
transform 1 0 448 0 1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1486834041
transform 1 0 2240 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_37
timestamp 1486834041
transform 1 0 2408 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_51
timestamp 1486834041
transform 1 0 3192 0 1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_67
timestamp 1486834041
transform 1 0 4088 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_71
timestamp 1486834041
transform 1 0 4312 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_73
timestamp 1486834041
transform 1 0 4424 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_84
timestamp 1486834041
transform 1 0 5040 0 1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_100
timestamp 1486834041
transform 1 0 5936 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_104
timestamp 1486834041
transform 1 0 6160 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_107
timestamp 1486834041
transform 1 0 6328 0 1 3528
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_171
timestamp 1486834041
transform 1 0 9912 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_187
timestamp 1486834041
transform 1 0 10808 0 1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_219
timestamp 1486834041
transform 1 0 12600 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_221
timestamp 1486834041
transform 1 0 12712 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_232
timestamp 1486834041
transform 1 0 13328 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_240
timestamp 1486834041
transform 1 0 13776 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_244
timestamp 1486834041
transform 1 0 14000 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_247
timestamp 1486834041
transform 1 0 14168 0 1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_279
timestamp 1486834041
transform 1 0 15960 0 1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_295
timestamp 1486834041
transform 1 0 16856 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_303
timestamp 1486834041
transform 1 0 17304 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_314
timestamp 1486834041
transform 1 0 17920 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_317
timestamp 1486834041
transform 1 0 18088 0 1 3528
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_381
timestamp 1486834041
transform 1 0 21672 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_387
timestamp 1486834041
transform 1 0 22008 0 1 3528
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_451
timestamp 1486834041
transform 1 0 25592 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_457
timestamp 1486834041
transform 1 0 25928 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_465
timestamp 1486834041
transform 1 0 26376 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_469
timestamp 1486834041
transform 1 0 26600 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_2
timestamp 1486834041
transform 1 0 448 0 -1 4312
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_66
timestamp 1486834041
transform 1 0 4032 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_72
timestamp 1486834041
transform 1 0 4368 0 -1 4312
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_136
timestamp 1486834041
transform 1 0 7952 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_142
timestamp 1486834041
transform 1 0 8288 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_150
timestamp 1486834041
transform 1 0 8736 0 -1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_161
timestamp 1486834041
transform 1 0 9352 0 -1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_177
timestamp 1486834041
transform 1 0 10248 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_185
timestamp 1486834041
transform 1 0 10696 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_189
timestamp 1486834041
transform 1 0 10920 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_201
timestamp 1486834041
transform 1 0 11592 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_209
timestamp 1486834041
transform 1 0 12040 0 -1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_212
timestamp 1486834041
transform 1 0 12208 0 -1 4312
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_244
timestamp 1486834041
transform 1 0 14000 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_262
timestamp 1486834041
transform 1 0 15008 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_264
timestamp 1486834041
transform 1 0 15120 0 -1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_275
timestamp 1486834041
transform 1 0 15736 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_279
timestamp 1486834041
transform 1 0 15960 0 -1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_282
timestamp 1486834041
transform 1 0 16128 0 -1 4312
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_346
timestamp 1486834041
transform 1 0 19712 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_352
timestamp 1486834041
transform 1 0 20048 0 -1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_368
timestamp 1486834041
transform 1 0 20944 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_376
timestamp 1486834041
transform 1 0 21392 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_390
timestamp 1486834041
transform 1 0 22176 0 -1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_406
timestamp 1486834041
transform 1 0 23072 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_414
timestamp 1486834041
transform 1 0 23520 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_418
timestamp 1486834041
transform 1 0 23744 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_422
timestamp 1486834041
transform 1 0 23968 0 -1 4312
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_454
timestamp 1486834041
transform 1 0 25760 0 -1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_470
timestamp 1486834041
transform 1 0 26656 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_474
timestamp 1486834041
transform 1 0 26880 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_492
timestamp 1486834041
transform 1 0 27888 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_496
timestamp 1486834041
transform 1 0 28112 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_498
timestamp 1486834041
transform 1 0 28224 0 -1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_2
timestamp 1486834041
transform 1 0 448 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_10
timestamp 1486834041
transform 1 0 896 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_22
timestamp 1486834041
transform 1 0 1568 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_30
timestamp 1486834041
transform 1 0 2016 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1486834041
transform 1 0 2240 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_37
timestamp 1486834041
transform 1 0 2408 0 1 4312
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_101
timestamp 1486834041
transform 1 0 5992 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_107
timestamp 1486834041
transform 1 0 6328 0 1 4312
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_171
timestamp 1486834041
transform 1 0 9912 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_177
timestamp 1486834041
transform 1 0 10248 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_203
timestamp 1486834041
transform 1 0 11704 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_229
timestamp 1486834041
transform 1 0 13160 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_237
timestamp 1486834041
transform 1 0 13608 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_241
timestamp 1486834041
transform 1 0 13832 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_255
timestamp 1486834041
transform 1 0 14616 0 1 4312
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_287
timestamp 1486834041
transform 1 0 16408 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_303
timestamp 1486834041
transform 1 0 17304 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_311
timestamp 1486834041
transform 1 0 17752 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_317
timestamp 1486834041
transform 1 0 18088 0 1 4312
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_349
timestamp 1486834041
transform 1 0 19880 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_357
timestamp 1486834041
transform 1 0 20328 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_368
timestamp 1486834041
transform 1 0 20944 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_376
timestamp 1486834041
transform 1 0 21392 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_380
timestamp 1486834041
transform 1 0 21616 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_382
timestamp 1486834041
transform 1 0 21728 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_395
timestamp 1486834041
transform 1 0 22456 0 1 4312
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_427
timestamp 1486834041
transform 1 0 24248 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_443
timestamp 1486834041
transform 1 0 25144 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_451
timestamp 1486834041
transform 1 0 25592 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_457
timestamp 1486834041
transform 1 0 25928 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_465
timestamp 1486834041
transform 1 0 26376 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_469
timestamp 1486834041
transform 1 0 26600 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_2
timestamp 1486834041
transform 1 0 448 0 -1 5096
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_66
timestamp 1486834041
transform 1 0 4032 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_72
timestamp 1486834041
transform 1 0 4368 0 -1 5096
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_136
timestamp 1486834041
transform 1 0 7952 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_142
timestamp 1486834041
transform 1 0 8288 0 -1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_158
timestamp 1486834041
transform 1 0 9184 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_162
timestamp 1486834041
transform 1 0 9408 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_174
timestamp 1486834041
transform 1 0 10080 0 -1 5096
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_206
timestamp 1486834041
transform 1 0 11872 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_212
timestamp 1486834041
transform 1 0 12208 0 -1 5096
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_276
timestamp 1486834041
transform 1 0 15792 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_282
timestamp 1486834041
transform 1 0 16128 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_294
timestamp 1486834041
transform 1 0 16800 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_298
timestamp 1486834041
transform 1 0 17024 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_310
timestamp 1486834041
transform 1 0 17696 0 -1 5096
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_342
timestamp 1486834041
transform 1 0 19488 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_352
timestamp 1486834041
transform 1 0 20048 0 -1 5096
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_416
timestamp 1486834041
transform 1 0 23632 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_422
timestamp 1486834041
transform 1 0 23968 0 -1 5096
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_454
timestamp 1486834041
transform 1 0 25760 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_492
timestamp 1486834041
transform 1 0 27888 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_496
timestamp 1486834041
transform 1 0 28112 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_498
timestamp 1486834041
transform 1 0 28224 0 -1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_2
timestamp 1486834041
transform 1 0 448 0 1 5096
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1486834041
transform 1 0 2240 0 1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_37
timestamp 1486834041
transform 1 0 2408 0 1 5096
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_101
timestamp 1486834041
transform 1 0 5992 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_107
timestamp 1486834041
transform 1 0 6328 0 1 5096
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_171
timestamp 1486834041
transform 1 0 9912 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_177
timestamp 1486834041
transform 1 0 10248 0 1 5096
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_241
timestamp 1486834041
transform 1 0 13832 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_247
timestamp 1486834041
transform 1 0 14168 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_259
timestamp 1486834041
transform 1 0 14840 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_263
timestamp 1486834041
transform 1 0 15064 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_265
timestamp 1486834041
transform 1 0 15176 0 1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_276
timestamp 1486834041
transform 1 0 15792 0 1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_292
timestamp 1486834041
transform 1 0 16688 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_296
timestamp 1486834041
transform 1 0 16912 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_298
timestamp 1486834041
transform 1 0 17024 0 1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_309
timestamp 1486834041
transform 1 0 17640 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_313
timestamp 1486834041
transform 1 0 17864 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_317
timestamp 1486834041
transform 1 0 18088 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_325
timestamp 1486834041
transform 1 0 18536 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_329
timestamp 1486834041
transform 1 0 18760 0 1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_340
timestamp 1486834041
transform 1 0 19376 0 1 5096
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_372
timestamp 1486834041
transform 1 0 21168 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_380
timestamp 1486834041
transform 1 0 21616 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_384
timestamp 1486834041
transform 1 0 21840 0 1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_387
timestamp 1486834041
transform 1 0 22008 0 1 5096
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_451
timestamp 1486834041
transform 1 0 25592 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_2
timestamp 1486834041
transform 1 0 448 0 -1 5880
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_66
timestamp 1486834041
transform 1 0 4032 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_72
timestamp 1486834041
transform 1 0 4368 0 -1 5880
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_104
timestamp 1486834041
transform 1 0 6160 0 -1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_130
timestamp 1486834041
transform 1 0 7616 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_138
timestamp 1486834041
transform 1 0 8064 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_142
timestamp 1486834041
transform 1 0 8288 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_150
timestamp 1486834041
transform 1 0 8736 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_154
timestamp 1486834041
transform 1 0 8960 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_165
timestamp 1486834041
transform 1 0 9576 0 -1 5880
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_197
timestamp 1486834041
transform 1 0 11368 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_199
timestamp 1486834041
transform 1 0 11480 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_202
timestamp 1486834041
transform 1 0 11648 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_206
timestamp 1486834041
transform 1 0 11872 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_220
timestamp 1486834041
transform 1 0 12656 0 -1 5880
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_252
timestamp 1486834041
transform 1 0 14448 0 -1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_268
timestamp 1486834041
transform 1 0 15344 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_276
timestamp 1486834041
transform 1 0 15792 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_282
timestamp 1486834041
transform 1 0 16128 0 -1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_298
timestamp 1486834041
transform 1 0 17024 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_302
timestamp 1486834041
transform 1 0 17248 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_314
timestamp 1486834041
transform 1 0 17920 0 -1 5880
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_346
timestamp 1486834041
transform 1 0 19712 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_352
timestamp 1486834041
transform 1 0 20048 0 -1 5880
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_384
timestamp 1486834041
transform 1 0 21840 0 -1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_400
timestamp 1486834041
transform 1 0 22736 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_408
timestamp 1486834041
transform 1 0 23184 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_424
timestamp 1486834041
transform 1 0 24080 0 -1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_440
timestamp 1486834041
transform 1 0 24976 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_492
timestamp 1486834041
transform 1 0 27888 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_496
timestamp 1486834041
transform 1 0 28112 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_498
timestamp 1486834041
transform 1 0 28224 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_2
timestamp 1486834041
transform 1 0 448 0 1 5880
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1486834041
transform 1 0 2240 0 1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_37
timestamp 1486834041
transform 1 0 2408 0 1 5880
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_69
timestamp 1486834041
transform 1 0 4200 0 1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_85
timestamp 1486834041
transform 1 0 5096 0 1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_96
timestamp 1486834041
transform 1 0 5712 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_104
timestamp 1486834041
transform 1 0 6160 0 1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_107
timestamp 1486834041
transform 1 0 6328 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_115
timestamp 1486834041
transform 1 0 6776 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_119
timestamp 1486834041
transform 1 0 7000 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_145
timestamp 1486834041
transform 1 0 8456 0 1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_161
timestamp 1486834041
transform 1 0 9352 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_169
timestamp 1486834041
transform 1 0 9800 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_173
timestamp 1486834041
transform 1 0 10024 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_187
timestamp 1486834041
transform 1 0 10808 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_191
timestamp 1486834041
transform 1 0 11032 0 1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_210
timestamp 1486834041
transform 1 0 12096 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_218
timestamp 1486834041
transform 1 0 12544 0 1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_239
timestamp 1486834041
transform 1 0 13720 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_255
timestamp 1486834041
transform 1 0 14616 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_259
timestamp 1486834041
transform 1 0 14840 0 1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_270
timestamp 1486834041
transform 1 0 15456 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_278
timestamp 1486834041
transform 1 0 15904 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_290
timestamp 1486834041
transform 1 0 16576 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_298
timestamp 1486834041
transform 1 0 17024 0 1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_313
timestamp 1486834041
transform 1 0 17864 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_317
timestamp 1486834041
transform 1 0 18088 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_321
timestamp 1486834041
transform 1 0 18312 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_323
timestamp 1486834041
transform 1 0 18424 0 1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_334
timestamp 1486834041
transform 1 0 19040 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_342
timestamp 1486834041
transform 1 0 19488 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_346
timestamp 1486834041
transform 1 0 19712 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_348
timestamp 1486834041
transform 1 0 19824 0 1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_359
timestamp 1486834041
transform 1 0 20440 0 1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_375
timestamp 1486834041
transform 1 0 21336 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_383
timestamp 1486834041
transform 1 0 21784 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_387
timestamp 1486834041
transform 1 0 22008 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_399
timestamp 1486834041
transform 1 0 22680 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_407
timestamp 1486834041
transform 1 0 23128 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_419
timestamp 1486834041
transform 1 0 23800 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_427
timestamp 1486834041
transform 1 0 24248 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_431
timestamp 1486834041
transform 1 0 24472 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_443
timestamp 1486834041
transform 1 0 25144 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_451
timestamp 1486834041
transform 1 0 25592 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_2
timestamp 1486834041
transform 1 0 448 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_10
timestamp 1486834041
transform 1 0 896 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_17
timestamp 1486834041
transform 1 0 1288 0 -1 6664
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_33
timestamp 1486834041
transform 1 0 2184 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_50
timestamp 1486834041
transform 1 0 3136 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_70
timestamp 1486834041
transform 1 0 4256 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_78
timestamp 1486834041
transform 1 0 4704 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_82
timestamp 1486834041
transform 1 0 4928 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_97
timestamp 1486834041
transform 1 0 5768 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_101
timestamp 1486834041
transform 1 0 5992 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_104
timestamp 1486834041
transform 1 0 6160 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_106
timestamp 1486834041
transform 1 0 6272 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_121
timestamp 1486834041
transform 1 0 7112 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_129
timestamp 1486834041
transform 1 0 7560 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_133
timestamp 1486834041
transform 1 0 7784 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_135
timestamp 1486834041
transform 1 0 7896 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_138
timestamp 1486834041
transform 1 0 8064 0 -1 6664
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_154
timestamp 1486834041
transform 1 0 8960 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_169
timestamp 1486834041
transform 1 0 9800 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_172
timestamp 1486834041
transform 1 0 9968 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_176
timestamp 1486834041
transform 1 0 10192 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_178
timestamp 1486834041
transform 1 0 10304 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_193
timestamp 1486834041
transform 1 0 11144 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_201
timestamp 1486834041
transform 1 0 11592 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_203
timestamp 1486834041
transform 1 0 11704 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_220
timestamp 1486834041
transform 1 0 12656 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_240
timestamp 1486834041
transform 1 0 13776 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_248
timestamp 1486834041
transform 1 0 14224 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_250
timestamp 1486834041
transform 1 0 14336 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_265
timestamp 1486834041
transform 1 0 15176 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_269
timestamp 1486834041
transform 1 0 15400 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_271
timestamp 1486834041
transform 1 0 15512 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_274
timestamp 1486834041
transform 1 0 15680 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_289
timestamp 1486834041
transform 1 0 16520 0 -1 6664
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_305
timestamp 1486834041
transform 1 0 17416 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_308
timestamp 1486834041
transform 1 0 17584 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_316
timestamp 1486834041
transform 1 0 18032 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_320
timestamp 1486834041
transform 1 0 18256 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_322
timestamp 1486834041
transform 1 0 18368 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_337
timestamp 1486834041
transform 1 0 19208 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_339
timestamp 1486834041
transform 1 0 19320 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_342
timestamp 1486834041
transform 1 0 19488 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_346
timestamp 1486834041
transform 1 0 19712 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_361
timestamp 1486834041
transform 1 0 20552 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_369
timestamp 1486834041
transform 1 0 21000 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_373
timestamp 1486834041
transform 1 0 21224 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_390
timestamp 1486834041
transform 1 0 22176 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_410
timestamp 1486834041
transform 1 0 23296 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_418
timestamp 1486834041
transform 1 0 23744 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_433
timestamp 1486834041
transform 1 0 24584 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_441
timestamp 1486834041
transform 1 0 25032 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_458
timestamp 1486834041
transform 1 0 25984 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_478
timestamp 1486834041
transform 1 0 27104 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_482
timestamp 1486834041
transform 1 0 27328 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_484
timestamp 1486834041
transform 1 0 27440 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output1
timestamp 1486834041
transform 1 0 25928 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output2
timestamp 1486834041
transform 1 0 26712 0 1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output3
timestamp 1486834041
transform 1 0 26992 0 -1 2744
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output4
timestamp 1486834041
transform 1 0 27496 0 1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output5
timestamp 1486834041
transform 1 0 26712 0 1 2744
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output6
timestamp 1486834041
transform 1 0 26992 0 -1 3528
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output7
timestamp 1486834041
transform 1 0 27496 0 1 2744
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output8
timestamp 1486834041
transform 1 0 26712 0 1 3528
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output9
timestamp 1486834041
transform 1 0 27496 0 1 3528
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output10
timestamp 1486834041
transform 1 0 27496 0 1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output11
timestamp 1486834041
transform 1 0 26712 0 1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output12
timestamp 1486834041
transform 1 0 26208 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output13
timestamp 1486834041
transform 1 0 27496 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output14
timestamp 1486834041
transform 1 0 26992 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output15
timestamp 1486834041
transform 1 0 26712 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output16
timestamp 1486834041
transform 1 0 27496 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output17
timestamp 1486834041
transform 1 0 26992 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output18
timestamp 1486834041
transform 1 0 27496 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output19
timestamp 1486834041
transform 1 0 26712 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output20
timestamp 1486834041
transform 1 0 26208 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output21
timestamp 1486834041
transform 1 0 25928 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output22
timestamp 1486834041
transform 1 0 26992 0 -1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output23
timestamp 1486834041
transform 1 0 25424 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output24
timestamp 1486834041
transform 1 0 26208 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output25
timestamp 1486834041
transform 1 0 25424 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output26
timestamp 1486834041
transform 1 0 26208 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output27
timestamp 1486834041
transform 1 0 26208 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output28
timestamp 1486834041
transform 1 0 26992 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output29
timestamp 1486834041
transform 1 0 27496 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output30
timestamp 1486834041
transform 1 0 26712 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output31
timestamp 1486834041
transform 1 0 26992 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output32
timestamp 1486834041
transform 1 0 27496 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output33
timestamp 1486834041
transform -1 0 3136 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output34
timestamp 1486834041
transform -1 0 16520 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output35
timestamp 1486834041
transform -1 0 17864 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output36
timestamp 1486834041
transform -1 0 19208 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output37
timestamp 1486834041
transform -1 0 20552 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output38
timestamp 1486834041
transform -1 0 22176 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output39
timestamp 1486834041
transform -1 0 23184 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output40
timestamp 1486834041
transform -1 0 24584 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output41
timestamp 1486834041
transform -1 0 25984 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output42
timestamp 1486834041
transform 1 0 26208 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output43
timestamp 1486834041
transform 1 0 25928 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output44
timestamp 1486834041
transform -1 0 4144 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output45
timestamp 1486834041
transform 1 0 4984 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output46
timestamp 1486834041
transform -1 0 7112 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output47
timestamp 1486834041
transform -1 0 8456 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output48
timestamp 1486834041
transform -1 0 9800 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output49
timestamp 1486834041
transform -1 0 11144 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output50
timestamp 1486834041
transform -1 0 12656 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output51
timestamp 1486834041
transform -1 0 13664 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output52
timestamp 1486834041
transform -1 0 15176 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output53
timestamp 1486834041
transform 1 0 11312 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output54
timestamp 1486834041
transform 1 0 10976 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output55
timestamp 1486834041
transform 1 0 12488 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output56
timestamp 1486834041
transform 1 0 12936 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output57
timestamp 1486834041
transform 1 0 12096 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output58
timestamp 1486834041
transform 1 0 13272 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output59
timestamp 1486834041
transform 1 0 12936 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output60
timestamp 1486834041
transform 1 0 12880 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output61
timestamp 1486834041
transform -1 0 14504 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output62
timestamp 1486834041
transform -1 0 14728 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output63
timestamp 1486834041
transform -1 0 15288 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output64
timestamp 1486834041
transform 1 0 14728 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output65
timestamp 1486834041
transform 1 0 15680 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output66
timestamp 1486834041
transform 1 0 15176 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output67
timestamp 1486834041
transform 1 0 16464 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output68
timestamp 1486834041
transform 1 0 16128 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output69
timestamp 1486834041
transform 1 0 15960 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output70
timestamp 1486834041
transform -1 0 16912 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output71
timestamp 1486834041
transform -1 0 17696 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output72
timestamp 1486834041
transform -1 0 17528 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output73
timestamp 1486834041
transform 1 0 17584 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output74
timestamp 1486834041
transform -1 0 21056 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output75
timestamp 1486834041
transform -1 0 20440 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output76
timestamp 1486834041
transform -1 0 20832 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output77
timestamp 1486834041
transform -1 0 21616 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output78
timestamp 1486834041
transform -1 0 20832 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output79
timestamp 1486834041
transform -1 0 21224 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output80
timestamp 1486834041
transform -1 0 18480 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output81
timestamp 1486834041
transform -1 0 17976 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output82
timestamp 1486834041
transform 1 0 18368 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output83
timestamp 1486834041
transform 1 0 18088 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output84
timestamp 1486834041
transform -1 0 19264 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output85
timestamp 1486834041
transform -1 0 18872 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output86
timestamp 1486834041
transform -1 0 20272 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output87
timestamp 1486834041
transform -1 0 19656 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output88
timestamp 1486834041
transform -1 0 19656 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output89
timestamp 1486834041
transform -1 0 22176 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output90
timestamp 1486834041
transform 1 0 24080 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output91
timestamp 1486834041
transform 1 0 23968 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output92
timestamp 1486834041
transform 1 0 23576 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output93
timestamp 1486834041
transform 1 0 23240 0 1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output94
timestamp 1486834041
transform 1 0 24360 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output95
timestamp 1486834041
transform 1 0 24752 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output96
timestamp 1486834041
transform 1 0 21616 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output97
timestamp 1486834041
transform 1 0 20832 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output98
timestamp 1486834041
transform 1 0 22176 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output99
timestamp 1486834041
transform 1 0 22400 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output100
timestamp 1486834041
transform 1 0 21616 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output101
timestamp 1486834041
transform 1 0 22008 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output102
timestamp 1486834041
transform 1 0 23296 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output103
timestamp 1486834041
transform 1 0 22792 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output104
timestamp 1486834041
transform 1 0 22400 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output105
timestamp 1486834041
transform -1 0 1288 0 -1 6664
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_16
timestamp 1486834041
transform 1 0 336 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1486834041
transform -1 0 28392 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_17
timestamp 1486834041
transform 1 0 336 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1486834041
transform -1 0 28392 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_18
timestamp 1486834041
transform 1 0 336 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1486834041
transform -1 0 28392 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_19
timestamp 1486834041
transform 1 0 336 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1486834041
transform -1 0 28392 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_20
timestamp 1486834041
transform 1 0 336 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1486834041
transform -1 0 28392 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_21
timestamp 1486834041
transform 1 0 336 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1486834041
transform -1 0 28392 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_22
timestamp 1486834041
transform 1 0 336 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1486834041
transform -1 0 28392 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_23
timestamp 1486834041
transform 1 0 336 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1486834041
transform -1 0 28392 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_24
timestamp 1486834041
transform 1 0 336 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1486834041
transform -1 0 28392 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_25
timestamp 1486834041
transform 1 0 336 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1486834041
transform -1 0 28392 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_26
timestamp 1486834041
transform 1 0 336 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1486834041
transform -1 0 28392 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_27
timestamp 1486834041
transform 1 0 336 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1486834041
transform -1 0 28392 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_28
timestamp 1486834041
transform 1 0 336 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1486834041
transform -1 0 28392 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_29
timestamp 1486834041
transform 1 0 336 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1486834041
transform -1 0 28392 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_30
timestamp 1486834041
transform 1 0 336 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1486834041
transform -1 0 28392 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_31
timestamp 1486834041
transform 1 0 336 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1486834041
transform -1 0 28392 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_32
timestamp 1486834041
transform 1 0 2240 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_33
timestamp 1486834041
transform 1 0 4144 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_34
timestamp 1486834041
transform 1 0 6048 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_35
timestamp 1486834041
transform 1 0 7952 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_36
timestamp 1486834041
transform 1 0 9856 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_37
timestamp 1486834041
transform 1 0 11760 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_38
timestamp 1486834041
transform 1 0 13664 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_39
timestamp 1486834041
transform 1 0 15568 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_40
timestamp 1486834041
transform 1 0 17472 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_41
timestamp 1486834041
transform 1 0 19376 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_42
timestamp 1486834041
transform 1 0 21280 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_43
timestamp 1486834041
transform 1 0 23184 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_44
timestamp 1486834041
transform 1 0 25088 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_45
timestamp 1486834041
transform 1 0 26992 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_46
timestamp 1486834041
transform 1 0 4256 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_47
timestamp 1486834041
transform 1 0 8176 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_48
timestamp 1486834041
transform 1 0 12096 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_49
timestamp 1486834041
transform 1 0 16016 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_50
timestamp 1486834041
transform 1 0 19936 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_51
timestamp 1486834041
transform 1 0 23856 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_52
timestamp 1486834041
transform 1 0 27776 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_53
timestamp 1486834041
transform 1 0 2296 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_54
timestamp 1486834041
transform 1 0 6216 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_55
timestamp 1486834041
transform 1 0 10136 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_56
timestamp 1486834041
transform 1 0 14056 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_57
timestamp 1486834041
transform 1 0 17976 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_58
timestamp 1486834041
transform 1 0 21896 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_59
timestamp 1486834041
transform 1 0 25816 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_60
timestamp 1486834041
transform 1 0 4256 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_61
timestamp 1486834041
transform 1 0 8176 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_62
timestamp 1486834041
transform 1 0 12096 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_63
timestamp 1486834041
transform 1 0 16016 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_64
timestamp 1486834041
transform 1 0 19936 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_65
timestamp 1486834041
transform 1 0 23856 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_66
timestamp 1486834041
transform 1 0 27776 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_67
timestamp 1486834041
transform 1 0 2296 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_68
timestamp 1486834041
transform 1 0 6216 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_69
timestamp 1486834041
transform 1 0 10136 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_70
timestamp 1486834041
transform 1 0 14056 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_71
timestamp 1486834041
transform 1 0 17976 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_72
timestamp 1486834041
transform 1 0 21896 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_73
timestamp 1486834041
transform 1 0 25816 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_74
timestamp 1486834041
transform 1 0 4256 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_75
timestamp 1486834041
transform 1 0 8176 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_76
timestamp 1486834041
transform 1 0 12096 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_77
timestamp 1486834041
transform 1 0 16016 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_78
timestamp 1486834041
transform 1 0 19936 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_79
timestamp 1486834041
transform 1 0 23856 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_80
timestamp 1486834041
transform 1 0 27776 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_81
timestamp 1486834041
transform 1 0 2296 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_82
timestamp 1486834041
transform 1 0 6216 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_83
timestamp 1486834041
transform 1 0 10136 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_84
timestamp 1486834041
transform 1 0 14056 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_85
timestamp 1486834041
transform 1 0 17976 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_86
timestamp 1486834041
transform 1 0 21896 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_87
timestamp 1486834041
transform 1 0 25816 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_88
timestamp 1486834041
transform 1 0 4256 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_89
timestamp 1486834041
transform 1 0 8176 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_90
timestamp 1486834041
transform 1 0 12096 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_91
timestamp 1486834041
transform 1 0 16016 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_92
timestamp 1486834041
transform 1 0 19936 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_93
timestamp 1486834041
transform 1 0 23856 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_94
timestamp 1486834041
transform 1 0 27776 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_95
timestamp 1486834041
transform 1 0 2296 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_96
timestamp 1486834041
transform 1 0 6216 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_97
timestamp 1486834041
transform 1 0 10136 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_98
timestamp 1486834041
transform 1 0 14056 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_99
timestamp 1486834041
transform 1 0 17976 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_100
timestamp 1486834041
transform 1 0 21896 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_101
timestamp 1486834041
transform 1 0 25816 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_102
timestamp 1486834041
transform 1 0 4256 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_103
timestamp 1486834041
transform 1 0 8176 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_104
timestamp 1486834041
transform 1 0 12096 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_105
timestamp 1486834041
transform 1 0 16016 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_106
timestamp 1486834041
transform 1 0 19936 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_107
timestamp 1486834041
transform 1 0 23856 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_108
timestamp 1486834041
transform 1 0 27776 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_109
timestamp 1486834041
transform 1 0 2296 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_110
timestamp 1486834041
transform 1 0 6216 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_111
timestamp 1486834041
transform 1 0 10136 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_112
timestamp 1486834041
transform 1 0 14056 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_113
timestamp 1486834041
transform 1 0 17976 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_114
timestamp 1486834041
transform 1 0 21896 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_115
timestamp 1486834041
transform 1 0 25816 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_116
timestamp 1486834041
transform 1 0 4256 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_117
timestamp 1486834041
transform 1 0 8176 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_118
timestamp 1486834041
transform 1 0 12096 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_119
timestamp 1486834041
transform 1 0 16016 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_120
timestamp 1486834041
transform 1 0 19936 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_121
timestamp 1486834041
transform 1 0 23856 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_122
timestamp 1486834041
transform 1 0 27776 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_123
timestamp 1486834041
transform 1 0 2296 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_124
timestamp 1486834041
transform 1 0 6216 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_125
timestamp 1486834041
transform 1 0 10136 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_126
timestamp 1486834041
transform 1 0 14056 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_127
timestamp 1486834041
transform 1 0 17976 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_128
timestamp 1486834041
transform 1 0 21896 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_129
timestamp 1486834041
transform 1 0 25816 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_130
timestamp 1486834041
transform 1 0 4256 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_131
timestamp 1486834041
transform 1 0 8176 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_132
timestamp 1486834041
transform 1 0 12096 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_133
timestamp 1486834041
transform 1 0 16016 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_134
timestamp 1486834041
transform 1 0 19936 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_135
timestamp 1486834041
transform 1 0 23856 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_136
timestamp 1486834041
transform 1 0 27776 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_137
timestamp 1486834041
transform 1 0 2296 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_138
timestamp 1486834041
transform 1 0 6216 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_139
timestamp 1486834041
transform 1 0 10136 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_140
timestamp 1486834041
transform 1 0 14056 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_141
timestamp 1486834041
transform 1 0 17976 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_142
timestamp 1486834041
transform 1 0 21896 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_143
timestamp 1486834041
transform 1 0 25816 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_144
timestamp 1486834041
transform 1 0 2240 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_145
timestamp 1486834041
transform 1 0 4144 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_146
timestamp 1486834041
transform 1 0 6048 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_147
timestamp 1486834041
transform 1 0 7952 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_148
timestamp 1486834041
transform 1 0 9856 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_149
timestamp 1486834041
transform 1 0 11760 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_150
timestamp 1486834041
transform 1 0 13664 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_151
timestamp 1486834041
transform 1 0 15568 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_152
timestamp 1486834041
transform 1 0 17472 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_153
timestamp 1486834041
transform 1 0 19376 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_154
timestamp 1486834041
transform 1 0 21280 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_155
timestamp 1486834041
transform 1 0 23184 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_156
timestamp 1486834041
transform 1 0 25088 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_157
timestamp 1486834041
transform 1 0 26992 0 -1 6664
box -43 -43 155 435
<< labels >>
flabel metal2 s 11984 0 12040 56 0 FreeSans 224 0 0 0 Ci
port 0 nsew signal input
flabel metal3 s 0 0 56 56 0 FreeSans 224 0 0 0 FrameData[0]
port 1 nsew signal input
flabel metal3 s 0 2240 56 2296 0 FreeSans 224 0 0 0 FrameData[10]
port 2 nsew signal input
flabel metal3 s 0 2464 56 2520 0 FreeSans 224 0 0 0 FrameData[11]
port 3 nsew signal input
flabel metal3 s 0 2688 56 2744 0 FreeSans 224 0 0 0 FrameData[12]
port 4 nsew signal input
flabel metal3 s 0 2912 56 2968 0 FreeSans 224 0 0 0 FrameData[13]
port 5 nsew signal input
flabel metal3 s 0 3136 56 3192 0 FreeSans 224 0 0 0 FrameData[14]
port 6 nsew signal input
flabel metal3 s 0 3360 56 3416 0 FreeSans 224 0 0 0 FrameData[15]
port 7 nsew signal input
flabel metal3 s 0 3584 56 3640 0 FreeSans 224 0 0 0 FrameData[16]
port 8 nsew signal input
flabel metal3 s 0 3808 56 3864 0 FreeSans 224 0 0 0 FrameData[17]
port 9 nsew signal input
flabel metal3 s 0 4032 56 4088 0 FreeSans 224 0 0 0 FrameData[18]
port 10 nsew signal input
flabel metal3 s 0 4256 56 4312 0 FreeSans 224 0 0 0 FrameData[19]
port 11 nsew signal input
flabel metal3 s 0 224 56 280 0 FreeSans 224 0 0 0 FrameData[1]
port 12 nsew signal input
flabel metal3 s 0 4480 56 4536 0 FreeSans 224 0 0 0 FrameData[20]
port 13 nsew signal input
flabel metal3 s 0 4704 56 4760 0 FreeSans 224 0 0 0 FrameData[21]
port 14 nsew signal input
flabel metal3 s 0 4928 56 4984 0 FreeSans 224 0 0 0 FrameData[22]
port 15 nsew signal input
flabel metal3 s 0 5152 56 5208 0 FreeSans 224 0 0 0 FrameData[23]
port 16 nsew signal input
flabel metal3 s 0 5376 56 5432 0 FreeSans 224 0 0 0 FrameData[24]
port 17 nsew signal input
flabel metal3 s 0 5600 56 5656 0 FreeSans 224 0 0 0 FrameData[25]
port 18 nsew signal input
flabel metal3 s 0 5824 56 5880 0 FreeSans 224 0 0 0 FrameData[26]
port 19 nsew signal input
flabel metal3 s 0 6048 56 6104 0 FreeSans 224 0 0 0 FrameData[27]
port 20 nsew signal input
flabel metal3 s 0 6272 56 6328 0 FreeSans 224 0 0 0 FrameData[28]
port 21 nsew signal input
flabel metal3 s 0 6496 56 6552 0 FreeSans 224 0 0 0 FrameData[29]
port 22 nsew signal input
flabel metal3 s 0 448 56 504 0 FreeSans 224 0 0 0 FrameData[2]
port 23 nsew signal input
flabel metal3 s 0 6720 56 6776 0 FreeSans 224 0 0 0 FrameData[30]
port 24 nsew signal input
flabel metal3 s 0 6944 56 7000 0 FreeSans 224 0 0 0 FrameData[31]
port 25 nsew signal input
flabel metal3 s 0 672 56 728 0 FreeSans 224 0 0 0 FrameData[3]
port 26 nsew signal input
flabel metal3 s 0 896 56 952 0 FreeSans 224 0 0 0 FrameData[4]
port 27 nsew signal input
flabel metal3 s 0 1120 56 1176 0 FreeSans 224 0 0 0 FrameData[5]
port 28 nsew signal input
flabel metal3 s 0 1344 56 1400 0 FreeSans 224 0 0 0 FrameData[6]
port 29 nsew signal input
flabel metal3 s 0 1568 56 1624 0 FreeSans 224 0 0 0 FrameData[7]
port 30 nsew signal input
flabel metal3 s 0 1792 56 1848 0 FreeSans 224 0 0 0 FrameData[8]
port 31 nsew signal input
flabel metal3 s 0 2016 56 2072 0 FreeSans 224 0 0 0 FrameData[9]
port 32 nsew signal input
flabel metal3 s 28672 0 28728 56 0 FreeSans 224 0 0 0 FrameData_O[0]
port 33 nsew signal output
flabel metal3 s 28672 2240 28728 2296 0 FreeSans 224 0 0 0 FrameData_O[10]
port 34 nsew signal output
flabel metal3 s 28672 2464 28728 2520 0 FreeSans 224 0 0 0 FrameData_O[11]
port 35 nsew signal output
flabel metal3 s 28672 2688 28728 2744 0 FreeSans 224 0 0 0 FrameData_O[12]
port 36 nsew signal output
flabel metal3 s 28672 2912 28728 2968 0 FreeSans 224 0 0 0 FrameData_O[13]
port 37 nsew signal output
flabel metal3 s 28672 3136 28728 3192 0 FreeSans 224 0 0 0 FrameData_O[14]
port 38 nsew signal output
flabel metal3 s 28672 3360 28728 3416 0 FreeSans 224 0 0 0 FrameData_O[15]
port 39 nsew signal output
flabel metal3 s 28672 3584 28728 3640 0 FreeSans 224 0 0 0 FrameData_O[16]
port 40 nsew signal output
flabel metal3 s 28672 3808 28728 3864 0 FreeSans 224 0 0 0 FrameData_O[17]
port 41 nsew signal output
flabel metal3 s 28672 4032 28728 4088 0 FreeSans 224 0 0 0 FrameData_O[18]
port 42 nsew signal output
flabel metal3 s 28672 4256 28728 4312 0 FreeSans 224 0 0 0 FrameData_O[19]
port 43 nsew signal output
flabel metal3 s 28672 224 28728 280 0 FreeSans 224 0 0 0 FrameData_O[1]
port 44 nsew signal output
flabel metal3 s 28672 4480 28728 4536 0 FreeSans 224 0 0 0 FrameData_O[20]
port 45 nsew signal output
flabel metal3 s 28672 4704 28728 4760 0 FreeSans 224 0 0 0 FrameData_O[21]
port 46 nsew signal output
flabel metal3 s 28672 4928 28728 4984 0 FreeSans 224 0 0 0 FrameData_O[22]
port 47 nsew signal output
flabel metal3 s 28672 5152 28728 5208 0 FreeSans 224 0 0 0 FrameData_O[23]
port 48 nsew signal output
flabel metal3 s 28672 5376 28728 5432 0 FreeSans 224 0 0 0 FrameData_O[24]
port 49 nsew signal output
flabel metal3 s 28672 5600 28728 5656 0 FreeSans 224 0 0 0 FrameData_O[25]
port 50 nsew signal output
flabel metal3 s 28672 5824 28728 5880 0 FreeSans 224 0 0 0 FrameData_O[26]
port 51 nsew signal output
flabel metal3 s 28672 6048 28728 6104 0 FreeSans 224 0 0 0 FrameData_O[27]
port 52 nsew signal output
flabel metal3 s 28672 6272 28728 6328 0 FreeSans 224 0 0 0 FrameData_O[28]
port 53 nsew signal output
flabel metal3 s 28672 6496 28728 6552 0 FreeSans 224 0 0 0 FrameData_O[29]
port 54 nsew signal output
flabel metal3 s 28672 448 28728 504 0 FreeSans 224 0 0 0 FrameData_O[2]
port 55 nsew signal output
flabel metal3 s 28672 6720 28728 6776 0 FreeSans 224 0 0 0 FrameData_O[30]
port 56 nsew signal output
flabel metal3 s 28672 6944 28728 7000 0 FreeSans 224 0 0 0 FrameData_O[31]
port 57 nsew signal output
flabel metal3 s 28672 672 28728 728 0 FreeSans 224 0 0 0 FrameData_O[3]
port 58 nsew signal output
flabel metal3 s 28672 896 28728 952 0 FreeSans 224 0 0 0 FrameData_O[4]
port 59 nsew signal output
flabel metal3 s 28672 1120 28728 1176 0 FreeSans 224 0 0 0 FrameData_O[5]
port 60 nsew signal output
flabel metal3 s 28672 1344 28728 1400 0 FreeSans 224 0 0 0 FrameData_O[6]
port 61 nsew signal output
flabel metal3 s 28672 1568 28728 1624 0 FreeSans 224 0 0 0 FrameData_O[7]
port 62 nsew signal output
flabel metal3 s 28672 1792 28728 1848 0 FreeSans 224 0 0 0 FrameData_O[8]
port 63 nsew signal output
flabel metal3 s 28672 2016 28728 2072 0 FreeSans 224 0 0 0 FrameData_O[9]
port 64 nsew signal output
flabel metal2 s 24080 0 24136 56 0 FreeSans 224 0 0 0 FrameStrobe[0]
port 65 nsew signal input
flabel metal2 s 26320 0 26376 56 0 FreeSans 224 0 0 0 FrameStrobe[10]
port 66 nsew signal input
flabel metal2 s 26544 0 26600 56 0 FreeSans 224 0 0 0 FrameStrobe[11]
port 67 nsew signal input
flabel metal2 s 26768 0 26824 56 0 FreeSans 224 0 0 0 FrameStrobe[12]
port 68 nsew signal input
flabel metal2 s 26992 0 27048 56 0 FreeSans 224 0 0 0 FrameStrobe[13]
port 69 nsew signal input
flabel metal2 s 27216 0 27272 56 0 FreeSans 224 0 0 0 FrameStrobe[14]
port 70 nsew signal input
flabel metal2 s 27440 0 27496 56 0 FreeSans 224 0 0 0 FrameStrobe[15]
port 71 nsew signal input
flabel metal2 s 27664 0 27720 56 0 FreeSans 224 0 0 0 FrameStrobe[16]
port 72 nsew signal input
flabel metal2 s 27888 0 27944 56 0 FreeSans 224 0 0 0 FrameStrobe[17]
port 73 nsew signal input
flabel metal2 s 28112 0 28168 56 0 FreeSans 224 0 0 0 FrameStrobe[18]
port 74 nsew signal input
flabel metal2 s 28336 0 28392 56 0 FreeSans 224 0 0 0 FrameStrobe[19]
port 75 nsew signal input
flabel metal2 s 24304 0 24360 56 0 FreeSans 224 0 0 0 FrameStrobe[1]
port 76 nsew signal input
flabel metal2 s 24528 0 24584 56 0 FreeSans 224 0 0 0 FrameStrobe[2]
port 77 nsew signal input
flabel metal2 s 24752 0 24808 56 0 FreeSans 224 0 0 0 FrameStrobe[3]
port 78 nsew signal input
flabel metal2 s 24976 0 25032 56 0 FreeSans 224 0 0 0 FrameStrobe[4]
port 79 nsew signal input
flabel metal2 s 25200 0 25256 56 0 FreeSans 224 0 0 0 FrameStrobe[5]
port 80 nsew signal input
flabel metal2 s 25424 0 25480 56 0 FreeSans 224 0 0 0 FrameStrobe[6]
port 81 nsew signal input
flabel metal2 s 25648 0 25704 56 0 FreeSans 224 0 0 0 FrameStrobe[7]
port 82 nsew signal input
flabel metal2 s 25872 0 25928 56 0 FreeSans 224 0 0 0 FrameStrobe[8]
port 83 nsew signal input
flabel metal2 s 26096 0 26152 56 0 FreeSans 224 0 0 0 FrameStrobe[9]
port 84 nsew signal input
flabel metal2 s 2240 7056 2296 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[0]
port 85 nsew signal output
flabel metal2 s 15680 7056 15736 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[10]
port 86 nsew signal output
flabel metal2 s 17024 7056 17080 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[11]
port 87 nsew signal output
flabel metal2 s 18368 7056 18424 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[12]
port 88 nsew signal output
flabel metal2 s 19712 7056 19768 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[13]
port 89 nsew signal output
flabel metal2 s 21056 7056 21112 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[14]
port 90 nsew signal output
flabel metal2 s 22400 7056 22456 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[15]
port 91 nsew signal output
flabel metal2 s 23744 7056 23800 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[16]
port 92 nsew signal output
flabel metal2 s 25088 7056 25144 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[17]
port 93 nsew signal output
flabel metal2 s 26432 7056 26488 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[18]
port 94 nsew signal output
flabel metal2 s 27776 7056 27832 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[19]
port 95 nsew signal output
flabel metal2 s 3584 7056 3640 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[1]
port 96 nsew signal output
flabel metal2 s 4928 7056 4984 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[2]
port 97 nsew signal output
flabel metal2 s 6272 7056 6328 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[3]
port 98 nsew signal output
flabel metal2 s 7616 7056 7672 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[4]
port 99 nsew signal output
flabel metal2 s 8960 7056 9016 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[5]
port 100 nsew signal output
flabel metal2 s 10304 7056 10360 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[6]
port 101 nsew signal output
flabel metal2 s 11648 7056 11704 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[7]
port 102 nsew signal output
flabel metal2 s 12992 7056 13048 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[8]
port 103 nsew signal output
flabel metal2 s 14336 7056 14392 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[9]
port 104 nsew signal output
flabel metal2 s 336 0 392 56 0 FreeSans 224 0 0 0 N1END[0]
port 105 nsew signal input
flabel metal2 s 560 0 616 56 0 FreeSans 224 0 0 0 N1END[1]
port 106 nsew signal input
flabel metal2 s 784 0 840 56 0 FreeSans 224 0 0 0 N1END[2]
port 107 nsew signal input
flabel metal2 s 1008 0 1064 56 0 FreeSans 224 0 0 0 N1END[3]
port 108 nsew signal input
flabel metal2 s 3024 0 3080 56 0 FreeSans 224 0 0 0 N2END[0]
port 109 nsew signal input
flabel metal2 s 3248 0 3304 56 0 FreeSans 224 0 0 0 N2END[1]
port 110 nsew signal input
flabel metal2 s 3472 0 3528 56 0 FreeSans 224 0 0 0 N2END[2]
port 111 nsew signal input
flabel metal2 s 3696 0 3752 56 0 FreeSans 224 0 0 0 N2END[3]
port 112 nsew signal input
flabel metal2 s 3920 0 3976 56 0 FreeSans 224 0 0 0 N2END[4]
port 113 nsew signal input
flabel metal2 s 4144 0 4200 56 0 FreeSans 224 0 0 0 N2END[5]
port 114 nsew signal input
flabel metal2 s 4368 0 4424 56 0 FreeSans 224 0 0 0 N2END[6]
port 115 nsew signal input
flabel metal2 s 4592 0 4648 56 0 FreeSans 224 0 0 0 N2END[7]
port 116 nsew signal input
flabel metal2 s 1232 0 1288 56 0 FreeSans 224 0 0 0 N2MID[0]
port 117 nsew signal input
flabel metal2 s 1456 0 1512 56 0 FreeSans 224 0 0 0 N2MID[1]
port 118 nsew signal input
flabel metal2 s 1680 0 1736 56 0 FreeSans 224 0 0 0 N2MID[2]
port 119 nsew signal input
flabel metal2 s 1904 0 1960 56 0 FreeSans 224 0 0 0 N2MID[3]
port 120 nsew signal input
flabel metal2 s 2128 0 2184 56 0 FreeSans 224 0 0 0 N2MID[4]
port 121 nsew signal input
flabel metal2 s 2352 0 2408 56 0 FreeSans 224 0 0 0 N2MID[5]
port 122 nsew signal input
flabel metal2 s 2576 0 2632 56 0 FreeSans 224 0 0 0 N2MID[6]
port 123 nsew signal input
flabel metal2 s 2800 0 2856 56 0 FreeSans 224 0 0 0 N2MID[7]
port 124 nsew signal input
flabel metal2 s 4816 0 4872 56 0 FreeSans 224 0 0 0 N4END[0]
port 125 nsew signal input
flabel metal2 s 7056 0 7112 56 0 FreeSans 224 0 0 0 N4END[10]
port 126 nsew signal input
flabel metal2 s 7280 0 7336 56 0 FreeSans 224 0 0 0 N4END[11]
port 127 nsew signal input
flabel metal2 s 7504 0 7560 56 0 FreeSans 224 0 0 0 N4END[12]
port 128 nsew signal input
flabel metal2 s 7728 0 7784 56 0 FreeSans 224 0 0 0 N4END[13]
port 129 nsew signal input
flabel metal2 s 7952 0 8008 56 0 FreeSans 224 0 0 0 N4END[14]
port 130 nsew signal input
flabel metal2 s 8176 0 8232 56 0 FreeSans 224 0 0 0 N4END[15]
port 131 nsew signal input
flabel metal2 s 5040 0 5096 56 0 FreeSans 224 0 0 0 N4END[1]
port 132 nsew signal input
flabel metal2 s 5264 0 5320 56 0 FreeSans 224 0 0 0 N4END[2]
port 133 nsew signal input
flabel metal2 s 5488 0 5544 56 0 FreeSans 224 0 0 0 N4END[3]
port 134 nsew signal input
flabel metal2 s 5712 0 5768 56 0 FreeSans 224 0 0 0 N4END[4]
port 135 nsew signal input
flabel metal2 s 5936 0 5992 56 0 FreeSans 224 0 0 0 N4END[5]
port 136 nsew signal input
flabel metal2 s 6160 0 6216 56 0 FreeSans 224 0 0 0 N4END[6]
port 137 nsew signal input
flabel metal2 s 6384 0 6440 56 0 FreeSans 224 0 0 0 N4END[7]
port 138 nsew signal input
flabel metal2 s 6608 0 6664 56 0 FreeSans 224 0 0 0 N4END[8]
port 139 nsew signal input
flabel metal2 s 6832 0 6888 56 0 FreeSans 224 0 0 0 N4END[9]
port 140 nsew signal input
flabel metal2 s 8400 0 8456 56 0 FreeSans 224 0 0 0 NN4END[0]
port 141 nsew signal input
flabel metal2 s 10640 0 10696 56 0 FreeSans 224 0 0 0 NN4END[10]
port 142 nsew signal input
flabel metal2 s 10864 0 10920 56 0 FreeSans 224 0 0 0 NN4END[11]
port 143 nsew signal input
flabel metal2 s 11088 0 11144 56 0 FreeSans 224 0 0 0 NN4END[12]
port 144 nsew signal input
flabel metal2 s 11312 0 11368 56 0 FreeSans 224 0 0 0 NN4END[13]
port 145 nsew signal input
flabel metal2 s 11536 0 11592 56 0 FreeSans 224 0 0 0 NN4END[14]
port 146 nsew signal input
flabel metal2 s 11760 0 11816 56 0 FreeSans 224 0 0 0 NN4END[15]
port 147 nsew signal input
flabel metal2 s 8624 0 8680 56 0 FreeSans 224 0 0 0 NN4END[1]
port 148 nsew signal input
flabel metal2 s 8848 0 8904 56 0 FreeSans 224 0 0 0 NN4END[2]
port 149 nsew signal input
flabel metal2 s 9072 0 9128 56 0 FreeSans 224 0 0 0 NN4END[3]
port 150 nsew signal input
flabel metal2 s 9296 0 9352 56 0 FreeSans 224 0 0 0 NN4END[4]
port 151 nsew signal input
flabel metal2 s 9520 0 9576 56 0 FreeSans 224 0 0 0 NN4END[5]
port 152 nsew signal input
flabel metal2 s 9744 0 9800 56 0 FreeSans 224 0 0 0 NN4END[6]
port 153 nsew signal input
flabel metal2 s 9968 0 10024 56 0 FreeSans 224 0 0 0 NN4END[7]
port 154 nsew signal input
flabel metal2 s 10192 0 10248 56 0 FreeSans 224 0 0 0 NN4END[8]
port 155 nsew signal input
flabel metal2 s 10416 0 10472 56 0 FreeSans 224 0 0 0 NN4END[9]
port 156 nsew signal input
flabel metal2 s 12208 0 12264 56 0 FreeSans 224 0 0 0 S1BEG[0]
port 157 nsew signal output
flabel metal2 s 12432 0 12488 56 0 FreeSans 224 0 0 0 S1BEG[1]
port 158 nsew signal output
flabel metal2 s 12656 0 12712 56 0 FreeSans 224 0 0 0 S1BEG[2]
port 159 nsew signal output
flabel metal2 s 12880 0 12936 56 0 FreeSans 224 0 0 0 S1BEG[3]
port 160 nsew signal output
flabel metal2 s 13104 0 13160 56 0 FreeSans 224 0 0 0 S2BEG[0]
port 161 nsew signal output
flabel metal2 s 13328 0 13384 56 0 FreeSans 224 0 0 0 S2BEG[1]
port 162 nsew signal output
flabel metal2 s 13552 0 13608 56 0 FreeSans 224 0 0 0 S2BEG[2]
port 163 nsew signal output
flabel metal2 s 13776 0 13832 56 0 FreeSans 224 0 0 0 S2BEG[3]
port 164 nsew signal output
flabel metal2 s 14000 0 14056 56 0 FreeSans 224 0 0 0 S2BEG[4]
port 165 nsew signal output
flabel metal2 s 14224 0 14280 56 0 FreeSans 224 0 0 0 S2BEG[5]
port 166 nsew signal output
flabel metal2 s 14448 0 14504 56 0 FreeSans 224 0 0 0 S2BEG[6]
port 167 nsew signal output
flabel metal2 s 14672 0 14728 56 0 FreeSans 224 0 0 0 S2BEG[7]
port 168 nsew signal output
flabel metal2 s 14896 0 14952 56 0 FreeSans 224 0 0 0 S2BEGb[0]
port 169 nsew signal output
flabel metal2 s 15120 0 15176 56 0 FreeSans 224 0 0 0 S2BEGb[1]
port 170 nsew signal output
flabel metal2 s 15344 0 15400 56 0 FreeSans 224 0 0 0 S2BEGb[2]
port 171 nsew signal output
flabel metal2 s 15568 0 15624 56 0 FreeSans 224 0 0 0 S2BEGb[3]
port 172 nsew signal output
flabel metal2 s 15792 0 15848 56 0 FreeSans 224 0 0 0 S2BEGb[4]
port 173 nsew signal output
flabel metal2 s 16016 0 16072 56 0 FreeSans 224 0 0 0 S2BEGb[5]
port 174 nsew signal output
flabel metal2 s 16240 0 16296 56 0 FreeSans 224 0 0 0 S2BEGb[6]
port 175 nsew signal output
flabel metal2 s 16464 0 16520 56 0 FreeSans 224 0 0 0 S2BEGb[7]
port 176 nsew signal output
flabel metal2 s 16688 0 16744 56 0 FreeSans 224 0 0 0 S4BEG[0]
port 177 nsew signal output
flabel metal2 s 18928 0 18984 56 0 FreeSans 224 0 0 0 S4BEG[10]
port 178 nsew signal output
flabel metal2 s 19152 0 19208 56 0 FreeSans 224 0 0 0 S4BEG[11]
port 179 nsew signal output
flabel metal2 s 19376 0 19432 56 0 FreeSans 224 0 0 0 S4BEG[12]
port 180 nsew signal output
flabel metal2 s 19600 0 19656 56 0 FreeSans 224 0 0 0 S4BEG[13]
port 181 nsew signal output
flabel metal2 s 19824 0 19880 56 0 FreeSans 224 0 0 0 S4BEG[14]
port 182 nsew signal output
flabel metal2 s 20048 0 20104 56 0 FreeSans 224 0 0 0 S4BEG[15]
port 183 nsew signal output
flabel metal2 s 16912 0 16968 56 0 FreeSans 224 0 0 0 S4BEG[1]
port 184 nsew signal output
flabel metal2 s 17136 0 17192 56 0 FreeSans 224 0 0 0 S4BEG[2]
port 185 nsew signal output
flabel metal2 s 17360 0 17416 56 0 FreeSans 224 0 0 0 S4BEG[3]
port 186 nsew signal output
flabel metal2 s 17584 0 17640 56 0 FreeSans 224 0 0 0 S4BEG[4]
port 187 nsew signal output
flabel metal2 s 17808 0 17864 56 0 FreeSans 224 0 0 0 S4BEG[5]
port 188 nsew signal output
flabel metal2 s 18032 0 18088 56 0 FreeSans 224 0 0 0 S4BEG[6]
port 189 nsew signal output
flabel metal2 s 18256 0 18312 56 0 FreeSans 224 0 0 0 S4BEG[7]
port 190 nsew signal output
flabel metal2 s 18480 0 18536 56 0 FreeSans 224 0 0 0 S4BEG[8]
port 191 nsew signal output
flabel metal2 s 18704 0 18760 56 0 FreeSans 224 0 0 0 S4BEG[9]
port 192 nsew signal output
flabel metal2 s 20272 0 20328 56 0 FreeSans 224 0 0 0 SS4BEG[0]
port 193 nsew signal output
flabel metal2 s 22512 0 22568 56 0 FreeSans 224 0 0 0 SS4BEG[10]
port 194 nsew signal output
flabel metal2 s 22736 0 22792 56 0 FreeSans 224 0 0 0 SS4BEG[11]
port 195 nsew signal output
flabel metal2 s 22960 0 23016 56 0 FreeSans 224 0 0 0 SS4BEG[12]
port 196 nsew signal output
flabel metal2 s 23184 0 23240 56 0 FreeSans 224 0 0 0 SS4BEG[13]
port 197 nsew signal output
flabel metal2 s 23408 0 23464 56 0 FreeSans 224 0 0 0 SS4BEG[14]
port 198 nsew signal output
flabel metal2 s 23632 0 23688 56 0 FreeSans 224 0 0 0 SS4BEG[15]
port 199 nsew signal output
flabel metal2 s 20496 0 20552 56 0 FreeSans 224 0 0 0 SS4BEG[1]
port 200 nsew signal output
flabel metal2 s 20720 0 20776 56 0 FreeSans 224 0 0 0 SS4BEG[2]
port 201 nsew signal output
flabel metal2 s 20944 0 21000 56 0 FreeSans 224 0 0 0 SS4BEG[3]
port 202 nsew signal output
flabel metal2 s 21168 0 21224 56 0 FreeSans 224 0 0 0 SS4BEG[4]
port 203 nsew signal output
flabel metal2 s 21392 0 21448 56 0 FreeSans 224 0 0 0 SS4BEG[5]
port 204 nsew signal output
flabel metal2 s 21616 0 21672 56 0 FreeSans 224 0 0 0 SS4BEG[6]
port 205 nsew signal output
flabel metal2 s 21840 0 21896 56 0 FreeSans 224 0 0 0 SS4BEG[7]
port 206 nsew signal output
flabel metal2 s 22064 0 22120 56 0 FreeSans 224 0 0 0 SS4BEG[8]
port 207 nsew signal output
flabel metal2 s 22288 0 22344 56 0 FreeSans 224 0 0 0 SS4BEG[9]
port 208 nsew signal output
flabel metal2 s 23856 0 23912 56 0 FreeSans 224 0 0 0 UserCLK
port 209 nsew signal input
flabel metal2 s 896 7056 952 7112 0 FreeSans 224 0 0 0 UserCLKo
port 210 nsew signal output
flabel metal4 s 1888 0 2048 7112 0 FreeSans 736 90 0 0 VDD
port 211 nsew power bidirectional
flabel metal4 s 1888 0 2048 28 0 FreeSans 184 0 0 0 VDD
port 211 nsew power bidirectional
flabel metal4 s 1888 7084 2048 7112 0 FreeSans 184 0 0 0 VDD
port 211 nsew power bidirectional
flabel metal4 s 11888 0 12048 7112 0 FreeSans 736 90 0 0 VDD
port 211 nsew power bidirectional
flabel metal4 s 11888 0 12048 28 0 FreeSans 184 0 0 0 VDD
port 211 nsew power bidirectional
flabel metal4 s 11888 7084 12048 7112 0 FreeSans 184 0 0 0 VDD
port 211 nsew power bidirectional
flabel metal4 s 21888 0 22048 7112 0 FreeSans 736 90 0 0 VDD
port 211 nsew power bidirectional
flabel metal4 s 21888 0 22048 28 0 FreeSans 184 0 0 0 VDD
port 211 nsew power bidirectional
flabel metal4 s 21888 7084 22048 7112 0 FreeSans 184 0 0 0 VDD
port 211 nsew power bidirectional
flabel metal4 s 2218 0 2378 7112 0 FreeSans 736 90 0 0 VSS
port 212 nsew ground bidirectional
flabel metal4 s 2218 0 2378 28 0 FreeSans 184 0 0 0 VSS
port 212 nsew ground bidirectional
flabel metal4 s 2218 7084 2378 7112 0 FreeSans 184 0 0 0 VSS
port 212 nsew ground bidirectional
flabel metal4 s 12218 0 12378 7112 0 FreeSans 736 90 0 0 VSS
port 212 nsew ground bidirectional
flabel metal4 s 12218 0 12378 28 0 FreeSans 184 0 0 0 VSS
port 212 nsew ground bidirectional
flabel metal4 s 12218 7084 12378 7112 0 FreeSans 184 0 0 0 VSS
port 212 nsew ground bidirectional
flabel metal4 s 22218 0 22378 7112 0 FreeSans 736 90 0 0 VSS
port 212 nsew ground bidirectional
flabel metal4 s 22218 0 22378 28 0 FreeSans 184 0 0 0 VSS
port 212 nsew ground bidirectional
flabel metal4 s 22218 7084 22378 7112 0 FreeSans 184 0 0 0 VSS
port 212 nsew ground bidirectional
rlabel metal1 14364 6272 14364 6272 0 VDD
rlabel metal1 14364 6664 14364 6664 0 VSS
rlabel metal3 259 28 259 28 0 FrameData[0]
rlabel metal3 1743 2268 1743 2268 0 FrameData[10]
rlabel metal3 11760 1036 11760 1036 0 FrameData[11]
rlabel metal3 63 2716 63 2716 0 FrameData[12]
rlabel metal3 1743 2940 1743 2940 0 FrameData[13]
rlabel metal3 119 3164 119 3164 0 FrameData[14]
rlabel metal3 399 3388 399 3388 0 FrameData[15]
rlabel metal3 1071 3612 1071 3612 0 FrameData[16]
rlabel metal2 10920 2268 10920 2268 0 FrameData[17]
rlabel metal2 10276 3500 10276 3500 0 FrameData[18]
rlabel metal2 11900 3556 11900 3556 0 FrameData[19]
rlabel metal2 14812 1064 14812 1064 0 FrameData[1]
rlabel metal2 14364 3346 14364 3346 0 FrameData[20]
rlabel metal3 11172 4172 11172 4172 0 FrameData[21]
rlabel metal3 2380 3724 2380 3724 0 FrameData[22]
rlabel metal3 427 5180 427 5180 0 FrameData[23]
rlabel metal3 11816 3780 11816 3780 0 FrameData[24]
rlabel metal3 1715 5628 1715 5628 0 FrameData[25]
rlabel metal3 1071 5852 1071 5852 0 FrameData[26]
rlabel metal3 231 6076 231 6076 0 FrameData[27]
rlabel metal3 931 6300 931 6300 0 FrameData[28]
rlabel metal3 427 6524 427 6524 0 FrameData[29]
rlabel metal3 175 476 175 476 0 FrameData[2]
rlabel metal2 11564 6440 11564 6440 0 FrameData[30]
rlabel metal3 11620 2380 11620 2380 0 FrameData[31]
rlabel metal3 1491 700 1491 700 0 FrameData[3]
rlabel metal3 567 924 567 924 0 FrameData[4]
rlabel metal3 1071 1148 1071 1148 0 FrameData[5]
rlabel metal3 287 1372 287 1372 0 FrameData[6]
rlabel metal3 203 1596 203 1596 0 FrameData[7]
rlabel metal3 1799 1820 1799 1820 0 FrameData[8]
rlabel metal3 2191 2044 2191 2044 0 FrameData[9]
rlabel metal3 28609 28 28609 28 0 FrameData_O[0]
rlabel metal3 27993 2268 27993 2268 0 FrameData_O[10]
rlabel metal3 27594 2548 27594 2548 0 FrameData_O[11]
rlabel metal2 28084 2492 28084 2492 0 FrameData_O[12]
rlabel metal2 27300 2968 27300 2968 0 FrameData_O[13]
rlabel metal2 27580 3192 27580 3192 0 FrameData_O[14]
rlabel metal2 28084 3220 28084 3220 0 FrameData_O[15]
rlabel metal2 27300 3696 27300 3696 0 FrameData_O[16]
rlabel metal3 28385 3836 28385 3836 0 FrameData_O[17]
rlabel metal3 28329 4060 28329 4060 0 FrameData_O[18]
rlabel metal2 27188 4368 27188 4368 0 FrameData_O[19]
rlabel metal3 28581 252 28581 252 0 FrameData_O[1]
rlabel metal3 28385 4508 28385 4508 0 FrameData_O[20]
rlabel metal2 27580 4760 27580 4760 0 FrameData_O[21]
rlabel metal2 27300 5208 27300 5208 0 FrameData_O[22]
rlabel metal3 28329 5180 28329 5180 0 FrameData_O[23]
rlabel metal2 27580 5488 27580 5488 0 FrameData_O[24]
rlabel metal3 28385 5628 28385 5628 0 FrameData_O[25]
rlabel metal3 27454 6020 27454 6020 0 FrameData_O[26]
rlabel metal2 26796 5544 26796 5544 0 FrameData_O[27]
rlabel metal2 26516 5432 26516 5432 0 FrameData_O[28]
rlabel metal3 28000 4172 28000 4172 0 FrameData_O[29]
rlabel metal2 26012 560 26012 560 0 FrameData_O[2]
rlabel metal3 28553 6748 28553 6748 0 FrameData_O[30]
rlabel metal3 28441 6972 28441 6972 0 FrameData_O[31]
rlabel metal3 27741 700 27741 700 0 FrameData_O[3]
rlabel metal3 27741 924 27741 924 0 FrameData_O[4]
rlabel metal2 27468 1092 27468 1092 0 FrameData_O[5]
rlabel metal2 28084 1036 28084 1036 0 FrameData_O[6]
rlabel metal2 27300 1540 27300 1540 0 FrameData_O[7]
rlabel metal3 28077 1820 28077 1820 0 FrameData_O[8]
rlabel metal2 28084 1764 28084 1764 0 FrameData_O[9]
rlabel metal2 24108 2121 24108 2121 0 FrameStrobe[0]
rlabel metal2 24444 1736 24444 1736 0 FrameStrobe[10]
rlabel metal2 26572 819 26572 819 0 FrameStrobe[11]
rlabel metal2 26796 315 26796 315 0 FrameStrobe[12]
rlabel metal2 26012 896 26012 896 0 FrameStrobe[13]
rlabel metal3 26684 1820 26684 1820 0 FrameStrobe[14]
rlabel metal3 25032 924 25032 924 0 FrameStrobe[15]
rlabel metal2 25004 1904 25004 1904 0 FrameStrobe[16]
rlabel metal3 26376 2044 26376 2044 0 FrameStrobe[17]
rlabel metal2 26628 2744 26628 2744 0 FrameStrobe[18]
rlabel metal2 25788 1904 25788 1904 0 FrameStrobe[19]
rlabel metal2 24332 847 24332 847 0 FrameStrobe[1]
rlabel metal2 24556 259 24556 259 0 FrameStrobe[2]
rlabel metal2 24780 791 24780 791 0 FrameStrobe[3]
rlabel metal2 25004 427 25004 427 0 FrameStrobe[4]
rlabel metal2 25228 63 25228 63 0 FrameStrobe[5]
rlabel metal2 25452 399 25452 399 0 FrameStrobe[6]
rlabel metal2 25676 847 25676 847 0 FrameStrobe[7]
rlabel metal2 25900 63 25900 63 0 FrameStrobe[8]
rlabel metal2 26124 371 26124 371 0 FrameStrobe[9]
rlabel metal2 2268 7049 2268 7049 0 FrameStrobe_O[0]
rlabel metal2 15932 6580 15932 6580 0 FrameStrobe_O[10]
rlabel metal2 17276 6384 17276 6384 0 FrameStrobe_O[11]
rlabel metal2 18396 6909 18396 6909 0 FrameStrobe_O[12]
rlabel metal2 19740 7049 19740 7049 0 FrameStrobe_O[13]
rlabel metal2 21084 6909 21084 6909 0 FrameStrobe_O[14]
rlabel metal2 22428 7049 22428 7049 0 FrameStrobe_O[15]
rlabel metal2 23772 7049 23772 7049 0 FrameStrobe_O[16]
rlabel metal2 25116 7049 25116 7049 0 FrameStrobe_O[17]
rlabel metal2 26460 6825 26460 6825 0 FrameStrobe_O[18]
rlabel metal2 27804 6629 27804 6629 0 FrameStrobe_O[19]
rlabel metal2 3612 6741 3612 6741 0 FrameStrobe_O[1]
rlabel metal2 4956 7049 4956 7049 0 FrameStrobe_O[2]
rlabel metal2 6300 7049 6300 7049 0 FrameStrobe_O[3]
rlabel metal2 7868 6356 7868 6356 0 FrameStrobe_O[4]
rlabel metal2 8988 7049 8988 7049 0 FrameStrobe_O[5]
rlabel metal2 10332 6909 10332 6909 0 FrameStrobe_O[6]
rlabel metal2 11676 6909 11676 6909 0 FrameStrobe_O[7]
rlabel metal2 13020 6741 13020 6741 0 FrameStrobe_O[8]
rlabel metal2 14364 6741 14364 6741 0 FrameStrobe_O[9]
rlabel metal2 364 1463 364 1463 0 N1END[0]
rlabel metal2 588 427 588 427 0 N1END[1]
rlabel metal2 812 679 812 679 0 N1END[2]
rlabel metal2 1036 1435 1036 1435 0 N1END[3]
rlabel metal2 3052 1379 3052 1379 0 N2END[0]
rlabel metal2 3276 259 3276 259 0 N2END[1]
rlabel metal2 12180 3724 12180 3724 0 N2END[2]
rlabel metal2 3724 735 3724 735 0 N2END[3]
rlabel metal2 3948 539 3948 539 0 N2END[4]
rlabel metal2 4172 623 4172 623 0 N2END[5]
rlabel metal2 6748 1260 6748 1260 0 N2END[6]
rlabel metal2 13804 1400 13804 1400 0 N2END[7]
rlabel metal2 1260 427 1260 427 0 N2MID[0]
rlabel metal2 1484 1099 1484 1099 0 N2MID[1]
rlabel metal2 1708 847 1708 847 0 N2MID[2]
rlabel metal2 1932 371 1932 371 0 N2MID[3]
rlabel metal2 2156 399 2156 399 0 N2MID[4]
rlabel metal2 2380 175 2380 175 0 N2MID[5]
rlabel metal2 2604 427 2604 427 0 N2MID[6]
rlabel metal2 2828 1015 2828 1015 0 N2MID[7]
rlabel metal3 23408 2660 23408 2660 0 N4END[0]
rlabel metal4 11172 5488 11172 5488 0 N4END[10]
rlabel metal3 12572 3360 12572 3360 0 N4END[11]
rlabel metal3 12180 3444 12180 3444 0 N4END[12]
rlabel metal2 12684 1568 12684 1568 0 N4END[13]
rlabel metal2 7980 819 7980 819 0 N4END[14]
rlabel metal2 1148 532 1148 532 0 N4END[15]
rlabel metal2 22260 3052 22260 3052 0 N4END[1]
rlabel metal2 23268 1988 23268 1988 0 N4END[2]
rlabel metal4 10948 3164 10948 3164 0 N4END[3]
rlabel metal2 10724 2156 10724 2156 0 N4END[4]
rlabel metal2 11788 5404 11788 5404 0 N4END[5]
rlabel metal2 12180 4508 12180 4508 0 N4END[6]
rlabel metal2 12068 2800 12068 2800 0 N4END[7]
rlabel metal2 6636 1043 6636 1043 0 N4END[8]
rlabel metal2 11228 308 11228 308 0 N4END[9]
rlabel metal2 1764 1904 1764 1904 0 NN4END[0]
rlabel metal2 10780 812 10780 812 0 NN4END[10]
rlabel metal2 11564 1288 11564 1288 0 NN4END[11]
rlabel metal2 12124 1232 12124 1232 0 NN4END[12]
rlabel metal3 11788 2548 11788 2548 0 NN4END[13]
rlabel metal3 12264 3276 12264 3276 0 NN4END[14]
rlabel metal2 11788 315 11788 315 0 NN4END[15]
rlabel metal3 3276 3612 3276 3612 0 NN4END[1]
rlabel metal3 6300 3612 6300 3612 0 NN4END[2]
rlabel metal2 5516 1232 5516 1232 0 NN4END[3]
rlabel metal3 6272 2548 6272 2548 0 NN4END[4]
rlabel metal2 6412 1372 6412 1372 0 NN4END[5]
rlabel metal2 7588 1792 7588 1792 0 NN4END[6]
rlabel metal3 9632 4060 9632 4060 0 NN4END[7]
rlabel metal2 10220 1043 10220 1043 0 NN4END[8]
rlabel metal3 10304 2548 10304 2548 0 NN4END[9]
rlabel metal2 12236 175 12236 175 0 S1BEG[0]
rlabel metal2 12460 287 12460 287 0 S1BEG[1]
rlabel metal2 12684 259 12684 259 0 S1BEG[2]
rlabel metal2 12908 343 12908 343 0 S1BEG[3]
rlabel metal2 13132 287 13132 287 0 S2BEG[0]
rlabel metal2 13356 287 13356 287 0 S2BEG[1]
rlabel metal2 13580 455 13580 455 0 S2BEG[2]
rlabel metal2 13804 343 13804 343 0 S2BEG[3]
rlabel metal2 14028 483 14028 483 0 S2BEG[4]
rlabel metal2 14252 287 14252 287 0 S2BEG[5]
rlabel metal2 14476 455 14476 455 0 S2BEG[6]
rlabel metal2 14700 259 14700 259 0 S2BEG[7]
rlabel metal2 14924 231 14924 231 0 S2BEGb[0]
rlabel metal2 15148 343 15148 343 0 S2BEGb[1]
rlabel metal2 15372 119 15372 119 0 S2BEGb[2]
rlabel metal2 15596 455 15596 455 0 S2BEGb[3]
rlabel metal2 15820 343 15820 343 0 S2BEGb[4]
rlabel metal2 16044 175 16044 175 0 S2BEGb[5]
rlabel metal2 16268 231 16268 231 0 S2BEGb[6]
rlabel metal2 16492 371 16492 371 0 S2BEGb[7]
rlabel metal2 16716 259 16716 259 0 S4BEG[0]
rlabel metal2 18956 147 18956 147 0 S4BEG[10]
rlabel metal2 19180 203 19180 203 0 S4BEG[11]
rlabel metal2 19404 175 19404 175 0 S4BEG[12]
rlabel metal2 19628 455 19628 455 0 S4BEG[13]
rlabel metal2 19852 427 19852 427 0 S4BEG[14]
rlabel metal2 20076 259 20076 259 0 S4BEG[15]
rlabel metal2 16940 203 16940 203 0 S4BEG[1]
rlabel metal2 17164 427 17164 427 0 S4BEG[2]
rlabel metal2 17388 231 17388 231 0 S4BEG[3]
rlabel metal2 17612 455 17612 455 0 S4BEG[4]
rlabel metal2 17836 119 17836 119 0 S4BEG[5]
rlabel metal2 18060 847 18060 847 0 S4BEG[6]
rlabel metal2 18284 287 18284 287 0 S4BEG[7]
rlabel metal2 18508 567 18508 567 0 S4BEG[8]
rlabel metal2 18732 203 18732 203 0 S4BEG[9]
rlabel metal2 20300 287 20300 287 0 SS4BEG[0]
rlabel metal2 22540 119 22540 119 0 SS4BEG[10]
rlabel metal2 22764 231 22764 231 0 SS4BEG[11]
rlabel metal2 22988 455 22988 455 0 SS4BEG[12]
rlabel metal2 23212 903 23212 903 0 SS4BEG[13]
rlabel metal2 23436 315 23436 315 0 SS4BEG[14]
rlabel metal2 23660 91 23660 91 0 SS4BEG[15]
rlabel metal3 21910 868 21910 868 0 SS4BEG[1]
rlabel metal2 20748 427 20748 427 0 SS4BEG[2]
rlabel metal2 20972 231 20972 231 0 SS4BEG[3]
rlabel metal2 22764 952 22764 952 0 SS4BEG[4]
rlabel metal2 22148 1064 22148 1064 0 SS4BEG[5]
rlabel metal2 22428 1064 22428 1064 0 SS4BEG[6]
rlabel metal2 21868 147 21868 147 0 SS4BEG[7]
rlabel metal2 22092 63 22092 63 0 SS4BEG[8]
rlabel metal2 22316 175 22316 175 0 SS4BEG[9]
rlabel metal2 23884 847 23884 847 0 UserCLK
rlabel metal2 1036 6692 1036 6692 0 UserCLKo
rlabel metal3 12180 1120 12180 1120 0 net1
rlabel metal2 10724 3640 10724 3640 0 net10
rlabel metal3 13580 2352 13580 2352 0 net100
rlabel metal2 21924 3556 21924 3556 0 net101
rlabel metal2 23380 336 23380 336 0 net102
rlabel metal2 11508 3416 11508 3416 0 net103
rlabel metal2 12852 2240 12852 2240 0 net104
rlabel metal3 12278 4172 12278 4172 0 net105
rlabel metal3 26012 4452 26012 4452 0 net11
rlabel metal2 15092 1204 15092 1204 0 net12
rlabel metal2 27636 5544 27636 5544 0 net13
rlabel metal3 12628 4396 12628 4396 0 net14
rlabel metal2 14924 3864 14924 3864 0 net15
rlabel metal2 25284 5208 25284 5208 0 net16
rlabel metal2 27076 5488 27076 5488 0 net17
rlabel metal2 27692 5516 27692 5516 0 net18
rlabel metal3 20664 6076 20664 6076 0 net19
rlabel metal2 23380 3080 23380 3080 0 net2
rlabel metal2 26404 5348 26404 5348 0 net20
rlabel metal2 26068 5236 26068 5236 0 net21
rlabel metal3 21868 3472 21868 3472 0 net22
rlabel metal2 25508 1568 25508 1568 0 net23
rlabel metal4 13412 4844 13412 4844 0 net24
rlabel metal2 25508 5880 25508 5880 0 net25
rlabel metal2 26404 1736 26404 1736 0 net26
rlabel metal2 26320 2100 26320 2100 0 net27
rlabel metal3 26404 1036 26404 1036 0 net28
rlabel metal2 21868 616 21868 616 0 net29
rlabel metal3 22428 4060 22428 4060 0 net3
rlabel metal2 24388 1820 24388 1820 0 net30
rlabel metal2 26236 5180 26236 5180 0 net31
rlabel metal2 27552 1372 27552 1372 0 net32
rlabel metal2 3052 6104 3052 6104 0 net33
rlabel metal2 24164 3220 24164 3220 0 net34
rlabel metal3 18172 6020 18172 6020 0 net35
rlabel metal3 19544 6132 19544 6132 0 net36
rlabel metal2 25620 1736 25620 1736 0 net37
rlabel metal3 25200 5348 25200 5348 0 net38
rlabel metal2 23380 924 23380 924 0 net39
rlabel metal2 27580 2184 27580 2184 0 net4
rlabel metal2 24584 1820 24584 1820 0 net40
rlabel metal3 26124 6468 26124 6468 0 net41
rlabel metal2 26236 6468 26236 6468 0 net42
rlabel metal2 25396 1848 25396 1848 0 net43
rlabel metal2 4060 6664 4060 6664 0 net44
rlabel metal2 5208 6132 5208 6132 0 net45
rlabel metal2 7140 6104 7140 6104 0 net46
rlabel metal3 8736 5740 8736 5740 0 net47
rlabel metal2 10332 6300 10332 6300 0 net48
rlabel metal2 11172 6300 11172 6300 0 net49
rlabel metal2 26796 2996 26796 2996 0 net5
rlabel metal3 12908 6132 12908 6132 0 net50
rlabel metal3 13972 5348 13972 5348 0 net51
rlabel metal2 15148 6048 15148 6048 0 net52
rlabel metal2 11396 1232 11396 1232 0 net53
rlabel metal2 8932 952 8932 952 0 net54
rlabel metal2 12628 1344 12628 1344 0 net55
rlabel metal2 10724 1204 10724 1204 0 net56
rlabel metal2 12180 1400 12180 1400 0 net57
rlabel metal2 13356 1120 13356 1120 0 net58
rlabel metal2 12964 1036 12964 1036 0 net59
rlabel metal3 11844 3192 11844 3192 0 net6
rlabel metal2 13076 896 13076 896 0 net60
rlabel metal2 14420 2618 14420 2618 0 net61
rlabel metal2 14700 588 14700 588 0 net62
rlabel metal2 15204 1792 15204 1792 0 net63
rlabel metal2 14868 1540 14868 1540 0 net64
rlabel metal2 15764 1148 15764 1148 0 net65
rlabel metal2 11508 1568 11508 1568 0 net66
rlabel metal2 12852 756 12852 756 0 net67
rlabel metal2 14644 1176 14644 1176 0 net68
rlabel metal2 15932 1176 15932 1176 0 net69
rlabel metal3 26376 2996 26376 2996 0 net7
rlabel metal2 16716 1932 16716 1932 0 net70
rlabel metal2 17892 1176 17892 1176 0 net71
rlabel metal2 17444 1736 17444 1736 0 net72
rlabel metal3 2240 1036 2240 1036 0 net73
rlabel metal2 20972 672 20972 672 0 net74
rlabel metal2 21868 3248 21868 3248 0 net75
rlabel metal2 22764 1932 22764 1932 0 net76
rlabel metal2 21476 1344 21476 1344 0 net77
rlabel metal2 20804 2576 20804 2576 0 net78
rlabel metal2 23772 2800 23772 2800 0 net79
rlabel metal2 12628 5628 12628 5628 0 net8
rlabel metal3 19012 980 19012 980 0 net80
rlabel metal2 18452 1960 18452 1960 0 net81
rlabel metal2 18592 588 18592 588 0 net82
rlabel metal3 18004 1372 18004 1372 0 net83
rlabel metal2 19040 980 19040 980 0 net84
rlabel metal2 19572 2492 19572 2492 0 net85
rlabel metal2 20048 588 20048 588 0 net86
rlabel metal2 19460 2128 19460 2128 0 net87
rlabel metal3 20272 2212 20272 2212 0 net88
rlabel metal2 22092 672 22092 672 0 net89
rlabel metal3 25284 3892 25284 3892 0 net9
rlabel metal3 13748 504 13748 504 0 net90
rlabel metal3 12180 2800 12180 2800 0 net91
rlabel metal2 23660 1400 23660 1400 0 net92
rlabel metal3 10948 1792 10948 1792 0 net93
rlabel metal2 2716 3612 2716 3612 0 net94
rlabel metal2 1316 1988 1316 1988 0 net95
rlabel metal3 13524 952 13524 952 0 net96
rlabel metal2 12684 3024 12684 3024 0 net97
rlabel metal2 14140 1232 14140 1232 0 net98
rlabel metal2 12516 1456 12516 1456 0 net99
<< properties >>
string FIXED_BBOX 0 0 28728 7112
<< end >>
