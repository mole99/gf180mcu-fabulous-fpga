magic
tech gf180mcuD
magscale 1 5
timestamp 1764324290
<< metal1 >>
rect 336 6677 26040 6694
rect 336 6651 2233 6677
rect 2259 6651 2285 6677
rect 2311 6651 2337 6677
rect 2363 6651 12233 6677
rect 12259 6651 12285 6677
rect 12311 6651 12337 6677
rect 12363 6651 22233 6677
rect 22259 6651 22285 6677
rect 22311 6651 22337 6677
rect 22363 6651 26040 6677
rect 336 6634 26040 6651
rect 19839 6593 19865 6599
rect 905 6567 911 6593
rect 937 6567 943 6593
rect 19839 6561 19865 6567
rect 22135 6593 22161 6599
rect 22135 6561 22161 6567
rect 23647 6593 23673 6599
rect 23647 6561 23673 6567
rect 24599 6593 24625 6599
rect 24599 6561 24625 6567
rect 2641 6511 2647 6537
rect 2673 6511 2679 6537
rect 3033 6511 3039 6537
rect 3065 6511 3071 6537
rect 6449 6511 6455 6537
rect 6481 6511 6487 6537
rect 1079 6481 1105 6487
rect 22807 6481 22833 6487
rect 3985 6455 3991 6481
rect 4017 6455 4023 6481
rect 5217 6455 5223 6481
rect 5249 6455 5255 6481
rect 6841 6455 6847 6481
rect 6873 6455 6879 6481
rect 7681 6455 7687 6481
rect 7713 6455 7719 6481
rect 8913 6455 8919 6481
rect 8945 6455 8951 6481
rect 9753 6455 9759 6481
rect 9785 6455 9791 6481
rect 11265 6455 11271 6481
rect 11297 6455 11303 6481
rect 12497 6455 12503 6481
rect 12529 6455 12535 6481
rect 13449 6455 13455 6481
rect 13481 6455 13487 6481
rect 14961 6455 14967 6481
rect 14993 6455 14999 6481
rect 16361 6455 16367 6481
rect 16393 6455 16399 6481
rect 17369 6455 17375 6481
rect 17401 6455 17407 6481
rect 18769 6455 18775 6481
rect 18801 6455 18807 6481
rect 19553 6455 19559 6481
rect 19585 6455 19591 6481
rect 21065 6455 21071 6481
rect 21097 6455 21103 6481
rect 21849 6455 21855 6481
rect 21881 6455 21887 6481
rect 1079 6449 1105 6455
rect 22807 6449 22833 6455
rect 23087 6481 23113 6487
rect 25271 6481 25297 6487
rect 23361 6455 23367 6481
rect 23393 6455 23399 6481
rect 24369 6455 24375 6481
rect 24401 6455 24407 6481
rect 23087 6449 23113 6455
rect 25271 6449 25297 6455
rect 3487 6425 3513 6431
rect 3487 6393 3513 6399
rect 4719 6425 4745 6431
rect 4719 6393 4745 6399
rect 7183 6425 7209 6431
rect 7183 6393 7209 6399
rect 8415 6425 8441 6431
rect 10879 6425 10905 6431
rect 9417 6399 9423 6425
rect 9449 6399 9455 6425
rect 8415 6393 8441 6399
rect 10879 6393 10905 6399
rect 12111 6425 12137 6431
rect 14575 6425 14601 6431
rect 13113 6399 13119 6425
rect 13145 6399 13151 6425
rect 12111 6393 12137 6399
rect 14575 6393 14601 6399
rect 15863 6425 15889 6431
rect 15863 6393 15889 6399
rect 16871 6425 16897 6431
rect 16871 6393 16897 6399
rect 18271 6425 18297 6431
rect 18271 6393 18297 6399
rect 20679 6425 20705 6431
rect 25489 6399 25495 6425
rect 25521 6399 25527 6425
rect 20679 6393 20705 6399
rect 336 6285 26040 6302
rect 336 6259 1903 6285
rect 1929 6259 1955 6285
rect 1981 6259 2007 6285
rect 2033 6259 11903 6285
rect 11929 6259 11955 6285
rect 11981 6259 12007 6285
rect 12033 6259 21903 6285
rect 21929 6259 21955 6285
rect 21981 6259 22007 6285
rect 22033 6259 26040 6285
rect 336 6242 26040 6259
rect 24039 6201 24065 6207
rect 24039 6169 24065 6175
rect 1359 6145 1385 6151
rect 15247 6145 15273 6151
rect 14849 6119 14855 6145
rect 14881 6119 14887 6145
rect 1359 6113 1385 6119
rect 15247 6113 15273 6119
rect 16591 6145 16617 6151
rect 16591 6113 16617 6119
rect 17039 6145 17065 6151
rect 20847 6145 20873 6151
rect 18825 6119 18831 6145
rect 18857 6119 18863 6145
rect 17039 6113 17065 6119
rect 20847 6113 20873 6119
rect 21295 6145 21321 6151
rect 24823 6145 24849 6151
rect 23025 6119 23031 6145
rect 23057 6119 23063 6145
rect 21295 6113 21321 6119
rect 24823 6113 24849 6119
rect 25607 6145 25633 6151
rect 25607 6113 25633 6119
rect 1129 6063 1135 6089
rect 1161 6063 1167 6089
rect 5049 6063 5055 6089
rect 5081 6063 5087 6089
rect 15017 6063 15023 6089
rect 15049 6063 15055 6089
rect 23305 6063 23311 6089
rect 23337 6063 23343 6089
rect 24369 6063 24375 6089
rect 24401 6063 24407 6089
rect 3767 6033 3793 6039
rect 3767 6001 3793 6007
rect 5279 6033 5305 6039
rect 5279 6001 5305 6007
rect 16871 6033 16897 6039
rect 16871 6001 16897 6007
rect 22359 6033 22385 6039
rect 23529 6007 23535 6033
rect 23561 6007 23567 6033
rect 25097 6007 25103 6033
rect 25129 6007 25135 6033
rect 22359 6001 22385 6007
rect 3487 5977 3513 5983
rect 3487 5945 3513 5951
rect 15527 5977 15553 5983
rect 16255 5977 16281 5983
rect 16081 5951 16087 5977
rect 16113 5951 16119 5977
rect 15527 5945 15553 5951
rect 16255 5945 16281 5951
rect 17319 5977 17345 5983
rect 17319 5945 17345 5951
rect 19055 5977 19081 5983
rect 19055 5945 19081 5951
rect 20567 5977 20593 5983
rect 20567 5945 20593 5951
rect 21015 5977 21041 5983
rect 21015 5945 21041 5951
rect 22079 5977 22105 5983
rect 22079 5945 22105 5951
rect 336 5893 26040 5910
rect 336 5867 2233 5893
rect 2259 5867 2285 5893
rect 2311 5867 2337 5893
rect 2363 5867 12233 5893
rect 12259 5867 12285 5893
rect 12311 5867 12337 5893
rect 12363 5867 22233 5893
rect 22259 5867 22285 5893
rect 22311 5867 22337 5893
rect 22363 5867 26040 5893
rect 336 5850 26040 5867
rect 7799 5809 7825 5815
rect 7799 5777 7825 5783
rect 9087 5809 9113 5815
rect 9087 5777 9113 5783
rect 22695 5809 22721 5815
rect 22695 5777 22721 5783
rect 8807 5753 8833 5759
rect 8807 5721 8833 5727
rect 19055 5753 19081 5759
rect 23137 5727 23143 5753
rect 23169 5727 23175 5753
rect 23529 5727 23535 5753
rect 23561 5727 23567 5753
rect 19055 5721 19081 5727
rect 12727 5697 12753 5703
rect 19273 5671 19279 5697
rect 19305 5671 19311 5697
rect 24481 5671 24487 5697
rect 24513 5671 24519 5697
rect 25265 5671 25271 5697
rect 25297 5671 25303 5697
rect 12727 5665 12753 5671
rect 22975 5641 23001 5647
rect 7569 5615 7575 5641
rect 7601 5615 7607 5641
rect 12497 5615 12503 5641
rect 12529 5615 12535 5641
rect 22975 5609 23001 5615
rect 24935 5641 24961 5647
rect 24935 5609 24961 5615
rect 25719 5585 25745 5591
rect 25719 5553 25745 5559
rect 336 5501 26040 5518
rect 336 5475 1903 5501
rect 1929 5475 1955 5501
rect 1981 5475 2007 5501
rect 2033 5475 11903 5501
rect 11929 5475 11955 5501
rect 11981 5475 12007 5501
rect 12033 5475 21903 5501
rect 21929 5475 21955 5501
rect 21981 5475 22007 5501
rect 22033 5475 26040 5501
rect 336 5458 26040 5475
rect 24039 5417 24065 5423
rect 24039 5385 24065 5391
rect 18719 5361 18745 5367
rect 11209 5335 11215 5361
rect 11241 5335 11247 5361
rect 13393 5335 13399 5361
rect 13425 5335 13431 5361
rect 17649 5335 17655 5361
rect 17681 5335 17687 5361
rect 18719 5329 18745 5335
rect 24823 5361 24849 5367
rect 24823 5329 24849 5335
rect 23087 5305 23113 5311
rect 24369 5279 24375 5305
rect 24401 5279 24407 5305
rect 23087 5273 23113 5279
rect 23367 5249 23393 5255
rect 23529 5223 23535 5249
rect 23561 5223 23567 5249
rect 25097 5223 25103 5249
rect 25129 5223 25135 5249
rect 25489 5223 25495 5249
rect 25521 5223 25527 5249
rect 23367 5217 23393 5223
rect 11439 5193 11465 5199
rect 11439 5161 11465 5167
rect 13623 5193 13649 5199
rect 13623 5161 13649 5167
rect 17879 5193 17905 5199
rect 17879 5161 17905 5167
rect 18999 5193 19025 5199
rect 18999 5161 19025 5167
rect 336 5109 26040 5126
rect 336 5083 2233 5109
rect 2259 5083 2285 5109
rect 2311 5083 2337 5109
rect 2363 5083 12233 5109
rect 12259 5083 12285 5109
rect 12311 5083 12337 5109
rect 12363 5083 22233 5109
rect 22259 5083 22285 5109
rect 22311 5083 22337 5109
rect 22363 5083 26040 5109
rect 336 5066 26040 5083
rect 2871 4969 2897 4975
rect 2871 4937 2897 4943
rect 1079 4913 1105 4919
rect 1079 4881 1105 4887
rect 2591 4913 2617 4919
rect 2591 4881 2617 4887
rect 3487 4913 3513 4919
rect 3487 4881 3513 4887
rect 7799 4913 7825 4919
rect 7799 4881 7825 4887
rect 9647 4913 9673 4919
rect 9647 4881 9673 4887
rect 16479 4913 16505 4919
rect 23759 4913 23785 4919
rect 23529 4887 23535 4913
rect 23561 4887 23567 4913
rect 24425 4887 24431 4913
rect 24457 4887 24463 4913
rect 25209 4887 25215 4913
rect 25241 4887 25247 4913
rect 16479 4881 16505 4887
rect 23759 4881 23785 4887
rect 3767 4857 3793 4863
rect 849 4831 855 4857
rect 881 4831 887 4857
rect 3767 4825 3793 4831
rect 8079 4857 8105 4863
rect 8079 4825 8105 4831
rect 9927 4857 9953 4863
rect 9927 4825 9953 4831
rect 16199 4857 16225 4863
rect 16199 4825 16225 4831
rect 24935 4857 24961 4863
rect 24935 4825 24961 4831
rect 25719 4801 25745 4807
rect 25719 4769 25745 4775
rect 336 4717 26040 4734
rect 336 4691 1903 4717
rect 1929 4691 1955 4717
rect 1981 4691 2007 4717
rect 2033 4691 11903 4717
rect 11929 4691 11955 4717
rect 11981 4691 12007 4717
rect 12033 4691 21903 4717
rect 21929 4691 21955 4717
rect 21981 4691 22007 4717
rect 22033 4691 26040 4717
rect 336 4674 26040 4691
rect 24823 4633 24849 4639
rect 24823 4601 24849 4607
rect 22751 4577 22777 4583
rect 2137 4551 2143 4577
rect 2169 4551 2175 4577
rect 22751 4545 22777 4551
rect 24151 4577 24177 4583
rect 24151 4545 24177 4551
rect 5279 4521 5305 4527
rect 5279 4489 5305 4495
rect 22471 4521 22497 4527
rect 24369 4495 24375 4521
rect 24401 4495 24407 4521
rect 25153 4495 25159 4521
rect 25185 4495 25191 4521
rect 22471 4489 22497 4495
rect 5559 4465 5585 4471
rect 5559 4433 5585 4439
rect 23871 4465 23897 4471
rect 25489 4439 25495 4465
rect 25521 4439 25527 4465
rect 23871 4433 23897 4439
rect 1919 4409 1945 4415
rect 1919 4377 1945 4383
rect 336 4325 26040 4342
rect 336 4299 2233 4325
rect 2259 4299 2285 4325
rect 2311 4299 2337 4325
rect 2363 4299 12233 4325
rect 12259 4299 12285 4325
rect 12311 4299 12337 4325
rect 12363 4299 22233 4325
rect 22259 4299 22285 4325
rect 22311 4299 22337 4325
rect 22363 4299 26040 4325
rect 336 4282 26040 4299
rect 15135 4185 15161 4191
rect 15135 4153 15161 4159
rect 23255 4185 23281 4191
rect 23255 4153 23281 4159
rect 25047 4185 25073 4191
rect 25047 4153 25073 4159
rect 15415 4129 15441 4135
rect 9249 4103 9255 4129
rect 9281 4103 9287 4129
rect 11769 4103 11775 4129
rect 11801 4103 11807 4129
rect 15415 4097 15441 4103
rect 21295 4129 21321 4135
rect 24599 4129 24625 4135
rect 24369 4103 24375 4129
rect 24401 4103 24407 4129
rect 21295 4097 21321 4103
rect 24599 4097 24625 4103
rect 24767 4129 24793 4135
rect 25209 4103 25215 4129
rect 25241 4103 25247 4129
rect 24767 4097 24793 4103
rect 9479 4073 9505 4079
rect 9479 4041 9505 4047
rect 11999 4073 12025 4079
rect 21513 4047 21519 4073
rect 21545 4047 21551 4073
rect 23473 4047 23479 4073
rect 23505 4047 23511 4073
rect 11999 4041 12025 4047
rect 25719 4017 25745 4023
rect 25719 3985 25745 3991
rect 336 3933 26040 3950
rect 336 3907 1903 3933
rect 1929 3907 1955 3933
rect 1981 3907 2007 3933
rect 2033 3907 11903 3933
rect 11929 3907 11955 3933
rect 11981 3907 12007 3933
rect 12033 3907 21903 3933
rect 21929 3907 21955 3933
rect 21981 3907 22007 3933
rect 22033 3907 26040 3933
rect 336 3890 26040 3907
rect 25607 3849 25633 3855
rect 25607 3817 25633 3823
rect 24151 3793 24177 3799
rect 24151 3761 24177 3767
rect 24823 3793 24849 3799
rect 24823 3761 24849 3767
rect 12279 3737 12305 3743
rect 24369 3711 24375 3737
rect 24401 3711 24407 3737
rect 25097 3711 25103 3737
rect 25129 3711 25135 3737
rect 12279 3705 12305 3711
rect 799 3681 825 3687
rect 799 3649 825 3655
rect 2871 3681 2897 3687
rect 2871 3649 2897 3655
rect 4215 3681 4241 3687
rect 4215 3649 4241 3655
rect 11271 3681 11297 3687
rect 11271 3649 11297 3655
rect 12559 3681 12585 3687
rect 12559 3649 12585 3655
rect 23871 3681 23897 3687
rect 23871 3649 23897 3655
rect 1079 3625 1105 3631
rect 1079 3593 1105 3599
rect 3151 3625 3177 3631
rect 3151 3593 3177 3599
rect 4495 3625 4521 3631
rect 4495 3593 4521 3599
rect 10991 3625 11017 3631
rect 10991 3593 11017 3599
rect 336 3541 26040 3558
rect 336 3515 2233 3541
rect 2259 3515 2285 3541
rect 2311 3515 2337 3541
rect 2363 3515 12233 3541
rect 12259 3515 12285 3541
rect 12311 3515 12337 3541
rect 12363 3515 22233 3541
rect 22259 3515 22285 3541
rect 22311 3515 22337 3541
rect 22363 3515 26040 3541
rect 336 3498 26040 3515
rect 16871 3457 16897 3463
rect 16871 3425 16897 3431
rect 4159 3345 4185 3351
rect 13623 3345 13649 3351
rect 7849 3319 7855 3345
rect 7881 3319 7887 3345
rect 8409 3319 8415 3345
rect 8441 3319 8447 3345
rect 4159 3313 4185 3319
rect 13623 3313 13649 3319
rect 15303 3345 15329 3351
rect 21071 3345 21097 3351
rect 17649 3319 17655 3345
rect 17681 3319 17687 3345
rect 15303 3313 15329 3319
rect 21071 3313 21097 3319
rect 22135 3345 22161 3351
rect 24425 3319 24431 3345
rect 24457 3319 24463 3345
rect 25209 3319 25215 3345
rect 25241 3319 25247 3345
rect 22135 3313 22161 3319
rect 8639 3289 8665 3295
rect 15583 3289 15609 3295
rect 3929 3263 3935 3289
rect 3961 3263 3967 3289
rect 8017 3263 8023 3289
rect 8049 3263 8055 3289
rect 13841 3263 13847 3289
rect 13873 3263 13879 3289
rect 8639 3257 8665 3263
rect 15583 3257 15609 3263
rect 17151 3289 17177 3295
rect 17151 3257 17177 3263
rect 17879 3289 17905 3295
rect 25719 3289 25745 3295
rect 21289 3263 21295 3289
rect 21321 3263 21327 3289
rect 22353 3263 22359 3289
rect 22385 3263 22391 3289
rect 24873 3263 24879 3289
rect 24905 3263 24911 3289
rect 17879 3257 17905 3263
rect 25719 3257 25745 3263
rect 336 3149 26040 3166
rect 336 3123 1903 3149
rect 1929 3123 1955 3149
rect 1981 3123 2007 3149
rect 2033 3123 11903 3149
rect 11929 3123 11955 3149
rect 11981 3123 12007 3149
rect 12033 3123 21903 3149
rect 21929 3123 21955 3149
rect 21981 3123 22007 3149
rect 22033 3123 26040 3149
rect 336 3106 26040 3123
rect 25607 3065 25633 3071
rect 25607 3033 25633 3039
rect 17375 3009 17401 3015
rect 849 2983 855 3009
rect 881 2983 887 3009
rect 5889 2983 5895 3009
rect 5921 2983 5927 3009
rect 6449 2983 6455 3009
rect 6481 2983 6487 3009
rect 15801 2983 15807 3009
rect 15833 2983 15839 3009
rect 18825 2983 18831 3009
rect 18857 2983 18863 3009
rect 17375 2977 17401 2983
rect 18607 2953 18633 2959
rect 2529 2927 2535 2953
rect 2561 2927 2567 2953
rect 15129 2927 15135 2953
rect 15161 2927 15167 2953
rect 15633 2927 15639 2953
rect 15665 2927 15671 2953
rect 18607 2921 18633 2927
rect 20511 2953 20537 2959
rect 20511 2921 20537 2927
rect 23143 2953 23169 2959
rect 23143 2921 23169 2927
rect 24207 2953 24233 2959
rect 24207 2921 24233 2927
rect 2759 2897 2785 2903
rect 2759 2865 2785 2871
rect 6119 2897 6145 2903
rect 6119 2865 6145 2871
rect 15359 2897 15385 2903
rect 15359 2865 15385 2871
rect 16311 2897 16337 2903
rect 18439 2897 18465 2903
rect 16473 2871 16479 2897
rect 16505 2871 16511 2897
rect 17873 2871 17879 2897
rect 17905 2871 17911 2897
rect 16311 2865 16337 2871
rect 18439 2865 18465 2871
rect 19335 2897 19361 2903
rect 19335 2865 19361 2871
rect 20791 2897 20817 2903
rect 20791 2865 20817 2871
rect 23423 2897 23449 2903
rect 23423 2865 23449 2871
rect 23591 2897 23617 2903
rect 23591 2865 23617 2871
rect 23871 2897 23897 2903
rect 23871 2865 23897 2871
rect 24487 2897 24513 2903
rect 24487 2865 24513 2871
rect 24935 2897 24961 2903
rect 25097 2871 25103 2897
rect 25129 2871 25135 2897
rect 24935 2865 24961 2871
rect 1079 2841 1105 2847
rect 1079 2809 1105 2815
rect 6679 2841 6705 2847
rect 6679 2809 6705 2815
rect 16031 2841 16057 2847
rect 16031 2809 16057 2815
rect 16759 2841 16785 2847
rect 16759 2809 16785 2815
rect 18159 2841 18185 2847
rect 18159 2809 18185 2815
rect 19055 2841 19081 2847
rect 19055 2809 19081 2815
rect 24655 2841 24681 2847
rect 24655 2809 24681 2815
rect 336 2757 26040 2774
rect 336 2731 2233 2757
rect 2259 2731 2285 2757
rect 2311 2731 2337 2757
rect 2363 2731 12233 2757
rect 12259 2731 12285 2757
rect 12311 2731 12337 2757
rect 12363 2731 22233 2757
rect 22259 2731 22285 2757
rect 22311 2731 22337 2757
rect 22363 2731 26040 2757
rect 336 2714 26040 2731
rect 12783 2673 12809 2679
rect 12783 2641 12809 2647
rect 2143 2617 2169 2623
rect 2143 2585 2169 2591
rect 7071 2617 7097 2623
rect 20399 2617 20425 2623
rect 15241 2591 15247 2617
rect 15273 2591 15279 2617
rect 17593 2591 17599 2617
rect 17625 2591 17631 2617
rect 18377 2591 18383 2617
rect 18409 2591 18415 2617
rect 19161 2591 19167 2617
rect 19193 2591 19199 2617
rect 25209 2591 25215 2617
rect 25241 2591 25247 2617
rect 25601 2591 25607 2617
rect 25633 2591 25639 2617
rect 7071 2585 7097 2591
rect 20399 2585 20425 2591
rect 2423 2561 2449 2567
rect 2423 2529 2449 2535
rect 7351 2561 7377 2567
rect 14799 2561 14825 2567
rect 8801 2535 8807 2561
rect 8833 2535 8839 2561
rect 7351 2529 7377 2535
rect 14799 2529 14825 2535
rect 15079 2561 15105 2567
rect 16193 2535 16199 2561
rect 16225 2535 16231 2561
rect 17985 2535 17991 2561
rect 18017 2535 18023 2561
rect 20169 2535 20175 2561
rect 20201 2535 20207 2561
rect 24425 2535 24431 2561
rect 24457 2535 24463 2561
rect 24817 2535 24823 2561
rect 24849 2535 24855 2561
rect 15079 2529 15105 2535
rect 13063 2505 13089 2511
rect 8969 2479 8975 2505
rect 9001 2479 9007 2505
rect 13063 2473 13089 2479
rect 15527 2449 15553 2455
rect 15527 2417 15553 2423
rect 16479 2449 16505 2455
rect 16479 2417 16505 2423
rect 17095 2449 17121 2455
rect 17095 2417 17121 2423
rect 18663 2449 18689 2455
rect 18663 2417 18689 2423
rect 336 2365 26040 2382
rect 336 2339 1903 2365
rect 1929 2339 1955 2365
rect 1981 2339 2007 2365
rect 2033 2339 11903 2365
rect 11929 2339 11955 2365
rect 11981 2339 12007 2365
rect 12033 2339 21903 2365
rect 21929 2339 21955 2365
rect 21981 2339 22007 2365
rect 22033 2339 26040 2365
rect 336 2322 26040 2339
rect 25439 2281 25465 2287
rect 25439 2249 25465 2255
rect 14519 2225 14545 2231
rect 18271 2225 18297 2231
rect 24095 2225 24121 2231
rect 16417 2199 16423 2225
rect 16449 2199 16455 2225
rect 18993 2199 18999 2225
rect 19025 2199 19031 2225
rect 14519 2193 14545 2199
rect 18271 2193 18297 2199
rect 24095 2193 24121 2199
rect 11831 2169 11857 2175
rect 12777 2143 12783 2169
rect 12809 2143 12815 2169
rect 14289 2143 14295 2169
rect 14321 2143 14327 2169
rect 14681 2143 14687 2169
rect 14713 2143 14719 2169
rect 15465 2143 15471 2169
rect 15497 2143 15503 2169
rect 17145 2143 17151 2169
rect 17177 2143 17183 2169
rect 18769 2143 18775 2169
rect 18801 2143 18807 2169
rect 24369 2143 24375 2169
rect 24401 2143 24407 2169
rect 25601 2143 25607 2169
rect 25633 2143 25639 2169
rect 11831 2137 11857 2143
rect 967 2113 993 2119
rect 967 2081 993 2087
rect 6399 2113 6425 2119
rect 22471 2113 22497 2119
rect 11993 2087 11999 2113
rect 12025 2087 12031 2113
rect 15857 2087 15863 2113
rect 15889 2087 15895 2113
rect 16865 2087 16871 2113
rect 16897 2087 16903 2113
rect 6399 2081 6425 2087
rect 22471 2081 22497 2087
rect 23815 2113 23841 2119
rect 24705 2087 24711 2113
rect 24737 2087 24743 2113
rect 23815 2081 23841 2087
rect 1247 2057 1273 2063
rect 1247 2025 1273 2031
rect 6679 2057 6705 2063
rect 6679 2025 6705 2031
rect 11551 2057 11577 2063
rect 11551 2025 11577 2031
rect 12279 2057 12305 2063
rect 12279 2025 12305 2031
rect 13063 2057 13089 2063
rect 13063 2025 13089 2031
rect 14967 2057 14993 2063
rect 14967 2025 14993 2031
rect 17319 2057 17345 2063
rect 17319 2025 17345 2031
rect 19223 2057 19249 2063
rect 19223 2025 19249 2031
rect 22191 2057 22217 2063
rect 22191 2025 22217 2031
rect 336 1973 26040 1990
rect 336 1947 2233 1973
rect 2259 1947 2285 1973
rect 2311 1947 2337 1973
rect 2363 1947 12233 1973
rect 12259 1947 12285 1973
rect 12311 1947 12337 1973
rect 12363 1947 22233 1973
rect 22259 1947 22285 1973
rect 22311 1947 22337 1973
rect 22363 1947 26040 1973
rect 336 1930 26040 1947
rect 5559 1833 5585 1839
rect 5559 1801 5585 1807
rect 9199 1833 9225 1839
rect 12839 1833 12865 1839
rect 11377 1807 11383 1833
rect 11409 1807 11415 1833
rect 13001 1807 13007 1833
rect 13033 1807 13039 1833
rect 14121 1807 14127 1833
rect 14153 1807 14159 1833
rect 14905 1807 14911 1833
rect 14937 1807 14943 1833
rect 17593 1807 17599 1833
rect 17625 1807 17631 1833
rect 18377 1807 18383 1833
rect 18409 1807 18415 1833
rect 19161 1807 19167 1833
rect 19193 1807 19199 1833
rect 25209 1807 25215 1833
rect 25241 1807 25247 1833
rect 9199 1801 9225 1807
rect 12839 1801 12865 1807
rect 5279 1777 5305 1783
rect 8969 1751 8975 1777
rect 9001 1751 9007 1777
rect 12609 1751 12615 1777
rect 12641 1751 12647 1777
rect 16193 1751 16199 1777
rect 16225 1751 16231 1777
rect 23529 1751 23535 1777
rect 23561 1751 23567 1777
rect 24425 1751 24431 1777
rect 24457 1751 24463 1777
rect 5279 1745 5305 1751
rect 16479 1721 16505 1727
rect 11825 1695 11831 1721
rect 11857 1695 11863 1721
rect 16479 1689 16505 1695
rect 17879 1721 17905 1727
rect 17879 1689 17905 1695
rect 18663 1721 18689 1727
rect 24935 1721 24961 1727
rect 23697 1695 23703 1721
rect 23729 1695 23735 1721
rect 18663 1689 18689 1695
rect 24935 1689 24961 1695
rect 25719 1721 25745 1727
rect 25719 1689 25745 1695
rect 13287 1665 13313 1671
rect 13287 1633 13313 1639
rect 14407 1665 14433 1671
rect 14407 1633 14433 1639
rect 15191 1665 15217 1671
rect 15191 1633 15217 1639
rect 17095 1665 17121 1671
rect 17095 1633 17121 1639
rect 336 1581 26040 1598
rect 336 1555 1903 1581
rect 1929 1555 1955 1581
rect 1981 1555 2007 1581
rect 2033 1555 11903 1581
rect 11929 1555 11955 1581
rect 11981 1555 12007 1581
rect 12033 1555 21903 1581
rect 21929 1555 21955 1581
rect 21981 1555 22007 1581
rect 22033 1555 26040 1581
rect 336 1538 26040 1555
rect 1751 1441 1777 1447
rect 1751 1409 1777 1415
rect 5223 1441 5249 1447
rect 5223 1409 5249 1415
rect 5671 1441 5697 1447
rect 24039 1441 24065 1447
rect 17593 1415 17599 1441
rect 17625 1415 17631 1441
rect 25545 1415 25551 1441
rect 25577 1415 25583 1441
rect 5671 1409 5697 1415
rect 24039 1409 24065 1415
rect 1471 1385 1497 1391
rect 23087 1385 23113 1391
rect 11769 1359 11775 1385
rect 11801 1359 11807 1385
rect 12609 1359 12615 1385
rect 12641 1359 12647 1385
rect 13337 1359 13343 1385
rect 13369 1359 13375 1385
rect 14345 1359 14351 1385
rect 14377 1359 14383 1385
rect 15017 1359 15023 1385
rect 15049 1359 15055 1385
rect 15801 1359 15807 1385
rect 15833 1359 15839 1385
rect 16585 1359 16591 1385
rect 16617 1359 16623 1385
rect 17425 1359 17431 1385
rect 17457 1359 17463 1385
rect 18769 1359 18775 1385
rect 18801 1359 18807 1385
rect 19553 1359 19559 1385
rect 19585 1359 19591 1385
rect 23529 1359 23535 1385
rect 23561 1359 23567 1385
rect 25097 1359 25103 1385
rect 25129 1359 25135 1385
rect 1471 1353 1497 1359
rect 23087 1353 23113 1359
rect 11607 1329 11633 1335
rect 20007 1329 20033 1335
rect 12161 1303 12167 1329
rect 12193 1303 12199 1329
rect 18377 1303 18383 1329
rect 18409 1303 18415 1329
rect 19161 1303 19167 1329
rect 19193 1303 19199 1329
rect 11607 1297 11633 1303
rect 20007 1297 20033 1303
rect 23367 1329 23393 1335
rect 24313 1303 24319 1329
rect 24345 1303 24351 1329
rect 24705 1303 24711 1329
rect 24737 1303 24743 1329
rect 23367 1297 23393 1303
rect 4943 1273 4969 1279
rect 4943 1241 4969 1247
rect 5391 1273 5417 1279
rect 5391 1241 5417 1247
rect 11327 1273 11353 1279
rect 11327 1241 11353 1247
rect 12839 1273 12865 1279
rect 12839 1241 12865 1247
rect 13623 1273 13649 1279
rect 13623 1241 13649 1247
rect 14519 1273 14545 1279
rect 14519 1241 14545 1247
rect 15303 1273 15329 1279
rect 15303 1241 15329 1247
rect 16087 1273 16113 1279
rect 16087 1241 16113 1247
rect 16871 1273 16897 1279
rect 16871 1241 16897 1247
rect 19727 1273 19753 1279
rect 19727 1241 19753 1247
rect 336 1189 26040 1206
rect 336 1163 2233 1189
rect 2259 1163 2285 1189
rect 2311 1163 2337 1189
rect 2363 1163 12233 1189
rect 12259 1163 12285 1189
rect 12311 1163 12337 1189
rect 12363 1163 22233 1189
rect 22259 1163 22285 1189
rect 22311 1163 22337 1189
rect 22363 1163 26040 1189
rect 336 1146 26040 1163
rect 2199 1105 2225 1111
rect 2199 1073 2225 1079
rect 19335 1105 19361 1111
rect 19335 1073 19361 1079
rect 2479 1049 2505 1055
rect 2479 1017 2505 1023
rect 9367 1049 9393 1055
rect 9367 1017 9393 1023
rect 10655 1049 10681 1055
rect 22471 1049 22497 1055
rect 11377 1023 11383 1049
rect 11409 1023 11415 1049
rect 12889 1023 12895 1049
rect 12921 1023 12927 1049
rect 13673 1023 13679 1049
rect 13705 1023 13711 1049
rect 14457 1023 14463 1049
rect 14489 1023 14495 1049
rect 15241 1023 15247 1049
rect 15273 1023 15279 1049
rect 16193 1023 16199 1049
rect 16225 1023 16231 1049
rect 16977 1023 16983 1049
rect 17009 1023 17015 1049
rect 10655 1017 10681 1023
rect 22471 1017 22497 1023
rect 22751 1049 22777 1055
rect 22751 1017 22777 1023
rect 10375 993 10401 999
rect 19615 993 19641 999
rect 23759 993 23785 999
rect 5833 967 5839 993
rect 5865 967 5871 993
rect 9137 967 9143 993
rect 9169 967 9175 993
rect 12497 967 12503 993
rect 12529 967 12535 993
rect 18377 967 18383 993
rect 18409 967 18415 993
rect 18545 967 18551 993
rect 18577 967 18583 993
rect 23529 967 23535 993
rect 23561 967 23567 993
rect 24481 967 24487 993
rect 24513 967 24519 993
rect 25209 967 25215 993
rect 25241 967 25247 993
rect 10375 961 10401 967
rect 19615 961 19641 967
rect 23759 961 23785 967
rect 12727 937 12753 943
rect 5665 911 5671 937
rect 5697 911 5703 937
rect 11769 911 11775 937
rect 11801 911 11807 937
rect 12727 905 12753 911
rect 24935 937 24961 943
rect 24935 905 24961 911
rect 25719 937 25745 943
rect 25719 905 25745 911
rect 13175 881 13201 887
rect 13175 849 13201 855
rect 13959 881 13985 887
rect 13959 849 13985 855
rect 14743 881 14769 887
rect 14743 849 14769 855
rect 15527 881 15553 887
rect 15527 849 15553 855
rect 16479 881 16505 887
rect 16479 849 16505 855
rect 17263 881 17289 887
rect 17263 849 17289 855
rect 17879 881 17905 887
rect 17879 849 17905 855
rect 18831 881 18857 887
rect 18831 849 18857 855
rect 336 797 26040 814
rect 336 771 1903 797
rect 1929 771 1955 797
rect 1981 771 2007 797
rect 2033 771 11903 797
rect 11929 771 11955 797
rect 11981 771 12007 797
rect 12033 771 21903 797
rect 21929 771 21955 797
rect 21981 771 22007 797
rect 22033 771 26040 797
rect 336 754 26040 771
rect 18943 713 18969 719
rect 18943 681 18969 687
rect 24879 713 24905 719
rect 24879 681 24905 687
rect 10767 657 10793 663
rect 19671 657 19697 663
rect 11489 631 11495 657
rect 11521 631 11527 657
rect 10767 625 10793 631
rect 19671 625 19697 631
rect 24095 657 24121 663
rect 24095 625 24121 631
rect 25551 657 25577 663
rect 25551 625 25577 631
rect 25271 601 25297 607
rect 10257 575 10263 601
rect 10289 575 10295 601
rect 11041 575 11047 601
rect 11073 575 11079 601
rect 13561 575 13567 601
rect 13593 575 13599 601
rect 13841 575 13847 601
rect 13873 575 13879 601
rect 14625 575 14631 601
rect 14657 575 14663 601
rect 16529 575 16535 601
rect 16561 575 16567 601
rect 17649 575 17655 601
rect 17681 575 17687 601
rect 18489 575 18495 601
rect 18521 575 18527 601
rect 20057 575 20063 601
rect 20089 575 20095 601
rect 23697 575 23703 601
rect 23729 575 23735 601
rect 24369 575 24375 601
rect 24401 575 24407 601
rect 25271 569 25297 575
rect 12161 519 12167 545
rect 12193 519 12199 545
rect 12553 519 12559 545
rect 12585 519 12591 545
rect 15745 519 15751 545
rect 15777 519 15783 545
rect 20561 519 20567 545
rect 20593 519 20599 545
rect 20953 519 20959 545
rect 20985 519 20991 545
rect 13287 489 13313 495
rect 13287 457 13313 463
rect 14127 489 14153 495
rect 14127 457 14153 463
rect 14911 489 14937 495
rect 14911 457 14937 463
rect 16031 489 16057 495
rect 16031 457 16057 463
rect 16815 489 16841 495
rect 16815 457 16841 463
rect 17935 489 17961 495
rect 17935 457 17961 463
rect 336 405 26040 422
rect 336 379 2233 405
rect 2259 379 2285 405
rect 2311 379 2337 405
rect 2363 379 12233 405
rect 12259 379 12285 405
rect 12311 379 12337 405
rect 12363 379 22233 405
rect 22259 379 22285 405
rect 22311 379 22337 405
rect 22363 379 26040 405
rect 336 362 26040 379
<< via1 >>
rect 2233 6651 2259 6677
rect 2285 6651 2311 6677
rect 2337 6651 2363 6677
rect 12233 6651 12259 6677
rect 12285 6651 12311 6677
rect 12337 6651 12363 6677
rect 22233 6651 22259 6677
rect 22285 6651 22311 6677
rect 22337 6651 22363 6677
rect 911 6567 937 6593
rect 19839 6567 19865 6593
rect 22135 6567 22161 6593
rect 23647 6567 23673 6593
rect 24599 6567 24625 6593
rect 2647 6511 2673 6537
rect 3039 6511 3065 6537
rect 6455 6511 6481 6537
rect 1079 6455 1105 6481
rect 3991 6455 4017 6481
rect 5223 6455 5249 6481
rect 6847 6455 6873 6481
rect 7687 6455 7713 6481
rect 8919 6455 8945 6481
rect 9759 6455 9785 6481
rect 11271 6455 11297 6481
rect 12503 6455 12529 6481
rect 13455 6455 13481 6481
rect 14967 6455 14993 6481
rect 16367 6455 16393 6481
rect 17375 6455 17401 6481
rect 18775 6455 18801 6481
rect 19559 6455 19585 6481
rect 21071 6455 21097 6481
rect 21855 6455 21881 6481
rect 22807 6455 22833 6481
rect 23087 6455 23113 6481
rect 23367 6455 23393 6481
rect 24375 6455 24401 6481
rect 25271 6455 25297 6481
rect 3487 6399 3513 6425
rect 4719 6399 4745 6425
rect 7183 6399 7209 6425
rect 8415 6399 8441 6425
rect 9423 6399 9449 6425
rect 10879 6399 10905 6425
rect 12111 6399 12137 6425
rect 13119 6399 13145 6425
rect 14575 6399 14601 6425
rect 15863 6399 15889 6425
rect 16871 6399 16897 6425
rect 18271 6399 18297 6425
rect 20679 6399 20705 6425
rect 25495 6399 25521 6425
rect 1903 6259 1929 6285
rect 1955 6259 1981 6285
rect 2007 6259 2033 6285
rect 11903 6259 11929 6285
rect 11955 6259 11981 6285
rect 12007 6259 12033 6285
rect 21903 6259 21929 6285
rect 21955 6259 21981 6285
rect 22007 6259 22033 6285
rect 24039 6175 24065 6201
rect 1359 6119 1385 6145
rect 14855 6119 14881 6145
rect 15247 6119 15273 6145
rect 16591 6119 16617 6145
rect 17039 6119 17065 6145
rect 18831 6119 18857 6145
rect 20847 6119 20873 6145
rect 21295 6119 21321 6145
rect 23031 6119 23057 6145
rect 24823 6119 24849 6145
rect 25607 6119 25633 6145
rect 1135 6063 1161 6089
rect 5055 6063 5081 6089
rect 15023 6063 15049 6089
rect 23311 6063 23337 6089
rect 24375 6063 24401 6089
rect 3767 6007 3793 6033
rect 5279 6007 5305 6033
rect 16871 6007 16897 6033
rect 22359 6007 22385 6033
rect 23535 6007 23561 6033
rect 25103 6007 25129 6033
rect 3487 5951 3513 5977
rect 15527 5951 15553 5977
rect 16087 5951 16113 5977
rect 16255 5951 16281 5977
rect 17319 5951 17345 5977
rect 19055 5951 19081 5977
rect 20567 5951 20593 5977
rect 21015 5951 21041 5977
rect 22079 5951 22105 5977
rect 2233 5867 2259 5893
rect 2285 5867 2311 5893
rect 2337 5867 2363 5893
rect 12233 5867 12259 5893
rect 12285 5867 12311 5893
rect 12337 5867 12363 5893
rect 22233 5867 22259 5893
rect 22285 5867 22311 5893
rect 22337 5867 22363 5893
rect 7799 5783 7825 5809
rect 9087 5783 9113 5809
rect 22695 5783 22721 5809
rect 8807 5727 8833 5753
rect 19055 5727 19081 5753
rect 23143 5727 23169 5753
rect 23535 5727 23561 5753
rect 12727 5671 12753 5697
rect 19279 5671 19305 5697
rect 24487 5671 24513 5697
rect 25271 5671 25297 5697
rect 7575 5615 7601 5641
rect 12503 5615 12529 5641
rect 22975 5615 23001 5641
rect 24935 5615 24961 5641
rect 25719 5559 25745 5585
rect 1903 5475 1929 5501
rect 1955 5475 1981 5501
rect 2007 5475 2033 5501
rect 11903 5475 11929 5501
rect 11955 5475 11981 5501
rect 12007 5475 12033 5501
rect 21903 5475 21929 5501
rect 21955 5475 21981 5501
rect 22007 5475 22033 5501
rect 24039 5391 24065 5417
rect 11215 5335 11241 5361
rect 13399 5335 13425 5361
rect 17655 5335 17681 5361
rect 18719 5335 18745 5361
rect 24823 5335 24849 5361
rect 23087 5279 23113 5305
rect 24375 5279 24401 5305
rect 23367 5223 23393 5249
rect 23535 5223 23561 5249
rect 25103 5223 25129 5249
rect 25495 5223 25521 5249
rect 11439 5167 11465 5193
rect 13623 5167 13649 5193
rect 17879 5167 17905 5193
rect 18999 5167 19025 5193
rect 2233 5083 2259 5109
rect 2285 5083 2311 5109
rect 2337 5083 2363 5109
rect 12233 5083 12259 5109
rect 12285 5083 12311 5109
rect 12337 5083 12363 5109
rect 22233 5083 22259 5109
rect 22285 5083 22311 5109
rect 22337 5083 22363 5109
rect 2871 4943 2897 4969
rect 1079 4887 1105 4913
rect 2591 4887 2617 4913
rect 3487 4887 3513 4913
rect 7799 4887 7825 4913
rect 9647 4887 9673 4913
rect 16479 4887 16505 4913
rect 23535 4887 23561 4913
rect 23759 4887 23785 4913
rect 24431 4887 24457 4913
rect 25215 4887 25241 4913
rect 855 4831 881 4857
rect 3767 4831 3793 4857
rect 8079 4831 8105 4857
rect 9927 4831 9953 4857
rect 16199 4831 16225 4857
rect 24935 4831 24961 4857
rect 25719 4775 25745 4801
rect 1903 4691 1929 4717
rect 1955 4691 1981 4717
rect 2007 4691 2033 4717
rect 11903 4691 11929 4717
rect 11955 4691 11981 4717
rect 12007 4691 12033 4717
rect 21903 4691 21929 4717
rect 21955 4691 21981 4717
rect 22007 4691 22033 4717
rect 24823 4607 24849 4633
rect 2143 4551 2169 4577
rect 22751 4551 22777 4577
rect 24151 4551 24177 4577
rect 5279 4495 5305 4521
rect 22471 4495 22497 4521
rect 24375 4495 24401 4521
rect 25159 4495 25185 4521
rect 5559 4439 5585 4465
rect 23871 4439 23897 4465
rect 25495 4439 25521 4465
rect 1919 4383 1945 4409
rect 2233 4299 2259 4325
rect 2285 4299 2311 4325
rect 2337 4299 2363 4325
rect 12233 4299 12259 4325
rect 12285 4299 12311 4325
rect 12337 4299 12363 4325
rect 22233 4299 22259 4325
rect 22285 4299 22311 4325
rect 22337 4299 22363 4325
rect 15135 4159 15161 4185
rect 23255 4159 23281 4185
rect 25047 4159 25073 4185
rect 9255 4103 9281 4129
rect 11775 4103 11801 4129
rect 15415 4103 15441 4129
rect 21295 4103 21321 4129
rect 24375 4103 24401 4129
rect 24599 4103 24625 4129
rect 24767 4103 24793 4129
rect 25215 4103 25241 4129
rect 9479 4047 9505 4073
rect 11999 4047 12025 4073
rect 21519 4047 21545 4073
rect 23479 4047 23505 4073
rect 25719 3991 25745 4017
rect 1903 3907 1929 3933
rect 1955 3907 1981 3933
rect 2007 3907 2033 3933
rect 11903 3907 11929 3933
rect 11955 3907 11981 3933
rect 12007 3907 12033 3933
rect 21903 3907 21929 3933
rect 21955 3907 21981 3933
rect 22007 3907 22033 3933
rect 25607 3823 25633 3849
rect 24151 3767 24177 3793
rect 24823 3767 24849 3793
rect 12279 3711 12305 3737
rect 24375 3711 24401 3737
rect 25103 3711 25129 3737
rect 799 3655 825 3681
rect 2871 3655 2897 3681
rect 4215 3655 4241 3681
rect 11271 3655 11297 3681
rect 12559 3655 12585 3681
rect 23871 3655 23897 3681
rect 1079 3599 1105 3625
rect 3151 3599 3177 3625
rect 4495 3599 4521 3625
rect 10991 3599 11017 3625
rect 2233 3515 2259 3541
rect 2285 3515 2311 3541
rect 2337 3515 2363 3541
rect 12233 3515 12259 3541
rect 12285 3515 12311 3541
rect 12337 3515 12363 3541
rect 22233 3515 22259 3541
rect 22285 3515 22311 3541
rect 22337 3515 22363 3541
rect 16871 3431 16897 3457
rect 4159 3319 4185 3345
rect 7855 3319 7881 3345
rect 8415 3319 8441 3345
rect 13623 3319 13649 3345
rect 15303 3319 15329 3345
rect 17655 3319 17681 3345
rect 21071 3319 21097 3345
rect 22135 3319 22161 3345
rect 24431 3319 24457 3345
rect 25215 3319 25241 3345
rect 3935 3263 3961 3289
rect 8023 3263 8049 3289
rect 8639 3263 8665 3289
rect 13847 3263 13873 3289
rect 15583 3263 15609 3289
rect 17151 3263 17177 3289
rect 17879 3263 17905 3289
rect 21295 3263 21321 3289
rect 22359 3263 22385 3289
rect 24879 3263 24905 3289
rect 25719 3263 25745 3289
rect 1903 3123 1929 3149
rect 1955 3123 1981 3149
rect 2007 3123 2033 3149
rect 11903 3123 11929 3149
rect 11955 3123 11981 3149
rect 12007 3123 12033 3149
rect 21903 3123 21929 3149
rect 21955 3123 21981 3149
rect 22007 3123 22033 3149
rect 25607 3039 25633 3065
rect 855 2983 881 3009
rect 5895 2983 5921 3009
rect 6455 2983 6481 3009
rect 15807 2983 15833 3009
rect 17375 2983 17401 3009
rect 18831 2983 18857 3009
rect 2535 2927 2561 2953
rect 15135 2927 15161 2953
rect 15639 2927 15665 2953
rect 18607 2927 18633 2953
rect 20511 2927 20537 2953
rect 23143 2927 23169 2953
rect 24207 2927 24233 2953
rect 2759 2871 2785 2897
rect 6119 2871 6145 2897
rect 15359 2871 15385 2897
rect 16311 2871 16337 2897
rect 16479 2871 16505 2897
rect 17879 2871 17905 2897
rect 18439 2871 18465 2897
rect 19335 2871 19361 2897
rect 20791 2871 20817 2897
rect 23423 2871 23449 2897
rect 23591 2871 23617 2897
rect 23871 2871 23897 2897
rect 24487 2871 24513 2897
rect 24935 2871 24961 2897
rect 25103 2871 25129 2897
rect 1079 2815 1105 2841
rect 6679 2815 6705 2841
rect 16031 2815 16057 2841
rect 16759 2815 16785 2841
rect 18159 2815 18185 2841
rect 19055 2815 19081 2841
rect 24655 2815 24681 2841
rect 2233 2731 2259 2757
rect 2285 2731 2311 2757
rect 2337 2731 2363 2757
rect 12233 2731 12259 2757
rect 12285 2731 12311 2757
rect 12337 2731 12363 2757
rect 22233 2731 22259 2757
rect 22285 2731 22311 2757
rect 22337 2731 22363 2757
rect 12783 2647 12809 2673
rect 2143 2591 2169 2617
rect 7071 2591 7097 2617
rect 15247 2591 15273 2617
rect 17599 2591 17625 2617
rect 18383 2591 18409 2617
rect 19167 2591 19193 2617
rect 20399 2591 20425 2617
rect 25215 2591 25241 2617
rect 25607 2591 25633 2617
rect 2423 2535 2449 2561
rect 7351 2535 7377 2561
rect 8807 2535 8833 2561
rect 14799 2535 14825 2561
rect 15079 2535 15105 2561
rect 16199 2535 16225 2561
rect 17991 2535 18017 2561
rect 20175 2535 20201 2561
rect 24431 2535 24457 2561
rect 24823 2535 24849 2561
rect 8975 2479 9001 2505
rect 13063 2479 13089 2505
rect 15527 2423 15553 2449
rect 16479 2423 16505 2449
rect 17095 2423 17121 2449
rect 18663 2423 18689 2449
rect 1903 2339 1929 2365
rect 1955 2339 1981 2365
rect 2007 2339 2033 2365
rect 11903 2339 11929 2365
rect 11955 2339 11981 2365
rect 12007 2339 12033 2365
rect 21903 2339 21929 2365
rect 21955 2339 21981 2365
rect 22007 2339 22033 2365
rect 25439 2255 25465 2281
rect 14519 2199 14545 2225
rect 16423 2199 16449 2225
rect 18271 2199 18297 2225
rect 18999 2199 19025 2225
rect 24095 2199 24121 2225
rect 11831 2143 11857 2169
rect 12783 2143 12809 2169
rect 14295 2143 14321 2169
rect 14687 2143 14713 2169
rect 15471 2143 15497 2169
rect 17151 2143 17177 2169
rect 18775 2143 18801 2169
rect 24375 2143 24401 2169
rect 25607 2143 25633 2169
rect 967 2087 993 2113
rect 6399 2087 6425 2113
rect 11999 2087 12025 2113
rect 15863 2087 15889 2113
rect 16871 2087 16897 2113
rect 22471 2087 22497 2113
rect 23815 2087 23841 2113
rect 24711 2087 24737 2113
rect 1247 2031 1273 2057
rect 6679 2031 6705 2057
rect 11551 2031 11577 2057
rect 12279 2031 12305 2057
rect 13063 2031 13089 2057
rect 14967 2031 14993 2057
rect 17319 2031 17345 2057
rect 19223 2031 19249 2057
rect 22191 2031 22217 2057
rect 2233 1947 2259 1973
rect 2285 1947 2311 1973
rect 2337 1947 2363 1973
rect 12233 1947 12259 1973
rect 12285 1947 12311 1973
rect 12337 1947 12363 1973
rect 22233 1947 22259 1973
rect 22285 1947 22311 1973
rect 22337 1947 22363 1973
rect 5559 1807 5585 1833
rect 9199 1807 9225 1833
rect 11383 1807 11409 1833
rect 12839 1807 12865 1833
rect 13007 1807 13033 1833
rect 14127 1807 14153 1833
rect 14911 1807 14937 1833
rect 17599 1807 17625 1833
rect 18383 1807 18409 1833
rect 19167 1807 19193 1833
rect 25215 1807 25241 1833
rect 5279 1751 5305 1777
rect 8975 1751 9001 1777
rect 12615 1751 12641 1777
rect 16199 1751 16225 1777
rect 23535 1751 23561 1777
rect 24431 1751 24457 1777
rect 11831 1695 11857 1721
rect 16479 1695 16505 1721
rect 17879 1695 17905 1721
rect 18663 1695 18689 1721
rect 23703 1695 23729 1721
rect 24935 1695 24961 1721
rect 25719 1695 25745 1721
rect 13287 1639 13313 1665
rect 14407 1639 14433 1665
rect 15191 1639 15217 1665
rect 17095 1639 17121 1665
rect 1903 1555 1929 1581
rect 1955 1555 1981 1581
rect 2007 1555 2033 1581
rect 11903 1555 11929 1581
rect 11955 1555 11981 1581
rect 12007 1555 12033 1581
rect 21903 1555 21929 1581
rect 21955 1555 21981 1581
rect 22007 1555 22033 1581
rect 1751 1415 1777 1441
rect 5223 1415 5249 1441
rect 5671 1415 5697 1441
rect 17599 1415 17625 1441
rect 24039 1415 24065 1441
rect 25551 1415 25577 1441
rect 1471 1359 1497 1385
rect 11775 1359 11801 1385
rect 12615 1359 12641 1385
rect 13343 1359 13369 1385
rect 14351 1359 14377 1385
rect 15023 1359 15049 1385
rect 15807 1359 15833 1385
rect 16591 1359 16617 1385
rect 17431 1359 17457 1385
rect 18775 1359 18801 1385
rect 19559 1359 19585 1385
rect 23087 1359 23113 1385
rect 23535 1359 23561 1385
rect 25103 1359 25129 1385
rect 11607 1303 11633 1329
rect 12167 1303 12193 1329
rect 18383 1303 18409 1329
rect 19167 1303 19193 1329
rect 20007 1303 20033 1329
rect 23367 1303 23393 1329
rect 24319 1303 24345 1329
rect 24711 1303 24737 1329
rect 4943 1247 4969 1273
rect 5391 1247 5417 1273
rect 11327 1247 11353 1273
rect 12839 1247 12865 1273
rect 13623 1247 13649 1273
rect 14519 1247 14545 1273
rect 15303 1247 15329 1273
rect 16087 1247 16113 1273
rect 16871 1247 16897 1273
rect 19727 1247 19753 1273
rect 2233 1163 2259 1189
rect 2285 1163 2311 1189
rect 2337 1163 2363 1189
rect 12233 1163 12259 1189
rect 12285 1163 12311 1189
rect 12337 1163 12363 1189
rect 22233 1163 22259 1189
rect 22285 1163 22311 1189
rect 22337 1163 22363 1189
rect 2199 1079 2225 1105
rect 19335 1079 19361 1105
rect 2479 1023 2505 1049
rect 9367 1023 9393 1049
rect 10655 1023 10681 1049
rect 11383 1023 11409 1049
rect 12895 1023 12921 1049
rect 13679 1023 13705 1049
rect 14463 1023 14489 1049
rect 15247 1023 15273 1049
rect 16199 1023 16225 1049
rect 16983 1023 17009 1049
rect 22471 1023 22497 1049
rect 22751 1023 22777 1049
rect 5839 967 5865 993
rect 9143 967 9169 993
rect 10375 967 10401 993
rect 12503 967 12529 993
rect 18383 967 18409 993
rect 18551 967 18577 993
rect 19615 967 19641 993
rect 23535 967 23561 993
rect 23759 967 23785 993
rect 24487 967 24513 993
rect 25215 967 25241 993
rect 5671 911 5697 937
rect 11775 911 11801 937
rect 12727 911 12753 937
rect 24935 911 24961 937
rect 25719 911 25745 937
rect 13175 855 13201 881
rect 13959 855 13985 881
rect 14743 855 14769 881
rect 15527 855 15553 881
rect 16479 855 16505 881
rect 17263 855 17289 881
rect 17879 855 17905 881
rect 18831 855 18857 881
rect 1903 771 1929 797
rect 1955 771 1981 797
rect 2007 771 2033 797
rect 11903 771 11929 797
rect 11955 771 11981 797
rect 12007 771 12033 797
rect 21903 771 21929 797
rect 21955 771 21981 797
rect 22007 771 22033 797
rect 18943 687 18969 713
rect 24879 687 24905 713
rect 10767 631 10793 657
rect 11495 631 11521 657
rect 19671 631 19697 657
rect 24095 631 24121 657
rect 25551 631 25577 657
rect 10263 575 10289 601
rect 11047 575 11073 601
rect 13567 575 13593 601
rect 13847 575 13873 601
rect 14631 575 14657 601
rect 16535 575 16561 601
rect 17655 575 17681 601
rect 18495 575 18521 601
rect 20063 575 20089 601
rect 23703 575 23729 601
rect 24375 575 24401 601
rect 25271 575 25297 601
rect 12167 519 12193 545
rect 12559 519 12585 545
rect 15751 519 15777 545
rect 20567 519 20593 545
rect 20959 519 20985 545
rect 13287 463 13313 489
rect 14127 463 14153 489
rect 14911 463 14937 489
rect 16031 463 16057 489
rect 16815 463 16841 489
rect 17935 463 17961 489
rect 2233 379 2259 405
rect 2285 379 2311 405
rect 2337 379 2363 405
rect 12233 379 12259 405
rect 12285 379 12311 405
rect 12337 379 12363 405
rect 22233 379 22259 405
rect 22285 379 22311 405
rect 22337 379 22363 405
<< metal2 >>
rect 784 7056 840 7112
rect 2016 7056 2072 7112
rect 3248 7056 3304 7112
rect 4480 7056 4536 7112
rect 5712 7056 5768 7112
rect 6944 7056 7000 7112
rect 8176 7056 8232 7112
rect 9408 7056 9464 7112
rect 10640 7056 10696 7112
rect 11872 7056 11928 7112
rect 13104 7056 13160 7112
rect 14336 7056 14392 7112
rect 15568 7056 15624 7112
rect 16800 7056 16856 7112
rect 18032 7056 18088 7112
rect 19264 7056 19320 7112
rect 20496 7056 20552 7112
rect 21728 7056 21784 7112
rect 798 6818 826 7056
rect 798 6790 938 6818
rect 910 6593 938 6790
rect 910 6567 911 6593
rect 937 6567 938 6593
rect 910 6561 938 6567
rect 1134 6762 1162 6767
rect 1078 6482 1106 6487
rect 1078 6435 1106 6454
rect 574 6314 602 6319
rect 350 6090 378 6095
rect 350 4858 378 6062
rect 574 5810 602 6286
rect 1134 6089 1162 6734
rect 1638 6538 1666 6543
rect 1358 6426 1386 6431
rect 1358 6145 1386 6398
rect 1358 6119 1359 6145
rect 1385 6119 1386 6145
rect 1358 6113 1386 6119
rect 1134 6063 1135 6089
rect 1161 6063 1162 6089
rect 1134 6057 1162 6063
rect 574 5777 602 5782
rect 1638 5026 1666 6510
rect 2030 6538 2058 7056
rect 3262 7042 3290 7056
rect 3262 7009 3290 7014
rect 3486 7042 3514 7047
rect 3038 6762 3066 6767
rect 2232 6678 2364 6683
rect 2260 6650 2284 6678
rect 2312 6650 2336 6678
rect 2232 6645 2364 6650
rect 2030 6505 2058 6510
rect 2646 6538 2674 6543
rect 2646 6491 2674 6510
rect 3038 6537 3066 6734
rect 3038 6511 3039 6537
rect 3065 6511 3066 6537
rect 3038 6505 3066 6511
rect 2478 6482 2506 6487
rect 1902 6286 2034 6291
rect 1930 6258 1954 6286
rect 1982 6258 2006 6286
rect 1902 6253 2034 6258
rect 2232 5894 2364 5899
rect 2260 5866 2284 5894
rect 2312 5866 2336 5894
rect 2232 5861 2364 5866
rect 1902 5502 2034 5507
rect 1930 5474 1954 5502
rect 1982 5474 2006 5502
rect 1902 5469 2034 5474
rect 2422 5418 2450 5423
rect 2232 5110 2364 5115
rect 2260 5082 2284 5110
rect 2312 5082 2336 5110
rect 2232 5077 2364 5082
rect 1638 4993 1666 4998
rect 1078 4913 1106 4919
rect 1078 4887 1079 4913
rect 1105 4887 1106 4913
rect 350 4825 378 4830
rect 854 4857 882 4863
rect 854 4831 855 4857
rect 881 4831 882 4857
rect 798 3681 826 3687
rect 798 3655 799 3681
rect 825 3655 826 3681
rect 798 3346 826 3655
rect 854 3458 882 4831
rect 1078 4018 1106 4887
rect 1902 4718 2034 4723
rect 1930 4690 1954 4718
rect 1982 4690 2006 4718
rect 1902 4685 2034 4690
rect 2142 4577 2170 4583
rect 2142 4551 2143 4577
rect 2169 4551 2170 4577
rect 1918 4409 1946 4415
rect 1918 4383 1919 4409
rect 1945 4383 1946 4409
rect 1918 4214 1946 4383
rect 1078 3985 1106 3990
rect 1806 4186 1946 4214
rect 1078 3626 1106 3631
rect 1078 3625 1162 3626
rect 1078 3599 1079 3625
rect 1105 3599 1162 3625
rect 1078 3598 1162 3599
rect 1078 3593 1106 3598
rect 854 3425 882 3430
rect 798 3318 938 3346
rect 854 3010 882 3015
rect 854 2963 882 2982
rect 910 1722 938 3318
rect 1078 2842 1106 2847
rect 1078 2795 1106 2814
rect 966 2114 994 2119
rect 966 2067 994 2086
rect 910 1689 938 1694
rect 1134 210 1162 3598
rect 1806 3402 1834 4186
rect 1902 3934 2034 3939
rect 1930 3906 1954 3934
rect 1982 3906 2006 3934
rect 1902 3901 2034 3906
rect 2142 3738 2170 4551
rect 2232 4326 2364 4331
rect 2260 4298 2284 4326
rect 2312 4298 2336 4326
rect 2232 4293 2364 4298
rect 2422 4214 2450 5390
rect 2478 5194 2506 6454
rect 3486 6425 3514 7014
rect 4494 7042 4522 7056
rect 4494 7009 4522 7014
rect 4718 7042 4746 7047
rect 3486 6399 3487 6425
rect 3513 6399 3514 6425
rect 3486 6393 3514 6399
rect 3990 6481 4018 6487
rect 3990 6455 3991 6481
rect 4017 6455 4018 6481
rect 3766 6033 3794 6039
rect 3766 6007 3767 6033
rect 3793 6007 3794 6033
rect 3486 5977 3514 5983
rect 3486 5951 3487 5977
rect 3513 5951 3514 5977
rect 3486 5642 3514 5951
rect 3486 5609 3514 5614
rect 3542 5922 3570 5927
rect 2478 5161 2506 5166
rect 2758 4970 2786 4975
rect 2590 4913 2618 4919
rect 2590 4887 2591 4913
rect 2617 4887 2618 4913
rect 2422 4186 2506 4214
rect 2142 3705 2170 3710
rect 2478 3570 2506 4186
rect 2590 3626 2618 4887
rect 2702 4914 2730 4919
rect 2702 3682 2730 4886
rect 2758 3794 2786 4942
rect 2870 4970 2898 4975
rect 2870 4923 2898 4942
rect 3542 4970 3570 5894
rect 3766 5530 3794 6007
rect 3990 5586 4018 6455
rect 4718 6425 4746 7014
rect 5726 6538 5754 7056
rect 6958 7042 6986 7056
rect 6958 7009 6986 7014
rect 7182 7042 7210 7047
rect 5726 6505 5754 6510
rect 6454 6538 6482 6543
rect 6454 6491 6482 6510
rect 4718 6399 4719 6425
rect 4745 6399 4746 6425
rect 4718 6393 4746 6399
rect 5222 6481 5250 6487
rect 5222 6455 5223 6481
rect 5249 6455 5250 6481
rect 3990 5553 4018 5558
rect 5054 6089 5082 6095
rect 5054 6063 5055 6089
rect 5081 6063 5082 6089
rect 3766 5497 3794 5502
rect 5054 5250 5082 6063
rect 5222 5642 5250 6455
rect 6846 6482 6874 6487
rect 6846 6435 6874 6454
rect 7182 6425 7210 7014
rect 8190 7042 8218 7056
rect 8190 7009 8218 7014
rect 8414 7042 8442 7047
rect 7182 6399 7183 6425
rect 7209 6399 7210 6425
rect 7182 6393 7210 6399
rect 7686 6481 7714 6487
rect 7686 6455 7687 6481
rect 7713 6455 7714 6481
rect 6454 6146 6482 6151
rect 5222 5609 5250 5614
rect 5278 6033 5306 6039
rect 5278 6007 5279 6033
rect 5305 6007 5306 6033
rect 5054 5217 5082 5222
rect 5278 5250 5306 6007
rect 5278 5217 5306 5222
rect 3542 4937 3570 4942
rect 4270 5194 4298 5199
rect 3486 4913 3514 4919
rect 3486 4887 3487 4913
rect 3513 4887 3514 4913
rect 3374 4858 3402 4863
rect 2926 4802 2954 4807
rect 2926 3850 2954 4774
rect 3038 4522 3066 4527
rect 2982 4242 3010 4247
rect 2982 3906 3010 4214
rect 2982 3873 3010 3878
rect 2926 3817 2954 3822
rect 2758 3761 2786 3766
rect 2870 3682 2898 3687
rect 2702 3654 2842 3682
rect 2590 3593 2618 3598
rect 2232 3542 2364 3547
rect 2260 3514 2284 3542
rect 2312 3514 2336 3542
rect 2478 3537 2506 3542
rect 2232 3509 2364 3514
rect 1806 3369 1834 3374
rect 1902 3150 2034 3155
rect 1930 3122 1954 3150
rect 1982 3122 2006 3150
rect 1902 3117 2034 3122
rect 2534 3066 2562 3071
rect 2086 2954 2114 2959
rect 1806 2730 1834 2735
rect 1134 177 1162 182
rect 1246 2057 1274 2063
rect 1246 2031 1247 2057
rect 1273 2031 1274 2057
rect 1246 98 1274 2031
rect 1470 2058 1498 2063
rect 1470 1385 1498 2030
rect 1750 1442 1778 1447
rect 1750 1395 1778 1414
rect 1470 1359 1471 1385
rect 1497 1359 1498 1385
rect 1470 1353 1498 1359
rect 1302 1330 1330 1335
rect 1302 490 1330 1302
rect 1302 457 1330 462
rect 1806 490 1834 2702
rect 1902 2366 2034 2371
rect 1930 2338 1954 2366
rect 1982 2338 2006 2366
rect 1902 2333 2034 2338
rect 1902 1582 2034 1587
rect 1930 1554 1954 1582
rect 1982 1554 2006 1582
rect 1902 1549 2034 1554
rect 2086 1106 2114 2926
rect 2534 2953 2562 3038
rect 2534 2927 2535 2953
rect 2561 2927 2562 2953
rect 2534 2921 2562 2927
rect 2646 3010 2674 3015
rect 2232 2758 2364 2763
rect 2260 2730 2284 2758
rect 2312 2730 2336 2758
rect 2232 2725 2364 2730
rect 2142 2618 2170 2623
rect 2142 2571 2170 2590
rect 2422 2562 2450 2567
rect 2422 2515 2450 2534
rect 2534 2338 2562 2343
rect 2232 1974 2364 1979
rect 2260 1946 2284 1974
rect 2312 1946 2336 1974
rect 2232 1941 2364 1946
rect 2478 1610 2506 1615
rect 2232 1190 2364 1195
rect 2260 1162 2284 1190
rect 2312 1162 2336 1190
rect 2232 1157 2364 1162
rect 2198 1106 2226 1111
rect 2086 1105 2226 1106
rect 2086 1079 2199 1105
rect 2225 1079 2226 1105
rect 2086 1078 2226 1079
rect 2198 1073 2226 1078
rect 2478 1049 2506 1582
rect 2534 1442 2562 2310
rect 2534 1409 2562 1414
rect 2590 2114 2618 2119
rect 2478 1023 2479 1049
rect 2505 1023 2506 1049
rect 2478 1017 2506 1023
rect 2590 1050 2618 2086
rect 2646 1834 2674 2982
rect 2758 2897 2786 2903
rect 2758 2871 2759 2897
rect 2785 2871 2786 2897
rect 2758 2786 2786 2871
rect 2758 2753 2786 2758
rect 2646 1801 2674 1806
rect 2702 2226 2730 2231
rect 2702 1330 2730 2198
rect 2702 1297 2730 1302
rect 2814 1106 2842 3654
rect 2870 3635 2898 3654
rect 2926 3626 2954 3631
rect 2870 3458 2898 3463
rect 2870 2170 2898 3430
rect 2926 2506 2954 3598
rect 3038 2954 3066 4494
rect 3038 2921 3066 2926
rect 3094 4242 3122 4247
rect 2926 2473 2954 2478
rect 3094 2282 3122 4214
rect 3374 4130 3402 4830
rect 3374 4097 3402 4102
rect 3486 4074 3514 4887
rect 3766 4857 3794 4863
rect 3766 4831 3767 4857
rect 3793 4831 3794 4857
rect 3766 4298 3794 4831
rect 3766 4265 3794 4270
rect 3486 4041 3514 4046
rect 3206 4018 3234 4023
rect 3094 2249 3122 2254
rect 3150 3625 3178 3631
rect 3150 3599 3151 3625
rect 3177 3599 3178 3625
rect 2870 2137 2898 2142
rect 2814 1073 2842 1078
rect 2590 1017 2618 1022
rect 3150 882 3178 3599
rect 3150 849 3178 854
rect 1902 798 2034 803
rect 1930 770 1954 798
rect 1982 770 2006 798
rect 1902 765 2034 770
rect 1806 457 1834 462
rect 2232 406 2364 411
rect 2260 378 2284 406
rect 2312 378 2336 406
rect 2232 373 2364 378
rect 3206 154 3234 3990
rect 3710 3682 3738 3687
rect 3318 3066 3346 3071
rect 3318 1610 3346 3038
rect 3318 1577 3346 1582
rect 3374 3010 3402 3015
rect 3374 882 3402 2982
rect 3318 854 3402 882
rect 3542 1722 3570 1727
rect 3318 714 3346 854
rect 3318 681 3346 686
rect 3542 602 3570 1694
rect 3710 1162 3738 3654
rect 4214 3681 4242 3687
rect 4214 3655 4215 3681
rect 4241 3655 4242 3681
rect 4158 3345 4186 3351
rect 4158 3319 4159 3345
rect 4185 3319 4186 3345
rect 3934 3289 3962 3295
rect 3934 3263 3935 3289
rect 3961 3263 3962 3289
rect 3934 2002 3962 3263
rect 4158 3290 4186 3319
rect 4158 3257 4186 3262
rect 3934 1969 3962 1974
rect 4214 1946 4242 3655
rect 4270 3346 4298 5166
rect 4326 5138 4354 5143
rect 4326 3626 4354 5110
rect 4326 3593 4354 3598
rect 4382 4970 4410 4975
rect 4270 3313 4298 3318
rect 4214 1913 4242 1918
rect 4382 1890 4410 4942
rect 6454 4970 6482 6118
rect 7126 5922 7154 5927
rect 6454 4937 6482 4942
rect 6958 5474 6986 5479
rect 6958 4802 6986 5446
rect 7126 4970 7154 5894
rect 7574 5642 7602 5647
rect 7574 5595 7602 5614
rect 7126 4937 7154 4942
rect 7462 5530 7490 5535
rect 6958 4769 6986 4774
rect 6174 4690 6202 4695
rect 5278 4634 5306 4639
rect 5278 4521 5306 4606
rect 5278 4495 5279 4521
rect 5305 4495 5306 4521
rect 5278 4489 5306 4495
rect 5558 4465 5586 4471
rect 5558 4439 5559 4465
rect 5585 4439 5586 4465
rect 5558 4354 5586 4439
rect 5558 4321 5586 4326
rect 4494 3626 4522 3631
rect 4494 3579 4522 3598
rect 5558 3514 5586 3519
rect 4382 1857 4410 1862
rect 4998 2842 5026 2847
rect 3710 1129 3738 1134
rect 4942 1273 4970 1279
rect 4942 1247 4943 1273
rect 4969 1247 4970 1273
rect 3542 569 3570 574
rect 3206 121 3234 126
rect 1246 65 1274 70
rect 4942 42 4970 1247
rect 4998 490 5026 2814
rect 5558 1833 5586 3486
rect 6006 3290 6034 3295
rect 5894 3009 5922 3015
rect 5894 2983 5895 3009
rect 5921 2983 5922 3009
rect 5894 2170 5922 2983
rect 5894 2137 5922 2142
rect 5558 1807 5559 1833
rect 5585 1807 5586 1833
rect 5558 1801 5586 1807
rect 5782 2002 5810 2007
rect 5278 1777 5306 1783
rect 5278 1751 5279 1777
rect 5305 1751 5306 1777
rect 5222 1554 5250 1559
rect 5222 1441 5250 1526
rect 5222 1415 5223 1441
rect 5249 1415 5250 1441
rect 5222 1409 5250 1415
rect 4998 457 5026 462
rect 5278 266 5306 1751
rect 5670 1442 5698 1447
rect 5670 1395 5698 1414
rect 5390 1273 5418 1279
rect 5390 1247 5391 1273
rect 5417 1247 5418 1273
rect 5390 938 5418 1247
rect 5390 905 5418 910
rect 5670 938 5698 943
rect 5670 891 5698 910
rect 5782 434 5810 1974
rect 5838 994 5866 999
rect 5838 947 5866 966
rect 6006 714 6034 3262
rect 6174 3066 6202 4662
rect 7070 3906 7098 3911
rect 6790 3794 6818 3799
rect 6174 3033 6202 3038
rect 6510 3122 6538 3127
rect 6454 3009 6482 3015
rect 6454 2983 6455 3009
rect 6481 2983 6482 3009
rect 6118 2898 6146 2903
rect 6118 2851 6146 2870
rect 6118 2730 6146 2735
rect 6118 2338 6146 2702
rect 6118 2305 6146 2310
rect 6342 2618 6370 2623
rect 6342 1498 6370 2590
rect 6454 2618 6482 2983
rect 6454 2585 6482 2590
rect 6342 1465 6370 1470
rect 6398 2113 6426 2119
rect 6398 2087 6399 2113
rect 6425 2087 6426 2113
rect 6006 681 6034 686
rect 6398 658 6426 2087
rect 6510 1386 6538 3094
rect 6622 2954 6650 2959
rect 6510 1353 6538 1358
rect 6566 2506 6594 2511
rect 6566 1274 6594 2478
rect 6622 2450 6650 2926
rect 6678 2842 6706 2847
rect 6678 2795 6706 2814
rect 6622 2417 6650 2422
rect 6734 2394 6762 2399
rect 6678 2057 6706 2063
rect 6678 2031 6679 2057
rect 6705 2031 6706 2057
rect 6566 1246 6650 1274
rect 6398 625 6426 630
rect 5782 401 5810 406
rect 6510 490 6538 495
rect 5278 233 5306 238
rect 6398 210 6426 215
rect 6286 154 6314 159
rect 6174 98 6202 103
rect 6174 56 6202 70
rect 6286 56 6314 126
rect 6398 56 6426 182
rect 6510 56 6538 462
rect 6622 56 6650 1246
rect 6678 826 6706 2031
rect 6734 1554 6762 2366
rect 6790 1666 6818 3766
rect 6790 1633 6818 1638
rect 6958 3626 6986 3631
rect 6734 1521 6762 1526
rect 6678 793 6706 798
rect 6734 770 6762 775
rect 6734 56 6762 742
rect 6846 714 6874 719
rect 6846 56 6874 686
rect 6958 56 6986 3598
rect 7070 3290 7098 3878
rect 7070 3257 7098 3262
rect 7126 3682 7154 3687
rect 7126 3010 7154 3654
rect 7462 3066 7490 5502
rect 7686 4802 7714 6455
rect 8414 6425 8442 7014
rect 9198 6874 9226 6879
rect 8862 6594 8890 6599
rect 8414 6399 8415 6425
rect 8441 6399 8442 6425
rect 8414 6393 8442 6399
rect 8806 6482 8834 6487
rect 7798 5866 7826 5871
rect 7798 5809 7826 5838
rect 7798 5783 7799 5809
rect 7825 5783 7826 5809
rect 7798 5777 7826 5783
rect 8806 5753 8834 6454
rect 8862 5810 8890 6566
rect 8918 6481 8946 6487
rect 8918 6455 8919 6481
rect 8945 6455 8946 6481
rect 8918 6426 8946 6455
rect 8918 6393 8946 6398
rect 8862 5777 8890 5782
rect 9086 5978 9114 5983
rect 9086 5809 9114 5950
rect 9086 5783 9087 5809
rect 9113 5783 9114 5809
rect 9086 5777 9114 5783
rect 8806 5727 8807 5753
rect 8833 5727 8834 5753
rect 8806 5721 8834 5727
rect 8358 5194 8386 5199
rect 7686 4769 7714 4774
rect 7798 4913 7826 4919
rect 7798 4887 7799 4913
rect 7825 4887 7826 4913
rect 7462 3033 7490 3038
rect 7126 2977 7154 2982
rect 7182 2898 7210 2903
rect 7070 2674 7098 2679
rect 7070 2617 7098 2646
rect 7070 2591 7071 2617
rect 7097 2591 7098 2617
rect 7070 2585 7098 2591
rect 7070 994 7098 999
rect 7070 56 7098 966
rect 7182 56 7210 2870
rect 7518 2842 7546 2847
rect 7350 2562 7378 2567
rect 7350 2515 7378 2534
rect 7294 826 7322 831
rect 7294 56 7322 798
rect 7406 826 7434 831
rect 7406 56 7434 798
rect 7518 56 7546 2814
rect 7630 2562 7658 2567
rect 7630 56 7658 2534
rect 7798 1694 7826 4887
rect 8358 4914 8386 5166
rect 8358 4881 8386 4886
rect 8078 4857 8106 4863
rect 8078 4831 8079 4857
rect 8105 4831 8106 4857
rect 8078 4634 8106 4831
rect 8078 4601 8106 4606
rect 8302 4466 8330 4471
rect 7966 3514 7994 3519
rect 7742 1666 7826 1694
rect 7854 3345 7882 3351
rect 7854 3319 7855 3345
rect 7881 3319 7882 3345
rect 7742 56 7770 1666
rect 7854 56 7882 3319
rect 7966 56 7994 3486
rect 8022 3289 8050 3295
rect 8022 3263 8023 3289
rect 8049 3263 8050 3289
rect 8022 1162 8050 3263
rect 8190 2954 8218 2959
rect 8022 1129 8050 1134
rect 8078 2898 8106 2903
rect 8078 56 8106 2870
rect 8190 56 8218 2926
rect 8302 1722 8330 4438
rect 8750 4354 8778 4359
rect 8358 4242 8386 4247
rect 8358 3850 8386 4214
rect 8358 3817 8386 3822
rect 8414 3345 8442 3351
rect 8414 3319 8415 3345
rect 8441 3319 8442 3345
rect 8358 2450 8386 2455
rect 8358 2338 8386 2422
rect 8358 2305 8386 2310
rect 8302 1689 8330 1694
rect 8414 1694 8442 3319
rect 8638 3289 8666 3295
rect 8638 3263 8639 3289
rect 8665 3263 8666 3289
rect 8526 2842 8554 2847
rect 8414 1666 8498 1694
rect 8470 826 8498 1666
rect 8470 793 8498 798
rect 8414 490 8442 495
rect 8302 98 8330 103
rect 8302 56 8330 70
rect 8414 56 8442 462
rect 8526 56 8554 2814
rect 8638 1386 8666 3263
rect 8638 1353 8666 1358
rect 8694 1218 8722 1223
rect 8638 826 8666 831
rect 8638 56 8666 798
rect 8694 714 8722 1190
rect 8750 882 8778 4326
rect 9198 3122 9226 6846
rect 9422 6425 9450 7056
rect 10654 7042 10682 7056
rect 10654 7009 10682 7014
rect 10878 7042 10906 7047
rect 9758 6482 9786 6487
rect 9758 6435 9786 6454
rect 9422 6399 9423 6425
rect 9449 6399 9450 6425
rect 9422 6393 9450 6399
rect 10878 6425 10906 7014
rect 11886 7042 11914 7056
rect 11886 7009 11914 7014
rect 12110 7042 12138 7047
rect 10878 6399 10879 6425
rect 10905 6399 10906 6425
rect 10878 6393 10906 6399
rect 11270 6481 11298 6487
rect 11270 6455 11271 6481
rect 11297 6455 11298 6481
rect 10934 6090 10962 6095
rect 10150 6034 10178 6039
rect 9534 5642 9562 5647
rect 9310 4578 9338 4583
rect 9198 3089 9226 3094
rect 9254 4129 9282 4135
rect 9254 4103 9255 4129
rect 9281 4103 9282 4129
rect 9254 2898 9282 4103
rect 9310 4130 9338 4550
rect 9310 4097 9338 4102
rect 9478 4073 9506 4079
rect 9478 4047 9479 4073
rect 9505 4047 9506 4073
rect 9478 4018 9506 4047
rect 9478 3985 9506 3990
rect 9254 2865 9282 2870
rect 9366 3178 9394 3183
rect 8806 2561 8834 2567
rect 8806 2535 8807 2561
rect 8833 2535 8834 2561
rect 8806 938 8834 2535
rect 8974 2506 9002 2511
rect 8918 2505 9002 2506
rect 8918 2479 8975 2505
rect 9001 2479 9002 2505
rect 8918 2478 9002 2479
rect 8918 1274 8946 2478
rect 8974 2473 9002 2478
rect 9198 2058 9226 2063
rect 9198 1833 9226 2030
rect 9198 1807 9199 1833
rect 9225 1807 9226 1833
rect 9198 1801 9226 1807
rect 9254 2002 9282 2007
rect 8974 1777 9002 1783
rect 8974 1751 8975 1777
rect 9001 1751 9002 1777
rect 8974 1694 9002 1751
rect 8974 1666 9114 1694
rect 8918 1246 9058 1274
rect 8806 910 9002 938
rect 8750 854 8890 882
rect 8694 686 8778 714
rect 8750 56 8778 686
rect 8862 56 8890 854
rect 8974 56 9002 910
rect 9030 770 9058 1246
rect 9030 737 9058 742
rect 9086 56 9114 1666
rect 9142 994 9170 999
rect 9142 993 9226 994
rect 9142 967 9143 993
rect 9169 967 9226 993
rect 9142 966 9226 967
rect 9142 961 9170 966
rect 9198 56 9226 966
rect 9254 546 9282 1974
rect 9366 1049 9394 3150
rect 9366 1023 9367 1049
rect 9393 1023 9394 1049
rect 9366 1017 9394 1023
rect 9422 1274 9450 1279
rect 9254 513 9282 518
rect 9310 322 9338 327
rect 9310 56 9338 294
rect 9422 56 9450 1246
rect 9534 56 9562 5614
rect 10094 5026 10122 5031
rect 9646 4913 9674 4919
rect 9646 4887 9647 4913
rect 9673 4887 9674 4913
rect 9646 3514 9674 4887
rect 9926 4857 9954 4863
rect 9926 4831 9927 4857
rect 9953 4831 9954 4857
rect 9646 3481 9674 3486
rect 9870 3626 9898 3631
rect 9646 3346 9674 3351
rect 9646 56 9674 3318
rect 9758 1946 9786 1951
rect 9758 56 9786 1918
rect 9870 56 9898 3598
rect 9926 546 9954 4831
rect 10038 3962 10066 3967
rect 9982 3514 10010 3519
rect 9982 2506 10010 3486
rect 9982 2473 10010 2478
rect 10038 1694 10066 3934
rect 10094 3402 10122 4998
rect 10150 4466 10178 6006
rect 10150 4433 10178 4438
rect 10262 5586 10290 5591
rect 10094 3369 10122 3374
rect 10150 3794 10178 3799
rect 10150 1694 10178 3766
rect 9926 513 9954 518
rect 9982 1666 10066 1694
rect 10094 1666 10178 1694
rect 10206 2506 10234 2511
rect 9982 56 10010 1666
rect 10094 56 10122 1666
rect 10206 56 10234 2478
rect 10262 1442 10290 5558
rect 10710 5362 10738 5367
rect 10486 5082 10514 5087
rect 10486 4858 10514 5054
rect 10486 4825 10514 4830
rect 10654 3906 10682 3911
rect 10598 3010 10626 3015
rect 10486 2450 10514 2455
rect 10486 2282 10514 2422
rect 10486 2249 10514 2254
rect 10262 1409 10290 1414
rect 10318 994 10346 999
rect 10262 602 10290 607
rect 10262 555 10290 574
rect 10318 56 10346 966
rect 10374 993 10402 999
rect 10374 967 10375 993
rect 10401 967 10402 993
rect 10374 322 10402 967
rect 10486 546 10514 551
rect 10374 289 10402 294
rect 10430 518 10486 546
rect 10430 56 10458 518
rect 10486 513 10514 518
rect 10598 378 10626 2982
rect 10654 1049 10682 3878
rect 10654 1023 10655 1049
rect 10681 1023 10682 1049
rect 10654 1017 10682 1023
rect 10710 882 10738 5334
rect 10934 4690 10962 6062
rect 11214 5362 11242 5367
rect 11270 5362 11298 6455
rect 12110 6425 12138 7014
rect 12232 6678 12364 6683
rect 12260 6650 12284 6678
rect 12312 6650 12336 6678
rect 12232 6645 12364 6650
rect 12110 6399 12111 6425
rect 12137 6399 12138 6425
rect 12110 6393 12138 6399
rect 12502 6481 12530 6487
rect 12502 6455 12503 6481
rect 12529 6455 12530 6481
rect 11494 6370 11522 6375
rect 11494 5866 11522 6342
rect 11902 6286 12034 6291
rect 11930 6258 11954 6286
rect 11982 6258 12006 6286
rect 11902 6253 12034 6258
rect 11494 5833 11522 5838
rect 11550 6202 11578 6207
rect 11214 5361 11298 5362
rect 11214 5335 11215 5361
rect 11241 5335 11298 5361
rect 11214 5334 11298 5335
rect 11214 5329 11242 5334
rect 10934 4657 10962 4662
rect 11046 5306 11074 5311
rect 10934 4522 10962 4527
rect 10934 3682 10962 4494
rect 10934 3649 10962 3654
rect 10990 3626 11018 3631
rect 10990 3579 11018 3598
rect 10934 2674 10962 2679
rect 10934 2282 10962 2646
rect 11046 2338 11074 5278
rect 11438 5193 11466 5199
rect 11438 5167 11439 5193
rect 11465 5167 11466 5193
rect 11438 4970 11466 5167
rect 11438 4937 11466 4942
rect 11270 3682 11298 3687
rect 11270 3635 11298 3654
rect 11550 3458 11578 6174
rect 12232 5894 12364 5899
rect 12260 5866 12284 5894
rect 12312 5866 12336 5894
rect 12232 5861 12364 5866
rect 12110 5642 12138 5647
rect 12110 5530 12138 5614
rect 12502 5641 12530 6455
rect 12614 6482 12642 6487
rect 12502 5615 12503 5641
rect 12529 5615 12530 5641
rect 12502 5609 12530 5615
rect 12558 5642 12586 5647
rect 11902 5502 12034 5507
rect 11930 5474 11954 5502
rect 11982 5474 12006 5502
rect 12110 5497 12138 5502
rect 11902 5469 12034 5474
rect 12558 5306 12586 5614
rect 12502 5278 12586 5306
rect 12614 5306 12642 6454
rect 13118 6425 13146 7056
rect 14350 7042 14378 7056
rect 14350 7009 14378 7014
rect 14574 7042 14602 7047
rect 14126 6594 14154 6599
rect 13118 6399 13119 6425
rect 13145 6399 13146 6425
rect 13118 6393 13146 6399
rect 13454 6481 13482 6487
rect 13454 6455 13455 6481
rect 13481 6455 13482 6481
rect 11718 5138 11746 5143
rect 12446 5138 12474 5143
rect 11606 4466 11634 4471
rect 11606 3906 11634 4438
rect 11718 4186 11746 5110
rect 12232 5110 12364 5115
rect 12260 5082 12284 5110
rect 12312 5082 12336 5110
rect 12232 5077 12364 5082
rect 11902 4718 12034 4723
rect 11930 4690 11954 4718
rect 11982 4690 12006 4718
rect 11902 4685 12034 4690
rect 12446 4578 12474 5110
rect 12446 4545 12474 4550
rect 11718 4153 11746 4158
rect 12110 4354 12138 4359
rect 11606 3873 11634 3878
rect 11662 4130 11690 4135
rect 11494 3430 11578 3458
rect 11046 2305 11074 2310
rect 11102 2674 11130 2679
rect 10934 2249 10962 2254
rect 10990 1442 11018 1447
rect 10542 350 10626 378
rect 10654 854 10738 882
rect 10878 882 10906 887
rect 10542 56 10570 350
rect 10654 56 10682 854
rect 10766 658 10794 663
rect 10766 657 10850 658
rect 10766 631 10767 657
rect 10793 631 10850 657
rect 10766 630 10850 631
rect 10766 625 10794 630
rect 10822 154 10850 630
rect 10822 121 10850 126
rect 10766 98 10794 103
rect 10766 56 10794 70
rect 10878 56 10906 854
rect 10990 56 11018 1414
rect 11046 658 11074 663
rect 11046 601 11074 630
rect 11046 575 11047 601
rect 11073 575 11074 601
rect 11046 569 11074 575
rect 11102 56 11130 2646
rect 11270 2618 11298 2623
rect 11214 2562 11242 2567
rect 11158 1330 11186 1335
rect 11158 826 11186 1302
rect 11158 793 11186 798
rect 11214 56 11242 2534
rect 11270 378 11298 2590
rect 11382 1834 11410 1839
rect 11382 1787 11410 1806
rect 11438 1778 11466 1783
rect 11438 1386 11466 1750
rect 11382 1358 11466 1386
rect 11326 1274 11354 1279
rect 11326 1227 11354 1246
rect 11382 1162 11410 1358
rect 11494 1330 11522 3430
rect 11662 3234 11690 4102
rect 11774 4129 11802 4135
rect 11774 4103 11775 4129
rect 11801 4103 11802 4129
rect 11774 3962 11802 4103
rect 11998 4074 12026 4079
rect 11998 4027 12026 4046
rect 11774 3929 11802 3934
rect 11902 3934 12034 3939
rect 11930 3906 11954 3934
rect 11982 3906 12006 3934
rect 11902 3901 12034 3906
rect 12110 3906 12138 4326
rect 12232 4326 12364 4331
rect 12260 4298 12284 4326
rect 12312 4298 12336 4326
rect 12232 4293 12364 4298
rect 12110 3873 12138 3878
rect 12502 3850 12530 5278
rect 12614 5273 12642 5278
rect 12670 5978 12698 5983
rect 12558 5194 12586 5199
rect 12558 4802 12586 5166
rect 12558 4769 12586 4774
rect 12670 4522 12698 5950
rect 12726 5698 12754 5703
rect 12726 5651 12754 5670
rect 13342 5586 13370 5591
rect 12726 5362 12754 5367
rect 12726 4634 12754 5334
rect 13342 5250 13370 5558
rect 13398 5362 13426 5367
rect 13454 5362 13482 6455
rect 13398 5361 13482 5362
rect 13398 5335 13399 5361
rect 13425 5335 13482 5361
rect 13398 5334 13482 5335
rect 13790 6370 13818 6375
rect 13398 5329 13426 5334
rect 13342 5222 13426 5250
rect 13398 4746 13426 5222
rect 13622 5194 13650 5199
rect 13622 5147 13650 5166
rect 13398 4713 13426 4718
rect 12726 4601 12754 4606
rect 12670 4489 12698 4494
rect 13678 4298 13706 4303
rect 13678 4186 13706 4270
rect 13678 4153 13706 4158
rect 13790 4186 13818 6342
rect 13902 5866 13930 5871
rect 13902 5586 13930 5838
rect 14126 5698 14154 6566
rect 14574 6425 14602 7014
rect 15582 7042 15610 7056
rect 15582 7009 15610 7014
rect 15862 7042 15890 7047
rect 14574 6399 14575 6425
rect 14601 6399 14602 6425
rect 14574 6393 14602 6399
rect 14742 6874 14770 6879
rect 14126 5665 14154 5670
rect 13902 5553 13930 5558
rect 13790 4153 13818 4158
rect 14014 5474 14042 5479
rect 13678 4018 13706 4023
rect 12502 3817 12530 3822
rect 13398 3906 13426 3911
rect 12278 3794 12306 3799
rect 12278 3737 12306 3766
rect 12278 3711 12279 3737
rect 12305 3711 12306 3737
rect 12278 3705 12306 3711
rect 12558 3681 12586 3687
rect 12558 3655 12559 3681
rect 12585 3655 12586 3681
rect 12232 3542 12364 3547
rect 12260 3514 12284 3542
rect 12312 3514 12336 3542
rect 12232 3509 12364 3514
rect 12558 3402 12586 3655
rect 12670 3626 12698 3631
rect 12558 3369 12586 3374
rect 12614 3514 12642 3519
rect 11662 3201 11690 3206
rect 11902 3150 12034 3155
rect 11930 3122 11954 3150
rect 11982 3122 12006 3150
rect 11902 3117 12034 3122
rect 12614 3066 12642 3486
rect 12614 3033 12642 3038
rect 12166 2786 12194 2791
rect 12670 2786 12698 3598
rect 13006 3402 13034 3407
rect 12166 2394 12194 2758
rect 12232 2758 12364 2763
rect 12260 2730 12284 2758
rect 12312 2730 12336 2758
rect 12670 2753 12698 2758
rect 12782 2954 12810 2959
rect 12232 2725 12364 2730
rect 12782 2673 12810 2926
rect 12782 2647 12783 2673
rect 12809 2647 12810 2673
rect 12782 2641 12810 2647
rect 12894 2898 12922 2903
rect 12670 2506 12698 2511
rect 11902 2366 12034 2371
rect 11930 2338 11954 2366
rect 11982 2338 12006 2366
rect 12166 2361 12194 2366
rect 12558 2394 12586 2399
rect 11902 2333 12034 2338
rect 12110 2338 12138 2343
rect 11830 2170 11858 2175
rect 11830 2123 11858 2142
rect 11998 2114 12026 2119
rect 12110 2114 12138 2310
rect 11998 2067 12026 2086
rect 12054 2086 12138 2114
rect 11550 2057 11578 2063
rect 11550 2031 11551 2057
rect 11577 2031 11578 2057
rect 11550 1946 11578 2031
rect 12054 2002 12082 2086
rect 12278 2058 12306 2063
rect 12054 1969 12082 1974
rect 12110 2057 12306 2058
rect 12110 2031 12279 2057
rect 12305 2031 12306 2057
rect 12110 2030 12306 2031
rect 11550 1913 11578 1918
rect 11494 1297 11522 1302
rect 11550 1834 11578 1839
rect 11494 1162 11522 1167
rect 11382 1134 11466 1162
rect 11382 1050 11410 1055
rect 11382 1003 11410 1022
rect 11270 350 11354 378
rect 11326 56 11354 350
rect 11438 56 11466 1134
rect 11494 1050 11522 1134
rect 11494 1017 11522 1022
rect 11494 657 11522 663
rect 11494 631 11495 657
rect 11521 631 11522 657
rect 11494 266 11522 631
rect 11494 233 11522 238
rect 11550 56 11578 1806
rect 11830 1721 11858 1727
rect 11830 1695 11831 1721
rect 11857 1695 11858 1721
rect 11774 1386 11802 1391
rect 11774 1339 11802 1358
rect 11606 1330 11634 1335
rect 11606 1283 11634 1302
rect 11774 1274 11802 1279
rect 11774 1050 11802 1246
rect 11718 1022 11802 1050
rect 11718 602 11746 1022
rect 11662 574 11746 602
rect 11774 937 11802 943
rect 11774 911 11775 937
rect 11801 911 11802 937
rect 11662 56 11690 574
rect 11774 322 11802 911
rect 11830 714 11858 1695
rect 11902 1582 12034 1587
rect 11930 1554 11954 1582
rect 11982 1554 12006 1582
rect 11902 1549 12034 1554
rect 11998 1442 12026 1447
rect 11998 1218 12026 1414
rect 11998 1185 12026 1190
rect 11902 798 12034 803
rect 11930 770 11954 798
rect 11982 770 12006 798
rect 11902 765 12034 770
rect 11830 686 12026 714
rect 11774 289 11802 294
rect 11886 490 11914 495
rect 11774 210 11802 215
rect 11774 56 11802 182
rect 11886 56 11914 462
rect 11998 56 12026 686
rect 12110 322 12138 2030
rect 12278 2025 12306 2030
rect 12232 1974 12364 1979
rect 12260 1946 12284 1974
rect 12312 1946 12336 1974
rect 12232 1941 12364 1946
rect 12558 1694 12586 2366
rect 12670 2394 12698 2478
rect 12670 2361 12698 2366
rect 12782 2226 12810 2231
rect 12782 2169 12810 2198
rect 12894 2226 12922 2870
rect 13006 2394 13034 3374
rect 13398 3290 13426 3878
rect 13398 3257 13426 3262
rect 13622 3345 13650 3351
rect 13622 3319 13623 3345
rect 13649 3319 13650 3345
rect 13230 3178 13258 3183
rect 13062 2506 13090 2511
rect 13062 2459 13090 2478
rect 13006 2366 13146 2394
rect 12894 2193 12922 2198
rect 12782 2143 12783 2169
rect 12809 2143 12810 2169
rect 12782 2137 12810 2143
rect 13062 2058 13090 2063
rect 12894 2057 13090 2058
rect 12894 2031 13063 2057
rect 13089 2031 13090 2057
rect 12894 2030 13090 2031
rect 12838 2002 12866 2007
rect 12838 1833 12866 1974
rect 12838 1807 12839 1833
rect 12865 1807 12866 1833
rect 12838 1801 12866 1807
rect 12614 1778 12642 1797
rect 12614 1745 12642 1750
rect 12894 1694 12922 2030
rect 13062 2025 13090 2030
rect 13006 1890 13034 1895
rect 13006 1833 13034 1862
rect 13006 1807 13007 1833
rect 13033 1807 13034 1833
rect 13006 1801 13034 1807
rect 13118 1694 13146 2366
rect 12558 1666 12642 1694
rect 12614 1633 12642 1638
rect 12670 1666 12922 1694
rect 13062 1666 13146 1694
rect 12614 1385 12642 1391
rect 12614 1359 12615 1385
rect 12641 1359 12642 1385
rect 12166 1329 12194 1335
rect 12166 1303 12167 1329
rect 12193 1303 12194 1329
rect 12166 658 12194 1303
rect 12232 1190 12364 1195
rect 12260 1162 12284 1190
rect 12312 1162 12336 1190
rect 12232 1157 12364 1162
rect 12502 993 12530 999
rect 12502 967 12503 993
rect 12529 967 12530 993
rect 12166 630 12474 658
rect 12166 545 12194 551
rect 12166 519 12167 545
rect 12193 519 12194 545
rect 12166 434 12194 519
rect 12166 401 12194 406
rect 12232 406 12364 411
rect 12260 378 12284 406
rect 12312 378 12336 406
rect 12232 373 12364 378
rect 12334 322 12362 327
rect 12110 294 12250 322
rect 12110 154 12138 159
rect 12110 56 12138 126
rect 12222 56 12250 294
rect 12334 56 12362 294
rect 12446 56 12474 630
rect 12502 210 12530 967
rect 12614 938 12642 1359
rect 12614 905 12642 910
rect 12558 546 12586 551
rect 12558 499 12586 518
rect 12502 177 12530 182
rect 12558 266 12586 271
rect 12558 56 12586 238
rect 12670 56 12698 1666
rect 12950 1554 12978 1559
rect 12838 1274 12866 1279
rect 12782 1273 12866 1274
rect 12782 1247 12839 1273
rect 12865 1247 12866 1273
rect 12782 1246 12866 1247
rect 12726 938 12754 943
rect 12726 891 12754 910
rect 12782 56 12810 1246
rect 12838 1241 12866 1246
rect 12894 1106 12922 1111
rect 12894 1049 12922 1078
rect 12894 1023 12895 1049
rect 12921 1023 12922 1049
rect 12894 1017 12922 1023
rect 12838 994 12866 999
rect 12838 882 12866 966
rect 12838 849 12866 854
rect 12894 602 12922 607
rect 12894 56 12922 574
rect 12950 154 12978 1526
rect 12950 121 12978 126
rect 13006 546 13034 551
rect 13006 56 13034 518
rect 13062 266 13090 1666
rect 13230 1106 13258 3150
rect 13398 2506 13426 2511
rect 13230 1073 13258 1078
rect 13286 1665 13314 1671
rect 13286 1639 13287 1665
rect 13313 1639 13314 1665
rect 13174 882 13202 887
rect 13062 233 13090 238
rect 13118 881 13202 882
rect 13118 855 13175 881
rect 13201 855 13202 881
rect 13118 854 13202 855
rect 13118 56 13146 854
rect 13174 849 13202 854
rect 13230 714 13258 719
rect 13230 56 13258 686
rect 13286 602 13314 1639
rect 13342 1498 13370 1503
rect 13342 1385 13370 1470
rect 13342 1359 13343 1385
rect 13369 1359 13370 1385
rect 13342 1353 13370 1359
rect 13286 569 13314 574
rect 13398 602 13426 2478
rect 13454 1778 13482 1783
rect 13454 826 13482 1750
rect 13622 1554 13650 3319
rect 13622 1521 13650 1526
rect 13454 793 13482 798
rect 13510 1498 13538 1503
rect 13510 658 13538 1470
rect 13622 1273 13650 1279
rect 13622 1247 13623 1273
rect 13649 1247 13650 1273
rect 13622 714 13650 1247
rect 13678 1049 13706 3990
rect 13902 3626 13930 3631
rect 13846 3290 13874 3295
rect 13678 1023 13679 1049
rect 13705 1023 13706 1049
rect 13678 1017 13706 1023
rect 13734 3289 13874 3290
rect 13734 3263 13847 3289
rect 13873 3263 13874 3289
rect 13734 3262 13874 3263
rect 13622 681 13650 686
rect 13510 625 13538 630
rect 13398 569 13426 574
rect 13566 602 13594 607
rect 13734 602 13762 3262
rect 13846 3257 13874 3262
rect 13790 2786 13818 2791
rect 13790 1554 13818 2758
rect 13790 1521 13818 1526
rect 13902 1218 13930 3598
rect 14014 2450 14042 5446
rect 14238 5138 14266 5143
rect 14126 4802 14154 4807
rect 14126 4522 14154 4774
rect 14238 4802 14266 5110
rect 14350 5138 14378 5143
rect 14350 4970 14378 5110
rect 14350 4937 14378 4942
rect 14238 4769 14266 4774
rect 14686 4746 14714 4751
rect 14126 4489 14154 4494
rect 14350 4690 14378 4695
rect 14014 2417 14042 2422
rect 14238 3794 14266 3799
rect 14238 1946 14266 3766
rect 14294 2169 14322 2175
rect 14294 2143 14295 2169
rect 14321 2143 14322 2169
rect 14294 2058 14322 2143
rect 14294 2025 14322 2030
rect 14238 1918 14322 1946
rect 14126 1834 14154 1839
rect 14238 1834 14266 1839
rect 14126 1787 14154 1806
rect 14182 1806 14238 1834
rect 14182 1694 14210 1806
rect 14238 1801 14266 1806
rect 14294 1722 14322 1918
rect 13902 1185 13930 1190
rect 14070 1666 14210 1694
rect 14238 1694 14322 1722
rect 13958 882 13986 887
rect 13566 601 13762 602
rect 13566 575 13567 601
rect 13593 575 13762 601
rect 13566 574 13762 575
rect 13790 881 13986 882
rect 13790 855 13959 881
rect 13985 855 13986 881
rect 13790 854 13986 855
rect 13566 569 13594 574
rect 13286 490 13314 495
rect 13454 490 13482 495
rect 13286 489 13370 490
rect 13286 463 13287 489
rect 13313 463 13370 489
rect 13286 462 13370 463
rect 13286 457 13314 462
rect 13342 56 13370 462
rect 13454 56 13482 462
rect 13510 434 13538 439
rect 13790 434 13818 854
rect 13958 849 13986 854
rect 14014 826 14042 831
rect 13902 658 13930 663
rect 13846 602 13874 607
rect 13846 555 13874 574
rect 13510 322 13538 406
rect 13510 289 13538 294
rect 13566 406 13818 434
rect 13566 56 13594 406
rect 13790 322 13818 327
rect 13678 266 13706 271
rect 13678 56 13706 238
rect 13790 56 13818 294
rect 13902 56 13930 630
rect 14014 56 14042 798
rect 14070 434 14098 1666
rect 14238 602 14266 1694
rect 14350 1385 14378 4662
rect 14518 2506 14546 2511
rect 14518 2225 14546 2478
rect 14686 2338 14714 4718
rect 14686 2305 14714 2310
rect 14518 2199 14519 2225
rect 14545 2199 14546 2225
rect 14518 2193 14546 2199
rect 14686 2170 14714 2175
rect 14686 2123 14714 2142
rect 14574 2058 14602 2063
rect 14350 1359 14351 1385
rect 14377 1359 14378 1385
rect 14350 1353 14378 1359
rect 14406 1665 14434 1671
rect 14406 1639 14407 1665
rect 14433 1639 14434 1665
rect 14406 1274 14434 1639
rect 14350 1246 14434 1274
rect 14518 1273 14546 1279
rect 14518 1247 14519 1273
rect 14545 1247 14546 1273
rect 14350 826 14378 1246
rect 14350 793 14378 798
rect 14406 1162 14434 1167
rect 14182 574 14266 602
rect 14350 602 14378 607
rect 14126 490 14154 495
rect 14126 443 14154 462
rect 14070 401 14098 406
rect 14182 378 14210 574
rect 14182 345 14210 350
rect 14238 490 14266 495
rect 14126 210 14154 215
rect 14126 56 14154 182
rect 14238 56 14266 462
rect 14350 56 14378 574
rect 14406 546 14434 1134
rect 14462 1050 14490 1055
rect 14462 1003 14490 1022
rect 14406 513 14434 518
rect 14462 714 14490 719
rect 14462 56 14490 686
rect 14518 658 14546 1247
rect 14518 625 14546 630
rect 14574 56 14602 2030
rect 14742 1106 14770 6846
rect 15246 6762 15274 6767
rect 14966 6482 14994 6487
rect 14854 6481 14994 6482
rect 14854 6455 14967 6481
rect 14993 6455 14994 6481
rect 14854 6454 14994 6455
rect 14854 6145 14882 6454
rect 14966 6449 14994 6454
rect 14854 6119 14855 6145
rect 14881 6119 14882 6145
rect 14854 6113 14882 6119
rect 15246 6145 15274 6734
rect 15862 6425 15890 7014
rect 15862 6399 15863 6425
rect 15889 6399 15890 6425
rect 15862 6393 15890 6399
rect 16366 6481 16394 6487
rect 16366 6455 16367 6481
rect 16393 6455 16394 6481
rect 15246 6119 15247 6145
rect 15273 6119 15274 6145
rect 15246 6113 15274 6119
rect 16366 6146 16394 6455
rect 16366 6113 16394 6118
rect 16590 6426 16618 6431
rect 16814 6426 16842 7056
rect 18046 7042 18074 7056
rect 18046 7009 18074 7014
rect 18270 7042 18298 7047
rect 17374 6481 17402 6487
rect 17374 6455 17375 6481
rect 17401 6455 17402 6481
rect 16870 6426 16898 6431
rect 16814 6425 16898 6426
rect 16814 6399 16871 6425
rect 16897 6399 16898 6425
rect 16814 6398 16898 6399
rect 16590 6145 16618 6398
rect 16870 6393 16898 6398
rect 16590 6119 16591 6145
rect 16617 6119 16618 6145
rect 16590 6113 16618 6119
rect 17038 6146 17066 6151
rect 17038 6099 17066 6118
rect 15022 6090 15050 6095
rect 14966 6089 15050 6090
rect 14966 6063 15023 6089
rect 15049 6063 15050 6089
rect 14966 6062 15050 6063
rect 14798 6034 14826 6039
rect 14798 5642 14826 6006
rect 14798 5609 14826 5614
rect 14854 5922 14882 5927
rect 14854 4970 14882 5894
rect 14854 4937 14882 4942
rect 14910 5754 14938 5759
rect 14910 4466 14938 5726
rect 14910 4433 14938 4438
rect 14966 4354 14994 6062
rect 15022 6057 15050 6062
rect 15918 6090 15946 6095
rect 15526 5977 15554 5983
rect 15526 5951 15527 5977
rect 15553 5951 15554 5977
rect 15134 5810 15162 5815
rect 14966 4321 14994 4326
rect 15022 5418 15050 5423
rect 14910 4298 14938 4303
rect 14910 4242 14938 4270
rect 14910 4214 14994 4242
rect 14854 4074 14882 4079
rect 14798 2561 14826 2567
rect 14798 2535 14799 2561
rect 14825 2535 14826 2561
rect 14798 1162 14826 2535
rect 14854 1694 14882 4046
rect 14910 3682 14938 3687
rect 14910 1833 14938 3654
rect 14966 3346 14994 4214
rect 15022 3850 15050 5390
rect 15078 5362 15106 5367
rect 15078 4522 15106 5334
rect 15078 4489 15106 4494
rect 15134 4185 15162 5782
rect 15134 4159 15135 4185
rect 15161 4159 15162 4185
rect 15134 4153 15162 4159
rect 15190 5530 15218 5535
rect 15022 3817 15050 3822
rect 15078 4018 15106 4023
rect 14966 3313 14994 3318
rect 15078 3010 15106 3990
rect 15078 2977 15106 2982
rect 15134 2954 15162 2959
rect 15190 2954 15218 5502
rect 15526 5082 15554 5951
rect 15918 5810 15946 6062
rect 16870 6034 16898 6039
rect 16870 5987 16898 6006
rect 15918 5777 15946 5782
rect 16086 5977 16114 5983
rect 16086 5951 16087 5977
rect 16113 5951 16114 5977
rect 15526 5049 15554 5054
rect 15974 5418 16002 5423
rect 15470 4578 15498 4583
rect 15246 4186 15274 4191
rect 15246 3178 15274 4158
rect 15414 4129 15442 4135
rect 15414 4103 15415 4129
rect 15441 4103 15442 4129
rect 15414 3402 15442 4103
rect 15414 3369 15442 3374
rect 15302 3345 15330 3351
rect 15302 3319 15303 3345
rect 15329 3319 15330 3345
rect 15302 3290 15330 3319
rect 15302 3257 15330 3262
rect 15246 3150 15330 3178
rect 15134 2953 15218 2954
rect 15134 2927 15135 2953
rect 15161 2927 15218 2953
rect 15134 2926 15218 2927
rect 15134 2921 15162 2926
rect 15246 2898 15274 2903
rect 15246 2617 15274 2870
rect 15246 2591 15247 2617
rect 15273 2591 15274 2617
rect 15246 2585 15274 2591
rect 15078 2562 15106 2567
rect 15078 2515 15106 2534
rect 15134 2450 15162 2455
rect 14966 2058 14994 2063
rect 14966 2011 14994 2030
rect 14910 1807 14911 1833
rect 14937 1807 14938 1833
rect 14910 1801 14938 1807
rect 14854 1666 14938 1694
rect 14910 1638 15050 1666
rect 15022 1385 15050 1638
rect 15022 1359 15023 1385
rect 15049 1359 15050 1385
rect 15022 1353 15050 1359
rect 14798 1129 14826 1134
rect 14742 1073 14770 1078
rect 15022 1050 15050 1055
rect 14742 881 14770 887
rect 14742 855 14743 881
rect 14769 855 14770 881
rect 14630 770 14658 775
rect 14630 601 14658 742
rect 14630 575 14631 601
rect 14657 575 14658 601
rect 14630 569 14658 575
rect 14686 546 14714 551
rect 14686 56 14714 518
rect 14742 322 14770 855
rect 14742 289 14770 294
rect 14798 658 14826 663
rect 14798 56 14826 630
rect 14910 490 14938 495
rect 14854 489 14938 490
rect 14854 463 14911 489
rect 14937 463 14938 489
rect 14854 462 14938 463
rect 14854 266 14882 462
rect 14910 457 14938 462
rect 14854 233 14882 238
rect 14910 378 14938 383
rect 14910 56 14938 350
rect 15022 56 15050 1022
rect 15134 56 15162 2422
rect 15190 1665 15218 1671
rect 15190 1639 15191 1665
rect 15217 1639 15218 1665
rect 15190 714 15218 1639
rect 15246 1666 15274 1671
rect 15246 1049 15274 1638
rect 15302 1386 15330 3150
rect 15358 2898 15386 2903
rect 15358 2897 15442 2898
rect 15358 2871 15359 2897
rect 15385 2871 15442 2897
rect 15358 2870 15442 2871
rect 15358 2865 15386 2870
rect 15358 2618 15386 2623
rect 15358 1946 15386 2590
rect 15414 2002 15442 2870
rect 15470 2169 15498 4550
rect 15862 4298 15890 4303
rect 15582 3289 15610 3295
rect 15582 3263 15583 3289
rect 15609 3263 15610 3289
rect 15582 2730 15610 3263
rect 15638 3234 15666 3239
rect 15638 2953 15666 3206
rect 15638 2927 15639 2953
rect 15665 2927 15666 2953
rect 15638 2921 15666 2927
rect 15750 3010 15778 3015
rect 15582 2697 15610 2702
rect 15526 2450 15554 2455
rect 15526 2403 15554 2422
rect 15470 2143 15471 2169
rect 15497 2143 15498 2169
rect 15470 2137 15498 2143
rect 15694 2226 15722 2231
rect 15694 2002 15722 2198
rect 15414 1974 15498 2002
rect 15358 1918 15442 1946
rect 15302 1353 15330 1358
rect 15358 1722 15386 1727
rect 15246 1023 15247 1049
rect 15273 1023 15274 1049
rect 15246 1017 15274 1023
rect 15302 1273 15330 1279
rect 15302 1247 15303 1273
rect 15329 1247 15330 1273
rect 15190 681 15218 686
rect 15302 602 15330 1247
rect 15302 569 15330 574
rect 15246 322 15274 327
rect 15246 56 15274 294
rect 15358 56 15386 1694
rect 15414 1442 15442 1918
rect 15470 1610 15498 1974
rect 15694 1969 15722 1974
rect 15750 1834 15778 2982
rect 15750 1801 15778 1806
rect 15806 3009 15834 3015
rect 15806 2983 15807 3009
rect 15833 2983 15834 3009
rect 15806 1694 15834 2983
rect 15862 2450 15890 4270
rect 15974 3514 16002 5390
rect 16086 5026 16114 5951
rect 16254 5977 16282 5983
rect 16254 5951 16255 5977
rect 16281 5951 16282 5977
rect 16086 4993 16114 4998
rect 16142 5642 16170 5647
rect 15974 3481 16002 3486
rect 16030 4578 16058 4583
rect 16030 3402 16058 4550
rect 15862 2417 15890 2422
rect 15918 3374 16058 3402
rect 16086 3794 16114 3799
rect 15918 2282 15946 3374
rect 16086 3290 16114 3766
rect 16086 3257 16114 3262
rect 16030 2841 16058 2847
rect 16030 2815 16031 2841
rect 16057 2815 16058 2841
rect 16030 2618 16058 2815
rect 16030 2585 16058 2590
rect 15918 2249 15946 2254
rect 15974 2338 16002 2343
rect 15470 1577 15498 1582
rect 15750 1666 15834 1694
rect 15862 2113 15890 2119
rect 15862 2087 15863 2113
rect 15889 2087 15890 2113
rect 15414 1409 15442 1414
rect 15750 994 15778 1666
rect 15806 1610 15834 1615
rect 15806 1385 15834 1582
rect 15806 1359 15807 1385
rect 15833 1359 15834 1385
rect 15806 1353 15834 1359
rect 15862 1050 15890 2087
rect 15862 1017 15890 1022
rect 15918 1666 15946 1671
rect 15750 966 15834 994
rect 15806 938 15834 966
rect 15806 910 15890 938
rect 15526 881 15554 887
rect 15526 855 15527 881
rect 15553 855 15554 881
rect 15470 714 15498 719
rect 15470 56 15498 686
rect 15526 210 15554 855
rect 15750 882 15778 887
rect 15778 854 15834 882
rect 15750 849 15778 854
rect 15694 826 15722 831
rect 15526 177 15554 182
rect 15582 266 15610 271
rect 15582 56 15610 238
rect 15694 56 15722 798
rect 15750 545 15778 551
rect 15750 519 15751 545
rect 15777 519 15778 545
rect 15750 154 15778 519
rect 15750 121 15778 126
rect 15806 56 15834 854
rect 15862 602 15890 910
rect 15862 569 15890 574
rect 15918 56 15946 1638
rect 15974 1610 16002 2310
rect 16142 2282 16170 5614
rect 16198 4858 16226 4863
rect 16198 4811 16226 4830
rect 16254 3850 16282 5951
rect 17318 5978 17346 5983
rect 17318 5931 17346 5950
rect 16814 5586 16842 5591
rect 16702 5082 16730 5087
rect 16478 4913 16506 4919
rect 16478 4887 16479 4913
rect 16505 4887 16506 4913
rect 16478 4298 16506 4887
rect 16478 4265 16506 4270
rect 16646 4634 16674 4639
rect 16254 3817 16282 3822
rect 16310 2897 16338 2903
rect 16310 2871 16311 2897
rect 16337 2871 16338 2897
rect 16310 2618 16338 2871
rect 16310 2585 16338 2590
rect 16478 2897 16506 2903
rect 16478 2871 16479 2897
rect 16505 2871 16506 2897
rect 16198 2562 16226 2567
rect 16198 2515 16226 2534
rect 16478 2562 16506 2871
rect 16478 2529 16506 2534
rect 16534 2898 16562 2903
rect 16478 2450 16506 2455
rect 16142 2249 16170 2254
rect 16254 2449 16506 2450
rect 16254 2423 16479 2449
rect 16505 2423 16506 2449
rect 16254 2422 16506 2423
rect 16198 1778 16226 1783
rect 16198 1731 16226 1750
rect 15974 1577 16002 1582
rect 16198 1330 16226 1335
rect 16086 1273 16114 1279
rect 16086 1247 16087 1273
rect 16113 1247 16114 1273
rect 16086 658 16114 1247
rect 16198 1049 16226 1302
rect 16198 1023 16199 1049
rect 16225 1023 16226 1049
rect 16198 1017 16226 1023
rect 16086 625 16114 630
rect 16030 490 16058 495
rect 16030 443 16058 462
rect 16254 322 16282 2422
rect 16478 2417 16506 2422
rect 16534 2338 16562 2870
rect 16366 2310 16562 2338
rect 16590 2730 16618 2735
rect 16030 294 16282 322
rect 16310 2058 16338 2063
rect 16030 56 16058 294
rect 16310 266 16338 2030
rect 16254 238 16338 266
rect 16142 210 16170 215
rect 16142 56 16170 182
rect 16254 56 16282 238
rect 16366 56 16394 2310
rect 16422 2225 16450 2231
rect 16422 2199 16423 2225
rect 16449 2199 16450 2225
rect 16422 826 16450 2199
rect 16478 1722 16506 1741
rect 16478 1689 16506 1694
rect 16590 1385 16618 2702
rect 16646 2506 16674 4606
rect 16646 2473 16674 2478
rect 16590 1359 16591 1385
rect 16617 1359 16618 1385
rect 16590 1353 16618 1359
rect 16646 1722 16674 1727
rect 16422 793 16450 798
rect 16478 881 16506 887
rect 16478 855 16479 881
rect 16505 855 16506 881
rect 16478 434 16506 855
rect 16646 826 16674 1694
rect 16702 1498 16730 5054
rect 16814 4186 16842 5558
rect 17374 5362 17402 6455
rect 18270 6425 18298 7014
rect 19278 6594 19306 7056
rect 20510 7042 20538 7056
rect 20510 7009 20538 7014
rect 20678 7042 20706 7047
rect 19278 6561 19306 6566
rect 19838 6594 19866 6599
rect 19838 6547 19866 6566
rect 18774 6482 18802 6487
rect 18774 6481 19026 6482
rect 18774 6455 18775 6481
rect 18801 6455 19026 6481
rect 18774 6454 19026 6455
rect 18774 6449 18802 6454
rect 18270 6399 18271 6425
rect 18297 6399 18298 6425
rect 18270 6393 18298 6399
rect 17374 5329 17402 5334
rect 17430 6314 17458 6319
rect 16814 4153 16842 4158
rect 16870 3682 16898 3687
rect 16870 3457 16898 3654
rect 16870 3431 16871 3457
rect 16897 3431 16898 3457
rect 16870 3425 16898 3431
rect 17150 3289 17178 3295
rect 17150 3263 17151 3289
rect 17177 3263 17178 3289
rect 16758 2898 16786 2903
rect 16758 2841 16786 2870
rect 16758 2815 16759 2841
rect 16785 2815 16786 2841
rect 16758 2809 16786 2815
rect 17094 2450 17122 2455
rect 16926 2449 17122 2450
rect 16926 2423 17095 2449
rect 17121 2423 17122 2449
rect 16926 2422 17122 2423
rect 16870 2113 16898 2119
rect 16870 2087 16871 2113
rect 16897 2087 16898 2113
rect 16702 1470 16786 1498
rect 16590 798 16674 826
rect 16702 1330 16730 1335
rect 16534 602 16562 607
rect 16534 555 16562 574
rect 16478 401 16506 406
rect 16534 490 16562 495
rect 16534 322 16562 462
rect 16478 294 16562 322
rect 16478 56 16506 294
rect 16590 56 16618 798
rect 16702 56 16730 1302
rect 16758 154 16786 1470
rect 16870 1442 16898 2087
rect 16870 1409 16898 1414
rect 16870 1273 16898 1279
rect 16870 1247 16871 1273
rect 16897 1247 16898 1273
rect 16870 714 16898 1247
rect 16870 681 16898 686
rect 16814 546 16842 551
rect 16814 489 16842 518
rect 16814 463 16815 489
rect 16841 463 16842 489
rect 16814 457 16842 463
rect 16926 378 16954 2422
rect 17094 2417 17122 2422
rect 16982 2170 17010 2175
rect 16982 1049 17010 2142
rect 17150 2169 17178 3263
rect 17374 3010 17402 3015
rect 17150 2143 17151 2169
rect 17177 2143 17178 2169
rect 17150 2137 17178 2143
rect 17206 3009 17402 3010
rect 17206 2983 17375 3009
rect 17401 2983 17402 3009
rect 17206 2982 17402 2983
rect 17094 1666 17122 1671
rect 17094 1619 17122 1638
rect 17206 1442 17234 2982
rect 17374 2977 17402 2982
rect 17374 2562 17402 2567
rect 17318 2058 17346 2063
rect 17318 2011 17346 2030
rect 16982 1023 16983 1049
rect 17009 1023 17010 1049
rect 16982 1017 17010 1023
rect 17038 1414 17234 1442
rect 17262 1778 17290 1783
rect 16758 121 16786 126
rect 16814 350 16954 378
rect 16814 56 16842 350
rect 16926 154 16954 159
rect 16926 56 16954 126
rect 17038 56 17066 1414
rect 17262 994 17290 1750
rect 17150 966 17290 994
rect 17150 56 17178 966
rect 17262 881 17290 887
rect 17262 855 17263 881
rect 17289 855 17290 881
rect 17262 322 17290 855
rect 17262 289 17290 294
rect 17374 210 17402 2534
rect 17430 1385 17458 6286
rect 18494 6202 18522 6207
rect 17654 5922 17682 5927
rect 17654 5642 17682 5894
rect 17654 5609 17682 5614
rect 17654 5361 17682 5367
rect 17654 5335 17655 5361
rect 17681 5335 17682 5361
rect 17654 5306 17682 5335
rect 17654 5273 17682 5278
rect 18494 5306 18522 6174
rect 18830 6146 18858 6151
rect 18830 6099 18858 6118
rect 18494 5273 18522 5278
rect 18662 6034 18690 6039
rect 17878 5193 17906 5199
rect 17878 5167 17879 5193
rect 17905 5167 17906 5193
rect 17822 3850 17850 3855
rect 17654 3345 17682 3351
rect 17654 3319 17655 3345
rect 17681 3319 17682 3345
rect 17654 3178 17682 3319
rect 17654 3145 17682 3150
rect 17766 3346 17794 3351
rect 17598 2898 17626 2903
rect 17598 2617 17626 2870
rect 17598 2591 17599 2617
rect 17625 2591 17626 2617
rect 17598 2585 17626 2591
rect 17654 2618 17682 2623
rect 17598 1834 17626 1839
rect 17598 1787 17626 1806
rect 17598 1442 17626 1447
rect 17598 1395 17626 1414
rect 17430 1359 17431 1385
rect 17457 1359 17458 1385
rect 17430 1353 17458 1359
rect 17262 182 17402 210
rect 17430 1106 17458 1111
rect 17262 56 17290 182
rect 17430 154 17458 1078
rect 17374 126 17458 154
rect 17486 826 17514 831
rect 17374 56 17402 126
rect 17486 56 17514 798
rect 17654 601 17682 2590
rect 17654 575 17655 601
rect 17681 575 17682 601
rect 17654 569 17682 575
rect 17710 770 17738 775
rect 17598 546 17626 551
rect 17598 56 17626 518
rect 17710 56 17738 742
rect 17766 602 17794 3318
rect 17766 569 17794 574
rect 17822 56 17850 3822
rect 17878 3458 17906 5167
rect 17878 3425 17906 3430
rect 18102 5138 18130 5143
rect 18046 3402 18074 3407
rect 17878 3290 17906 3295
rect 17878 3289 17962 3290
rect 17878 3263 17879 3289
rect 17905 3263 17962 3289
rect 17878 3262 17962 3263
rect 17878 3257 17906 3262
rect 17878 2897 17906 2903
rect 17878 2871 17879 2897
rect 17905 2871 17906 2897
rect 17878 2730 17906 2871
rect 17878 2697 17906 2702
rect 17934 1834 17962 3262
rect 17990 2562 18018 2567
rect 17990 2515 18018 2534
rect 17934 1801 17962 1806
rect 17878 1722 17906 1741
rect 17878 1689 17906 1694
rect 17878 882 17906 887
rect 17878 835 17906 854
rect 17934 489 17962 495
rect 17934 463 17935 489
rect 17961 463 17962 489
rect 17934 266 17962 463
rect 17934 233 17962 238
rect 17934 98 17962 103
rect 17934 56 17962 70
rect 18046 56 18074 3374
rect 18102 378 18130 5110
rect 18326 4298 18354 4303
rect 18158 2841 18186 2847
rect 18158 2815 18159 2841
rect 18185 2815 18186 2841
rect 18158 2674 18186 2815
rect 18158 2641 18186 2646
rect 18270 2225 18298 2231
rect 18270 2199 18271 2225
rect 18297 2199 18298 2225
rect 18102 345 18130 350
rect 18158 1386 18186 1391
rect 18158 56 18186 1358
rect 18270 826 18298 2199
rect 18326 882 18354 4270
rect 18662 3850 18690 6006
rect 18998 5754 19026 6454
rect 19558 6481 19586 6487
rect 19558 6455 19559 6481
rect 19585 6455 19586 6481
rect 19558 6146 19586 6455
rect 20678 6425 20706 7014
rect 21742 6986 21770 7056
rect 21826 6986 21882 7098
rect 22960 7056 23016 7112
rect 24192 7056 24248 7112
rect 25424 7056 25480 7112
rect 21742 6958 21882 6986
rect 21854 6594 21882 6958
rect 22232 6678 22364 6683
rect 22260 6650 22284 6678
rect 22312 6650 22336 6678
rect 22232 6645 22364 6650
rect 21854 6561 21882 6566
rect 22134 6594 22162 6599
rect 22134 6547 22162 6566
rect 22974 6594 23002 7056
rect 23478 6986 23506 6991
rect 22974 6561 23002 6566
rect 23030 6930 23058 6935
rect 21126 6538 21154 6543
rect 21070 6482 21098 6487
rect 20678 6399 20679 6425
rect 20705 6399 20706 6425
rect 20678 6393 20706 6399
rect 20846 6481 21098 6482
rect 20846 6455 21071 6481
rect 21097 6455 21098 6481
rect 20846 6454 21098 6455
rect 19558 6113 19586 6118
rect 20846 6145 20874 6454
rect 21070 6449 21098 6454
rect 20846 6119 20847 6145
rect 20873 6119 20874 6145
rect 20846 6113 20874 6119
rect 19334 6090 19362 6095
rect 19054 5977 19082 5983
rect 19054 5951 19055 5977
rect 19081 5951 19082 5977
rect 19054 5866 19082 5951
rect 19054 5833 19082 5838
rect 19054 5754 19082 5759
rect 18998 5753 19082 5754
rect 18998 5727 19055 5753
rect 19081 5727 19082 5753
rect 18998 5726 19082 5727
rect 19054 5721 19082 5726
rect 19278 5697 19306 5703
rect 19278 5671 19279 5697
rect 19305 5671 19306 5697
rect 18718 5362 18746 5367
rect 18718 5315 18746 5334
rect 18942 5194 18970 5199
rect 18886 4186 18914 4191
rect 18662 3822 18746 3850
rect 18550 3458 18578 3463
rect 18382 3290 18410 3295
rect 18382 2617 18410 3262
rect 18382 2591 18383 2617
rect 18409 2591 18410 2617
rect 18382 2585 18410 2591
rect 18438 2897 18466 2903
rect 18438 2871 18439 2897
rect 18465 2871 18466 2897
rect 18382 1834 18410 1839
rect 18438 1834 18466 2871
rect 18382 1833 18466 1834
rect 18382 1807 18383 1833
rect 18409 1807 18466 1833
rect 18382 1806 18466 1807
rect 18494 2114 18522 2119
rect 18382 1801 18410 1806
rect 18382 1330 18410 1335
rect 18382 1283 18410 1302
rect 18494 1050 18522 2086
rect 18550 1218 18578 3430
rect 18606 2954 18634 2959
rect 18606 2907 18634 2926
rect 18662 2450 18690 2455
rect 18550 1185 18578 1190
rect 18606 2449 18690 2450
rect 18606 2423 18663 2449
rect 18689 2423 18690 2449
rect 18606 2422 18690 2423
rect 18494 1022 18578 1050
rect 18382 994 18410 999
rect 18382 947 18410 966
rect 18550 993 18578 1022
rect 18550 967 18551 993
rect 18577 967 18578 993
rect 18550 961 18578 967
rect 18494 938 18522 943
rect 18326 854 18410 882
rect 18270 793 18298 798
rect 18270 658 18298 663
rect 18270 56 18298 630
rect 18382 56 18410 854
rect 18494 601 18522 910
rect 18606 770 18634 2422
rect 18662 2417 18690 2422
rect 18662 1778 18690 1783
rect 18662 1721 18690 1750
rect 18662 1695 18663 1721
rect 18689 1695 18690 1721
rect 18662 1689 18690 1695
rect 18606 737 18634 742
rect 18718 658 18746 3822
rect 18830 3009 18858 3015
rect 18830 2983 18831 3009
rect 18857 2983 18858 3009
rect 18774 2170 18802 2175
rect 18774 2123 18802 2142
rect 18774 1386 18802 1391
rect 18830 1386 18858 2983
rect 18774 1385 18858 1386
rect 18774 1359 18775 1385
rect 18801 1359 18858 1385
rect 18774 1358 18858 1359
rect 18774 1353 18802 1358
rect 18494 575 18495 601
rect 18521 575 18522 601
rect 18494 569 18522 575
rect 18550 630 18746 658
rect 18774 1218 18802 1223
rect 18550 490 18578 630
rect 18774 546 18802 1190
rect 18494 462 18578 490
rect 18606 518 18802 546
rect 18830 881 18858 887
rect 18830 855 18831 881
rect 18857 855 18858 881
rect 18494 56 18522 462
rect 18606 56 18634 518
rect 18830 490 18858 855
rect 18830 457 18858 462
rect 18718 378 18746 383
rect 18886 378 18914 4158
rect 18942 1694 18970 5166
rect 18998 5194 19026 5199
rect 18998 5193 19138 5194
rect 18998 5167 18999 5193
rect 19025 5167 19138 5193
rect 18998 5166 19138 5167
rect 18998 5161 19026 5166
rect 18998 4354 19026 4359
rect 18998 2674 19026 4326
rect 19054 2841 19082 2847
rect 19054 2815 19055 2841
rect 19081 2815 19082 2841
rect 19054 2786 19082 2815
rect 19054 2753 19082 2758
rect 18998 2646 19082 2674
rect 18998 2338 19026 2343
rect 18998 2225 19026 2310
rect 18998 2199 18999 2225
rect 19025 2199 19026 2225
rect 18998 2193 19026 2199
rect 18942 1666 19026 1694
rect 18942 714 18970 733
rect 18942 681 18970 686
rect 18998 602 19026 1666
rect 18718 56 18746 350
rect 18830 350 18914 378
rect 18942 574 19026 602
rect 18830 56 18858 350
rect 18942 56 18970 574
rect 19054 56 19082 2646
rect 19110 1694 19138 5166
rect 19166 2674 19194 2679
rect 19166 2617 19194 2646
rect 19166 2591 19167 2617
rect 19193 2591 19194 2617
rect 19166 2585 19194 2591
rect 19278 2562 19306 5671
rect 19334 5082 19362 6062
rect 20566 5977 20594 5983
rect 20566 5951 20567 5977
rect 20593 5951 20594 5977
rect 20230 5922 20258 5927
rect 19334 5049 19362 5054
rect 19502 5866 19530 5871
rect 19334 2898 19362 2903
rect 19334 2851 19362 2870
rect 19278 2534 19418 2562
rect 19222 2058 19250 2063
rect 19222 2011 19250 2030
rect 19334 2002 19362 2007
rect 19166 1834 19194 1839
rect 19166 1787 19194 1806
rect 19110 1666 19306 1694
rect 19278 1386 19306 1666
rect 19222 1358 19306 1386
rect 19166 1329 19194 1335
rect 19166 1303 19167 1329
rect 19193 1303 19194 1329
rect 19166 1106 19194 1303
rect 19222 1162 19250 1358
rect 19222 1134 19306 1162
rect 19166 1073 19194 1078
rect 19166 714 19194 719
rect 19110 658 19138 663
rect 19110 210 19138 630
rect 19110 177 19138 182
rect 19166 56 19194 686
rect 19278 56 19306 1134
rect 19334 1105 19362 1974
rect 19334 1079 19335 1105
rect 19361 1079 19362 1105
rect 19334 1073 19362 1079
rect 19390 56 19418 2534
rect 19446 1722 19474 1727
rect 19446 770 19474 1694
rect 19446 737 19474 742
rect 19502 56 19530 5838
rect 20062 2954 20090 2959
rect 20062 2170 20090 2926
rect 20062 2137 20090 2142
rect 20174 2561 20202 2567
rect 20174 2535 20175 2561
rect 20201 2535 20202 2561
rect 19670 2058 19698 2063
rect 19558 1386 19586 1391
rect 19558 1339 19586 1358
rect 19670 1050 19698 2030
rect 20174 1498 20202 2535
rect 20174 1465 20202 1470
rect 20006 1329 20034 1335
rect 20006 1303 20007 1329
rect 20033 1303 20034 1329
rect 19726 1274 19754 1279
rect 19726 1227 19754 1246
rect 19670 1022 19754 1050
rect 19614 994 19642 999
rect 19614 947 19642 966
rect 19614 826 19642 831
rect 19614 56 19642 798
rect 19670 657 19698 663
rect 19670 631 19671 657
rect 19697 631 19698 657
rect 19670 154 19698 631
rect 19670 121 19698 126
rect 19726 56 19754 1022
rect 19838 770 19866 775
rect 19838 56 19866 742
rect 19950 658 19978 663
rect 19950 56 19978 630
rect 20006 602 20034 1303
rect 20230 714 20258 5894
rect 20286 3626 20314 3631
rect 20286 1498 20314 3598
rect 20510 3010 20538 3015
rect 20510 2953 20538 2982
rect 20510 2927 20511 2953
rect 20537 2927 20538 2953
rect 20510 2921 20538 2927
rect 20342 2898 20370 2903
rect 20342 1722 20370 2870
rect 20398 2730 20426 2735
rect 20398 2617 20426 2702
rect 20398 2591 20399 2617
rect 20425 2591 20426 2617
rect 20398 2585 20426 2591
rect 20342 1689 20370 1694
rect 20286 1465 20314 1470
rect 20342 1554 20370 1559
rect 20230 681 20258 686
rect 20342 714 20370 1526
rect 20566 826 20594 5951
rect 21014 5977 21042 5983
rect 21014 5951 21015 5977
rect 21041 5951 21042 5977
rect 20902 5474 20930 5479
rect 20622 4970 20650 4975
rect 20622 3066 20650 4942
rect 20622 3033 20650 3038
rect 20790 2897 20818 2903
rect 20790 2871 20791 2897
rect 20817 2871 20818 2897
rect 20790 1834 20818 2871
rect 20790 1801 20818 1806
rect 20902 1834 20930 5446
rect 20902 1801 20930 1806
rect 20566 793 20594 798
rect 21014 770 21042 5951
rect 21126 5754 21154 6510
rect 21462 6482 21490 6487
rect 21294 6146 21322 6151
rect 21294 6099 21322 6118
rect 21126 5721 21154 5726
rect 21406 5978 21434 5983
rect 21126 5642 21154 5647
rect 21070 3345 21098 3351
rect 21070 3319 21071 3345
rect 21097 3319 21098 3345
rect 21070 2506 21098 3319
rect 21070 2473 21098 2478
rect 21126 2114 21154 5614
rect 21294 4129 21322 4135
rect 21294 4103 21295 4129
rect 21321 4103 21322 4129
rect 21294 4018 21322 4103
rect 21294 3985 21322 3990
rect 21294 3290 21322 3295
rect 21294 3243 21322 3262
rect 21126 2081 21154 2086
rect 21014 737 21042 742
rect 20342 681 20370 686
rect 20062 602 20090 607
rect 20006 601 20090 602
rect 20006 575 20063 601
rect 20089 575 20090 601
rect 20006 574 20090 575
rect 20062 569 20090 574
rect 20566 546 20594 551
rect 20566 499 20594 518
rect 20958 546 20986 551
rect 20958 499 20986 518
rect 20062 490 20090 495
rect 20062 56 20090 462
rect 21406 490 21434 5950
rect 21462 2338 21490 6454
rect 21854 6482 21882 6487
rect 21854 6435 21882 6454
rect 22806 6481 22834 6487
rect 22806 6455 22807 6481
rect 22833 6455 22834 6481
rect 21902 6286 22034 6291
rect 21930 6258 21954 6286
rect 21982 6258 22006 6286
rect 21902 6253 22034 6258
rect 22358 6034 22386 6039
rect 22358 5987 22386 6006
rect 22078 5978 22106 5983
rect 22078 5931 22106 5950
rect 21686 5922 21714 5927
rect 21462 2305 21490 2310
rect 21518 4073 21546 4079
rect 21518 4047 21519 4073
rect 21545 4047 21546 4073
rect 21518 1386 21546 4047
rect 21686 3402 21714 5894
rect 22232 5894 22364 5899
rect 22260 5866 22284 5894
rect 22312 5866 22336 5894
rect 22232 5861 22364 5866
rect 22694 5810 22722 5815
rect 22694 5763 22722 5782
rect 21902 5502 22034 5507
rect 21930 5474 21954 5502
rect 21982 5474 22006 5502
rect 21902 5469 22034 5474
rect 22232 5110 22364 5115
rect 22260 5082 22284 5110
rect 22312 5082 22336 5110
rect 22232 5077 22364 5082
rect 21902 4718 22034 4723
rect 21930 4690 21954 4718
rect 21982 4690 22006 4718
rect 21902 4685 22034 4690
rect 22750 4578 22778 4583
rect 22750 4531 22778 4550
rect 22470 4522 22498 4527
rect 22470 4475 22498 4494
rect 22232 4326 22364 4331
rect 22260 4298 22284 4326
rect 22312 4298 22336 4326
rect 22232 4293 22364 4298
rect 21902 3934 22034 3939
rect 21930 3906 21954 3934
rect 21982 3906 22006 3934
rect 21902 3901 22034 3906
rect 22232 3542 22364 3547
rect 22260 3514 22284 3542
rect 22312 3514 22336 3542
rect 22232 3509 22364 3514
rect 21686 3369 21714 3374
rect 22134 3346 22162 3351
rect 22134 3299 22162 3318
rect 22358 3289 22386 3295
rect 22358 3263 22359 3289
rect 22385 3263 22386 3289
rect 21902 3150 22034 3155
rect 21930 3122 21954 3150
rect 21982 3122 22006 3150
rect 21902 3117 22034 3122
rect 22358 2954 22386 3263
rect 22358 2921 22386 2926
rect 22232 2758 22364 2763
rect 22260 2730 22284 2758
rect 22312 2730 22336 2758
rect 22232 2725 22364 2730
rect 21902 2366 22034 2371
rect 21930 2338 21954 2366
rect 21982 2338 22006 2366
rect 21902 2333 22034 2338
rect 22470 2113 22498 2119
rect 22470 2087 22471 2113
rect 22497 2087 22498 2113
rect 22190 2058 22218 2077
rect 22190 2025 22218 2030
rect 22232 1974 22364 1979
rect 22260 1946 22284 1974
rect 22312 1946 22336 1974
rect 22232 1941 22364 1946
rect 22470 1778 22498 2087
rect 22470 1745 22498 1750
rect 21902 1582 22034 1587
rect 21930 1554 21954 1582
rect 21982 1554 22006 1582
rect 21902 1549 22034 1554
rect 21518 1353 21546 1358
rect 22750 1274 22778 1279
rect 22232 1190 22364 1195
rect 22260 1162 22284 1190
rect 22312 1162 22336 1190
rect 22232 1157 22364 1162
rect 22470 1050 22498 1055
rect 22470 1003 22498 1022
rect 22750 1049 22778 1246
rect 22750 1023 22751 1049
rect 22777 1023 22778 1049
rect 22750 1017 22778 1023
rect 21902 798 22034 803
rect 21930 770 21954 798
rect 21982 770 22006 798
rect 21902 765 22034 770
rect 22806 658 22834 6455
rect 23030 6145 23058 6902
rect 23086 6482 23114 6487
rect 23086 6435 23114 6454
rect 23366 6481 23394 6487
rect 23366 6455 23367 6481
rect 23393 6455 23394 6481
rect 23030 6119 23031 6145
rect 23057 6119 23058 6145
rect 23030 6113 23058 6119
rect 23366 6146 23394 6455
rect 23366 6113 23394 6118
rect 23310 6090 23338 6095
rect 23310 6043 23338 6062
rect 23478 5866 23506 6958
rect 23646 6594 23674 6599
rect 23646 6547 23674 6566
rect 24206 6594 24234 7056
rect 25214 6762 25242 6767
rect 24206 6561 24234 6566
rect 24598 6594 24626 6599
rect 24598 6547 24626 6566
rect 24374 6482 24402 6487
rect 24374 6435 24402 6454
rect 24038 6202 24066 6207
rect 24038 6155 24066 6174
rect 24822 6145 24850 6151
rect 24822 6119 24823 6145
rect 24849 6119 24850 6145
rect 24374 6089 24402 6095
rect 24374 6063 24375 6089
rect 24401 6063 24402 6089
rect 23534 6034 23562 6039
rect 23534 5987 23562 6006
rect 23478 5833 23506 5838
rect 23142 5754 23170 5759
rect 23142 5707 23170 5726
rect 23534 5754 23562 5759
rect 23534 5707 23562 5726
rect 22974 5641 23002 5647
rect 22974 5615 22975 5641
rect 23001 5615 23002 5641
rect 22974 5082 23002 5615
rect 24038 5474 24066 5479
rect 24038 5417 24066 5446
rect 24038 5391 24039 5417
rect 24065 5391 24066 5417
rect 24038 5385 24066 5391
rect 24374 5418 24402 6063
rect 24822 5922 24850 6119
rect 25102 6034 25130 6039
rect 24822 5889 24850 5894
rect 25046 6033 25130 6034
rect 25046 6007 25103 6033
rect 25129 6007 25130 6033
rect 25046 6006 25130 6007
rect 24486 5697 24514 5703
rect 24486 5671 24487 5697
rect 24513 5671 24514 5697
rect 24486 5418 24514 5671
rect 24934 5642 24962 5647
rect 24934 5595 24962 5614
rect 24374 5390 24458 5418
rect 23086 5306 23114 5311
rect 23086 5259 23114 5278
rect 24374 5305 24402 5311
rect 24374 5279 24375 5305
rect 24401 5279 24402 5305
rect 23366 5250 23394 5255
rect 23534 5250 23562 5255
rect 23366 5249 23562 5250
rect 23366 5223 23367 5249
rect 23393 5223 23535 5249
rect 23561 5223 23562 5249
rect 23366 5222 23562 5223
rect 23366 5217 23394 5222
rect 23534 5217 23562 5222
rect 24374 5250 24402 5279
rect 24374 5217 24402 5222
rect 22974 5049 23002 5054
rect 24374 5082 24402 5087
rect 23142 5026 23170 5031
rect 23142 2953 23170 4998
rect 24150 5026 24178 5031
rect 23534 4913 23562 4919
rect 23534 4887 23535 4913
rect 23561 4887 23562 4913
rect 23534 4802 23562 4887
rect 23758 4914 23786 4919
rect 23758 4867 23786 4886
rect 23534 4769 23562 4774
rect 24150 4577 24178 4998
rect 24150 4551 24151 4577
rect 24177 4551 24178 4577
rect 24150 4545 24178 4551
rect 24206 4522 24234 4527
rect 23870 4466 23898 4471
rect 23870 4419 23898 4438
rect 23254 4186 23282 4191
rect 23254 4139 23282 4158
rect 23478 4074 23506 4079
rect 23478 4027 23506 4046
rect 24150 3794 24178 3799
rect 24150 3747 24178 3766
rect 23870 3682 23898 3687
rect 23870 3635 23898 3654
rect 23142 2927 23143 2953
rect 23169 2927 23170 2953
rect 23142 2921 23170 2927
rect 24206 2953 24234 4494
rect 24374 4521 24402 5054
rect 24430 5026 24458 5390
rect 24486 5385 24514 5390
rect 24822 5361 24850 5367
rect 24822 5335 24823 5361
rect 24849 5335 24850 5361
rect 24822 5194 24850 5335
rect 24822 5161 24850 5166
rect 24430 4993 24458 4998
rect 24430 4914 24458 4919
rect 24430 4867 24458 4886
rect 24934 4858 24962 4863
rect 24934 4811 24962 4830
rect 24822 4634 24850 4639
rect 24822 4587 24850 4606
rect 24374 4495 24375 4521
rect 24401 4495 24402 4521
rect 24374 4489 24402 4495
rect 25046 4185 25074 6006
rect 25102 6001 25130 6006
rect 25214 5754 25242 6734
rect 25382 6538 25410 6543
rect 25270 6481 25298 6487
rect 25270 6455 25271 6481
rect 25297 6455 25298 6481
rect 25270 5866 25298 6455
rect 25270 5833 25298 5838
rect 25326 6314 25354 6319
rect 25214 5721 25242 5726
rect 25270 5697 25298 5703
rect 25270 5671 25271 5697
rect 25297 5671 25298 5697
rect 25102 5249 25130 5255
rect 25102 5223 25103 5249
rect 25129 5223 25130 5249
rect 25102 4410 25130 5223
rect 25214 4913 25242 4919
rect 25214 4887 25215 4913
rect 25241 4887 25242 4913
rect 25214 4578 25242 4887
rect 25214 4545 25242 4550
rect 25102 4377 25130 4382
rect 25158 4521 25186 4527
rect 25158 4495 25159 4521
rect 25185 4495 25186 4521
rect 25046 4159 25047 4185
rect 25073 4159 25074 4185
rect 25046 4153 25074 4159
rect 25102 4242 25130 4247
rect 24374 4130 24402 4135
rect 24598 4130 24626 4135
rect 24374 4129 24458 4130
rect 24374 4103 24375 4129
rect 24401 4103 24458 4129
rect 24374 4102 24458 4103
rect 24374 4097 24402 4102
rect 24374 3738 24402 3743
rect 24374 3691 24402 3710
rect 24430 3626 24458 4102
rect 24598 4083 24626 4102
rect 24766 4129 24794 4135
rect 24766 4103 24767 4129
rect 24793 4103 24794 4129
rect 24766 4018 24794 4103
rect 24766 3985 24794 3990
rect 24430 3593 24458 3598
rect 24822 3793 24850 3799
rect 24822 3767 24823 3793
rect 24849 3767 24850 3793
rect 24822 3402 24850 3767
rect 25102 3737 25130 4214
rect 25158 4074 25186 4495
rect 25214 4130 25242 4135
rect 25214 4083 25242 4102
rect 25158 4041 25186 4046
rect 25270 3794 25298 5671
rect 25326 4634 25354 6286
rect 25382 5474 25410 6510
rect 25438 6202 25466 7056
rect 25438 6169 25466 6174
rect 25494 6425 25522 6431
rect 25494 6399 25495 6425
rect 25521 6399 25522 6425
rect 25494 6090 25522 6399
rect 25494 6057 25522 6062
rect 25606 6145 25634 6151
rect 25606 6119 25607 6145
rect 25633 6119 25634 6145
rect 25382 5441 25410 5446
rect 25606 5418 25634 6119
rect 25606 5385 25634 5390
rect 25662 6090 25690 6095
rect 25494 5249 25522 5255
rect 25494 5223 25495 5249
rect 25521 5223 25522 5249
rect 25494 4746 25522 5223
rect 25662 4858 25690 6062
rect 25718 5585 25746 5591
rect 25718 5559 25719 5585
rect 25745 5559 25746 5585
rect 25718 4970 25746 5559
rect 25718 4937 25746 4942
rect 25662 4825 25690 4830
rect 25494 4713 25522 4718
rect 25718 4801 25746 4807
rect 25718 4775 25719 4801
rect 25745 4775 25746 4801
rect 25326 4601 25354 4606
rect 25718 4522 25746 4775
rect 25718 4489 25746 4494
rect 25494 4465 25522 4471
rect 25494 4439 25495 4465
rect 25521 4439 25522 4465
rect 25494 4298 25522 4439
rect 25494 4265 25522 4270
rect 25606 4074 25634 4079
rect 25606 3849 25634 4046
rect 25606 3823 25607 3849
rect 25633 3823 25634 3849
rect 25606 3817 25634 3823
rect 25718 4017 25746 4023
rect 25718 3991 25719 4017
rect 25745 3991 25746 4017
rect 25718 3850 25746 3991
rect 25718 3817 25746 3822
rect 25270 3761 25298 3766
rect 25102 3711 25103 3737
rect 25129 3711 25130 3737
rect 25102 3705 25130 3711
rect 24822 3369 24850 3374
rect 25718 3626 25746 3631
rect 24430 3346 24458 3351
rect 24430 3299 24458 3318
rect 25214 3345 25242 3351
rect 25214 3319 25215 3345
rect 25241 3319 25242 3345
rect 24206 2927 24207 2953
rect 24233 2927 24234 2953
rect 24206 2921 24234 2927
rect 24878 3289 24906 3295
rect 24878 3263 24879 3289
rect 24905 3263 24906 3289
rect 24878 2954 24906 3263
rect 25214 3066 25242 3319
rect 25718 3289 25746 3598
rect 25718 3263 25719 3289
rect 25745 3263 25746 3289
rect 25718 3257 25746 3263
rect 25214 3033 25242 3038
rect 25606 3178 25634 3183
rect 25606 3065 25634 3150
rect 25606 3039 25607 3065
rect 25633 3039 25634 3065
rect 25606 3033 25634 3039
rect 24878 2921 24906 2926
rect 23422 2897 23450 2903
rect 23422 2871 23423 2897
rect 23449 2871 23450 2897
rect 23422 2562 23450 2871
rect 23590 2898 23618 2903
rect 23590 2851 23618 2870
rect 23870 2897 23898 2903
rect 23870 2871 23871 2897
rect 23897 2871 23898 2897
rect 23422 2529 23450 2534
rect 23814 2114 23842 2119
rect 23814 2067 23842 2086
rect 23534 1834 23562 1839
rect 23534 1777 23562 1806
rect 23534 1751 23535 1777
rect 23561 1751 23562 1777
rect 23534 1745 23562 1751
rect 23702 1721 23730 1727
rect 23702 1695 23703 1721
rect 23729 1695 23730 1721
rect 23534 1498 23562 1503
rect 23086 1442 23114 1447
rect 23086 1385 23114 1414
rect 23086 1359 23087 1385
rect 23113 1359 23114 1385
rect 23086 1353 23114 1359
rect 23534 1385 23562 1470
rect 23534 1359 23535 1385
rect 23561 1359 23562 1385
rect 23534 1353 23562 1359
rect 23366 1330 23394 1335
rect 23366 1283 23394 1302
rect 23534 1106 23562 1111
rect 23534 993 23562 1078
rect 23534 967 23535 993
rect 23561 967 23562 993
rect 23534 961 23562 967
rect 22806 625 22834 630
rect 23702 601 23730 1695
rect 23758 994 23786 999
rect 23758 947 23786 966
rect 23702 575 23703 601
rect 23729 575 23730 601
rect 23702 569 23730 575
rect 23870 546 23898 2871
rect 24486 2897 24514 2903
rect 24486 2871 24487 2897
rect 24513 2871 24514 2897
rect 24486 2618 24514 2871
rect 24934 2897 24962 2903
rect 24934 2871 24935 2897
rect 24961 2871 24962 2897
rect 24486 2585 24514 2590
rect 24654 2841 24682 2847
rect 24654 2815 24655 2841
rect 24681 2815 24682 2841
rect 24374 2562 24402 2567
rect 24094 2226 24122 2231
rect 24094 2179 24122 2198
rect 24374 2169 24402 2534
rect 24430 2561 24458 2567
rect 24430 2535 24431 2561
rect 24457 2535 24458 2561
rect 24430 2226 24458 2535
rect 24654 2450 24682 2815
rect 24934 2674 24962 2871
rect 25102 2897 25130 2903
rect 25102 2871 25103 2897
rect 25129 2871 25130 2897
rect 25102 2842 25130 2871
rect 25102 2809 25130 2814
rect 24934 2641 24962 2646
rect 25606 2730 25634 2735
rect 25214 2618 25242 2623
rect 25214 2571 25242 2590
rect 25606 2617 25634 2702
rect 25606 2591 25607 2617
rect 25633 2591 25634 2617
rect 25606 2585 25634 2591
rect 24822 2562 24850 2567
rect 24822 2515 24850 2534
rect 25550 2562 25578 2567
rect 24654 2417 24682 2422
rect 25438 2506 25466 2511
rect 25438 2281 25466 2478
rect 25438 2255 25439 2281
rect 25465 2255 25466 2281
rect 25438 2249 25466 2255
rect 25550 2282 25578 2534
rect 25550 2249 25578 2254
rect 24430 2193 24458 2198
rect 24374 2143 24375 2169
rect 24401 2143 24402 2169
rect 24374 2137 24402 2143
rect 25606 2169 25634 2175
rect 25606 2143 25607 2169
rect 25633 2143 25634 2169
rect 24710 2113 24738 2119
rect 24710 2087 24711 2113
rect 24737 2087 24738 2113
rect 24710 1834 24738 2087
rect 24710 1801 24738 1806
rect 25214 1890 25242 1895
rect 25214 1833 25242 1862
rect 25214 1807 25215 1833
rect 25241 1807 25242 1833
rect 25214 1801 25242 1807
rect 24430 1777 24458 1783
rect 24430 1751 24431 1777
rect 24457 1751 24458 1777
rect 24038 1442 24066 1447
rect 24038 1395 24066 1414
rect 24318 1329 24346 1335
rect 24318 1303 24319 1329
rect 24345 1303 24346 1329
rect 24318 714 24346 1303
rect 24318 681 24346 686
rect 24374 1330 24402 1335
rect 23870 513 23898 518
rect 24094 657 24122 663
rect 24094 631 24095 657
rect 24121 631 24122 657
rect 21406 457 21434 462
rect 24094 490 24122 631
rect 24374 601 24402 1302
rect 24430 1274 24458 1751
rect 25102 1778 25130 1783
rect 24934 1722 24962 1727
rect 24934 1675 24962 1694
rect 24430 1241 24458 1246
rect 24486 1666 24514 1671
rect 24486 993 24514 1638
rect 25102 1385 25130 1750
rect 25494 1722 25522 1727
rect 25102 1359 25103 1385
rect 25129 1359 25130 1385
rect 25102 1353 25130 1359
rect 25326 1442 25354 1447
rect 24710 1330 24738 1335
rect 24710 1283 24738 1302
rect 24486 967 24487 993
rect 24513 967 24514 993
rect 24486 961 24514 967
rect 25214 994 25242 999
rect 25214 947 25242 966
rect 24934 938 24962 943
rect 24934 891 24962 910
rect 24878 714 24906 719
rect 24878 667 24906 686
rect 24374 575 24375 601
rect 24401 575 24402 601
rect 24374 569 24402 575
rect 25270 602 25298 607
rect 25270 555 25298 574
rect 24094 457 24122 462
rect 22232 406 22364 411
rect 22260 378 22284 406
rect 22312 378 22336 406
rect 22232 373 22364 378
rect 25326 266 25354 1414
rect 25494 1386 25522 1694
rect 25550 1610 25578 1615
rect 25550 1441 25578 1582
rect 25550 1415 25551 1441
rect 25577 1415 25578 1441
rect 25550 1409 25578 1415
rect 25494 1353 25522 1358
rect 25326 233 25354 238
rect 25438 1330 25466 1335
rect 4942 9 4970 14
rect 6160 0 6216 56
rect 6272 0 6328 56
rect 6384 0 6440 56
rect 6496 0 6552 56
rect 6608 0 6664 56
rect 6720 0 6776 56
rect 6832 0 6888 56
rect 6944 0 7000 56
rect 7056 0 7112 56
rect 7168 0 7224 56
rect 7280 0 7336 56
rect 7392 0 7448 56
rect 7504 0 7560 56
rect 7616 0 7672 56
rect 7728 0 7784 56
rect 7840 0 7896 56
rect 7952 0 8008 56
rect 8064 0 8120 56
rect 8176 0 8232 56
rect 8288 0 8344 56
rect 8400 0 8456 56
rect 8512 0 8568 56
rect 8624 0 8680 56
rect 8736 0 8792 56
rect 8848 0 8904 56
rect 8960 0 9016 56
rect 9072 0 9128 56
rect 9184 0 9240 56
rect 9296 0 9352 56
rect 9408 0 9464 56
rect 9520 0 9576 56
rect 9632 0 9688 56
rect 9744 0 9800 56
rect 9856 0 9912 56
rect 9968 0 10024 56
rect 10080 0 10136 56
rect 10192 0 10248 56
rect 10304 0 10360 56
rect 10416 0 10472 56
rect 10528 0 10584 56
rect 10640 0 10696 56
rect 10752 0 10808 56
rect 10864 0 10920 56
rect 10976 0 11032 56
rect 11088 0 11144 56
rect 11200 0 11256 56
rect 11312 0 11368 56
rect 11424 0 11480 56
rect 11536 0 11592 56
rect 11648 0 11704 56
rect 11760 0 11816 56
rect 11872 0 11928 56
rect 11984 0 12040 56
rect 12096 0 12152 56
rect 12208 0 12264 56
rect 12320 0 12376 56
rect 12432 0 12488 56
rect 12544 0 12600 56
rect 12656 0 12712 56
rect 12768 0 12824 56
rect 12880 0 12936 56
rect 12992 0 13048 56
rect 13104 0 13160 56
rect 13216 0 13272 56
rect 13328 0 13384 56
rect 13440 0 13496 56
rect 13552 0 13608 56
rect 13664 0 13720 56
rect 13776 0 13832 56
rect 13888 0 13944 56
rect 14000 0 14056 56
rect 14112 0 14168 56
rect 14224 0 14280 56
rect 14336 0 14392 56
rect 14448 0 14504 56
rect 14560 0 14616 56
rect 14672 0 14728 56
rect 14784 0 14840 56
rect 14896 0 14952 56
rect 15008 0 15064 56
rect 15120 0 15176 56
rect 15232 0 15288 56
rect 15344 0 15400 56
rect 15456 0 15512 56
rect 15568 0 15624 56
rect 15680 0 15736 56
rect 15792 0 15848 56
rect 15904 0 15960 56
rect 16016 0 16072 56
rect 16128 0 16184 56
rect 16240 0 16296 56
rect 16352 0 16408 56
rect 16464 0 16520 56
rect 16576 0 16632 56
rect 16688 0 16744 56
rect 16800 0 16856 56
rect 16912 0 16968 56
rect 17024 0 17080 56
rect 17136 0 17192 56
rect 17248 0 17304 56
rect 17360 0 17416 56
rect 17472 0 17528 56
rect 17584 0 17640 56
rect 17696 0 17752 56
rect 17808 0 17864 56
rect 17920 0 17976 56
rect 18032 0 18088 56
rect 18144 0 18200 56
rect 18256 0 18312 56
rect 18368 0 18424 56
rect 18480 0 18536 56
rect 18592 0 18648 56
rect 18704 0 18760 56
rect 18816 0 18872 56
rect 18928 0 18984 56
rect 19040 0 19096 56
rect 19152 0 19208 56
rect 19264 0 19320 56
rect 19376 0 19432 56
rect 19488 0 19544 56
rect 19600 0 19656 56
rect 19712 0 19768 56
rect 19824 0 19880 56
rect 19936 0 19992 56
rect 20048 0 20104 56
rect 25438 42 25466 1302
rect 25550 658 25578 663
rect 25606 658 25634 2143
rect 25718 2058 25746 2063
rect 25718 1721 25746 2030
rect 25718 1695 25719 1721
rect 25745 1695 25746 1721
rect 25718 1689 25746 1695
rect 25718 1162 25746 1167
rect 25718 937 25746 1134
rect 25718 911 25719 937
rect 25745 911 25746 937
rect 25718 905 25746 911
rect 25550 657 25634 658
rect 25550 631 25551 657
rect 25577 631 25634 657
rect 25550 630 25634 631
rect 25550 625 25578 630
rect 25438 9 25466 14
<< via2 >>
rect 1134 6734 1162 6762
rect 1078 6481 1106 6482
rect 1078 6455 1079 6481
rect 1079 6455 1105 6481
rect 1105 6455 1106 6481
rect 1078 6454 1106 6455
rect 574 6286 602 6314
rect 350 6062 378 6090
rect 1638 6510 1666 6538
rect 1358 6398 1386 6426
rect 574 5782 602 5810
rect 3262 7014 3290 7042
rect 3486 7014 3514 7042
rect 3038 6734 3066 6762
rect 2232 6677 2260 6678
rect 2232 6651 2233 6677
rect 2233 6651 2259 6677
rect 2259 6651 2260 6677
rect 2232 6650 2260 6651
rect 2284 6677 2312 6678
rect 2284 6651 2285 6677
rect 2285 6651 2311 6677
rect 2311 6651 2312 6677
rect 2284 6650 2312 6651
rect 2336 6677 2364 6678
rect 2336 6651 2337 6677
rect 2337 6651 2363 6677
rect 2363 6651 2364 6677
rect 2336 6650 2364 6651
rect 2030 6510 2058 6538
rect 2646 6537 2674 6538
rect 2646 6511 2647 6537
rect 2647 6511 2673 6537
rect 2673 6511 2674 6537
rect 2646 6510 2674 6511
rect 2478 6454 2506 6482
rect 1902 6285 1930 6286
rect 1902 6259 1903 6285
rect 1903 6259 1929 6285
rect 1929 6259 1930 6285
rect 1902 6258 1930 6259
rect 1954 6285 1982 6286
rect 1954 6259 1955 6285
rect 1955 6259 1981 6285
rect 1981 6259 1982 6285
rect 1954 6258 1982 6259
rect 2006 6285 2034 6286
rect 2006 6259 2007 6285
rect 2007 6259 2033 6285
rect 2033 6259 2034 6285
rect 2006 6258 2034 6259
rect 2232 5893 2260 5894
rect 2232 5867 2233 5893
rect 2233 5867 2259 5893
rect 2259 5867 2260 5893
rect 2232 5866 2260 5867
rect 2284 5893 2312 5894
rect 2284 5867 2285 5893
rect 2285 5867 2311 5893
rect 2311 5867 2312 5893
rect 2284 5866 2312 5867
rect 2336 5893 2364 5894
rect 2336 5867 2337 5893
rect 2337 5867 2363 5893
rect 2363 5867 2364 5893
rect 2336 5866 2364 5867
rect 1902 5501 1930 5502
rect 1902 5475 1903 5501
rect 1903 5475 1929 5501
rect 1929 5475 1930 5501
rect 1902 5474 1930 5475
rect 1954 5501 1982 5502
rect 1954 5475 1955 5501
rect 1955 5475 1981 5501
rect 1981 5475 1982 5501
rect 1954 5474 1982 5475
rect 2006 5501 2034 5502
rect 2006 5475 2007 5501
rect 2007 5475 2033 5501
rect 2033 5475 2034 5501
rect 2006 5474 2034 5475
rect 2422 5390 2450 5418
rect 2232 5109 2260 5110
rect 2232 5083 2233 5109
rect 2233 5083 2259 5109
rect 2259 5083 2260 5109
rect 2232 5082 2260 5083
rect 2284 5109 2312 5110
rect 2284 5083 2285 5109
rect 2285 5083 2311 5109
rect 2311 5083 2312 5109
rect 2284 5082 2312 5083
rect 2336 5109 2364 5110
rect 2336 5083 2337 5109
rect 2337 5083 2363 5109
rect 2363 5083 2364 5109
rect 2336 5082 2364 5083
rect 1638 4998 1666 5026
rect 350 4830 378 4858
rect 1902 4717 1930 4718
rect 1902 4691 1903 4717
rect 1903 4691 1929 4717
rect 1929 4691 1930 4717
rect 1902 4690 1930 4691
rect 1954 4717 1982 4718
rect 1954 4691 1955 4717
rect 1955 4691 1981 4717
rect 1981 4691 1982 4717
rect 1954 4690 1982 4691
rect 2006 4717 2034 4718
rect 2006 4691 2007 4717
rect 2007 4691 2033 4717
rect 2033 4691 2034 4717
rect 2006 4690 2034 4691
rect 1078 3990 1106 4018
rect 854 3430 882 3458
rect 854 3009 882 3010
rect 854 2983 855 3009
rect 855 2983 881 3009
rect 881 2983 882 3009
rect 854 2982 882 2983
rect 1078 2841 1106 2842
rect 1078 2815 1079 2841
rect 1079 2815 1105 2841
rect 1105 2815 1106 2841
rect 1078 2814 1106 2815
rect 966 2113 994 2114
rect 966 2087 967 2113
rect 967 2087 993 2113
rect 993 2087 994 2113
rect 966 2086 994 2087
rect 910 1694 938 1722
rect 1902 3933 1930 3934
rect 1902 3907 1903 3933
rect 1903 3907 1929 3933
rect 1929 3907 1930 3933
rect 1902 3906 1930 3907
rect 1954 3933 1982 3934
rect 1954 3907 1955 3933
rect 1955 3907 1981 3933
rect 1981 3907 1982 3933
rect 1954 3906 1982 3907
rect 2006 3933 2034 3934
rect 2006 3907 2007 3933
rect 2007 3907 2033 3933
rect 2033 3907 2034 3933
rect 2006 3906 2034 3907
rect 2232 4325 2260 4326
rect 2232 4299 2233 4325
rect 2233 4299 2259 4325
rect 2259 4299 2260 4325
rect 2232 4298 2260 4299
rect 2284 4325 2312 4326
rect 2284 4299 2285 4325
rect 2285 4299 2311 4325
rect 2311 4299 2312 4325
rect 2284 4298 2312 4299
rect 2336 4325 2364 4326
rect 2336 4299 2337 4325
rect 2337 4299 2363 4325
rect 2363 4299 2364 4325
rect 2336 4298 2364 4299
rect 4494 7014 4522 7042
rect 4718 7014 4746 7042
rect 3486 5614 3514 5642
rect 3542 5894 3570 5922
rect 2478 5166 2506 5194
rect 2758 4942 2786 4970
rect 2142 3710 2170 3738
rect 2702 4886 2730 4914
rect 2870 4969 2898 4970
rect 2870 4943 2871 4969
rect 2871 4943 2897 4969
rect 2897 4943 2898 4969
rect 2870 4942 2898 4943
rect 6958 7014 6986 7042
rect 7182 7014 7210 7042
rect 5726 6510 5754 6538
rect 6454 6537 6482 6538
rect 6454 6511 6455 6537
rect 6455 6511 6481 6537
rect 6481 6511 6482 6537
rect 6454 6510 6482 6511
rect 3990 5558 4018 5586
rect 3766 5502 3794 5530
rect 6846 6481 6874 6482
rect 6846 6455 6847 6481
rect 6847 6455 6873 6481
rect 6873 6455 6874 6481
rect 6846 6454 6874 6455
rect 8190 7014 8218 7042
rect 8414 7014 8442 7042
rect 6454 6118 6482 6146
rect 5222 5614 5250 5642
rect 5054 5222 5082 5250
rect 5278 5222 5306 5250
rect 3542 4942 3570 4970
rect 4270 5166 4298 5194
rect 3374 4830 3402 4858
rect 2926 4774 2954 4802
rect 3038 4494 3066 4522
rect 2982 4214 3010 4242
rect 2982 3878 3010 3906
rect 2926 3822 2954 3850
rect 2758 3766 2786 3794
rect 2590 3598 2618 3626
rect 2232 3541 2260 3542
rect 2232 3515 2233 3541
rect 2233 3515 2259 3541
rect 2259 3515 2260 3541
rect 2232 3514 2260 3515
rect 2284 3541 2312 3542
rect 2284 3515 2285 3541
rect 2285 3515 2311 3541
rect 2311 3515 2312 3541
rect 2284 3514 2312 3515
rect 2336 3541 2364 3542
rect 2336 3515 2337 3541
rect 2337 3515 2363 3541
rect 2363 3515 2364 3541
rect 2478 3542 2506 3570
rect 2336 3514 2364 3515
rect 1806 3374 1834 3402
rect 1902 3149 1930 3150
rect 1902 3123 1903 3149
rect 1903 3123 1929 3149
rect 1929 3123 1930 3149
rect 1902 3122 1930 3123
rect 1954 3149 1982 3150
rect 1954 3123 1955 3149
rect 1955 3123 1981 3149
rect 1981 3123 1982 3149
rect 1954 3122 1982 3123
rect 2006 3149 2034 3150
rect 2006 3123 2007 3149
rect 2007 3123 2033 3149
rect 2033 3123 2034 3149
rect 2006 3122 2034 3123
rect 2534 3038 2562 3066
rect 2086 2926 2114 2954
rect 1806 2702 1834 2730
rect 1134 182 1162 210
rect 1470 2030 1498 2058
rect 1750 1441 1778 1442
rect 1750 1415 1751 1441
rect 1751 1415 1777 1441
rect 1777 1415 1778 1441
rect 1750 1414 1778 1415
rect 1302 1302 1330 1330
rect 1302 462 1330 490
rect 1902 2365 1930 2366
rect 1902 2339 1903 2365
rect 1903 2339 1929 2365
rect 1929 2339 1930 2365
rect 1902 2338 1930 2339
rect 1954 2365 1982 2366
rect 1954 2339 1955 2365
rect 1955 2339 1981 2365
rect 1981 2339 1982 2365
rect 1954 2338 1982 2339
rect 2006 2365 2034 2366
rect 2006 2339 2007 2365
rect 2007 2339 2033 2365
rect 2033 2339 2034 2365
rect 2006 2338 2034 2339
rect 1902 1581 1930 1582
rect 1902 1555 1903 1581
rect 1903 1555 1929 1581
rect 1929 1555 1930 1581
rect 1902 1554 1930 1555
rect 1954 1581 1982 1582
rect 1954 1555 1955 1581
rect 1955 1555 1981 1581
rect 1981 1555 1982 1581
rect 1954 1554 1982 1555
rect 2006 1581 2034 1582
rect 2006 1555 2007 1581
rect 2007 1555 2033 1581
rect 2033 1555 2034 1581
rect 2006 1554 2034 1555
rect 2646 2982 2674 3010
rect 2232 2757 2260 2758
rect 2232 2731 2233 2757
rect 2233 2731 2259 2757
rect 2259 2731 2260 2757
rect 2232 2730 2260 2731
rect 2284 2757 2312 2758
rect 2284 2731 2285 2757
rect 2285 2731 2311 2757
rect 2311 2731 2312 2757
rect 2284 2730 2312 2731
rect 2336 2757 2364 2758
rect 2336 2731 2337 2757
rect 2337 2731 2363 2757
rect 2363 2731 2364 2757
rect 2336 2730 2364 2731
rect 2142 2617 2170 2618
rect 2142 2591 2143 2617
rect 2143 2591 2169 2617
rect 2169 2591 2170 2617
rect 2142 2590 2170 2591
rect 2422 2561 2450 2562
rect 2422 2535 2423 2561
rect 2423 2535 2449 2561
rect 2449 2535 2450 2561
rect 2422 2534 2450 2535
rect 2534 2310 2562 2338
rect 2232 1973 2260 1974
rect 2232 1947 2233 1973
rect 2233 1947 2259 1973
rect 2259 1947 2260 1973
rect 2232 1946 2260 1947
rect 2284 1973 2312 1974
rect 2284 1947 2285 1973
rect 2285 1947 2311 1973
rect 2311 1947 2312 1973
rect 2284 1946 2312 1947
rect 2336 1973 2364 1974
rect 2336 1947 2337 1973
rect 2337 1947 2363 1973
rect 2363 1947 2364 1973
rect 2336 1946 2364 1947
rect 2478 1582 2506 1610
rect 2232 1189 2260 1190
rect 2232 1163 2233 1189
rect 2233 1163 2259 1189
rect 2259 1163 2260 1189
rect 2232 1162 2260 1163
rect 2284 1189 2312 1190
rect 2284 1163 2285 1189
rect 2285 1163 2311 1189
rect 2311 1163 2312 1189
rect 2284 1162 2312 1163
rect 2336 1189 2364 1190
rect 2336 1163 2337 1189
rect 2337 1163 2363 1189
rect 2363 1163 2364 1189
rect 2336 1162 2364 1163
rect 2534 1414 2562 1442
rect 2590 2086 2618 2114
rect 2758 2758 2786 2786
rect 2646 1806 2674 1834
rect 2702 2198 2730 2226
rect 2702 1302 2730 1330
rect 2870 3681 2898 3682
rect 2870 3655 2871 3681
rect 2871 3655 2897 3681
rect 2897 3655 2898 3681
rect 2870 3654 2898 3655
rect 2926 3598 2954 3626
rect 2870 3430 2898 3458
rect 3038 2926 3066 2954
rect 3094 4214 3122 4242
rect 2926 2478 2954 2506
rect 3374 4102 3402 4130
rect 3766 4270 3794 4298
rect 3486 4046 3514 4074
rect 3206 3990 3234 4018
rect 3094 2254 3122 2282
rect 2870 2142 2898 2170
rect 2814 1078 2842 1106
rect 2590 1022 2618 1050
rect 3150 854 3178 882
rect 1902 797 1930 798
rect 1902 771 1903 797
rect 1903 771 1929 797
rect 1929 771 1930 797
rect 1902 770 1930 771
rect 1954 797 1982 798
rect 1954 771 1955 797
rect 1955 771 1981 797
rect 1981 771 1982 797
rect 1954 770 1982 771
rect 2006 797 2034 798
rect 2006 771 2007 797
rect 2007 771 2033 797
rect 2033 771 2034 797
rect 2006 770 2034 771
rect 1806 462 1834 490
rect 2232 405 2260 406
rect 2232 379 2233 405
rect 2233 379 2259 405
rect 2259 379 2260 405
rect 2232 378 2260 379
rect 2284 405 2312 406
rect 2284 379 2285 405
rect 2285 379 2311 405
rect 2311 379 2312 405
rect 2284 378 2312 379
rect 2336 405 2364 406
rect 2336 379 2337 405
rect 2337 379 2363 405
rect 2363 379 2364 405
rect 2336 378 2364 379
rect 3710 3654 3738 3682
rect 3318 3038 3346 3066
rect 3318 1582 3346 1610
rect 3374 2982 3402 3010
rect 3542 1694 3570 1722
rect 3318 686 3346 714
rect 4158 3262 4186 3290
rect 3934 1974 3962 2002
rect 4326 5110 4354 5138
rect 4326 3598 4354 3626
rect 4382 4942 4410 4970
rect 4270 3318 4298 3346
rect 4214 1918 4242 1946
rect 7126 5894 7154 5922
rect 6454 4942 6482 4970
rect 6958 5446 6986 5474
rect 7574 5641 7602 5642
rect 7574 5615 7575 5641
rect 7575 5615 7601 5641
rect 7601 5615 7602 5641
rect 7574 5614 7602 5615
rect 7126 4942 7154 4970
rect 7462 5502 7490 5530
rect 6958 4774 6986 4802
rect 6174 4662 6202 4690
rect 5278 4606 5306 4634
rect 5558 4326 5586 4354
rect 4494 3625 4522 3626
rect 4494 3599 4495 3625
rect 4495 3599 4521 3625
rect 4521 3599 4522 3625
rect 4494 3598 4522 3599
rect 5558 3486 5586 3514
rect 4382 1862 4410 1890
rect 4998 2814 5026 2842
rect 3710 1134 3738 1162
rect 3542 574 3570 602
rect 3206 126 3234 154
rect 1246 70 1274 98
rect 6006 3262 6034 3290
rect 5894 2142 5922 2170
rect 5782 1974 5810 2002
rect 5222 1526 5250 1554
rect 4998 462 5026 490
rect 5670 1441 5698 1442
rect 5670 1415 5671 1441
rect 5671 1415 5697 1441
rect 5697 1415 5698 1441
rect 5670 1414 5698 1415
rect 5390 910 5418 938
rect 5670 937 5698 938
rect 5670 911 5671 937
rect 5671 911 5697 937
rect 5697 911 5698 937
rect 5670 910 5698 911
rect 5838 993 5866 994
rect 5838 967 5839 993
rect 5839 967 5865 993
rect 5865 967 5866 993
rect 5838 966 5866 967
rect 7070 3878 7098 3906
rect 6790 3766 6818 3794
rect 6174 3038 6202 3066
rect 6510 3094 6538 3122
rect 6118 2897 6146 2898
rect 6118 2871 6119 2897
rect 6119 2871 6145 2897
rect 6145 2871 6146 2897
rect 6118 2870 6146 2871
rect 6118 2702 6146 2730
rect 6118 2310 6146 2338
rect 6342 2590 6370 2618
rect 6454 2590 6482 2618
rect 6342 1470 6370 1498
rect 6006 686 6034 714
rect 6622 2926 6650 2954
rect 6510 1358 6538 1386
rect 6566 2478 6594 2506
rect 6678 2841 6706 2842
rect 6678 2815 6679 2841
rect 6679 2815 6705 2841
rect 6705 2815 6706 2841
rect 6678 2814 6706 2815
rect 6622 2422 6650 2450
rect 6734 2366 6762 2394
rect 6398 630 6426 658
rect 5782 406 5810 434
rect 6510 462 6538 490
rect 5278 238 5306 266
rect 6398 182 6426 210
rect 6286 126 6314 154
rect 6174 70 6202 98
rect 6790 1638 6818 1666
rect 6958 3598 6986 3626
rect 6734 1526 6762 1554
rect 6678 798 6706 826
rect 6734 742 6762 770
rect 6846 686 6874 714
rect 7070 3262 7098 3290
rect 7126 3654 7154 3682
rect 9198 6846 9226 6874
rect 8862 6566 8890 6594
rect 8806 6454 8834 6482
rect 7798 5838 7826 5866
rect 8918 6398 8946 6426
rect 8862 5782 8890 5810
rect 9086 5950 9114 5978
rect 8358 5166 8386 5194
rect 7686 4774 7714 4802
rect 7462 3038 7490 3066
rect 7126 2982 7154 3010
rect 7182 2870 7210 2898
rect 7070 2646 7098 2674
rect 7070 966 7098 994
rect 7518 2814 7546 2842
rect 7350 2561 7378 2562
rect 7350 2535 7351 2561
rect 7351 2535 7377 2561
rect 7377 2535 7378 2561
rect 7350 2534 7378 2535
rect 7294 798 7322 826
rect 7406 798 7434 826
rect 7630 2534 7658 2562
rect 8358 4886 8386 4914
rect 8078 4606 8106 4634
rect 8302 4438 8330 4466
rect 7966 3486 7994 3514
rect 8190 2926 8218 2954
rect 8022 1134 8050 1162
rect 8078 2870 8106 2898
rect 8750 4326 8778 4354
rect 8358 4214 8386 4242
rect 8358 3822 8386 3850
rect 8358 2422 8386 2450
rect 8358 2310 8386 2338
rect 8302 1694 8330 1722
rect 8526 2814 8554 2842
rect 8470 798 8498 826
rect 8414 462 8442 490
rect 8302 70 8330 98
rect 8638 1358 8666 1386
rect 8694 1190 8722 1218
rect 8638 798 8666 826
rect 10654 7014 10682 7042
rect 10878 7014 10906 7042
rect 9758 6481 9786 6482
rect 9758 6455 9759 6481
rect 9759 6455 9785 6481
rect 9785 6455 9786 6481
rect 9758 6454 9786 6455
rect 11886 7014 11914 7042
rect 12110 7014 12138 7042
rect 10934 6062 10962 6090
rect 10150 6006 10178 6034
rect 9534 5614 9562 5642
rect 9310 4550 9338 4578
rect 9198 3094 9226 3122
rect 9310 4102 9338 4130
rect 9478 3990 9506 4018
rect 9254 2870 9282 2898
rect 9366 3150 9394 3178
rect 9198 2030 9226 2058
rect 9254 1974 9282 2002
rect 9030 742 9058 770
rect 9422 1246 9450 1274
rect 9254 518 9282 546
rect 9310 294 9338 322
rect 10094 4998 10122 5026
rect 9646 3486 9674 3514
rect 9870 3598 9898 3626
rect 9646 3318 9674 3346
rect 9758 1918 9786 1946
rect 10038 3934 10066 3962
rect 9982 3486 10010 3514
rect 9982 2478 10010 2506
rect 10150 4438 10178 4466
rect 10262 5558 10290 5586
rect 10094 3374 10122 3402
rect 10150 3766 10178 3794
rect 9926 518 9954 546
rect 10206 2478 10234 2506
rect 10710 5334 10738 5362
rect 10486 5054 10514 5082
rect 10486 4830 10514 4858
rect 10654 3878 10682 3906
rect 10598 2982 10626 3010
rect 10486 2422 10514 2450
rect 10486 2254 10514 2282
rect 10262 1414 10290 1442
rect 10318 966 10346 994
rect 10262 601 10290 602
rect 10262 575 10263 601
rect 10263 575 10289 601
rect 10289 575 10290 601
rect 10262 574 10290 575
rect 10374 294 10402 322
rect 10486 518 10514 546
rect 12232 6677 12260 6678
rect 12232 6651 12233 6677
rect 12233 6651 12259 6677
rect 12259 6651 12260 6677
rect 12232 6650 12260 6651
rect 12284 6677 12312 6678
rect 12284 6651 12285 6677
rect 12285 6651 12311 6677
rect 12311 6651 12312 6677
rect 12284 6650 12312 6651
rect 12336 6677 12364 6678
rect 12336 6651 12337 6677
rect 12337 6651 12363 6677
rect 12363 6651 12364 6677
rect 12336 6650 12364 6651
rect 11494 6342 11522 6370
rect 11902 6285 11930 6286
rect 11902 6259 11903 6285
rect 11903 6259 11929 6285
rect 11929 6259 11930 6285
rect 11902 6258 11930 6259
rect 11954 6285 11982 6286
rect 11954 6259 11955 6285
rect 11955 6259 11981 6285
rect 11981 6259 11982 6285
rect 11954 6258 11982 6259
rect 12006 6285 12034 6286
rect 12006 6259 12007 6285
rect 12007 6259 12033 6285
rect 12033 6259 12034 6285
rect 12006 6258 12034 6259
rect 11494 5838 11522 5866
rect 11550 6174 11578 6202
rect 10934 4662 10962 4690
rect 11046 5278 11074 5306
rect 10934 4494 10962 4522
rect 10934 3654 10962 3682
rect 10990 3625 11018 3626
rect 10990 3599 10991 3625
rect 10991 3599 11017 3625
rect 11017 3599 11018 3625
rect 10990 3598 11018 3599
rect 10934 2646 10962 2674
rect 11438 4942 11466 4970
rect 11270 3681 11298 3682
rect 11270 3655 11271 3681
rect 11271 3655 11297 3681
rect 11297 3655 11298 3681
rect 11270 3654 11298 3655
rect 12232 5893 12260 5894
rect 12232 5867 12233 5893
rect 12233 5867 12259 5893
rect 12259 5867 12260 5893
rect 12232 5866 12260 5867
rect 12284 5893 12312 5894
rect 12284 5867 12285 5893
rect 12285 5867 12311 5893
rect 12311 5867 12312 5893
rect 12284 5866 12312 5867
rect 12336 5893 12364 5894
rect 12336 5867 12337 5893
rect 12337 5867 12363 5893
rect 12363 5867 12364 5893
rect 12336 5866 12364 5867
rect 12110 5614 12138 5642
rect 12614 6454 12642 6482
rect 12558 5614 12586 5642
rect 11902 5501 11930 5502
rect 11902 5475 11903 5501
rect 11903 5475 11929 5501
rect 11929 5475 11930 5501
rect 11902 5474 11930 5475
rect 11954 5501 11982 5502
rect 11954 5475 11955 5501
rect 11955 5475 11981 5501
rect 11981 5475 11982 5501
rect 11954 5474 11982 5475
rect 12006 5501 12034 5502
rect 12006 5475 12007 5501
rect 12007 5475 12033 5501
rect 12033 5475 12034 5501
rect 12110 5502 12138 5530
rect 12006 5474 12034 5475
rect 14350 7014 14378 7042
rect 14574 7014 14602 7042
rect 14126 6566 14154 6594
rect 12614 5278 12642 5306
rect 11718 5110 11746 5138
rect 11606 4438 11634 4466
rect 12232 5109 12260 5110
rect 12232 5083 12233 5109
rect 12233 5083 12259 5109
rect 12259 5083 12260 5109
rect 12232 5082 12260 5083
rect 12284 5109 12312 5110
rect 12284 5083 12285 5109
rect 12285 5083 12311 5109
rect 12311 5083 12312 5109
rect 12284 5082 12312 5083
rect 12336 5109 12364 5110
rect 12336 5083 12337 5109
rect 12337 5083 12363 5109
rect 12363 5083 12364 5109
rect 12336 5082 12364 5083
rect 12446 5110 12474 5138
rect 11902 4717 11930 4718
rect 11902 4691 11903 4717
rect 11903 4691 11929 4717
rect 11929 4691 11930 4717
rect 11902 4690 11930 4691
rect 11954 4717 11982 4718
rect 11954 4691 11955 4717
rect 11955 4691 11981 4717
rect 11981 4691 11982 4717
rect 11954 4690 11982 4691
rect 12006 4717 12034 4718
rect 12006 4691 12007 4717
rect 12007 4691 12033 4717
rect 12033 4691 12034 4717
rect 12006 4690 12034 4691
rect 12446 4550 12474 4578
rect 11718 4158 11746 4186
rect 12110 4326 12138 4354
rect 11606 3878 11634 3906
rect 11662 4102 11690 4130
rect 11046 2310 11074 2338
rect 11102 2646 11130 2674
rect 10934 2254 10962 2282
rect 10990 1414 11018 1442
rect 10878 854 10906 882
rect 10822 126 10850 154
rect 10766 70 10794 98
rect 11046 630 11074 658
rect 11270 2590 11298 2618
rect 11214 2534 11242 2562
rect 11158 1302 11186 1330
rect 11158 798 11186 826
rect 11382 1833 11410 1834
rect 11382 1807 11383 1833
rect 11383 1807 11409 1833
rect 11409 1807 11410 1833
rect 11382 1806 11410 1807
rect 11438 1750 11466 1778
rect 11326 1273 11354 1274
rect 11326 1247 11327 1273
rect 11327 1247 11353 1273
rect 11353 1247 11354 1273
rect 11326 1246 11354 1247
rect 11998 4073 12026 4074
rect 11998 4047 11999 4073
rect 11999 4047 12025 4073
rect 12025 4047 12026 4073
rect 11998 4046 12026 4047
rect 11774 3934 11802 3962
rect 11902 3933 11930 3934
rect 11902 3907 11903 3933
rect 11903 3907 11929 3933
rect 11929 3907 11930 3933
rect 11902 3906 11930 3907
rect 11954 3933 11982 3934
rect 11954 3907 11955 3933
rect 11955 3907 11981 3933
rect 11981 3907 11982 3933
rect 11954 3906 11982 3907
rect 12006 3933 12034 3934
rect 12006 3907 12007 3933
rect 12007 3907 12033 3933
rect 12033 3907 12034 3933
rect 12006 3906 12034 3907
rect 12232 4325 12260 4326
rect 12232 4299 12233 4325
rect 12233 4299 12259 4325
rect 12259 4299 12260 4325
rect 12232 4298 12260 4299
rect 12284 4325 12312 4326
rect 12284 4299 12285 4325
rect 12285 4299 12311 4325
rect 12311 4299 12312 4325
rect 12284 4298 12312 4299
rect 12336 4325 12364 4326
rect 12336 4299 12337 4325
rect 12337 4299 12363 4325
rect 12363 4299 12364 4325
rect 12336 4298 12364 4299
rect 12110 3878 12138 3906
rect 12670 5950 12698 5978
rect 12558 5166 12586 5194
rect 12558 4774 12586 4802
rect 12726 5697 12754 5698
rect 12726 5671 12727 5697
rect 12727 5671 12753 5697
rect 12753 5671 12754 5697
rect 12726 5670 12754 5671
rect 13342 5558 13370 5586
rect 12726 5334 12754 5362
rect 13790 6342 13818 6370
rect 13622 5193 13650 5194
rect 13622 5167 13623 5193
rect 13623 5167 13649 5193
rect 13649 5167 13650 5193
rect 13622 5166 13650 5167
rect 13398 4718 13426 4746
rect 12726 4606 12754 4634
rect 12670 4494 12698 4522
rect 13678 4270 13706 4298
rect 13678 4158 13706 4186
rect 13902 5838 13930 5866
rect 15582 7014 15610 7042
rect 15862 7014 15890 7042
rect 14742 6846 14770 6874
rect 14126 5670 14154 5698
rect 13902 5558 13930 5586
rect 13790 4158 13818 4186
rect 14014 5446 14042 5474
rect 13678 3990 13706 4018
rect 12502 3822 12530 3850
rect 13398 3878 13426 3906
rect 12278 3766 12306 3794
rect 12232 3541 12260 3542
rect 12232 3515 12233 3541
rect 12233 3515 12259 3541
rect 12259 3515 12260 3541
rect 12232 3514 12260 3515
rect 12284 3541 12312 3542
rect 12284 3515 12285 3541
rect 12285 3515 12311 3541
rect 12311 3515 12312 3541
rect 12284 3514 12312 3515
rect 12336 3541 12364 3542
rect 12336 3515 12337 3541
rect 12337 3515 12363 3541
rect 12363 3515 12364 3541
rect 12336 3514 12364 3515
rect 12670 3598 12698 3626
rect 12558 3374 12586 3402
rect 12614 3486 12642 3514
rect 11662 3206 11690 3234
rect 11902 3149 11930 3150
rect 11902 3123 11903 3149
rect 11903 3123 11929 3149
rect 11929 3123 11930 3149
rect 11902 3122 11930 3123
rect 11954 3149 11982 3150
rect 11954 3123 11955 3149
rect 11955 3123 11981 3149
rect 11981 3123 11982 3149
rect 11954 3122 11982 3123
rect 12006 3149 12034 3150
rect 12006 3123 12007 3149
rect 12007 3123 12033 3149
rect 12033 3123 12034 3149
rect 12006 3122 12034 3123
rect 12614 3038 12642 3066
rect 12166 2758 12194 2786
rect 13006 3374 13034 3402
rect 12232 2757 12260 2758
rect 12232 2731 12233 2757
rect 12233 2731 12259 2757
rect 12259 2731 12260 2757
rect 12232 2730 12260 2731
rect 12284 2757 12312 2758
rect 12284 2731 12285 2757
rect 12285 2731 12311 2757
rect 12311 2731 12312 2757
rect 12284 2730 12312 2731
rect 12336 2757 12364 2758
rect 12336 2731 12337 2757
rect 12337 2731 12363 2757
rect 12363 2731 12364 2757
rect 12670 2758 12698 2786
rect 12782 2926 12810 2954
rect 12336 2730 12364 2731
rect 12894 2870 12922 2898
rect 12670 2478 12698 2506
rect 11902 2365 11930 2366
rect 11902 2339 11903 2365
rect 11903 2339 11929 2365
rect 11929 2339 11930 2365
rect 11902 2338 11930 2339
rect 11954 2365 11982 2366
rect 11954 2339 11955 2365
rect 11955 2339 11981 2365
rect 11981 2339 11982 2365
rect 11954 2338 11982 2339
rect 12006 2365 12034 2366
rect 12006 2339 12007 2365
rect 12007 2339 12033 2365
rect 12033 2339 12034 2365
rect 12166 2366 12194 2394
rect 12558 2366 12586 2394
rect 12006 2338 12034 2339
rect 12110 2310 12138 2338
rect 11830 2169 11858 2170
rect 11830 2143 11831 2169
rect 11831 2143 11857 2169
rect 11857 2143 11858 2169
rect 11830 2142 11858 2143
rect 11998 2113 12026 2114
rect 11998 2087 11999 2113
rect 11999 2087 12025 2113
rect 12025 2087 12026 2113
rect 11998 2086 12026 2087
rect 12054 1974 12082 2002
rect 11550 1918 11578 1946
rect 11494 1302 11522 1330
rect 11550 1806 11578 1834
rect 11382 1049 11410 1050
rect 11382 1023 11383 1049
rect 11383 1023 11409 1049
rect 11409 1023 11410 1049
rect 11382 1022 11410 1023
rect 11494 1134 11522 1162
rect 11494 1022 11522 1050
rect 11494 238 11522 266
rect 11774 1385 11802 1386
rect 11774 1359 11775 1385
rect 11775 1359 11801 1385
rect 11801 1359 11802 1385
rect 11774 1358 11802 1359
rect 11606 1329 11634 1330
rect 11606 1303 11607 1329
rect 11607 1303 11633 1329
rect 11633 1303 11634 1329
rect 11606 1302 11634 1303
rect 11774 1246 11802 1274
rect 11902 1581 11930 1582
rect 11902 1555 11903 1581
rect 11903 1555 11929 1581
rect 11929 1555 11930 1581
rect 11902 1554 11930 1555
rect 11954 1581 11982 1582
rect 11954 1555 11955 1581
rect 11955 1555 11981 1581
rect 11981 1555 11982 1581
rect 11954 1554 11982 1555
rect 12006 1581 12034 1582
rect 12006 1555 12007 1581
rect 12007 1555 12033 1581
rect 12033 1555 12034 1581
rect 12006 1554 12034 1555
rect 11998 1414 12026 1442
rect 11998 1190 12026 1218
rect 11902 797 11930 798
rect 11902 771 11903 797
rect 11903 771 11929 797
rect 11929 771 11930 797
rect 11902 770 11930 771
rect 11954 797 11982 798
rect 11954 771 11955 797
rect 11955 771 11981 797
rect 11981 771 11982 797
rect 11954 770 11982 771
rect 12006 797 12034 798
rect 12006 771 12007 797
rect 12007 771 12033 797
rect 12033 771 12034 797
rect 12006 770 12034 771
rect 11774 294 11802 322
rect 11886 462 11914 490
rect 11774 182 11802 210
rect 12232 1973 12260 1974
rect 12232 1947 12233 1973
rect 12233 1947 12259 1973
rect 12259 1947 12260 1973
rect 12232 1946 12260 1947
rect 12284 1973 12312 1974
rect 12284 1947 12285 1973
rect 12285 1947 12311 1973
rect 12311 1947 12312 1973
rect 12284 1946 12312 1947
rect 12336 1973 12364 1974
rect 12336 1947 12337 1973
rect 12337 1947 12363 1973
rect 12363 1947 12364 1973
rect 12336 1946 12364 1947
rect 12670 2366 12698 2394
rect 12782 2198 12810 2226
rect 13398 3262 13426 3290
rect 13230 3150 13258 3178
rect 13062 2505 13090 2506
rect 13062 2479 13063 2505
rect 13063 2479 13089 2505
rect 13089 2479 13090 2505
rect 13062 2478 13090 2479
rect 12894 2198 12922 2226
rect 12838 1974 12866 2002
rect 12614 1777 12642 1778
rect 12614 1751 12615 1777
rect 12615 1751 12641 1777
rect 12641 1751 12642 1777
rect 12614 1750 12642 1751
rect 13006 1862 13034 1890
rect 12614 1638 12642 1666
rect 12232 1189 12260 1190
rect 12232 1163 12233 1189
rect 12233 1163 12259 1189
rect 12259 1163 12260 1189
rect 12232 1162 12260 1163
rect 12284 1189 12312 1190
rect 12284 1163 12285 1189
rect 12285 1163 12311 1189
rect 12311 1163 12312 1189
rect 12284 1162 12312 1163
rect 12336 1189 12364 1190
rect 12336 1163 12337 1189
rect 12337 1163 12363 1189
rect 12363 1163 12364 1189
rect 12336 1162 12364 1163
rect 12166 406 12194 434
rect 12232 405 12260 406
rect 12232 379 12233 405
rect 12233 379 12259 405
rect 12259 379 12260 405
rect 12232 378 12260 379
rect 12284 405 12312 406
rect 12284 379 12285 405
rect 12285 379 12311 405
rect 12311 379 12312 405
rect 12284 378 12312 379
rect 12336 405 12364 406
rect 12336 379 12337 405
rect 12337 379 12363 405
rect 12363 379 12364 405
rect 12336 378 12364 379
rect 12110 126 12138 154
rect 12334 294 12362 322
rect 12614 910 12642 938
rect 12558 545 12586 546
rect 12558 519 12559 545
rect 12559 519 12585 545
rect 12585 519 12586 545
rect 12558 518 12586 519
rect 12502 182 12530 210
rect 12558 238 12586 266
rect 12950 1526 12978 1554
rect 12726 937 12754 938
rect 12726 911 12727 937
rect 12727 911 12753 937
rect 12753 911 12754 937
rect 12726 910 12754 911
rect 12894 1078 12922 1106
rect 12838 966 12866 994
rect 12838 854 12866 882
rect 12894 574 12922 602
rect 12950 126 12978 154
rect 13006 518 13034 546
rect 13398 2478 13426 2506
rect 13230 1078 13258 1106
rect 13062 238 13090 266
rect 13230 686 13258 714
rect 13342 1470 13370 1498
rect 13286 574 13314 602
rect 13454 1750 13482 1778
rect 13622 1526 13650 1554
rect 13454 798 13482 826
rect 13510 1470 13538 1498
rect 13902 3598 13930 3626
rect 13622 686 13650 714
rect 13510 630 13538 658
rect 13398 574 13426 602
rect 13790 2758 13818 2786
rect 13790 1526 13818 1554
rect 14238 5110 14266 5138
rect 14126 4774 14154 4802
rect 14350 5110 14378 5138
rect 14350 4942 14378 4970
rect 14238 4774 14266 4802
rect 14686 4718 14714 4746
rect 14126 4494 14154 4522
rect 14350 4662 14378 4690
rect 14014 2422 14042 2450
rect 14238 3766 14266 3794
rect 14294 2030 14322 2058
rect 14126 1833 14154 1834
rect 14126 1807 14127 1833
rect 14127 1807 14153 1833
rect 14153 1807 14154 1833
rect 14126 1806 14154 1807
rect 14238 1806 14266 1834
rect 13902 1190 13930 1218
rect 13454 462 13482 490
rect 14014 798 14042 826
rect 13902 630 13930 658
rect 13846 601 13874 602
rect 13846 575 13847 601
rect 13847 575 13873 601
rect 13873 575 13874 601
rect 13846 574 13874 575
rect 13510 406 13538 434
rect 13510 294 13538 322
rect 13790 294 13818 322
rect 13678 238 13706 266
rect 14518 2478 14546 2506
rect 14686 2310 14714 2338
rect 14686 2169 14714 2170
rect 14686 2143 14687 2169
rect 14687 2143 14713 2169
rect 14713 2143 14714 2169
rect 14686 2142 14714 2143
rect 14574 2030 14602 2058
rect 14350 798 14378 826
rect 14406 1134 14434 1162
rect 14350 574 14378 602
rect 14126 489 14154 490
rect 14126 463 14127 489
rect 14127 463 14153 489
rect 14153 463 14154 489
rect 14126 462 14154 463
rect 14070 406 14098 434
rect 14182 350 14210 378
rect 14238 462 14266 490
rect 14126 182 14154 210
rect 14462 1049 14490 1050
rect 14462 1023 14463 1049
rect 14463 1023 14489 1049
rect 14489 1023 14490 1049
rect 14462 1022 14490 1023
rect 14406 518 14434 546
rect 14462 686 14490 714
rect 14518 630 14546 658
rect 15246 6734 15274 6762
rect 16366 6118 16394 6146
rect 16590 6398 16618 6426
rect 18046 7014 18074 7042
rect 18270 7014 18298 7042
rect 17038 6145 17066 6146
rect 17038 6119 17039 6145
rect 17039 6119 17065 6145
rect 17065 6119 17066 6145
rect 17038 6118 17066 6119
rect 14798 6006 14826 6034
rect 14798 5614 14826 5642
rect 14854 5894 14882 5922
rect 14854 4942 14882 4970
rect 14910 5726 14938 5754
rect 14910 4438 14938 4466
rect 15918 6062 15946 6090
rect 15134 5782 15162 5810
rect 14966 4326 14994 4354
rect 15022 5390 15050 5418
rect 14910 4270 14938 4298
rect 14854 4046 14882 4074
rect 14910 3654 14938 3682
rect 15078 5334 15106 5362
rect 15078 4494 15106 4522
rect 15190 5502 15218 5530
rect 15022 3822 15050 3850
rect 15078 3990 15106 4018
rect 14966 3318 14994 3346
rect 15078 2982 15106 3010
rect 16870 6033 16898 6034
rect 16870 6007 16871 6033
rect 16871 6007 16897 6033
rect 16897 6007 16898 6033
rect 16870 6006 16898 6007
rect 15918 5782 15946 5810
rect 15526 5054 15554 5082
rect 15974 5390 16002 5418
rect 15470 4550 15498 4578
rect 15246 4158 15274 4186
rect 15414 3374 15442 3402
rect 15302 3262 15330 3290
rect 15246 2870 15274 2898
rect 15078 2561 15106 2562
rect 15078 2535 15079 2561
rect 15079 2535 15105 2561
rect 15105 2535 15106 2561
rect 15078 2534 15106 2535
rect 15134 2422 15162 2450
rect 14966 2057 14994 2058
rect 14966 2031 14967 2057
rect 14967 2031 14993 2057
rect 14993 2031 14994 2057
rect 14966 2030 14994 2031
rect 14798 1134 14826 1162
rect 14742 1078 14770 1106
rect 15022 1022 15050 1050
rect 14630 742 14658 770
rect 14686 518 14714 546
rect 14742 294 14770 322
rect 14798 630 14826 658
rect 14854 238 14882 266
rect 14910 350 14938 378
rect 15246 1638 15274 1666
rect 15358 2590 15386 2618
rect 15862 4270 15890 4298
rect 15638 3206 15666 3234
rect 15750 2982 15778 3010
rect 15582 2702 15610 2730
rect 15526 2449 15554 2450
rect 15526 2423 15527 2449
rect 15527 2423 15553 2449
rect 15553 2423 15554 2449
rect 15526 2422 15554 2423
rect 15694 2198 15722 2226
rect 15302 1358 15330 1386
rect 15358 1694 15386 1722
rect 15190 686 15218 714
rect 15302 574 15330 602
rect 15246 294 15274 322
rect 15694 1974 15722 2002
rect 15750 1806 15778 1834
rect 16086 4998 16114 5026
rect 16142 5614 16170 5642
rect 15974 3486 16002 3514
rect 16030 4550 16058 4578
rect 15862 2422 15890 2450
rect 16086 3766 16114 3794
rect 16086 3262 16114 3290
rect 16030 2590 16058 2618
rect 15918 2254 15946 2282
rect 15974 2310 16002 2338
rect 15470 1582 15498 1610
rect 15414 1414 15442 1442
rect 15806 1582 15834 1610
rect 15862 1022 15890 1050
rect 15918 1638 15946 1666
rect 15470 686 15498 714
rect 15750 854 15778 882
rect 15694 798 15722 826
rect 15526 182 15554 210
rect 15582 238 15610 266
rect 15750 126 15778 154
rect 15862 574 15890 602
rect 16198 4857 16226 4858
rect 16198 4831 16199 4857
rect 16199 4831 16225 4857
rect 16225 4831 16226 4857
rect 16198 4830 16226 4831
rect 17318 5977 17346 5978
rect 17318 5951 17319 5977
rect 17319 5951 17345 5977
rect 17345 5951 17346 5977
rect 17318 5950 17346 5951
rect 16814 5558 16842 5586
rect 16702 5054 16730 5082
rect 16478 4270 16506 4298
rect 16646 4606 16674 4634
rect 16254 3822 16282 3850
rect 16310 2590 16338 2618
rect 16198 2561 16226 2562
rect 16198 2535 16199 2561
rect 16199 2535 16225 2561
rect 16225 2535 16226 2561
rect 16198 2534 16226 2535
rect 16478 2534 16506 2562
rect 16534 2870 16562 2898
rect 16142 2254 16170 2282
rect 16198 1777 16226 1778
rect 16198 1751 16199 1777
rect 16199 1751 16225 1777
rect 16225 1751 16226 1777
rect 16198 1750 16226 1751
rect 15974 1582 16002 1610
rect 16198 1302 16226 1330
rect 16086 630 16114 658
rect 16030 489 16058 490
rect 16030 463 16031 489
rect 16031 463 16057 489
rect 16057 463 16058 489
rect 16030 462 16058 463
rect 16590 2702 16618 2730
rect 16310 2030 16338 2058
rect 16142 182 16170 210
rect 16478 1721 16506 1722
rect 16478 1695 16479 1721
rect 16479 1695 16505 1721
rect 16505 1695 16506 1721
rect 16478 1694 16506 1695
rect 16646 2478 16674 2506
rect 16646 1694 16674 1722
rect 16422 798 16450 826
rect 20510 7014 20538 7042
rect 20678 7014 20706 7042
rect 19278 6566 19306 6594
rect 19838 6593 19866 6594
rect 19838 6567 19839 6593
rect 19839 6567 19865 6593
rect 19865 6567 19866 6593
rect 19838 6566 19866 6567
rect 17374 5334 17402 5362
rect 17430 6286 17458 6314
rect 16814 4158 16842 4186
rect 16870 3654 16898 3682
rect 16758 2870 16786 2898
rect 16702 1302 16730 1330
rect 16534 601 16562 602
rect 16534 575 16535 601
rect 16535 575 16561 601
rect 16561 575 16562 601
rect 16534 574 16562 575
rect 16478 406 16506 434
rect 16534 462 16562 490
rect 16870 1414 16898 1442
rect 16870 686 16898 714
rect 16814 518 16842 546
rect 16982 2142 17010 2170
rect 17094 1665 17122 1666
rect 17094 1639 17095 1665
rect 17095 1639 17121 1665
rect 17121 1639 17122 1665
rect 17094 1638 17122 1639
rect 17374 2534 17402 2562
rect 17318 2057 17346 2058
rect 17318 2031 17319 2057
rect 17319 2031 17345 2057
rect 17345 2031 17346 2057
rect 17318 2030 17346 2031
rect 17262 1750 17290 1778
rect 16758 126 16786 154
rect 16926 126 16954 154
rect 17262 294 17290 322
rect 18494 6174 18522 6202
rect 17654 5894 17682 5922
rect 17654 5614 17682 5642
rect 17654 5278 17682 5306
rect 18830 6145 18858 6146
rect 18830 6119 18831 6145
rect 18831 6119 18857 6145
rect 18857 6119 18858 6145
rect 18830 6118 18858 6119
rect 18494 5278 18522 5306
rect 18662 6006 18690 6034
rect 17822 3822 17850 3850
rect 17654 3150 17682 3178
rect 17766 3318 17794 3346
rect 17598 2870 17626 2898
rect 17654 2590 17682 2618
rect 17598 1833 17626 1834
rect 17598 1807 17599 1833
rect 17599 1807 17625 1833
rect 17625 1807 17626 1833
rect 17598 1806 17626 1807
rect 17598 1441 17626 1442
rect 17598 1415 17599 1441
rect 17599 1415 17625 1441
rect 17625 1415 17626 1441
rect 17598 1414 17626 1415
rect 17430 1078 17458 1106
rect 17486 798 17514 826
rect 17710 742 17738 770
rect 17598 518 17626 546
rect 17766 574 17794 602
rect 17878 3430 17906 3458
rect 18102 5110 18130 5138
rect 18046 3374 18074 3402
rect 17878 2702 17906 2730
rect 17990 2561 18018 2562
rect 17990 2535 17991 2561
rect 17991 2535 18017 2561
rect 18017 2535 18018 2561
rect 17990 2534 18018 2535
rect 17934 1806 17962 1834
rect 17878 1721 17906 1722
rect 17878 1695 17879 1721
rect 17879 1695 17905 1721
rect 17905 1695 17906 1721
rect 17878 1694 17906 1695
rect 17878 881 17906 882
rect 17878 855 17879 881
rect 17879 855 17905 881
rect 17905 855 17906 881
rect 17878 854 17906 855
rect 17934 238 17962 266
rect 17934 70 17962 98
rect 18326 4270 18354 4298
rect 18158 2646 18186 2674
rect 18102 350 18130 378
rect 18158 1358 18186 1386
rect 22232 6677 22260 6678
rect 22232 6651 22233 6677
rect 22233 6651 22259 6677
rect 22259 6651 22260 6677
rect 22232 6650 22260 6651
rect 22284 6677 22312 6678
rect 22284 6651 22285 6677
rect 22285 6651 22311 6677
rect 22311 6651 22312 6677
rect 22284 6650 22312 6651
rect 22336 6677 22364 6678
rect 22336 6651 22337 6677
rect 22337 6651 22363 6677
rect 22363 6651 22364 6677
rect 22336 6650 22364 6651
rect 21854 6566 21882 6594
rect 22134 6593 22162 6594
rect 22134 6567 22135 6593
rect 22135 6567 22161 6593
rect 22161 6567 22162 6593
rect 22134 6566 22162 6567
rect 23478 6958 23506 6986
rect 22974 6566 23002 6594
rect 23030 6902 23058 6930
rect 21126 6510 21154 6538
rect 19558 6118 19586 6146
rect 19334 6062 19362 6090
rect 19054 5838 19082 5866
rect 18718 5361 18746 5362
rect 18718 5335 18719 5361
rect 18719 5335 18745 5361
rect 18745 5335 18746 5361
rect 18718 5334 18746 5335
rect 18942 5166 18970 5194
rect 18886 4158 18914 4186
rect 18550 3430 18578 3458
rect 18382 3262 18410 3290
rect 18494 2086 18522 2114
rect 18382 1329 18410 1330
rect 18382 1303 18383 1329
rect 18383 1303 18409 1329
rect 18409 1303 18410 1329
rect 18382 1302 18410 1303
rect 18606 2953 18634 2954
rect 18606 2927 18607 2953
rect 18607 2927 18633 2953
rect 18633 2927 18634 2953
rect 18606 2926 18634 2927
rect 18550 1190 18578 1218
rect 18382 993 18410 994
rect 18382 967 18383 993
rect 18383 967 18409 993
rect 18409 967 18410 993
rect 18382 966 18410 967
rect 18494 910 18522 938
rect 18270 798 18298 826
rect 18270 630 18298 658
rect 18662 1750 18690 1778
rect 18606 742 18634 770
rect 18774 2169 18802 2170
rect 18774 2143 18775 2169
rect 18775 2143 18801 2169
rect 18801 2143 18802 2169
rect 18774 2142 18802 2143
rect 18774 1190 18802 1218
rect 18830 462 18858 490
rect 18998 4326 19026 4354
rect 19054 2758 19082 2786
rect 18998 2310 19026 2338
rect 18942 713 18970 714
rect 18942 687 18943 713
rect 18943 687 18969 713
rect 18969 687 18970 713
rect 18942 686 18970 687
rect 18718 350 18746 378
rect 19166 2646 19194 2674
rect 20230 5894 20258 5922
rect 19334 5054 19362 5082
rect 19502 5838 19530 5866
rect 19334 2897 19362 2898
rect 19334 2871 19335 2897
rect 19335 2871 19361 2897
rect 19361 2871 19362 2897
rect 19334 2870 19362 2871
rect 19222 2057 19250 2058
rect 19222 2031 19223 2057
rect 19223 2031 19249 2057
rect 19249 2031 19250 2057
rect 19222 2030 19250 2031
rect 19334 1974 19362 2002
rect 19166 1833 19194 1834
rect 19166 1807 19167 1833
rect 19167 1807 19193 1833
rect 19193 1807 19194 1833
rect 19166 1806 19194 1807
rect 19166 1078 19194 1106
rect 19166 686 19194 714
rect 19110 630 19138 658
rect 19110 182 19138 210
rect 19446 1694 19474 1722
rect 19446 742 19474 770
rect 20062 2926 20090 2954
rect 20062 2142 20090 2170
rect 19670 2030 19698 2058
rect 19558 1385 19586 1386
rect 19558 1359 19559 1385
rect 19559 1359 19585 1385
rect 19585 1359 19586 1385
rect 19558 1358 19586 1359
rect 20174 1470 20202 1498
rect 19726 1273 19754 1274
rect 19726 1247 19727 1273
rect 19727 1247 19753 1273
rect 19753 1247 19754 1273
rect 19726 1246 19754 1247
rect 19614 993 19642 994
rect 19614 967 19615 993
rect 19615 967 19641 993
rect 19641 967 19642 993
rect 19614 966 19642 967
rect 19614 798 19642 826
rect 19670 126 19698 154
rect 19838 742 19866 770
rect 19950 630 19978 658
rect 20286 3598 20314 3626
rect 20510 2982 20538 3010
rect 20342 2870 20370 2898
rect 20398 2702 20426 2730
rect 20342 1694 20370 1722
rect 20286 1470 20314 1498
rect 20342 1526 20370 1554
rect 20230 686 20258 714
rect 20902 5446 20930 5474
rect 20622 4942 20650 4970
rect 20622 3038 20650 3066
rect 20790 1806 20818 1834
rect 20902 1806 20930 1834
rect 20566 798 20594 826
rect 21462 6454 21490 6482
rect 21294 6145 21322 6146
rect 21294 6119 21295 6145
rect 21295 6119 21321 6145
rect 21321 6119 21322 6145
rect 21294 6118 21322 6119
rect 21126 5726 21154 5754
rect 21406 5950 21434 5978
rect 21126 5614 21154 5642
rect 21070 2478 21098 2506
rect 21294 3990 21322 4018
rect 21294 3289 21322 3290
rect 21294 3263 21295 3289
rect 21295 3263 21321 3289
rect 21321 3263 21322 3289
rect 21294 3262 21322 3263
rect 21126 2086 21154 2114
rect 21014 742 21042 770
rect 20342 686 20370 714
rect 20566 545 20594 546
rect 20566 519 20567 545
rect 20567 519 20593 545
rect 20593 519 20594 545
rect 20566 518 20594 519
rect 20958 545 20986 546
rect 20958 519 20959 545
rect 20959 519 20985 545
rect 20985 519 20986 545
rect 20958 518 20986 519
rect 20062 462 20090 490
rect 21854 6481 21882 6482
rect 21854 6455 21855 6481
rect 21855 6455 21881 6481
rect 21881 6455 21882 6481
rect 21854 6454 21882 6455
rect 21902 6285 21930 6286
rect 21902 6259 21903 6285
rect 21903 6259 21929 6285
rect 21929 6259 21930 6285
rect 21902 6258 21930 6259
rect 21954 6285 21982 6286
rect 21954 6259 21955 6285
rect 21955 6259 21981 6285
rect 21981 6259 21982 6285
rect 21954 6258 21982 6259
rect 22006 6285 22034 6286
rect 22006 6259 22007 6285
rect 22007 6259 22033 6285
rect 22033 6259 22034 6285
rect 22006 6258 22034 6259
rect 22358 6033 22386 6034
rect 22358 6007 22359 6033
rect 22359 6007 22385 6033
rect 22385 6007 22386 6033
rect 22358 6006 22386 6007
rect 22078 5977 22106 5978
rect 22078 5951 22079 5977
rect 22079 5951 22105 5977
rect 22105 5951 22106 5977
rect 22078 5950 22106 5951
rect 21686 5894 21714 5922
rect 21462 2310 21490 2338
rect 22232 5893 22260 5894
rect 22232 5867 22233 5893
rect 22233 5867 22259 5893
rect 22259 5867 22260 5893
rect 22232 5866 22260 5867
rect 22284 5893 22312 5894
rect 22284 5867 22285 5893
rect 22285 5867 22311 5893
rect 22311 5867 22312 5893
rect 22284 5866 22312 5867
rect 22336 5893 22364 5894
rect 22336 5867 22337 5893
rect 22337 5867 22363 5893
rect 22363 5867 22364 5893
rect 22336 5866 22364 5867
rect 22694 5809 22722 5810
rect 22694 5783 22695 5809
rect 22695 5783 22721 5809
rect 22721 5783 22722 5809
rect 22694 5782 22722 5783
rect 21902 5501 21930 5502
rect 21902 5475 21903 5501
rect 21903 5475 21929 5501
rect 21929 5475 21930 5501
rect 21902 5474 21930 5475
rect 21954 5501 21982 5502
rect 21954 5475 21955 5501
rect 21955 5475 21981 5501
rect 21981 5475 21982 5501
rect 21954 5474 21982 5475
rect 22006 5501 22034 5502
rect 22006 5475 22007 5501
rect 22007 5475 22033 5501
rect 22033 5475 22034 5501
rect 22006 5474 22034 5475
rect 22232 5109 22260 5110
rect 22232 5083 22233 5109
rect 22233 5083 22259 5109
rect 22259 5083 22260 5109
rect 22232 5082 22260 5083
rect 22284 5109 22312 5110
rect 22284 5083 22285 5109
rect 22285 5083 22311 5109
rect 22311 5083 22312 5109
rect 22284 5082 22312 5083
rect 22336 5109 22364 5110
rect 22336 5083 22337 5109
rect 22337 5083 22363 5109
rect 22363 5083 22364 5109
rect 22336 5082 22364 5083
rect 21902 4717 21930 4718
rect 21902 4691 21903 4717
rect 21903 4691 21929 4717
rect 21929 4691 21930 4717
rect 21902 4690 21930 4691
rect 21954 4717 21982 4718
rect 21954 4691 21955 4717
rect 21955 4691 21981 4717
rect 21981 4691 21982 4717
rect 21954 4690 21982 4691
rect 22006 4717 22034 4718
rect 22006 4691 22007 4717
rect 22007 4691 22033 4717
rect 22033 4691 22034 4717
rect 22006 4690 22034 4691
rect 22750 4577 22778 4578
rect 22750 4551 22751 4577
rect 22751 4551 22777 4577
rect 22777 4551 22778 4577
rect 22750 4550 22778 4551
rect 22470 4521 22498 4522
rect 22470 4495 22471 4521
rect 22471 4495 22497 4521
rect 22497 4495 22498 4521
rect 22470 4494 22498 4495
rect 22232 4325 22260 4326
rect 22232 4299 22233 4325
rect 22233 4299 22259 4325
rect 22259 4299 22260 4325
rect 22232 4298 22260 4299
rect 22284 4325 22312 4326
rect 22284 4299 22285 4325
rect 22285 4299 22311 4325
rect 22311 4299 22312 4325
rect 22284 4298 22312 4299
rect 22336 4325 22364 4326
rect 22336 4299 22337 4325
rect 22337 4299 22363 4325
rect 22363 4299 22364 4325
rect 22336 4298 22364 4299
rect 21902 3933 21930 3934
rect 21902 3907 21903 3933
rect 21903 3907 21929 3933
rect 21929 3907 21930 3933
rect 21902 3906 21930 3907
rect 21954 3933 21982 3934
rect 21954 3907 21955 3933
rect 21955 3907 21981 3933
rect 21981 3907 21982 3933
rect 21954 3906 21982 3907
rect 22006 3933 22034 3934
rect 22006 3907 22007 3933
rect 22007 3907 22033 3933
rect 22033 3907 22034 3933
rect 22006 3906 22034 3907
rect 22232 3541 22260 3542
rect 22232 3515 22233 3541
rect 22233 3515 22259 3541
rect 22259 3515 22260 3541
rect 22232 3514 22260 3515
rect 22284 3541 22312 3542
rect 22284 3515 22285 3541
rect 22285 3515 22311 3541
rect 22311 3515 22312 3541
rect 22284 3514 22312 3515
rect 22336 3541 22364 3542
rect 22336 3515 22337 3541
rect 22337 3515 22363 3541
rect 22363 3515 22364 3541
rect 22336 3514 22364 3515
rect 21686 3374 21714 3402
rect 22134 3345 22162 3346
rect 22134 3319 22135 3345
rect 22135 3319 22161 3345
rect 22161 3319 22162 3345
rect 22134 3318 22162 3319
rect 21902 3149 21930 3150
rect 21902 3123 21903 3149
rect 21903 3123 21929 3149
rect 21929 3123 21930 3149
rect 21902 3122 21930 3123
rect 21954 3149 21982 3150
rect 21954 3123 21955 3149
rect 21955 3123 21981 3149
rect 21981 3123 21982 3149
rect 21954 3122 21982 3123
rect 22006 3149 22034 3150
rect 22006 3123 22007 3149
rect 22007 3123 22033 3149
rect 22033 3123 22034 3149
rect 22006 3122 22034 3123
rect 22358 2926 22386 2954
rect 22232 2757 22260 2758
rect 22232 2731 22233 2757
rect 22233 2731 22259 2757
rect 22259 2731 22260 2757
rect 22232 2730 22260 2731
rect 22284 2757 22312 2758
rect 22284 2731 22285 2757
rect 22285 2731 22311 2757
rect 22311 2731 22312 2757
rect 22284 2730 22312 2731
rect 22336 2757 22364 2758
rect 22336 2731 22337 2757
rect 22337 2731 22363 2757
rect 22363 2731 22364 2757
rect 22336 2730 22364 2731
rect 21902 2365 21930 2366
rect 21902 2339 21903 2365
rect 21903 2339 21929 2365
rect 21929 2339 21930 2365
rect 21902 2338 21930 2339
rect 21954 2365 21982 2366
rect 21954 2339 21955 2365
rect 21955 2339 21981 2365
rect 21981 2339 21982 2365
rect 21954 2338 21982 2339
rect 22006 2365 22034 2366
rect 22006 2339 22007 2365
rect 22007 2339 22033 2365
rect 22033 2339 22034 2365
rect 22006 2338 22034 2339
rect 22190 2057 22218 2058
rect 22190 2031 22191 2057
rect 22191 2031 22217 2057
rect 22217 2031 22218 2057
rect 22190 2030 22218 2031
rect 22232 1973 22260 1974
rect 22232 1947 22233 1973
rect 22233 1947 22259 1973
rect 22259 1947 22260 1973
rect 22232 1946 22260 1947
rect 22284 1973 22312 1974
rect 22284 1947 22285 1973
rect 22285 1947 22311 1973
rect 22311 1947 22312 1973
rect 22284 1946 22312 1947
rect 22336 1973 22364 1974
rect 22336 1947 22337 1973
rect 22337 1947 22363 1973
rect 22363 1947 22364 1973
rect 22336 1946 22364 1947
rect 22470 1750 22498 1778
rect 21902 1581 21930 1582
rect 21902 1555 21903 1581
rect 21903 1555 21929 1581
rect 21929 1555 21930 1581
rect 21902 1554 21930 1555
rect 21954 1581 21982 1582
rect 21954 1555 21955 1581
rect 21955 1555 21981 1581
rect 21981 1555 21982 1581
rect 21954 1554 21982 1555
rect 22006 1581 22034 1582
rect 22006 1555 22007 1581
rect 22007 1555 22033 1581
rect 22033 1555 22034 1581
rect 22006 1554 22034 1555
rect 21518 1358 21546 1386
rect 22750 1246 22778 1274
rect 22232 1189 22260 1190
rect 22232 1163 22233 1189
rect 22233 1163 22259 1189
rect 22259 1163 22260 1189
rect 22232 1162 22260 1163
rect 22284 1189 22312 1190
rect 22284 1163 22285 1189
rect 22285 1163 22311 1189
rect 22311 1163 22312 1189
rect 22284 1162 22312 1163
rect 22336 1189 22364 1190
rect 22336 1163 22337 1189
rect 22337 1163 22363 1189
rect 22363 1163 22364 1189
rect 22336 1162 22364 1163
rect 22470 1049 22498 1050
rect 22470 1023 22471 1049
rect 22471 1023 22497 1049
rect 22497 1023 22498 1049
rect 22470 1022 22498 1023
rect 21902 797 21930 798
rect 21902 771 21903 797
rect 21903 771 21929 797
rect 21929 771 21930 797
rect 21902 770 21930 771
rect 21954 797 21982 798
rect 21954 771 21955 797
rect 21955 771 21981 797
rect 21981 771 21982 797
rect 21954 770 21982 771
rect 22006 797 22034 798
rect 22006 771 22007 797
rect 22007 771 22033 797
rect 22033 771 22034 797
rect 22006 770 22034 771
rect 23086 6481 23114 6482
rect 23086 6455 23087 6481
rect 23087 6455 23113 6481
rect 23113 6455 23114 6481
rect 23086 6454 23114 6455
rect 23366 6118 23394 6146
rect 23310 6089 23338 6090
rect 23310 6063 23311 6089
rect 23311 6063 23337 6089
rect 23337 6063 23338 6089
rect 23310 6062 23338 6063
rect 23646 6593 23674 6594
rect 23646 6567 23647 6593
rect 23647 6567 23673 6593
rect 23673 6567 23674 6593
rect 23646 6566 23674 6567
rect 25214 6734 25242 6762
rect 24206 6566 24234 6594
rect 24598 6593 24626 6594
rect 24598 6567 24599 6593
rect 24599 6567 24625 6593
rect 24625 6567 24626 6593
rect 24598 6566 24626 6567
rect 24374 6481 24402 6482
rect 24374 6455 24375 6481
rect 24375 6455 24401 6481
rect 24401 6455 24402 6481
rect 24374 6454 24402 6455
rect 24038 6201 24066 6202
rect 24038 6175 24039 6201
rect 24039 6175 24065 6201
rect 24065 6175 24066 6201
rect 24038 6174 24066 6175
rect 23534 6033 23562 6034
rect 23534 6007 23535 6033
rect 23535 6007 23561 6033
rect 23561 6007 23562 6033
rect 23534 6006 23562 6007
rect 23478 5838 23506 5866
rect 23142 5753 23170 5754
rect 23142 5727 23143 5753
rect 23143 5727 23169 5753
rect 23169 5727 23170 5753
rect 23142 5726 23170 5727
rect 23534 5753 23562 5754
rect 23534 5727 23535 5753
rect 23535 5727 23561 5753
rect 23561 5727 23562 5753
rect 23534 5726 23562 5727
rect 24038 5446 24066 5474
rect 24822 5894 24850 5922
rect 24934 5641 24962 5642
rect 24934 5615 24935 5641
rect 24935 5615 24961 5641
rect 24961 5615 24962 5641
rect 24934 5614 24962 5615
rect 23086 5305 23114 5306
rect 23086 5279 23087 5305
rect 23087 5279 23113 5305
rect 23113 5279 23114 5305
rect 23086 5278 23114 5279
rect 24374 5222 24402 5250
rect 22974 5054 23002 5082
rect 24374 5054 24402 5082
rect 23142 4998 23170 5026
rect 24150 4998 24178 5026
rect 23758 4913 23786 4914
rect 23758 4887 23759 4913
rect 23759 4887 23785 4913
rect 23785 4887 23786 4913
rect 23758 4886 23786 4887
rect 23534 4774 23562 4802
rect 24206 4494 24234 4522
rect 23870 4465 23898 4466
rect 23870 4439 23871 4465
rect 23871 4439 23897 4465
rect 23897 4439 23898 4465
rect 23870 4438 23898 4439
rect 23254 4185 23282 4186
rect 23254 4159 23255 4185
rect 23255 4159 23281 4185
rect 23281 4159 23282 4185
rect 23254 4158 23282 4159
rect 23478 4073 23506 4074
rect 23478 4047 23479 4073
rect 23479 4047 23505 4073
rect 23505 4047 23506 4073
rect 23478 4046 23506 4047
rect 24150 3793 24178 3794
rect 24150 3767 24151 3793
rect 24151 3767 24177 3793
rect 24177 3767 24178 3793
rect 24150 3766 24178 3767
rect 23870 3681 23898 3682
rect 23870 3655 23871 3681
rect 23871 3655 23897 3681
rect 23897 3655 23898 3681
rect 23870 3654 23898 3655
rect 24486 5390 24514 5418
rect 24822 5166 24850 5194
rect 24430 4998 24458 5026
rect 24430 4913 24458 4914
rect 24430 4887 24431 4913
rect 24431 4887 24457 4913
rect 24457 4887 24458 4913
rect 24430 4886 24458 4887
rect 24934 4857 24962 4858
rect 24934 4831 24935 4857
rect 24935 4831 24961 4857
rect 24961 4831 24962 4857
rect 24934 4830 24962 4831
rect 24822 4633 24850 4634
rect 24822 4607 24823 4633
rect 24823 4607 24849 4633
rect 24849 4607 24850 4633
rect 24822 4606 24850 4607
rect 25382 6510 25410 6538
rect 25270 5838 25298 5866
rect 25326 6286 25354 6314
rect 25214 5726 25242 5754
rect 25214 4550 25242 4578
rect 25102 4382 25130 4410
rect 25102 4214 25130 4242
rect 24374 3737 24402 3738
rect 24374 3711 24375 3737
rect 24375 3711 24401 3737
rect 24401 3711 24402 3737
rect 24374 3710 24402 3711
rect 24598 4129 24626 4130
rect 24598 4103 24599 4129
rect 24599 4103 24625 4129
rect 24625 4103 24626 4129
rect 24598 4102 24626 4103
rect 24766 3990 24794 4018
rect 24430 3598 24458 3626
rect 25214 4129 25242 4130
rect 25214 4103 25215 4129
rect 25215 4103 25241 4129
rect 25241 4103 25242 4129
rect 25214 4102 25242 4103
rect 25158 4046 25186 4074
rect 25438 6174 25466 6202
rect 25494 6062 25522 6090
rect 25382 5446 25410 5474
rect 25606 5390 25634 5418
rect 25662 6062 25690 6090
rect 25718 4942 25746 4970
rect 25662 4830 25690 4858
rect 25494 4718 25522 4746
rect 25326 4606 25354 4634
rect 25718 4494 25746 4522
rect 25494 4270 25522 4298
rect 25606 4046 25634 4074
rect 25718 3822 25746 3850
rect 25270 3766 25298 3794
rect 24822 3374 24850 3402
rect 25718 3598 25746 3626
rect 24430 3345 24458 3346
rect 24430 3319 24431 3345
rect 24431 3319 24457 3345
rect 24457 3319 24458 3345
rect 24430 3318 24458 3319
rect 25214 3038 25242 3066
rect 25606 3150 25634 3178
rect 24878 2926 24906 2954
rect 23590 2897 23618 2898
rect 23590 2871 23591 2897
rect 23591 2871 23617 2897
rect 23617 2871 23618 2897
rect 23590 2870 23618 2871
rect 23422 2534 23450 2562
rect 23814 2113 23842 2114
rect 23814 2087 23815 2113
rect 23815 2087 23841 2113
rect 23841 2087 23842 2113
rect 23814 2086 23842 2087
rect 23534 1806 23562 1834
rect 23534 1470 23562 1498
rect 23086 1414 23114 1442
rect 23366 1329 23394 1330
rect 23366 1303 23367 1329
rect 23367 1303 23393 1329
rect 23393 1303 23394 1329
rect 23366 1302 23394 1303
rect 23534 1078 23562 1106
rect 22806 630 22834 658
rect 23758 993 23786 994
rect 23758 967 23759 993
rect 23759 967 23785 993
rect 23785 967 23786 993
rect 23758 966 23786 967
rect 24486 2590 24514 2618
rect 24374 2534 24402 2562
rect 24094 2225 24122 2226
rect 24094 2199 24095 2225
rect 24095 2199 24121 2225
rect 24121 2199 24122 2225
rect 24094 2198 24122 2199
rect 25102 2814 25130 2842
rect 24934 2646 24962 2674
rect 25606 2702 25634 2730
rect 25214 2617 25242 2618
rect 25214 2591 25215 2617
rect 25215 2591 25241 2617
rect 25241 2591 25242 2617
rect 25214 2590 25242 2591
rect 24822 2561 24850 2562
rect 24822 2535 24823 2561
rect 24823 2535 24849 2561
rect 24849 2535 24850 2561
rect 24822 2534 24850 2535
rect 25550 2534 25578 2562
rect 24654 2422 24682 2450
rect 25438 2478 25466 2506
rect 25550 2254 25578 2282
rect 24430 2198 24458 2226
rect 24710 1806 24738 1834
rect 25214 1862 25242 1890
rect 24038 1441 24066 1442
rect 24038 1415 24039 1441
rect 24039 1415 24065 1441
rect 24065 1415 24066 1441
rect 24038 1414 24066 1415
rect 24318 686 24346 714
rect 24374 1302 24402 1330
rect 23870 518 23898 546
rect 21406 462 21434 490
rect 25102 1750 25130 1778
rect 24934 1721 24962 1722
rect 24934 1695 24935 1721
rect 24935 1695 24961 1721
rect 24961 1695 24962 1721
rect 24934 1694 24962 1695
rect 24430 1246 24458 1274
rect 24486 1638 24514 1666
rect 25494 1694 25522 1722
rect 25326 1414 25354 1442
rect 24710 1329 24738 1330
rect 24710 1303 24711 1329
rect 24711 1303 24737 1329
rect 24737 1303 24738 1329
rect 24710 1302 24738 1303
rect 25214 993 25242 994
rect 25214 967 25215 993
rect 25215 967 25241 993
rect 25241 967 25242 993
rect 25214 966 25242 967
rect 24934 937 24962 938
rect 24934 911 24935 937
rect 24935 911 24961 937
rect 24961 911 24962 937
rect 24934 910 24962 911
rect 24878 713 24906 714
rect 24878 687 24879 713
rect 24879 687 24905 713
rect 24905 687 24906 713
rect 24878 686 24906 687
rect 25270 601 25298 602
rect 25270 575 25271 601
rect 25271 575 25297 601
rect 25297 575 25298 601
rect 25270 574 25298 575
rect 24094 462 24122 490
rect 22232 405 22260 406
rect 22232 379 22233 405
rect 22233 379 22259 405
rect 22259 379 22260 405
rect 22232 378 22260 379
rect 22284 405 22312 406
rect 22284 379 22285 405
rect 22285 379 22311 405
rect 22311 379 22312 405
rect 22284 378 22312 379
rect 22336 405 22364 406
rect 22336 379 22337 405
rect 22337 379 22363 405
rect 22363 379 22364 405
rect 22336 378 22364 379
rect 25550 1582 25578 1610
rect 25494 1358 25522 1386
rect 25326 238 25354 266
rect 25438 1302 25466 1330
rect 4942 14 4970 42
rect 25718 2030 25746 2058
rect 25718 1134 25746 1162
rect 25438 14 25466 42
<< metal3 >>
rect 3257 7014 3262 7042
rect 3290 7014 3486 7042
rect 3514 7014 3519 7042
rect 4489 7014 4494 7042
rect 4522 7014 4718 7042
rect 4746 7014 4751 7042
rect 6953 7014 6958 7042
rect 6986 7014 7182 7042
rect 7210 7014 7215 7042
rect 8185 7014 8190 7042
rect 8218 7014 8414 7042
rect 8442 7014 8447 7042
rect 10649 7014 10654 7042
rect 10682 7014 10878 7042
rect 10906 7014 10911 7042
rect 11881 7014 11886 7042
rect 11914 7014 12110 7042
rect 12138 7014 12143 7042
rect 14345 7014 14350 7042
rect 14378 7014 14574 7042
rect 14602 7014 14607 7042
rect 15577 7014 15582 7042
rect 15610 7014 15862 7042
rect 15890 7014 15895 7042
rect 18041 7014 18046 7042
rect 18074 7014 18270 7042
rect 18298 7014 18303 7042
rect 20505 7014 20510 7042
rect 20538 7014 20678 7042
rect 20706 7014 20711 7042
rect 0 6986 56 7000
rect 26320 6986 26376 7000
rect 0 6958 23478 6986
rect 23506 6958 23511 6986
rect 25046 6958 26376 6986
rect 0 6944 56 6958
rect 25046 6930 25074 6958
rect 26320 6944 26376 6958
rect 23025 6902 23030 6930
rect 23058 6902 25074 6930
rect 9193 6846 9198 6874
rect 9226 6846 14742 6874
rect 14770 6846 14775 6874
rect 0 6762 56 6776
rect 26320 6762 26376 6776
rect 0 6734 1134 6762
rect 1162 6734 1167 6762
rect 3033 6734 3038 6762
rect 3066 6734 15246 6762
rect 15274 6734 15279 6762
rect 25209 6734 25214 6762
rect 25242 6734 26376 6762
rect 0 6720 56 6734
rect 26320 6720 26376 6734
rect 2227 6650 2232 6678
rect 2260 6650 2284 6678
rect 2312 6650 2336 6678
rect 2364 6650 2369 6678
rect 12227 6650 12232 6678
rect 12260 6650 12284 6678
rect 12312 6650 12336 6678
rect 12364 6650 12369 6678
rect 22227 6650 22232 6678
rect 22260 6650 22284 6678
rect 22312 6650 22336 6678
rect 22364 6650 22369 6678
rect 8857 6566 8862 6594
rect 8890 6566 14126 6594
rect 14154 6566 14159 6594
rect 19273 6566 19278 6594
rect 19306 6566 19838 6594
rect 19866 6566 19871 6594
rect 21849 6566 21854 6594
rect 21882 6566 22134 6594
rect 22162 6566 22167 6594
rect 22969 6566 22974 6594
rect 23002 6566 23646 6594
rect 23674 6566 23679 6594
rect 24201 6566 24206 6594
rect 24234 6566 24598 6594
rect 24626 6566 24631 6594
rect 0 6538 56 6552
rect 26320 6538 26376 6552
rect 0 6510 1638 6538
rect 1666 6510 1671 6538
rect 2025 6510 2030 6538
rect 2058 6510 2646 6538
rect 2674 6510 2679 6538
rect 5721 6510 5726 6538
rect 5754 6510 6454 6538
rect 6482 6510 6487 6538
rect 6734 6510 21126 6538
rect 21154 6510 21159 6538
rect 25377 6510 25382 6538
rect 25410 6510 26376 6538
rect 0 6496 56 6510
rect 1073 6454 1078 6482
rect 1106 6454 2478 6482
rect 2506 6454 2511 6482
rect 6734 6426 6762 6510
rect 26320 6496 26376 6510
rect 6841 6454 6846 6482
rect 6874 6454 8806 6482
rect 8834 6454 8839 6482
rect 9753 6454 9758 6482
rect 9786 6454 12614 6482
rect 12642 6454 12647 6482
rect 21457 6454 21462 6482
rect 21490 6454 21854 6482
rect 21882 6454 21887 6482
rect 23081 6454 23086 6482
rect 23114 6454 24374 6482
rect 24402 6454 24407 6482
rect 1353 6398 1358 6426
rect 1386 6398 6762 6426
rect 8913 6398 8918 6426
rect 8946 6398 16590 6426
rect 16618 6398 16623 6426
rect 11489 6342 11494 6370
rect 11522 6342 13790 6370
rect 13818 6342 13823 6370
rect 0 6314 56 6328
rect 26320 6314 26376 6328
rect 0 6286 574 6314
rect 602 6286 607 6314
rect 12110 6286 17430 6314
rect 17458 6286 17463 6314
rect 25321 6286 25326 6314
rect 25354 6286 26376 6314
rect 0 6272 56 6286
rect 1897 6258 1902 6286
rect 1930 6258 1954 6286
rect 1982 6258 2006 6286
rect 2034 6258 2039 6286
rect 11897 6258 11902 6286
rect 11930 6258 11954 6286
rect 11982 6258 12006 6286
rect 12034 6258 12039 6286
rect 12110 6202 12138 6286
rect 21897 6258 21902 6286
rect 21930 6258 21954 6286
rect 21982 6258 22006 6286
rect 22034 6258 22039 6286
rect 26320 6272 26376 6286
rect 11545 6174 11550 6202
rect 11578 6174 12138 6202
rect 13337 6174 13342 6202
rect 13370 6174 18494 6202
rect 18522 6174 18527 6202
rect 24033 6174 24038 6202
rect 24066 6174 25438 6202
rect 25466 6174 25471 6202
rect 6449 6118 6454 6146
rect 6482 6118 16282 6146
rect 16361 6118 16366 6146
rect 16394 6118 17038 6146
rect 17066 6118 17071 6146
rect 18825 6118 18830 6146
rect 18858 6118 19558 6146
rect 19586 6118 19591 6146
rect 21289 6118 21294 6146
rect 21322 6118 23366 6146
rect 23394 6118 23399 6146
rect 0 6090 56 6104
rect 16254 6090 16282 6118
rect 26320 6090 26376 6104
rect 0 6062 350 6090
rect 378 6062 383 6090
rect 10929 6062 10934 6090
rect 10962 6062 15918 6090
rect 15946 6062 15951 6090
rect 16254 6062 19334 6090
rect 19362 6062 19367 6090
rect 23305 6062 23310 6090
rect 23338 6062 25494 6090
rect 25522 6062 25527 6090
rect 25657 6062 25662 6090
rect 25690 6062 26376 6090
rect 0 6048 56 6062
rect 26320 6048 26376 6062
rect 10145 6006 10150 6034
rect 10178 6006 14798 6034
rect 14826 6006 14831 6034
rect 16865 6006 16870 6034
rect 16898 6006 18662 6034
rect 18690 6006 18695 6034
rect 22353 6006 22358 6034
rect 22386 6006 23534 6034
rect 23562 6006 23567 6034
rect 9081 5950 9086 5978
rect 9114 5950 12586 5978
rect 12665 5950 12670 5978
rect 12698 5950 16310 5978
rect 16338 5950 16343 5978
rect 17313 5950 17318 5978
rect 17346 5950 18354 5978
rect 19217 5950 19222 5978
rect 19250 5950 20370 5978
rect 21401 5950 21406 5978
rect 21434 5950 22078 5978
rect 22106 5950 22111 5978
rect 3537 5894 3542 5922
rect 3570 5894 7126 5922
rect 7154 5894 7159 5922
rect 0 5866 56 5880
rect 2227 5866 2232 5894
rect 2260 5866 2284 5894
rect 2312 5866 2336 5894
rect 2364 5866 2369 5894
rect 12227 5866 12232 5894
rect 12260 5866 12284 5894
rect 12312 5866 12336 5894
rect 12364 5866 12369 5894
rect 12558 5866 12586 5950
rect 18326 5922 18354 5950
rect 20342 5922 20370 5950
rect 13342 5894 14854 5922
rect 14882 5894 14887 5922
rect 15974 5894 17654 5922
rect 17682 5894 17687 5922
rect 18326 5894 20230 5922
rect 20258 5894 20263 5922
rect 20342 5894 21686 5922
rect 21714 5894 21719 5922
rect 24817 5894 24822 5922
rect 24850 5894 25522 5922
rect 13342 5866 13370 5894
rect 15974 5866 16002 5894
rect 22227 5866 22232 5894
rect 22260 5866 22284 5894
rect 22312 5866 22336 5894
rect 22364 5866 22369 5894
rect 25494 5866 25522 5894
rect 26320 5866 26376 5880
rect 0 5838 490 5866
rect 7793 5838 7798 5866
rect 7826 5838 11494 5866
rect 11522 5838 11527 5866
rect 12558 5838 13370 5866
rect 13897 5838 13902 5866
rect 13930 5838 16002 5866
rect 19049 5838 19054 5866
rect 19082 5838 19502 5866
rect 19530 5838 19535 5866
rect 23473 5838 23478 5866
rect 23506 5838 25270 5866
rect 25298 5838 25303 5866
rect 25494 5838 26376 5866
rect 0 5824 56 5838
rect 462 5754 490 5838
rect 26320 5824 26376 5838
rect 569 5782 574 5810
rect 602 5782 8862 5810
rect 8890 5782 8895 5810
rect 9025 5782 9030 5810
rect 9058 5782 15134 5810
rect 15162 5782 15167 5810
rect 15913 5782 15918 5810
rect 15946 5782 19222 5810
rect 19250 5782 19255 5810
rect 19306 5782 22694 5810
rect 22722 5782 22727 5810
rect 462 5726 14910 5754
rect 14938 5726 14943 5754
rect 19306 5698 19334 5782
rect 21121 5726 21126 5754
rect 21154 5726 23142 5754
rect 23170 5726 23175 5754
rect 23529 5726 23534 5754
rect 23562 5726 25214 5754
rect 25242 5726 25247 5754
rect 12721 5670 12726 5698
rect 12754 5670 14042 5698
rect 14121 5670 14126 5698
rect 14154 5670 19334 5698
rect 0 5642 56 5656
rect 0 5614 3486 5642
rect 3514 5614 3519 5642
rect 5217 5614 5222 5642
rect 5250 5614 7574 5642
rect 7602 5614 7607 5642
rect 9529 5614 9534 5642
rect 9562 5614 12110 5642
rect 12138 5614 12143 5642
rect 12553 5614 12558 5642
rect 12586 5614 13482 5642
rect 0 5600 56 5614
rect 13454 5586 13482 5614
rect 14014 5586 14042 5670
rect 26320 5642 26376 5656
rect 14793 5614 14798 5642
rect 14826 5614 16142 5642
rect 16170 5614 16175 5642
rect 17649 5614 17654 5642
rect 17682 5614 21126 5642
rect 21154 5614 21159 5642
rect 24929 5614 24934 5642
rect 24962 5614 26376 5642
rect 26320 5600 26376 5614
rect 3985 5558 3990 5586
rect 4018 5558 9030 5586
rect 9058 5558 9063 5586
rect 10257 5558 10262 5586
rect 10290 5558 13342 5586
rect 13370 5558 13375 5586
rect 13454 5558 13902 5586
rect 13930 5558 13935 5586
rect 14014 5558 16814 5586
rect 16842 5558 16847 5586
rect 3761 5502 3766 5530
rect 3794 5502 7462 5530
rect 7490 5502 7495 5530
rect 12105 5502 12110 5530
rect 12138 5502 15190 5530
rect 15218 5502 15223 5530
rect 1897 5474 1902 5502
rect 1930 5474 1954 5502
rect 1982 5474 2006 5502
rect 2034 5474 2039 5502
rect 11897 5474 11902 5502
rect 11930 5474 11954 5502
rect 11982 5474 12006 5502
rect 12034 5474 12039 5502
rect 21897 5474 21902 5502
rect 21930 5474 21954 5502
rect 21982 5474 22006 5502
rect 22034 5474 22039 5502
rect 6953 5446 6958 5474
rect 6986 5446 7574 5474
rect 14009 5446 14014 5474
rect 14042 5446 20902 5474
rect 20930 5446 20935 5474
rect 24033 5446 24038 5474
rect 24066 5446 25382 5474
rect 25410 5446 25415 5474
rect 0 5418 56 5432
rect 7546 5418 7574 5446
rect 26320 5418 26376 5432
rect 0 5390 2422 5418
rect 2450 5390 2455 5418
rect 7546 5390 15022 5418
rect 15050 5390 15055 5418
rect 15969 5390 15974 5418
rect 16002 5390 24486 5418
rect 24514 5390 24519 5418
rect 25601 5390 25606 5418
rect 25634 5390 26376 5418
rect 0 5376 56 5390
rect 26320 5376 26376 5390
rect 10705 5334 10710 5362
rect 10738 5334 12726 5362
rect 12754 5334 12759 5362
rect 12833 5334 12838 5362
rect 12866 5334 15078 5362
rect 15106 5334 15111 5362
rect 17369 5334 17374 5362
rect 17402 5334 18718 5362
rect 18746 5334 18751 5362
rect 11041 5278 11046 5306
rect 11074 5278 12502 5306
rect 12530 5278 12535 5306
rect 12609 5278 12614 5306
rect 12642 5278 17654 5306
rect 17682 5278 17687 5306
rect 18489 5278 18494 5306
rect 18522 5278 23086 5306
rect 23114 5278 23119 5306
rect 2086 5222 5054 5250
rect 5082 5222 5087 5250
rect 5273 5222 5278 5250
rect 5306 5222 24374 5250
rect 24402 5222 24407 5250
rect 0 5194 56 5208
rect 2086 5194 2114 5222
rect 26320 5194 26376 5208
rect 0 5166 2114 5194
rect 2473 5166 2478 5194
rect 2506 5166 4270 5194
rect 4298 5166 4303 5194
rect 8353 5166 8358 5194
rect 8386 5166 12558 5194
rect 12586 5166 12591 5194
rect 13617 5166 13622 5194
rect 13650 5166 18942 5194
rect 18970 5166 18975 5194
rect 24817 5166 24822 5194
rect 24850 5166 26376 5194
rect 0 5152 56 5166
rect 26320 5152 26376 5166
rect 4321 5110 4326 5138
rect 4354 5110 11718 5138
rect 11746 5110 11751 5138
rect 12441 5110 12446 5138
rect 12474 5110 14238 5138
rect 14266 5110 14271 5138
rect 14345 5110 14350 5138
rect 14378 5110 18102 5138
rect 18130 5110 18135 5138
rect 2227 5082 2232 5110
rect 2260 5082 2284 5110
rect 2312 5082 2336 5110
rect 2364 5082 2369 5110
rect 12227 5082 12232 5110
rect 12260 5082 12284 5110
rect 12312 5082 12336 5110
rect 12364 5082 12369 5110
rect 22227 5082 22232 5110
rect 22260 5082 22284 5110
rect 22312 5082 22336 5110
rect 22364 5082 22369 5110
rect 7546 5054 10486 5082
rect 10514 5054 10519 5082
rect 12446 5054 14770 5082
rect 15521 5054 15526 5082
rect 15554 5054 16702 5082
rect 16730 5054 16735 5082
rect 19329 5054 19334 5082
rect 19362 5054 21854 5082
rect 22969 5054 22974 5082
rect 23002 5054 24374 5082
rect 24402 5054 24407 5082
rect 7546 5026 7574 5054
rect 12446 5026 12474 5054
rect 1633 4998 1638 5026
rect 1666 4998 7574 5026
rect 10089 4998 10094 5026
rect 10122 4998 12474 5026
rect 14742 5026 14770 5054
rect 21826 5026 21854 5054
rect 14742 4998 16086 5026
rect 16114 4998 16119 5026
rect 21826 4998 23142 5026
rect 23170 4998 23175 5026
rect 24145 4998 24150 5026
rect 24178 4998 24430 5026
rect 24458 4998 24463 5026
rect 0 4970 56 4984
rect 26320 4970 26376 4984
rect 0 4942 2758 4970
rect 2786 4942 2791 4970
rect 2865 4942 2870 4970
rect 2898 4942 3542 4970
rect 3570 4942 3575 4970
rect 4377 4942 4382 4970
rect 4410 4942 6454 4970
rect 6482 4942 6487 4970
rect 7121 4942 7126 4970
rect 7154 4942 10066 4970
rect 11433 4942 11438 4970
rect 11466 4942 14350 4970
rect 14378 4942 14383 4970
rect 14849 4942 14854 4970
rect 14882 4942 16590 4970
rect 16618 4942 16623 4970
rect 19306 4942 20622 4970
rect 20650 4942 20655 4970
rect 25713 4942 25718 4970
rect 25746 4942 26376 4970
rect 0 4928 56 4942
rect 10038 4914 10066 4942
rect 19306 4914 19334 4942
rect 26320 4928 26376 4942
rect 2697 4886 2702 4914
rect 2730 4886 8358 4914
rect 8386 4886 8391 4914
rect 10038 4886 19334 4914
rect 23753 4886 23758 4914
rect 23786 4886 24430 4914
rect 24458 4886 24463 4914
rect 345 4830 350 4858
rect 378 4830 3374 4858
rect 3402 4830 3407 4858
rect 10481 4830 10486 4858
rect 10514 4830 13342 4858
rect 13370 4830 13375 4858
rect 13449 4830 13454 4858
rect 13482 4830 16198 4858
rect 16226 4830 16231 4858
rect 24929 4830 24934 4858
rect 24962 4830 25662 4858
rect 25690 4830 25695 4858
rect 2921 4774 2926 4802
rect 2954 4774 6958 4802
rect 6986 4774 6991 4802
rect 7681 4774 7686 4802
rect 7714 4774 12474 4802
rect 12553 4774 12558 4802
rect 12586 4774 14126 4802
rect 14154 4774 14159 4802
rect 14233 4774 14238 4802
rect 14266 4774 23534 4802
rect 23562 4774 23567 4802
rect 0 4746 56 4760
rect 12446 4746 12474 4774
rect 26320 4746 26376 4760
rect 0 4718 1834 4746
rect 12446 4718 13286 4746
rect 13314 4718 13319 4746
rect 13393 4718 13398 4746
rect 13426 4718 14686 4746
rect 14714 4718 14719 4746
rect 25489 4718 25494 4746
rect 25522 4718 26376 4746
rect 0 4704 56 4718
rect 1806 4634 1834 4718
rect 1897 4690 1902 4718
rect 1930 4690 1954 4718
rect 1982 4690 2006 4718
rect 2034 4690 2039 4718
rect 11897 4690 11902 4718
rect 11930 4690 11954 4718
rect 11982 4690 12006 4718
rect 12034 4690 12039 4718
rect 21897 4690 21902 4718
rect 21930 4690 21954 4718
rect 21982 4690 22006 4718
rect 22034 4690 22039 4718
rect 26320 4704 26376 4718
rect 6169 4662 6174 4690
rect 6202 4662 10934 4690
rect 10962 4662 10967 4690
rect 12110 4662 14350 4690
rect 14378 4662 14383 4690
rect 12110 4634 12138 4662
rect 1806 4606 5278 4634
rect 5306 4606 5311 4634
rect 8073 4606 8078 4634
rect 8106 4606 12138 4634
rect 12721 4606 12726 4634
rect 12754 4606 16646 4634
rect 16674 4606 16679 4634
rect 24817 4606 24822 4634
rect 24850 4606 25326 4634
rect 25354 4606 25359 4634
rect 9305 4550 9310 4578
rect 9338 4550 12446 4578
rect 12474 4550 12479 4578
rect 13426 4550 15470 4578
rect 15498 4550 15503 4578
rect 16025 4550 16030 4578
rect 16058 4550 22666 4578
rect 22745 4550 22750 4578
rect 22778 4550 25214 4578
rect 25242 4550 25247 4578
rect 0 4522 56 4536
rect 0 4494 3038 4522
rect 3066 4494 3071 4522
rect 10929 4494 10934 4522
rect 10962 4494 12670 4522
rect 12698 4494 12703 4522
rect 0 4480 56 4494
rect 13426 4466 13454 4550
rect 22638 4522 22666 4550
rect 26320 4522 26376 4536
rect 14121 4494 14126 4522
rect 14154 4494 14966 4522
rect 14994 4494 14999 4522
rect 15073 4494 15078 4522
rect 15106 4494 22470 4522
rect 22498 4494 22503 4522
rect 22638 4494 24206 4522
rect 24234 4494 24239 4522
rect 25713 4494 25718 4522
rect 25746 4494 26376 4522
rect 26320 4480 26376 4494
rect 8297 4438 8302 4466
rect 8330 4438 10150 4466
rect 10178 4438 10183 4466
rect 11601 4438 11606 4466
rect 11634 4438 13454 4466
rect 14905 4438 14910 4466
rect 14938 4438 23870 4466
rect 23898 4438 23903 4466
rect 7546 4382 25102 4410
rect 25130 4382 25135 4410
rect 7546 4354 7574 4382
rect 5553 4326 5558 4354
rect 5586 4326 7574 4354
rect 8745 4326 8750 4354
rect 8778 4326 12110 4354
rect 12138 4326 12143 4354
rect 14961 4326 14966 4354
rect 14994 4326 18998 4354
rect 19026 4326 19031 4354
rect 0 4298 56 4312
rect 2227 4298 2232 4326
rect 2260 4298 2284 4326
rect 2312 4298 2336 4326
rect 2364 4298 2369 4326
rect 12227 4298 12232 4326
rect 12260 4298 12284 4326
rect 12312 4298 12336 4326
rect 12364 4298 12369 4326
rect 22227 4298 22232 4326
rect 22260 4298 22284 4326
rect 22312 4298 22336 4326
rect 22364 4298 22369 4326
rect 26320 4298 26376 4312
rect 0 4270 1218 4298
rect 3761 4270 3766 4298
rect 3794 4270 10514 4298
rect 13673 4270 13678 4298
rect 13706 4270 14910 4298
rect 14938 4270 14943 4298
rect 15017 4270 15022 4298
rect 15050 4270 15862 4298
rect 15890 4270 15895 4298
rect 16473 4270 16478 4298
rect 16506 4270 18326 4298
rect 18354 4270 18359 4298
rect 25489 4270 25494 4298
rect 25522 4270 26376 4298
rect 0 4256 56 4270
rect 1190 4242 1218 4270
rect 10486 4242 10514 4270
rect 26320 4256 26376 4270
rect 1190 4214 2982 4242
rect 3010 4214 3015 4242
rect 3089 4214 3094 4242
rect 3122 4214 8358 4242
rect 8386 4214 8391 4242
rect 10486 4214 25102 4242
rect 25130 4214 25135 4242
rect 11713 4158 11718 4186
rect 11746 4158 13678 4186
rect 13706 4158 13711 4186
rect 13785 4158 13790 4186
rect 13818 4158 15246 4186
rect 15274 4158 15279 4186
rect 16809 4158 16814 4186
rect 16842 4158 18886 4186
rect 18914 4158 18919 4186
rect 19306 4158 23254 4186
rect 23282 4158 23287 4186
rect 19306 4130 19334 4158
rect 3369 4102 3374 4130
rect 3402 4102 9310 4130
rect 9338 4102 9343 4130
rect 11657 4102 11662 4130
rect 11690 4102 19334 4130
rect 24593 4102 24598 4130
rect 24626 4102 25214 4130
rect 25242 4102 25247 4130
rect 0 4074 56 4088
rect 26320 4074 26376 4088
rect 0 4046 3486 4074
rect 3514 4046 3519 4074
rect 11993 4046 11998 4074
rect 12026 4046 14854 4074
rect 14882 4046 14887 4074
rect 23473 4046 23478 4074
rect 23506 4046 25158 4074
rect 25186 4046 25191 4074
rect 25601 4046 25606 4074
rect 25634 4046 26376 4074
rect 0 4032 56 4046
rect 26320 4032 26376 4046
rect 1073 3990 1078 4018
rect 1106 3990 3206 4018
rect 3234 3990 3239 4018
rect 9473 3990 9478 4018
rect 9506 3990 13678 4018
rect 13706 3990 13711 4018
rect 15073 3990 15078 4018
rect 15106 3990 21294 4018
rect 21322 3990 21327 4018
rect 21826 3990 24766 4018
rect 24794 3990 24799 4018
rect 21826 3962 21854 3990
rect 10033 3934 10038 3962
rect 10066 3934 11774 3962
rect 11802 3934 11807 3962
rect 14177 3934 14182 3962
rect 14210 3934 21854 3962
rect 1897 3906 1902 3934
rect 1930 3906 1954 3934
rect 1982 3906 2006 3934
rect 2034 3906 2039 3934
rect 11897 3906 11902 3934
rect 11930 3906 11954 3934
rect 11982 3906 12006 3934
rect 12034 3906 12039 3934
rect 21897 3906 21902 3934
rect 21930 3906 21954 3934
rect 21982 3906 22006 3934
rect 22034 3906 22039 3934
rect 2977 3878 2982 3906
rect 3010 3878 7070 3906
rect 7098 3878 7103 3906
rect 10649 3878 10654 3906
rect 10682 3878 11606 3906
rect 11634 3878 11639 3906
rect 12105 3878 12110 3906
rect 12138 3878 13398 3906
rect 13426 3878 13431 3906
rect 13505 3878 13510 3906
rect 13538 3878 16982 3906
rect 17010 3878 17015 3906
rect 0 3850 56 3864
rect 26320 3850 26376 3864
rect 0 3822 2926 3850
rect 2954 3822 2959 3850
rect 8353 3822 8358 3850
rect 8386 3822 12502 3850
rect 12530 3822 12535 3850
rect 15017 3822 15022 3850
rect 15050 3822 16142 3850
rect 16170 3822 16175 3850
rect 16249 3822 16254 3850
rect 16282 3822 17822 3850
rect 17850 3822 17855 3850
rect 25713 3822 25718 3850
rect 25746 3822 26376 3850
rect 0 3808 56 3822
rect 26320 3808 26376 3822
rect 2753 3766 2758 3794
rect 2786 3766 6790 3794
rect 6818 3766 6823 3794
rect 10145 3766 10150 3794
rect 10178 3766 12278 3794
rect 12306 3766 12311 3794
rect 14233 3766 14238 3794
rect 14266 3766 16086 3794
rect 16114 3766 16119 3794
rect 24145 3766 24150 3794
rect 24178 3766 25270 3794
rect 25298 3766 25303 3794
rect 2137 3710 2142 3738
rect 2170 3710 24374 3738
rect 24402 3710 24407 3738
rect 2865 3654 2870 3682
rect 2898 3654 3710 3682
rect 3738 3654 3743 3682
rect 7121 3654 7126 3682
rect 7154 3654 10934 3682
rect 10962 3654 10967 3682
rect 11265 3654 11270 3682
rect 11298 3654 14910 3682
rect 14938 3654 14943 3682
rect 15022 3654 16870 3682
rect 16898 3654 16903 3682
rect 16977 3654 16982 3682
rect 17010 3654 23870 3682
rect 23898 3654 23903 3682
rect 0 3626 56 3640
rect 15022 3626 15050 3654
rect 26320 3626 26376 3640
rect 0 3598 2590 3626
rect 2618 3598 2623 3626
rect 2921 3598 2926 3626
rect 2954 3598 4326 3626
rect 4354 3598 4359 3626
rect 4489 3598 4494 3626
rect 4522 3598 6958 3626
rect 6986 3598 6991 3626
rect 9865 3598 9870 3626
rect 9898 3598 10990 3626
rect 11018 3598 11023 3626
rect 11102 3598 12670 3626
rect 12698 3598 12703 3626
rect 13897 3598 13902 3626
rect 13930 3598 15050 3626
rect 16086 3598 20286 3626
rect 20314 3598 20319 3626
rect 21826 3598 24430 3626
rect 24458 3598 24463 3626
rect 25713 3598 25718 3626
rect 25746 3598 26376 3626
rect 0 3584 56 3598
rect 2473 3542 2478 3570
rect 2506 3542 10486 3570
rect 10514 3542 10519 3570
rect 2227 3514 2232 3542
rect 2260 3514 2284 3542
rect 2312 3514 2336 3542
rect 2364 3514 2369 3542
rect 11102 3514 11130 3598
rect 12227 3514 12232 3542
rect 12260 3514 12284 3542
rect 12312 3514 12336 3542
rect 12364 3514 12369 3542
rect 5553 3486 5558 3514
rect 5586 3486 7574 3514
rect 7961 3486 7966 3514
rect 7994 3486 9646 3514
rect 9674 3486 9679 3514
rect 9977 3486 9982 3514
rect 10010 3486 11130 3514
rect 12609 3486 12614 3514
rect 12642 3486 15974 3514
rect 16002 3486 16007 3514
rect 7546 3458 7574 3486
rect 16086 3458 16114 3598
rect 21826 3570 21854 3598
rect 26320 3584 26376 3598
rect 16193 3542 16198 3570
rect 16226 3542 21854 3570
rect 22227 3514 22232 3542
rect 22260 3514 22284 3542
rect 22312 3514 22336 3542
rect 22364 3514 22369 3542
rect 849 3430 854 3458
rect 882 3430 2870 3458
rect 2898 3430 2903 3458
rect 7546 3430 16114 3458
rect 17873 3430 17878 3458
rect 17906 3430 18550 3458
rect 18578 3430 18583 3458
rect 0 3402 56 3416
rect 26320 3402 26376 3416
rect 0 3374 1806 3402
rect 1834 3374 1839 3402
rect 6734 3374 10094 3402
rect 10122 3374 10127 3402
rect 12553 3374 12558 3402
rect 12586 3374 13006 3402
rect 13034 3374 13039 3402
rect 13426 3374 14182 3402
rect 14210 3374 14215 3402
rect 15409 3374 15414 3402
rect 15442 3374 18046 3402
rect 18074 3374 18079 3402
rect 21681 3374 21686 3402
rect 21714 3374 22666 3402
rect 24817 3374 24822 3402
rect 24850 3374 26376 3402
rect 0 3360 56 3374
rect 6734 3346 6762 3374
rect 13426 3346 13454 3374
rect 22638 3346 22666 3374
rect 26320 3360 26376 3374
rect 4265 3318 4270 3346
rect 4298 3318 6762 3346
rect 9641 3318 9646 3346
rect 9674 3318 10290 3346
rect 10481 3318 10486 3346
rect 10514 3318 13454 3346
rect 14961 3318 14966 3346
rect 14994 3318 17766 3346
rect 17794 3318 17799 3346
rect 17878 3318 22134 3346
rect 22162 3318 22167 3346
rect 22638 3318 24430 3346
rect 24458 3318 24463 3346
rect 10262 3290 10290 3318
rect 17878 3290 17906 3318
rect 4153 3262 4158 3290
rect 4186 3262 6006 3290
rect 6034 3262 6039 3290
rect 7065 3262 7070 3290
rect 7098 3262 7574 3290
rect 10262 3262 13146 3290
rect 13393 3262 13398 3290
rect 13426 3262 15302 3290
rect 15330 3262 15335 3290
rect 16081 3262 16086 3290
rect 16114 3262 17906 3290
rect 18377 3262 18382 3290
rect 18410 3262 21294 3290
rect 21322 3262 21327 3290
rect 7546 3234 7574 3262
rect 13118 3234 13146 3262
rect 7546 3206 11662 3234
rect 11690 3206 11695 3234
rect 11774 3206 13006 3234
rect 13034 3206 13039 3234
rect 13118 3206 15638 3234
rect 15666 3206 15671 3234
rect 0 3178 56 3192
rect 11774 3178 11802 3206
rect 26320 3178 26376 3192
rect 0 3150 1834 3178
rect 9361 3150 9366 3178
rect 9394 3150 11802 3178
rect 13225 3150 13230 3178
rect 13258 3150 17654 3178
rect 17682 3150 17687 3178
rect 25601 3150 25606 3178
rect 25634 3150 26376 3178
rect 0 3136 56 3150
rect 1806 3066 1834 3150
rect 1897 3122 1902 3150
rect 1930 3122 1954 3150
rect 1982 3122 2006 3150
rect 2034 3122 2039 3150
rect 11897 3122 11902 3150
rect 11930 3122 11954 3150
rect 11982 3122 12006 3150
rect 12034 3122 12039 3150
rect 21897 3122 21902 3150
rect 21930 3122 21954 3150
rect 21982 3122 22006 3150
rect 22034 3122 22039 3150
rect 26320 3136 26376 3150
rect 6505 3094 6510 3122
rect 6538 3094 9198 3122
rect 9226 3094 9231 3122
rect 1806 3038 2534 3066
rect 2562 3038 2567 3066
rect 3313 3038 3318 3066
rect 3346 3038 6174 3066
rect 6202 3038 6207 3066
rect 7457 3038 7462 3066
rect 7490 3038 12614 3066
rect 12642 3038 12647 3066
rect 20617 3038 20622 3066
rect 20650 3038 25214 3066
rect 25242 3038 25247 3066
rect 849 2982 854 3010
rect 882 2982 2646 3010
rect 2674 2982 2679 3010
rect 3369 2982 3374 3010
rect 3402 2982 7126 3010
rect 7154 2982 7159 3010
rect 10593 2982 10598 3010
rect 10626 2982 15078 3010
rect 15106 2982 15111 3010
rect 15745 2982 15750 3010
rect 15778 2982 20510 3010
rect 20538 2982 20543 3010
rect 0 2954 56 2968
rect 26320 2954 26376 2968
rect 0 2926 2086 2954
rect 2114 2926 2119 2954
rect 3033 2926 3038 2954
rect 3066 2926 6622 2954
rect 6650 2926 6655 2954
rect 8185 2926 8190 2954
rect 8218 2926 12782 2954
rect 12810 2926 12815 2954
rect 14961 2926 14966 2954
rect 14994 2926 18606 2954
rect 18634 2926 18639 2954
rect 20057 2926 20062 2954
rect 20090 2926 22358 2954
rect 22386 2926 22391 2954
rect 24873 2926 24878 2954
rect 24906 2926 26376 2954
rect 0 2912 56 2926
rect 26320 2912 26376 2926
rect 6113 2870 6118 2898
rect 6146 2870 7182 2898
rect 7210 2870 7215 2898
rect 8073 2870 8078 2898
rect 8106 2870 9254 2898
rect 9282 2870 9287 2898
rect 9422 2870 12894 2898
rect 12922 2870 12927 2898
rect 13001 2870 13006 2898
rect 13034 2870 15246 2898
rect 15274 2870 15279 2898
rect 16529 2870 16534 2898
rect 16562 2870 16758 2898
rect 16786 2870 16791 2898
rect 17593 2870 17598 2898
rect 17626 2870 19334 2898
rect 19362 2870 19367 2898
rect 20337 2870 20342 2898
rect 20370 2870 23590 2898
rect 23618 2870 23623 2898
rect 9422 2842 9450 2870
rect 1073 2814 1078 2842
rect 1106 2814 4998 2842
rect 5026 2814 5031 2842
rect 6673 2814 6678 2842
rect 6706 2814 7518 2842
rect 7546 2814 7551 2842
rect 8521 2814 8526 2842
rect 8554 2814 9450 2842
rect 10486 2814 25102 2842
rect 25130 2814 25135 2842
rect 10486 2786 10514 2814
rect 2753 2758 2758 2786
rect 2786 2758 10514 2786
rect 10593 2758 10598 2786
rect 10626 2758 12166 2786
rect 12194 2758 12199 2786
rect 12665 2758 12670 2786
rect 12698 2758 13790 2786
rect 13818 2758 13823 2786
rect 15190 2758 19054 2786
rect 19082 2758 19087 2786
rect 0 2730 56 2744
rect 2227 2730 2232 2758
rect 2260 2730 2284 2758
rect 2312 2730 2336 2758
rect 2364 2730 2369 2758
rect 12227 2730 12232 2758
rect 12260 2730 12284 2758
rect 12312 2730 12336 2758
rect 12364 2730 12369 2758
rect 0 2702 1806 2730
rect 1834 2702 1839 2730
rect 6113 2702 6118 2730
rect 6146 2702 11718 2730
rect 11746 2702 11751 2730
rect 0 2688 56 2702
rect 15190 2674 15218 2758
rect 22227 2730 22232 2758
rect 22260 2730 22284 2758
rect 22312 2730 22336 2758
rect 22364 2730 22369 2758
rect 26320 2730 26376 2744
rect 15577 2702 15582 2730
rect 15610 2702 16590 2730
rect 16618 2702 16623 2730
rect 17873 2702 17878 2730
rect 17906 2702 20398 2730
rect 20426 2702 20431 2730
rect 25601 2702 25606 2730
rect 25634 2702 26376 2730
rect 26320 2688 26376 2702
rect 7065 2646 7070 2674
rect 7098 2646 10934 2674
rect 10962 2646 10967 2674
rect 11097 2646 11102 2674
rect 11130 2646 15218 2674
rect 15246 2646 18158 2674
rect 18186 2646 18191 2674
rect 19161 2646 19166 2674
rect 19194 2646 24934 2674
rect 24962 2646 24967 2674
rect 15246 2618 15274 2646
rect 2137 2590 2142 2618
rect 2170 2590 6342 2618
rect 6370 2590 6375 2618
rect 6449 2590 6454 2618
rect 6482 2590 10598 2618
rect 10626 2590 10631 2618
rect 11265 2590 11270 2618
rect 11298 2590 15274 2618
rect 15353 2590 15358 2618
rect 15386 2590 16030 2618
rect 16058 2590 16063 2618
rect 16305 2590 16310 2618
rect 16338 2590 17654 2618
rect 17682 2590 17687 2618
rect 24481 2590 24486 2618
rect 24514 2590 25214 2618
rect 25242 2590 25247 2618
rect 2417 2534 2422 2562
rect 2450 2534 4214 2562
rect 7345 2534 7350 2562
rect 7378 2534 7630 2562
rect 7658 2534 7663 2562
rect 11209 2534 11214 2562
rect 11242 2534 14966 2562
rect 14994 2534 14999 2562
rect 15073 2534 15078 2562
rect 15106 2534 16198 2562
rect 16226 2534 16231 2562
rect 16473 2534 16478 2562
rect 16506 2534 16511 2562
rect 17369 2534 17374 2562
rect 17402 2534 17990 2562
rect 18018 2534 18023 2562
rect 23417 2534 23422 2562
rect 23450 2534 24374 2562
rect 24402 2534 24407 2562
rect 24817 2534 24822 2562
rect 24850 2534 25550 2562
rect 25578 2534 25583 2562
rect 0 2506 56 2520
rect 4186 2506 4214 2534
rect 16478 2506 16506 2534
rect 26320 2506 26376 2520
rect 0 2478 2926 2506
rect 2954 2478 2959 2506
rect 4186 2478 6566 2506
rect 6594 2478 6599 2506
rect 9142 2478 9982 2506
rect 10010 2478 10015 2506
rect 10201 2478 10206 2506
rect 10234 2478 12670 2506
rect 12698 2478 12703 2506
rect 13057 2478 13062 2506
rect 13090 2478 13398 2506
rect 13426 2478 13431 2506
rect 14513 2478 14518 2506
rect 14546 2478 16506 2506
rect 16641 2478 16646 2506
rect 16674 2478 21070 2506
rect 21098 2478 21103 2506
rect 25433 2478 25438 2506
rect 25466 2478 26376 2506
rect 0 2464 56 2478
rect 6617 2422 6622 2450
rect 6650 2422 8358 2450
rect 8386 2422 8391 2450
rect 9142 2394 9170 2478
rect 26320 2464 26376 2478
rect 10481 2422 10486 2450
rect 10514 2422 14014 2450
rect 14042 2422 14047 2450
rect 15129 2422 15134 2450
rect 15162 2422 15526 2450
rect 15554 2422 15559 2450
rect 15857 2422 15862 2450
rect 15890 2422 18662 2450
rect 18690 2422 18695 2450
rect 19306 2422 24654 2450
rect 24682 2422 24687 2450
rect 19306 2394 19334 2422
rect 6729 2366 6734 2394
rect 6762 2366 9170 2394
rect 12161 2366 12166 2394
rect 12194 2366 12558 2394
rect 12586 2366 12591 2394
rect 12665 2366 12670 2394
rect 12698 2366 19334 2394
rect 1897 2338 1902 2366
rect 1930 2338 1954 2366
rect 1982 2338 2006 2366
rect 2034 2338 2039 2366
rect 11897 2338 11902 2366
rect 11930 2338 11954 2366
rect 11982 2338 12006 2366
rect 12034 2338 12039 2366
rect 21897 2338 21902 2366
rect 21930 2338 21954 2366
rect 21982 2338 22006 2366
rect 22034 2338 22039 2366
rect 2529 2310 2534 2338
rect 2562 2310 6118 2338
rect 6146 2310 6151 2338
rect 8353 2310 8358 2338
rect 8386 2310 11046 2338
rect 11074 2310 11079 2338
rect 12105 2310 12110 2338
rect 12138 2310 13370 2338
rect 14681 2310 14686 2338
rect 14714 2310 15974 2338
rect 16002 2310 16007 2338
rect 18993 2310 18998 2338
rect 19026 2310 21462 2338
rect 21490 2310 21495 2338
rect 0 2282 56 2296
rect 13342 2282 13370 2310
rect 26320 2282 26376 2296
rect 0 2254 3094 2282
rect 3122 2254 3127 2282
rect 7546 2254 10486 2282
rect 10514 2254 10519 2282
rect 10929 2254 10934 2282
rect 10962 2254 13230 2282
rect 13258 2254 13263 2282
rect 13342 2254 15918 2282
rect 15946 2254 15951 2282
rect 16137 2254 16142 2282
rect 16170 2254 20202 2282
rect 25545 2254 25550 2282
rect 25578 2254 26376 2282
rect 0 2240 56 2254
rect 7546 2226 7574 2254
rect 2697 2198 2702 2226
rect 2730 2198 7574 2226
rect 10150 2198 12782 2226
rect 12810 2198 12815 2226
rect 12889 2198 12894 2226
rect 12922 2198 15694 2226
rect 15722 2198 15727 2226
rect 16305 2198 16310 2226
rect 16338 2198 19110 2226
rect 19138 2198 19143 2226
rect 10150 2170 10178 2198
rect 2865 2142 2870 2170
rect 2898 2142 4214 2170
rect 5889 2142 5894 2170
rect 5922 2142 10178 2170
rect 11825 2142 11830 2170
rect 11858 2142 14686 2170
rect 14714 2142 14719 2170
rect 15190 2142 16982 2170
rect 17010 2142 17015 2170
rect 18769 2142 18774 2170
rect 18802 2142 20062 2170
rect 20090 2142 20095 2170
rect 4186 2114 4214 2142
rect 15190 2114 15218 2142
rect 961 2086 966 2114
rect 994 2086 2590 2114
rect 2618 2086 2623 2114
rect 4186 2086 11998 2114
rect 12026 2086 12031 2114
rect 12614 2086 15218 2114
rect 15302 2086 18494 2114
rect 18522 2086 18527 2114
rect 0 2058 56 2072
rect 12614 2058 12642 2086
rect 0 2030 1470 2058
rect 1498 2030 1503 2058
rect 9193 2030 9198 2058
rect 9226 2030 12642 2058
rect 12721 2030 12726 2058
rect 12754 2030 14294 2058
rect 14322 2030 14327 2058
rect 14569 2030 14574 2058
rect 14602 2030 14966 2058
rect 14994 2030 14999 2058
rect 0 2016 56 2030
rect 15302 2002 15330 2086
rect 20174 2058 20202 2254
rect 26320 2240 26376 2254
rect 24089 2198 24094 2226
rect 24122 2198 24430 2226
rect 24458 2198 24463 2226
rect 21121 2086 21126 2114
rect 21154 2086 23814 2114
rect 23842 2086 23847 2114
rect 26320 2058 26376 2072
rect 16305 2030 16310 2058
rect 16338 2030 17318 2058
rect 17346 2030 17351 2058
rect 19217 2030 19222 2058
rect 19250 2030 19670 2058
rect 19698 2030 19703 2058
rect 20174 2030 22190 2058
rect 22218 2030 22223 2058
rect 25713 2030 25718 2058
rect 25746 2030 26376 2058
rect 26320 2016 26376 2030
rect 3929 1974 3934 2002
rect 3962 1974 5782 2002
rect 5810 1974 5815 2002
rect 9249 1974 9254 2002
rect 9282 1974 12054 2002
rect 12082 1974 12087 2002
rect 12833 1974 12838 2002
rect 12866 1974 15330 2002
rect 15689 1974 15694 2002
rect 15722 1974 19334 2002
rect 19362 1974 19367 2002
rect 2227 1946 2232 1974
rect 2260 1946 2284 1974
rect 2312 1946 2336 1974
rect 2364 1946 2369 1974
rect 12227 1946 12232 1974
rect 12260 1946 12284 1974
rect 12312 1946 12336 1974
rect 12364 1946 12369 1974
rect 22227 1946 22232 1974
rect 22260 1946 22284 1974
rect 22312 1946 22336 1974
rect 22364 1946 22369 1974
rect 4209 1918 4214 1946
rect 4242 1918 7574 1946
rect 9753 1918 9758 1946
rect 9786 1918 11550 1946
rect 11578 1918 11583 1946
rect 7546 1890 7574 1918
rect 1694 1862 4382 1890
rect 4410 1862 4415 1890
rect 7546 1862 13006 1890
rect 13034 1862 13039 1890
rect 13174 1862 25214 1890
rect 25242 1862 25247 1890
rect 0 1834 56 1848
rect 1694 1834 1722 1862
rect 0 1806 1722 1834
rect 2641 1806 2646 1834
rect 2674 1806 11382 1834
rect 11410 1806 11415 1834
rect 11545 1806 11550 1834
rect 11578 1806 12726 1834
rect 12754 1806 12759 1834
rect 0 1792 56 1806
rect 11433 1750 11438 1778
rect 11466 1750 12614 1778
rect 12642 1750 12647 1778
rect 13174 1722 13202 1862
rect 26320 1834 26376 1848
rect 13281 1806 13286 1834
rect 13314 1806 14126 1834
rect 14154 1806 14159 1834
rect 14233 1806 14238 1834
rect 14266 1806 15750 1834
rect 15778 1806 15783 1834
rect 17593 1806 17598 1834
rect 17626 1806 17934 1834
rect 17962 1806 17967 1834
rect 19161 1806 19166 1834
rect 19194 1806 20790 1834
rect 20818 1806 20823 1834
rect 20897 1806 20902 1834
rect 20930 1806 23534 1834
rect 23562 1806 23567 1834
rect 24705 1806 24710 1834
rect 24738 1806 26376 1834
rect 26320 1792 26376 1806
rect 13449 1750 13454 1778
rect 13482 1750 16198 1778
rect 16226 1750 16231 1778
rect 17257 1750 17262 1778
rect 17290 1750 18662 1778
rect 18690 1750 18695 1778
rect 22465 1750 22470 1778
rect 22498 1750 25102 1778
rect 25130 1750 25135 1778
rect 905 1694 910 1722
rect 938 1694 3542 1722
rect 3570 1694 3575 1722
rect 5838 1694 8302 1722
rect 8330 1694 8335 1722
rect 10066 1694 11634 1722
rect 11713 1694 11718 1722
rect 11746 1694 13202 1722
rect 15353 1694 15358 1722
rect 15386 1694 16478 1722
rect 16506 1694 16511 1722
rect 16641 1694 16646 1722
rect 16674 1694 17878 1722
rect 17906 1694 17911 1722
rect 19441 1694 19446 1722
rect 19474 1694 20342 1722
rect 20370 1694 20375 1722
rect 24929 1694 24934 1722
rect 24962 1694 25494 1722
rect 25522 1694 25527 1722
rect 5838 1666 5866 1694
rect 10066 1666 10094 1694
rect 1806 1638 5866 1666
rect 6785 1638 6790 1666
rect 6818 1638 10094 1666
rect 11606 1666 11634 1694
rect 11606 1638 12362 1666
rect 12609 1638 12614 1666
rect 12642 1638 15246 1666
rect 15274 1638 15279 1666
rect 15913 1638 15918 1666
rect 15946 1638 17094 1666
rect 17122 1638 17127 1666
rect 21826 1638 24486 1666
rect 24514 1638 24519 1666
rect 0 1610 56 1624
rect 1806 1610 1834 1638
rect 12334 1610 12362 1638
rect 21826 1610 21854 1638
rect 26320 1610 26376 1624
rect 0 1582 1834 1610
rect 2473 1582 2478 1610
rect 2506 1582 3318 1610
rect 3346 1582 3351 1610
rect 12334 1582 13510 1610
rect 13538 1582 13543 1610
rect 15465 1582 15470 1610
rect 15498 1582 15806 1610
rect 15834 1582 15839 1610
rect 15969 1582 15974 1610
rect 16002 1582 21854 1610
rect 25545 1582 25550 1610
rect 25578 1582 26376 1610
rect 0 1568 56 1582
rect 1897 1554 1902 1582
rect 1930 1554 1954 1582
rect 1982 1554 2006 1582
rect 2034 1554 2039 1582
rect 11897 1554 11902 1582
rect 11930 1554 11954 1582
rect 11982 1554 12006 1582
rect 12034 1554 12039 1582
rect 21897 1554 21902 1582
rect 21930 1554 21954 1582
rect 21982 1554 22006 1582
rect 22034 1554 22039 1582
rect 26320 1568 26376 1582
rect 5217 1526 5222 1554
rect 5250 1526 6734 1554
rect 6762 1526 6767 1554
rect 12945 1526 12950 1554
rect 12978 1526 13622 1554
rect 13650 1526 13655 1554
rect 13785 1526 13790 1554
rect 13818 1526 20342 1554
rect 20370 1526 20375 1554
rect 6337 1470 6342 1498
rect 6370 1470 13342 1498
rect 13370 1470 13375 1498
rect 13505 1470 13510 1498
rect 13538 1470 20174 1498
rect 20202 1470 20207 1498
rect 20281 1470 20286 1498
rect 20314 1470 23534 1498
rect 23562 1470 23567 1498
rect 1745 1414 1750 1442
rect 1778 1414 2534 1442
rect 2562 1414 2567 1442
rect 5665 1414 5670 1442
rect 5698 1414 10262 1442
rect 10290 1414 10295 1442
rect 10985 1414 10990 1442
rect 11018 1414 11914 1442
rect 11993 1414 11998 1442
rect 12026 1414 15414 1442
rect 15442 1414 15447 1442
rect 16865 1414 16870 1442
rect 16898 1414 17598 1442
rect 17626 1414 17631 1442
rect 19105 1414 19110 1442
rect 19138 1414 23086 1442
rect 23114 1414 23119 1442
rect 24033 1414 24038 1442
rect 24066 1414 25326 1442
rect 25354 1414 25359 1442
rect 0 1386 56 1400
rect 11886 1386 11914 1414
rect 26320 1386 26376 1400
rect 0 1358 6510 1386
rect 6538 1358 6543 1386
rect 8633 1358 8638 1386
rect 8666 1358 11774 1386
rect 11802 1358 11807 1386
rect 11886 1358 12642 1386
rect 12721 1358 12726 1386
rect 12754 1358 13454 1386
rect 15297 1358 15302 1386
rect 15330 1358 18158 1386
rect 18186 1358 18191 1386
rect 19553 1358 19558 1386
rect 19586 1358 21518 1386
rect 21546 1358 21551 1386
rect 25489 1358 25494 1386
rect 25522 1358 26376 1386
rect 0 1344 56 1358
rect 1297 1302 1302 1330
rect 1330 1302 2702 1330
rect 2730 1302 2735 1330
rect 11153 1302 11158 1330
rect 11186 1302 11494 1330
rect 11522 1302 11527 1330
rect 11601 1302 11606 1330
rect 11634 1302 12502 1330
rect 12530 1302 12535 1330
rect 12614 1274 12642 1358
rect 13426 1330 13454 1358
rect 26320 1344 26376 1358
rect 13426 1302 16198 1330
rect 16226 1302 16231 1330
rect 16697 1302 16702 1330
rect 16730 1302 18382 1330
rect 18410 1302 18415 1330
rect 23361 1302 23366 1330
rect 23394 1302 24374 1330
rect 24402 1302 24407 1330
rect 24705 1302 24710 1330
rect 24738 1302 25438 1330
rect 25466 1302 25471 1330
rect 9417 1246 9422 1274
rect 9450 1246 11326 1274
rect 11354 1246 11359 1274
rect 11769 1246 11774 1274
rect 11802 1246 12586 1274
rect 12614 1246 19726 1274
rect 19754 1246 19759 1274
rect 22745 1246 22750 1274
rect 22778 1246 24430 1274
rect 24458 1246 24463 1274
rect 12558 1218 12586 1246
rect 8689 1190 8694 1218
rect 8722 1190 11998 1218
rect 12026 1190 12031 1218
rect 12558 1190 13902 1218
rect 13930 1190 13935 1218
rect 18545 1190 18550 1218
rect 18578 1190 18774 1218
rect 18802 1190 18807 1218
rect 0 1162 56 1176
rect 2227 1162 2232 1190
rect 2260 1162 2284 1190
rect 2312 1162 2336 1190
rect 2364 1162 2369 1190
rect 12227 1162 12232 1190
rect 12260 1162 12284 1190
rect 12312 1162 12336 1190
rect 12364 1162 12369 1190
rect 22227 1162 22232 1190
rect 22260 1162 22284 1190
rect 22312 1162 22336 1190
rect 22364 1162 22369 1190
rect 26320 1162 26376 1176
rect 0 1134 1386 1162
rect 3705 1134 3710 1162
rect 3738 1134 7574 1162
rect 8017 1134 8022 1162
rect 8050 1134 11494 1162
rect 11522 1134 11527 1162
rect 14401 1134 14406 1162
rect 14434 1134 14798 1162
rect 14826 1134 14831 1162
rect 18657 1134 18662 1162
rect 18690 1134 21854 1162
rect 25713 1134 25718 1162
rect 25746 1134 26376 1162
rect 0 1120 56 1134
rect 1358 1106 1386 1134
rect 7546 1106 7574 1134
rect 21826 1106 21854 1134
rect 26320 1120 26376 1134
rect 1358 1078 2814 1106
rect 2842 1078 2847 1106
rect 7546 1078 12894 1106
rect 12922 1078 12927 1106
rect 13113 1078 13118 1106
rect 13146 1078 13230 1106
rect 13258 1078 13263 1106
rect 14737 1078 14742 1106
rect 14770 1078 15974 1106
rect 17425 1078 17430 1106
rect 17458 1078 19166 1106
rect 19194 1078 19199 1106
rect 21826 1078 23534 1106
rect 23562 1078 23567 1106
rect 15946 1050 15974 1078
rect 2585 1022 2590 1050
rect 2618 1022 11382 1050
rect 11410 1022 11415 1050
rect 11489 1022 11494 1050
rect 11522 1022 14462 1050
rect 14490 1022 14495 1050
rect 15017 1022 15022 1050
rect 15050 1022 15862 1050
rect 15890 1022 15895 1050
rect 15946 1022 22470 1050
rect 22498 1022 22503 1050
rect 5833 966 5838 994
rect 5866 966 7070 994
rect 7098 966 7103 994
rect 10313 966 10318 994
rect 10346 966 12838 994
rect 12866 966 12871 994
rect 18377 966 18382 994
rect 18410 966 19614 994
rect 19642 966 19647 994
rect 23753 966 23758 994
rect 23786 966 25214 994
rect 25242 966 25247 994
rect 0 938 56 952
rect 26320 938 26376 952
rect 0 910 5390 938
rect 5418 910 5423 938
rect 5665 910 5670 938
rect 5698 910 12614 938
rect 12642 910 12647 938
rect 12721 910 12726 938
rect 12754 910 18494 938
rect 18522 910 18527 938
rect 24929 910 24934 938
rect 24962 910 26376 938
rect 0 896 56 910
rect 26320 896 26376 910
rect 3145 854 3150 882
rect 3178 854 5474 882
rect 10873 854 10878 882
rect 10906 854 12446 882
rect 12474 854 12479 882
rect 12833 854 12838 882
rect 12866 854 14546 882
rect 15745 854 15750 882
rect 15778 854 17878 882
rect 17906 854 17911 882
rect 1897 770 1902 798
rect 1930 770 1954 798
rect 1982 770 2006 798
rect 2034 770 2039 798
rect 5446 770 5474 854
rect 14518 826 14546 854
rect 6673 798 6678 826
rect 6706 798 7294 826
rect 7322 798 7327 826
rect 7401 798 7406 826
rect 7434 798 8470 826
rect 8498 798 8503 826
rect 8633 798 8638 826
rect 8666 798 11158 826
rect 11186 798 11191 826
rect 12390 798 13454 826
rect 13482 798 13487 826
rect 14009 798 14014 826
rect 14042 798 14350 826
rect 14378 798 14383 826
rect 14518 798 14770 826
rect 15689 798 15694 826
rect 15722 798 16422 826
rect 16450 798 16455 826
rect 17481 798 17486 826
rect 17514 798 18270 826
rect 18298 798 18303 826
rect 19609 798 19614 826
rect 19642 798 20566 826
rect 20594 798 20599 826
rect 11897 770 11902 798
rect 11930 770 11954 798
rect 11982 770 12006 798
rect 12034 770 12039 798
rect 12390 770 12418 798
rect 14742 770 14770 798
rect 21897 770 21902 798
rect 21930 770 21954 798
rect 21982 770 22006 798
rect 22034 770 22039 798
rect 5446 742 6734 770
rect 6762 742 6767 770
rect 9025 742 9030 770
rect 9058 742 11298 770
rect 0 714 56 728
rect 11270 714 11298 742
rect 12110 742 12418 770
rect 12497 742 12502 770
rect 12530 742 14630 770
rect 14658 742 14663 770
rect 14742 742 17654 770
rect 17705 742 17710 770
rect 17738 742 18606 770
rect 18634 742 18639 770
rect 18718 742 19446 770
rect 19474 742 19479 770
rect 19833 742 19838 770
rect 19866 742 21014 770
rect 21042 742 21047 770
rect 12110 714 12138 742
rect 17626 714 17654 742
rect 18718 714 18746 742
rect 26320 714 26376 728
rect 0 686 3318 714
rect 3346 686 3351 714
rect 6001 686 6006 714
rect 6034 686 6846 714
rect 6874 686 6879 714
rect 11270 686 12138 714
rect 12166 686 13118 714
rect 13146 686 13151 714
rect 13225 686 13230 714
rect 13258 686 13622 714
rect 13650 686 13655 714
rect 14457 686 14462 714
rect 14490 686 15190 714
rect 15218 686 15223 714
rect 15465 686 15470 714
rect 15498 686 16870 714
rect 16898 686 16903 714
rect 17626 686 18746 714
rect 18937 686 18942 714
rect 18970 686 18975 714
rect 19161 686 19166 714
rect 19194 686 20230 714
rect 20258 686 20263 714
rect 20337 686 20342 714
rect 20370 686 24318 714
rect 24346 686 24351 714
rect 24873 686 24878 714
rect 24906 686 26376 714
rect 0 672 56 686
rect 12166 658 12194 686
rect 18942 658 18970 686
rect 26320 672 26376 686
rect 6393 630 6398 658
rect 6426 630 11046 658
rect 11074 630 11079 658
rect 11265 630 11270 658
rect 11298 630 12194 658
rect 12441 630 12446 658
rect 12474 630 13510 658
rect 13538 630 13543 658
rect 13897 630 13902 658
rect 13930 630 14518 658
rect 14546 630 14551 658
rect 14793 630 14798 658
rect 14826 630 16086 658
rect 16114 630 16119 658
rect 16585 630 16590 658
rect 16618 630 18270 658
rect 18298 630 18303 658
rect 18942 630 19110 658
rect 19138 630 19143 658
rect 19945 630 19950 658
rect 19978 630 22806 658
rect 22834 630 22839 658
rect 3537 574 3542 602
rect 3570 574 10262 602
rect 10290 574 10295 602
rect 10374 574 12502 602
rect 12530 574 12535 602
rect 12889 574 12894 602
rect 12922 574 13286 602
rect 13314 574 13319 602
rect 13393 574 13398 602
rect 13426 574 13846 602
rect 13874 574 13879 602
rect 14345 574 14350 602
rect 14378 574 15302 602
rect 15330 574 15335 602
rect 15857 574 15862 602
rect 15890 574 16534 602
rect 16562 574 16567 602
rect 17761 574 17766 602
rect 17794 574 25270 602
rect 25298 574 25303 602
rect 10374 546 10402 574
rect 4186 518 9254 546
rect 9282 518 9287 546
rect 9921 518 9926 546
rect 9954 518 10402 546
rect 10481 518 10486 546
rect 10514 518 12446 546
rect 12474 518 12479 546
rect 12553 518 12558 546
rect 12586 518 13006 546
rect 13034 518 13039 546
rect 13118 518 14406 546
rect 14434 518 14439 546
rect 14681 518 14686 546
rect 14714 518 16814 546
rect 16842 518 16847 546
rect 17593 518 17598 546
rect 17626 518 20566 546
rect 20594 518 20599 546
rect 20953 518 20958 546
rect 20986 518 23870 546
rect 23898 518 23903 546
rect 0 490 56 504
rect 4186 490 4214 518
rect 13118 490 13146 518
rect 26320 490 26376 504
rect 0 462 1302 490
rect 1330 462 1335 490
rect 1801 462 1806 490
rect 1834 462 4214 490
rect 4993 462 4998 490
rect 5026 462 6510 490
rect 6538 462 6543 490
rect 8409 462 8414 490
rect 8442 462 11270 490
rect 11298 462 11303 490
rect 11881 462 11886 490
rect 11914 462 13146 490
rect 13449 462 13454 490
rect 13482 462 14126 490
rect 14154 462 14159 490
rect 14233 462 14238 490
rect 14266 462 16030 490
rect 16058 462 16063 490
rect 16529 462 16534 490
rect 16562 462 18830 490
rect 18858 462 18863 490
rect 20057 462 20062 490
rect 20090 462 21406 490
rect 21434 462 21439 490
rect 24089 462 24094 490
rect 24122 462 26376 490
rect 0 448 56 462
rect 26320 448 26376 462
rect 5777 406 5782 434
rect 5810 406 12166 434
rect 12194 406 12199 434
rect 13505 406 13510 434
rect 13538 406 14070 434
rect 14098 406 14103 434
rect 14910 406 16478 434
rect 16506 406 16511 434
rect 2227 378 2232 406
rect 2260 378 2284 406
rect 2312 378 2336 406
rect 2364 378 2369 406
rect 12227 378 12232 406
rect 12260 378 12284 406
rect 12312 378 12336 406
rect 12364 378 12369 406
rect 14910 378 14938 406
rect 22227 378 22232 406
rect 22260 378 22284 406
rect 22312 378 22336 406
rect 22364 378 22369 406
rect 12441 350 12446 378
rect 12474 350 14182 378
rect 14210 350 14215 378
rect 14905 350 14910 378
rect 14938 350 14943 378
rect 18097 350 18102 378
rect 18130 350 18718 378
rect 18746 350 18751 378
rect 9305 294 9310 322
rect 9338 294 10374 322
rect 10402 294 10407 322
rect 11769 294 11774 322
rect 11802 294 12334 322
rect 12362 294 12367 322
rect 12670 294 13510 322
rect 13538 294 13543 322
rect 13785 294 13790 322
rect 13818 294 14742 322
rect 14770 294 14775 322
rect 15241 294 15246 322
rect 15274 294 17262 322
rect 17290 294 17295 322
rect 0 266 56 280
rect 0 238 5278 266
rect 5306 238 5311 266
rect 11489 238 11494 266
rect 11522 238 12558 266
rect 12586 238 12591 266
rect 0 224 56 238
rect 1129 182 1134 210
rect 1162 182 6398 210
rect 6426 182 6431 210
rect 11769 182 11774 210
rect 11802 182 12502 210
rect 12530 182 12535 210
rect 3201 126 3206 154
rect 3234 126 6286 154
rect 6314 126 6319 154
rect 10817 126 10822 154
rect 10850 126 12110 154
rect 12138 126 12143 154
rect 12670 98 12698 294
rect 26320 266 26376 280
rect 13057 238 13062 266
rect 13090 238 13594 266
rect 13673 238 13678 266
rect 13706 238 14854 266
rect 14882 238 14887 266
rect 15577 238 15582 266
rect 15610 238 17934 266
rect 17962 238 17967 266
rect 25321 238 25326 266
rect 25354 238 26376 266
rect 13566 154 13594 238
rect 26320 224 26376 238
rect 14121 182 14126 210
rect 14154 182 15526 210
rect 15554 182 15559 210
rect 16137 182 16142 210
rect 16170 182 19110 210
rect 19138 182 19143 210
rect 12945 126 12950 154
rect 12978 126 12983 154
rect 13566 126 15750 154
rect 15778 126 15783 154
rect 16753 126 16758 154
rect 16786 126 16791 154
rect 16921 126 16926 154
rect 16954 126 19670 154
rect 19698 126 19703 154
rect 1241 70 1246 98
rect 1274 70 6174 98
rect 6202 70 6207 98
rect 8297 70 8302 98
rect 8330 70 8335 98
rect 10761 70 10766 98
rect 10794 70 12698 98
rect 0 42 56 56
rect 8302 42 8330 70
rect 12950 42 12978 126
rect 16758 98 16786 126
rect 16758 70 17934 98
rect 17962 70 17967 98
rect 26320 42 26376 56
rect 0 14 4942 42
rect 4970 14 4975 42
rect 8302 14 12978 42
rect 25433 14 25438 42
rect 25466 14 26376 42
rect 0 0 56 14
rect 26320 0 26376 14
<< via3 >>
rect 2232 6650 2260 6678
rect 2284 6650 2312 6678
rect 2336 6650 2364 6678
rect 12232 6650 12260 6678
rect 12284 6650 12312 6678
rect 12336 6650 12364 6678
rect 22232 6650 22260 6678
rect 22284 6650 22312 6678
rect 22336 6650 22364 6678
rect 1902 6258 1930 6286
rect 1954 6258 1982 6286
rect 2006 6258 2034 6286
rect 11902 6258 11930 6286
rect 11954 6258 11982 6286
rect 12006 6258 12034 6286
rect 21902 6258 21930 6286
rect 21954 6258 21982 6286
rect 22006 6258 22034 6286
rect 13342 6174 13370 6202
rect 16310 5950 16338 5978
rect 19222 5950 19250 5978
rect 2232 5866 2260 5894
rect 2284 5866 2312 5894
rect 2336 5866 2364 5894
rect 12232 5866 12260 5894
rect 12284 5866 12312 5894
rect 12336 5866 12364 5894
rect 22232 5866 22260 5894
rect 22284 5866 22312 5894
rect 22336 5866 22364 5894
rect 9030 5782 9058 5810
rect 19222 5782 19250 5810
rect 9030 5558 9058 5586
rect 1902 5474 1930 5502
rect 1954 5474 1982 5502
rect 2006 5474 2034 5502
rect 11902 5474 11930 5502
rect 11954 5474 11982 5502
rect 12006 5474 12034 5502
rect 21902 5474 21930 5502
rect 21954 5474 21982 5502
rect 22006 5474 22034 5502
rect 12838 5334 12866 5362
rect 12502 5278 12530 5306
rect 2232 5082 2260 5110
rect 2284 5082 2312 5110
rect 2336 5082 2364 5110
rect 12232 5082 12260 5110
rect 12284 5082 12312 5110
rect 12336 5082 12364 5110
rect 22232 5082 22260 5110
rect 22284 5082 22312 5110
rect 22336 5082 22364 5110
rect 16590 4942 16618 4970
rect 13342 4830 13370 4858
rect 13454 4830 13482 4858
rect 13286 4718 13314 4746
rect 1902 4690 1930 4718
rect 1954 4690 1982 4718
rect 2006 4690 2034 4718
rect 11902 4690 11930 4718
rect 11954 4690 11982 4718
rect 12006 4690 12034 4718
rect 21902 4690 21930 4718
rect 21954 4690 21982 4718
rect 22006 4690 22034 4718
rect 14966 4494 14994 4522
rect 2232 4298 2260 4326
rect 2284 4298 2312 4326
rect 2336 4298 2364 4326
rect 12232 4298 12260 4326
rect 12284 4298 12312 4326
rect 12336 4298 12364 4326
rect 22232 4298 22260 4326
rect 22284 4298 22312 4326
rect 22336 4298 22364 4326
rect 15022 4270 15050 4298
rect 14182 3934 14210 3962
rect 1902 3906 1930 3934
rect 1954 3906 1982 3934
rect 2006 3906 2034 3934
rect 11902 3906 11930 3934
rect 11954 3906 11982 3934
rect 12006 3906 12034 3934
rect 21902 3906 21930 3934
rect 21954 3906 21982 3934
rect 22006 3906 22034 3934
rect 13510 3878 13538 3906
rect 16982 3878 17010 3906
rect 16142 3822 16170 3850
rect 16982 3654 17010 3682
rect 10486 3542 10514 3570
rect 2232 3514 2260 3542
rect 2284 3514 2312 3542
rect 2336 3514 2364 3542
rect 12232 3514 12260 3542
rect 12284 3514 12312 3542
rect 12336 3514 12364 3542
rect 16198 3542 16226 3570
rect 22232 3514 22260 3542
rect 22284 3514 22312 3542
rect 22336 3514 22364 3542
rect 14182 3374 14210 3402
rect 10486 3318 10514 3346
rect 13006 3206 13034 3234
rect 1902 3122 1930 3150
rect 1954 3122 1982 3150
rect 2006 3122 2034 3150
rect 11902 3122 11930 3150
rect 11954 3122 11982 3150
rect 12006 3122 12034 3150
rect 21902 3122 21930 3150
rect 21954 3122 21982 3150
rect 22006 3122 22034 3150
rect 14966 2926 14994 2954
rect 13006 2870 13034 2898
rect 10598 2758 10626 2786
rect 2232 2730 2260 2758
rect 2284 2730 2312 2758
rect 2336 2730 2364 2758
rect 12232 2730 12260 2758
rect 12284 2730 12312 2758
rect 12336 2730 12364 2758
rect 11718 2702 11746 2730
rect 22232 2730 22260 2758
rect 22284 2730 22312 2758
rect 22336 2730 22364 2758
rect 10598 2590 10626 2618
rect 14966 2534 14994 2562
rect 18662 2422 18690 2450
rect 1902 2338 1930 2366
rect 1954 2338 1982 2366
rect 2006 2338 2034 2366
rect 11902 2338 11930 2366
rect 11954 2338 11982 2366
rect 12006 2338 12034 2366
rect 21902 2338 21930 2366
rect 21954 2338 21982 2366
rect 22006 2338 22034 2366
rect 13230 2254 13258 2282
rect 16310 2198 16338 2226
rect 19110 2198 19138 2226
rect 12726 2030 12754 2058
rect 2232 1946 2260 1974
rect 2284 1946 2312 1974
rect 2336 1946 2364 1974
rect 12232 1946 12260 1974
rect 12284 1946 12312 1974
rect 12336 1946 12364 1974
rect 22232 1946 22260 1974
rect 22284 1946 22312 1974
rect 22336 1946 22364 1974
rect 12726 1806 12754 1834
rect 13286 1806 13314 1834
rect 11718 1694 11746 1722
rect 13510 1582 13538 1610
rect 1902 1554 1930 1582
rect 1954 1554 1982 1582
rect 2006 1554 2034 1582
rect 11902 1554 11930 1582
rect 11954 1554 11982 1582
rect 12006 1554 12034 1582
rect 21902 1554 21930 1582
rect 21954 1554 21982 1582
rect 22006 1554 22034 1582
rect 19110 1414 19138 1442
rect 12726 1358 12754 1386
rect 12502 1302 12530 1330
rect 2232 1162 2260 1190
rect 2284 1162 2312 1190
rect 2336 1162 2364 1190
rect 12232 1162 12260 1190
rect 12284 1162 12312 1190
rect 12336 1162 12364 1190
rect 22232 1162 22260 1190
rect 22284 1162 22312 1190
rect 22336 1162 22364 1190
rect 18662 1134 18690 1162
rect 13118 1078 13146 1106
rect 12446 854 12474 882
rect 1902 770 1930 798
rect 1954 770 1982 798
rect 2006 770 2034 798
rect 11902 770 11930 798
rect 11954 770 11982 798
rect 12006 770 12034 798
rect 21902 770 21930 798
rect 21954 770 21982 798
rect 22006 770 22034 798
rect 12502 742 12530 770
rect 13118 686 13146 714
rect 11270 630 11298 658
rect 12446 630 12474 658
rect 16590 630 16618 658
rect 12502 574 12530 602
rect 12446 518 12474 546
rect 11270 462 11298 490
rect 2232 378 2260 406
rect 2284 378 2312 406
rect 2336 378 2364 406
rect 12232 378 12260 406
rect 12284 378 12312 406
rect 12336 378 12364 406
rect 22232 378 22260 406
rect 22284 378 22312 406
rect 22336 378 22364 406
rect 12446 350 12474 378
<< metal4 >>
rect 1888 6286 2048 7112
rect 1888 6258 1902 6286
rect 1930 6258 1954 6286
rect 1982 6258 2006 6286
rect 2034 6258 2048 6286
rect 1888 5502 2048 6258
rect 1888 5474 1902 5502
rect 1930 5474 1954 5502
rect 1982 5474 2006 5502
rect 2034 5474 2048 5502
rect 1888 4718 2048 5474
rect 1888 4690 1902 4718
rect 1930 4690 1954 4718
rect 1982 4690 2006 4718
rect 2034 4690 2048 4718
rect 1888 3934 2048 4690
rect 1888 3906 1902 3934
rect 1930 3906 1954 3934
rect 1982 3906 2006 3934
rect 2034 3906 2048 3934
rect 1888 3150 2048 3906
rect 1888 3122 1902 3150
rect 1930 3122 1954 3150
rect 1982 3122 2006 3150
rect 2034 3122 2048 3150
rect 1888 2366 2048 3122
rect 1888 2338 1902 2366
rect 1930 2338 1954 2366
rect 1982 2338 2006 2366
rect 2034 2338 2048 2366
rect 1888 1582 2048 2338
rect 1888 1554 1902 1582
rect 1930 1554 1954 1582
rect 1982 1554 2006 1582
rect 2034 1554 2048 1582
rect 1888 798 2048 1554
rect 1888 770 1902 798
rect 1930 770 1954 798
rect 1982 770 2006 798
rect 2034 770 2048 798
rect 1888 0 2048 770
rect 2218 6678 2378 7112
rect 2218 6650 2232 6678
rect 2260 6650 2284 6678
rect 2312 6650 2336 6678
rect 2364 6650 2378 6678
rect 2218 5894 2378 6650
rect 2218 5866 2232 5894
rect 2260 5866 2284 5894
rect 2312 5866 2336 5894
rect 2364 5866 2378 5894
rect 2218 5110 2378 5866
rect 11888 6286 12048 7112
rect 11888 6258 11902 6286
rect 11930 6258 11954 6286
rect 11982 6258 12006 6286
rect 12034 6258 12048 6286
rect 9030 5810 9058 5815
rect 9030 5586 9058 5782
rect 9030 5553 9058 5558
rect 2218 5082 2232 5110
rect 2260 5082 2284 5110
rect 2312 5082 2336 5110
rect 2364 5082 2378 5110
rect 2218 4326 2378 5082
rect 2218 4298 2232 4326
rect 2260 4298 2284 4326
rect 2312 4298 2336 4326
rect 2364 4298 2378 4326
rect 2218 3542 2378 4298
rect 11888 5502 12048 6258
rect 11888 5474 11902 5502
rect 11930 5474 11954 5502
rect 11982 5474 12006 5502
rect 12034 5474 12048 5502
rect 11888 4718 12048 5474
rect 11888 4690 11902 4718
rect 11930 4690 11954 4718
rect 11982 4690 12006 4718
rect 12034 4690 12048 4718
rect 11888 3934 12048 4690
rect 11888 3906 11902 3934
rect 11930 3906 11954 3934
rect 11982 3906 12006 3934
rect 12034 3906 12048 3934
rect 2218 3514 2232 3542
rect 2260 3514 2284 3542
rect 2312 3514 2336 3542
rect 2364 3514 2378 3542
rect 2218 2758 2378 3514
rect 10486 3570 10514 3575
rect 10486 3346 10514 3542
rect 10486 3313 10514 3318
rect 11888 3150 12048 3906
rect 11888 3122 11902 3150
rect 11930 3122 11954 3150
rect 11982 3122 12006 3150
rect 12034 3122 12048 3150
rect 2218 2730 2232 2758
rect 2260 2730 2284 2758
rect 2312 2730 2336 2758
rect 2364 2730 2378 2758
rect 2218 1974 2378 2730
rect 10598 2786 10626 2791
rect 10598 2618 10626 2758
rect 10598 2585 10626 2590
rect 11718 2730 11746 2735
rect 2218 1946 2232 1974
rect 2260 1946 2284 1974
rect 2312 1946 2336 1974
rect 2364 1946 2378 1974
rect 2218 1190 2378 1946
rect 11718 1722 11746 2702
rect 11718 1689 11746 1694
rect 11888 2366 12048 3122
rect 11888 2338 11902 2366
rect 11930 2338 11954 2366
rect 11982 2338 12006 2366
rect 12034 2338 12048 2366
rect 2218 1162 2232 1190
rect 2260 1162 2284 1190
rect 2312 1162 2336 1190
rect 2364 1162 2378 1190
rect 2218 406 2378 1162
rect 11888 1582 12048 2338
rect 11888 1554 11902 1582
rect 11930 1554 11954 1582
rect 11982 1554 12006 1582
rect 12034 1554 12048 1582
rect 11888 798 12048 1554
rect 11888 770 11902 798
rect 11930 770 11954 798
rect 11982 770 12006 798
rect 12034 770 12048 798
rect 11270 658 11298 663
rect 11270 490 11298 630
rect 11270 457 11298 462
rect 2218 378 2232 406
rect 2260 378 2284 406
rect 2312 378 2336 406
rect 2364 378 2378 406
rect 2218 0 2378 378
rect 11888 0 12048 770
rect 12218 6678 12378 7112
rect 12218 6650 12232 6678
rect 12260 6650 12284 6678
rect 12312 6650 12336 6678
rect 12364 6650 12378 6678
rect 12218 5894 12378 6650
rect 21888 6286 22048 7112
rect 21888 6258 21902 6286
rect 21930 6258 21954 6286
rect 21982 6258 22006 6286
rect 22034 6258 22048 6286
rect 12218 5866 12232 5894
rect 12260 5866 12284 5894
rect 12312 5866 12336 5894
rect 12364 5866 12378 5894
rect 12218 5110 12378 5866
rect 13342 6202 13370 6207
rect 12502 5362 12866 5369
rect 12502 5341 12838 5362
rect 12502 5306 12530 5341
rect 12838 5329 12866 5334
rect 12502 5273 12530 5278
rect 12218 5082 12232 5110
rect 12260 5082 12284 5110
rect 12312 5082 12336 5110
rect 12364 5082 12378 5110
rect 12218 4326 12378 5082
rect 13342 4858 13370 6174
rect 16310 5978 16338 5983
rect 13342 4825 13370 4830
rect 13454 4858 13482 4863
rect 13454 4829 13482 4830
rect 13398 4801 13482 4829
rect 13286 4746 13314 4751
rect 13398 4739 13426 4801
rect 13314 4718 13426 4739
rect 13286 4711 13426 4718
rect 14966 4522 14994 4527
rect 14966 4469 14994 4494
rect 14966 4441 15050 4469
rect 12218 4298 12232 4326
rect 12260 4298 12284 4326
rect 12312 4298 12336 4326
rect 12364 4298 12378 4326
rect 12218 3542 12378 4298
rect 15022 4298 15050 4441
rect 15022 4265 15050 4270
rect 14182 3962 14210 3967
rect 12218 3514 12232 3542
rect 12260 3514 12284 3542
rect 12312 3514 12336 3542
rect 12364 3514 12378 3542
rect 12218 2758 12378 3514
rect 13510 3906 13538 3911
rect 13006 3234 13034 3239
rect 13006 2898 13034 3206
rect 13006 2865 13034 2870
rect 12218 2730 12232 2758
rect 12260 2730 12284 2758
rect 12312 2730 12336 2758
rect 12364 2730 12378 2758
rect 12218 1974 12378 2730
rect 13230 2282 13258 2287
rect 13230 2219 13258 2254
rect 13230 2191 13314 2219
rect 12218 1946 12232 1974
rect 12260 1946 12284 1974
rect 12312 1946 12336 1974
rect 12364 1946 12378 1974
rect 12218 1190 12378 1946
rect 12726 2058 12754 2063
rect 12726 1834 12754 2030
rect 12726 1801 12754 1806
rect 13286 1834 13314 2191
rect 13286 1801 13314 1806
rect 13510 1610 13538 3878
rect 14182 3402 14210 3934
rect 16142 3850 16170 3855
rect 16170 3822 16226 3839
rect 16142 3811 16226 3822
rect 16198 3570 16226 3811
rect 16198 3537 16226 3542
rect 14182 3369 14210 3374
rect 14966 2954 14994 2959
rect 14966 2562 14994 2926
rect 14966 2529 14994 2534
rect 16310 2226 16338 5950
rect 19222 5978 19250 5983
rect 19222 5810 19250 5950
rect 19222 5777 19250 5782
rect 21888 5502 22048 6258
rect 21888 5474 21902 5502
rect 21930 5474 21954 5502
rect 21982 5474 22006 5502
rect 22034 5474 22048 5502
rect 16310 2193 16338 2198
rect 16590 4970 16618 4975
rect 13510 1577 13538 1582
rect 12726 1386 12754 1391
rect 12502 1330 12530 1335
rect 12726 1319 12754 1358
rect 12530 1302 12754 1319
rect 12502 1291 12754 1302
rect 12218 1162 12232 1190
rect 12260 1162 12284 1190
rect 12312 1162 12336 1190
rect 12364 1162 12378 1190
rect 12218 406 12378 1162
rect 13118 1106 13146 1111
rect 12446 882 12474 887
rect 12446 658 12474 854
rect 12446 625 12474 630
rect 12502 770 12530 775
rect 12502 602 12530 742
rect 13118 714 13146 1078
rect 13118 681 13146 686
rect 16590 658 16618 4942
rect 21888 4718 22048 5474
rect 21888 4690 21902 4718
rect 21930 4690 21954 4718
rect 21982 4690 22006 4718
rect 22034 4690 22048 4718
rect 21888 3934 22048 4690
rect 16982 3906 17010 3911
rect 16982 3682 17010 3878
rect 16982 3649 17010 3654
rect 21888 3906 21902 3934
rect 21930 3906 21954 3934
rect 21982 3906 22006 3934
rect 22034 3906 22048 3934
rect 21888 3150 22048 3906
rect 21888 3122 21902 3150
rect 21930 3122 21954 3150
rect 21982 3122 22006 3150
rect 22034 3122 22048 3150
rect 18662 2450 18690 2455
rect 18662 1162 18690 2422
rect 21888 2366 22048 3122
rect 21888 2338 21902 2366
rect 21930 2338 21954 2366
rect 21982 2338 22006 2366
rect 22034 2338 22048 2366
rect 19110 2226 19138 2231
rect 19110 1442 19138 2198
rect 19110 1409 19138 1414
rect 21888 1582 22048 2338
rect 21888 1554 21902 1582
rect 21930 1554 21954 1582
rect 21982 1554 22006 1582
rect 22034 1554 22048 1582
rect 18662 1129 18690 1134
rect 16590 625 16618 630
rect 21888 798 22048 1554
rect 21888 770 21902 798
rect 21930 770 21954 798
rect 21982 770 22006 798
rect 22034 770 22048 798
rect 12502 569 12530 574
rect 12218 378 12232 406
rect 12260 378 12284 406
rect 12312 378 12336 406
rect 12364 378 12378 406
rect 12218 0 12378 378
rect 12446 546 12474 551
rect 12446 378 12474 518
rect 12446 345 12474 350
rect 21888 0 22048 770
rect 22218 6678 22378 7112
rect 22218 6650 22232 6678
rect 22260 6650 22284 6678
rect 22312 6650 22336 6678
rect 22364 6650 22378 6678
rect 22218 5894 22378 6650
rect 22218 5866 22232 5894
rect 22260 5866 22284 5894
rect 22312 5866 22336 5894
rect 22364 5866 22378 5894
rect 22218 5110 22378 5866
rect 22218 5082 22232 5110
rect 22260 5082 22284 5110
rect 22312 5082 22336 5110
rect 22364 5082 22378 5110
rect 22218 4326 22378 5082
rect 22218 4298 22232 4326
rect 22260 4298 22284 4326
rect 22312 4298 22336 4326
rect 22364 4298 22378 4326
rect 22218 3542 22378 4298
rect 22218 3514 22232 3542
rect 22260 3514 22284 3542
rect 22312 3514 22336 3542
rect 22364 3514 22378 3542
rect 22218 2758 22378 3514
rect 22218 2730 22232 2758
rect 22260 2730 22284 2758
rect 22312 2730 22336 2758
rect 22364 2730 22378 2758
rect 22218 1974 22378 2730
rect 22218 1946 22232 1974
rect 22260 1946 22284 1974
rect 22312 1946 22336 1974
rect 22364 1946 22378 1974
rect 22218 1190 22378 1946
rect 22218 1162 22232 1190
rect 22260 1162 22284 1190
rect 22312 1162 22336 1190
rect 22364 1162 22378 1190
rect 22218 406 22378 1162
rect 22218 378 22232 406
rect 22260 378 22284 406
rect 22312 378 22336 406
rect 22364 378 22378 406
rect 22218 0 22378 378
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _000_
timestamp 1486834041
transform 1 0 4872 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _001_
timestamp 1486834041
transform 1 0 5208 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _002_
timestamp 1486834041
transform 1 0 23408 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _003_
timestamp 1486834041
transform 1 0 23016 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _004_
timestamp 1486834041
transform 1 0 5320 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _005_
timestamp 1486834041
transform 1 0 23408 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _006_
timestamp 1486834041
transform 1 0 22400 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _007_
timestamp 1486834041
transform 1 0 22120 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _008_
timestamp 1486834041
transform 1 0 23072 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _009_
timestamp 1486834041
transform 1 0 1400 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _010_
timestamp 1486834041
transform 1 0 23744 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _011_
timestamp 1486834041
transform 1 0 25200 0 1 392
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _012_
timestamp 1486834041
transform 1 0 24136 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _013_
timestamp 1486834041
transform 1 0 2128 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _014_
timestamp 1486834041
transform 1 0 2408 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _015_
timestamp 1486834041
transform 1 0 1848 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _016_
timestamp 1486834041
transform 1 0 2520 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _017_
timestamp 1486834041
transform 1 0 24248 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _018_
timestamp 1486834041
transform 1 0 3416 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _019_
timestamp 1486834041
transform 1 0 23184 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _020_
timestamp 1486834041
transform 1 0 22400 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _021_
timestamp 1486834041
transform 1 0 5208 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _022_
timestamp 1486834041
transform 1 0 23800 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _023_
timestamp 1486834041
transform 1 0 4928 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _024_
timestamp 1486834041
transform 1 0 24696 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _025_
timestamp 1486834041
transform 1 0 3416 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _026_
timestamp 1486834041
transform 1 0 23800 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _027_
timestamp 1486834041
transform 1 0 23408 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _028_
timestamp 1486834041
transform 1 0 22624 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _029_
timestamp 1486834041
transform 1 0 23016 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _030_
timestamp 1486834041
transform 1 0 1008 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _031_
timestamp 1486834041
transform 1 0 25200 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _032_
timestamp 1486834041
transform -1 0 15624 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _033_
timestamp 1486834041
transform -1 0 15512 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _034_
timestamp 1486834041
transform -1 0 7896 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _035_
timestamp 1486834041
transform -1 0 9184 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _036_
timestamp 1486834041
transform -1 0 16576 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _037_
timestamp 1486834041
transform -1 0 16968 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _038_
timestamp 1486834041
transform -1 0 17976 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _039_
timestamp 1486834041
transform -1 0 11536 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _040_
timestamp 1486834041
transform -1 0 12824 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _041_
timestamp 1486834041
transform -1 0 13720 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _042_
timestamp 1486834041
transform -1 0 15176 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _043_
timestamp 1486834041
transform -1 0 17416 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _044_
timestamp 1486834041
transform -1 0 19096 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _045_
timestamp 1486834041
transform -1 0 19432 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _046_
timestamp 1486834041
transform -1 0 19152 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _047_
timestamp 1486834041
transform 1 0 20496 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _048_
timestamp 1486834041
transform -1 0 19320 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _049_
timestamp 1486834041
transform 1 0 20944 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _050_
timestamp 1486834041
transform 1 0 22736 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _051_
timestamp 1486834041
transform 1 0 22008 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _052_
timestamp 1486834041
transform -1 0 1176 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _053_
timestamp 1486834041
transform -1 0 1176 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _054_
timestamp 1486834041
transform -1 0 1176 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _055_
timestamp 1486834041
transform -1 0 1344 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _056_
timestamp 1486834041
transform 1 0 8288 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _057_
timestamp 1486834041
transform -1 0 6776 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _058_
timestamp 1486834041
transform -1 0 6216 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _059_
timestamp 1486834041
transform -1 0 5992 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _060_
timestamp 1486834041
transform -1 0 4592 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _061_
timestamp 1486834041
transform -1 0 4256 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _062_
timestamp 1486834041
transform -1 0 3248 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _063_
timestamp 1486834041
transform -1 0 2520 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _064_
timestamp 1486834041
transform 1 0 13552 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _065_
timestamp 1486834041
transform 1 0 12712 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _066_
timestamp 1486834041
transform 1 0 9128 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _067_
timestamp 1486834041
transform 1 0 9576 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _068_
timestamp 1486834041
transform 1 0 7728 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _069_
timestamp 1486834041
transform 1 0 7728 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _070_
timestamp 1486834041
transform -1 0 7448 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _071_
timestamp 1486834041
transform -1 0 6776 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _072_
timestamp 1486834041
transform 1 0 12208 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _073_
timestamp 1486834041
transform 1 0 11648 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _074_
timestamp 1486834041
transform 1 0 10920 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _075_
timestamp 1486834041
transform 1 0 11480 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _076_
timestamp 1486834041
transform 1 0 15512 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _077_
timestamp 1486834041
transform 1 0 15008 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _078_
timestamp 1486834041
transform 1 0 11256 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _079_
timestamp 1486834041
transform 1 0 10304 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _080_
timestamp 1486834041
transform 1 0 9016 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _081_
timestamp 1486834041
transform 1 0 8848 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _082_
timestamp 1486834041
transform 1 0 8680 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _083_
timestamp 1486834041
transform 1 0 15232 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _084_
timestamp 1486834041
transform 1 0 15960 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _085_
timestamp 1486834041
transform 1 0 17304 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _086_
timestamp 1486834041
transform 1 0 19264 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _087_
timestamp 1486834041
transform 1 0 17528 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _088_
timestamp 1486834041
transform 1 0 14728 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _089_
timestamp 1486834041
transform 1 0 12376 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _090_
timestamp 1486834041
transform 1 0 16800 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _091_
timestamp 1486834041
transform 1 0 14168 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _092_
timestamp 1486834041
transform 1 0 12488 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _093_
timestamp 1486834041
transform 1 0 18088 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _094_
timestamp 1486834041
transform 1 0 18536 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _095_
timestamp 1486834041
transform 1 0 18984 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _096_
timestamp 1486834041
transform 1 0 19656 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _097_
timestamp 1486834041
transform 1 0 20048 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _098_
timestamp 1486834041
transform 1 0 20440 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _099_
timestamp 1486834041
transform 1 0 21000 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _100_
timestamp 1486834041
transform 1 0 21224 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _101_
timestamp 1486834041
transform 1 0 22064 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _102_
timestamp 1486834041
transform 1 0 23520 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _103_
timestamp 1486834041
transform 1 0 24584 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _104_
timestamp 1486834041
transform -1 0 16352 0 1 5880
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2
timestamp 1486834041
transform 1 0 448 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36
timestamp 1486834041
transform 1 0 2352 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_70
timestamp 1486834041
transform 1 0 4256 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_104
timestamp 1486834041
transform 1 0 6160 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_138
timestamp 1486834041
transform 1 0 8064 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_172
timestamp 1486834041
transform 1 0 9968 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_206
timestamp 1486834041
transform 1 0 11872 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_268
timestamp 1486834041
transform 1 0 15344 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_302
timestamp 1486834041
transform 1 0 17248 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_336
timestamp 1486834041
transform 1 0 19152 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_370
timestamp 1486834041
transform 1 0 21056 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_376
timestamp 1486834041
transform 1 0 21392 0 1 392
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_410
timestamp 1486834041
transform 1 0 23296 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_452
timestamp 1486834041
transform 1 0 25648 0 1 392
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_456
timestamp 1486834041
transform 1 0 25872 0 1 392
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_2
timestamp 1486834041
transform 1 0 448 0 -1 1176
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_18
timestamp 1486834041
transform 1 0 1344 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_26
timestamp 1486834041
transform 1 0 1792 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_30
timestamp 1486834041
transform 1 0 2016 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_40
timestamp 1486834041
transform 1 0 2576 0 -1 1176
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_56
timestamp 1486834041
transform 1 0 3472 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_64
timestamp 1486834041
transform 1 0 3920 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_68
timestamp 1486834041
transform 1 0 4144 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_72
timestamp 1486834041
transform 1 0 4368 0 -1 1176
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_88
timestamp 1486834041
transform 1 0 5264 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_92
timestamp 1486834041
transform 1 0 5488 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_101
timestamp 1486834041
transform 1 0 5992 0 -1 1176
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_133
timestamp 1486834041
transform 1 0 7784 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_137
timestamp 1486834041
transform 1 0 8008 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_139
timestamp 1486834041
transform 1 0 8120 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_142
timestamp 1486834041
transform 1 0 8288 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_150
timestamp 1486834041
transform 1 0 8736 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_154
timestamp 1486834041
transform 1 0 8960 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_163
timestamp 1486834041
transform 1 0 9464 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_171
timestamp 1486834041
transform 1 0 9912 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_175
timestamp 1486834041
transform 1 0 10136 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_177
timestamp 1486834041
transform 1 0 10248 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_186
timestamp 1486834041
transform 1 0 10752 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_194
timestamp 1486834041
transform 1 0 11200 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_212
timestamp 1486834041
transform 1 0 12208 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_214
timestamp 1486834041
transform 1 0 12320 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_279
timestamp 1486834041
transform 1 0 15960 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_346
timestamp 1486834041
transform 1 0 19712 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_352
timestamp 1486834041
transform 1 0 20048 0 -1 1176
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_384
timestamp 1486834041
transform 1 0 21840 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_392
timestamp 1486834041
transform 1 0 22288 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_402
timestamp 1486834041
transform 1 0 22848 0 -1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_410
timestamp 1486834041
transform 1 0 23296 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_422
timestamp 1486834041
transform 1 0 23968 0 -1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_426
timestamp 1486834041
transform 1 0 24192 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_428
timestamp 1486834041
transform 1 0 24304 0 -1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_2
timestamp 1486834041
transform 1 0 448 0 1 1176
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_18
timestamp 1486834041
transform 1 0 1344 0 1 1176
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_27
timestamp 1486834041
transform 1 0 1848 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_37
timestamp 1486834041
transform 1 0 2408 0 1 1176
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_69
timestamp 1486834041
transform 1 0 4200 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_77
timestamp 1486834041
transform 1 0 4648 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_97
timestamp 1486834041
transform 1 0 5768 0 1 1176
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_107
timestamp 1486834041
transform 1 0 6328 0 1 1176
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_171
timestamp 1486834041
transform 1 0 9912 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_177
timestamp 1486834041
transform 1 0 10248 0 1 1176
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_193
timestamp 1486834041
transform 1 0 11144 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_311
timestamp 1486834041
transform 1 0 17752 0 1 1176
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_353
timestamp 1486834041
transform 1 0 20104 0 1 1176
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_387
timestamp 1486834041
transform 1 0 22008 0 1 1176
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_403
timestamp 1486834041
transform 1 0 22904 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_2
timestamp 1486834041
transform 1 0 448 0 -1 1960
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_66
timestamp 1486834041
transform 1 0 4032 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_72
timestamp 1486834041
transform 1 0 4368 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_80
timestamp 1486834041
transform 1 0 4816 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_84
timestamp 1486834041
transform 1 0 5040 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_86
timestamp 1486834041
transform 1 0 5152 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_95
timestamp 1486834041
transform 1 0 5656 0 -1 1960
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_127
timestamp 1486834041
transform 1 0 7448 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_135
timestamp 1486834041
transform 1 0 7896 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_139
timestamp 1486834041
transform 1 0 8120 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_142
timestamp 1486834041
transform 1 0 8288 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_150
timestamp 1486834041
transform 1 0 8736 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_160
timestamp 1486834041
transform 1 0 9296 0 -1 1960
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_192
timestamp 1486834041
transform 1 0 11088 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_212
timestamp 1486834041
transform 1 0 12208 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_216
timestamp 1486834041
transform 1 0 12432 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_239
timestamp 1486834041
transform 1 0 13720 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_243
timestamp 1486834041
transform 1 0 13944 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_273
timestamp 1486834041
transform 1 0 15624 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_277
timestamp 1486834041
transform 1 0 15848 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_279
timestamp 1486834041
transform 1 0 15960 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_338
timestamp 1486834041
transform 1 0 19264 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_346
timestamp 1486834041
transform 1 0 19712 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_352
timestamp 1486834041
transform 1 0 20048 0 -1 1960
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_384
timestamp 1486834041
transform 1 0 21840 0 -1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_400
timestamp 1486834041
transform 1 0 22736 0 -1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_408
timestamp 1486834041
transform 1 0 23184 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_422
timestamp 1486834041
transform 1 0 23968 0 -1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_426
timestamp 1486834041
transform 1 0 24192 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_428
timestamp 1486834041
transform 1 0 24304 0 -1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_2
timestamp 1486834041
transform 1 0 448 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_18
timestamp 1486834041
transform 1 0 1344 0 1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1486834041
transform 1 0 2240 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_37
timestamp 1486834041
transform 1 0 2408 0 1 1960
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_101
timestamp 1486834041
transform 1 0 5992 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_115
timestamp 1486834041
transform 1 0 6776 0 1 1960
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_147
timestamp 1486834041
transform 1 0 8568 0 1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_163
timestamp 1486834041
transform 1 0 9464 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_171
timestamp 1486834041
transform 1 0 9912 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_177
timestamp 1486834041
transform 1 0 10248 0 1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_193
timestamp 1486834041
transform 1 0 11144 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_197
timestamp 1486834041
transform 1 0 11368 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_235
timestamp 1486834041
transform 1 0 13496 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_243
timestamp 1486834041
transform 1 0 13944 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_311
timestamp 1486834041
transform 1 0 17752 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_339
timestamp 1486834041
transform 1 0 19320 0 1 1960
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_371
timestamp 1486834041
transform 1 0 21112 0 1 1960
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_379
timestamp 1486834041
transform 1 0 21560 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_383
timestamp 1486834041
transform 1 0 21784 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_387
timestamp 1486834041
transform 1 0 22008 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_397
timestamp 1486834041
transform 1 0 22568 0 1 1960
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_413
timestamp 1486834041
transform 1 0 23464 0 1 1960
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_417
timestamp 1486834041
transform 1 0 23688 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_426
timestamp 1486834041
transform 1 0 24192 0 1 1960
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_2
timestamp 1486834041
transform 1 0 448 0 -1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_18
timestamp 1486834041
transform 1 0 1344 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_26
timestamp 1486834041
transform 1 0 1792 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_30
timestamp 1486834041
transform 1 0 2016 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_39
timestamp 1486834041
transform 1 0 2520 0 -1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_55
timestamp 1486834041
transform 1 0 3416 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_63
timestamp 1486834041
transform 1 0 3864 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_67
timestamp 1486834041
transform 1 0 4088 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_69
timestamp 1486834041
transform 1 0 4200 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_72
timestamp 1486834041
transform 1 0 4368 0 -1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_104
timestamp 1486834041
transform 1 0 6160 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_112
timestamp 1486834041
transform 1 0 6608 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_116
timestamp 1486834041
transform 1 0 6832 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_118
timestamp 1486834041
transform 1 0 6944 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_127
timestamp 1486834041
transform 1 0 7448 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_135
timestamp 1486834041
transform 1 0 7896 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_139
timestamp 1486834041
transform 1 0 8120 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_142
timestamp 1486834041
transform 1 0 8288 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_146
timestamp 1486834041
transform 1 0 8512 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_148
timestamp 1486834041
transform 1 0 8624 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_157
timestamp 1486834041
transform 1 0 9128 0 -1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_189
timestamp 1486834041
transform 1 0 10920 0 -1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_205
timestamp 1486834041
transform 1 0 11816 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_209
timestamp 1486834041
transform 1 0 12040 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_212
timestamp 1486834041
transform 1 0 12208 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_220
timestamp 1486834041
transform 1 0 12656 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_229
timestamp 1486834041
transform 1 0 13160 0 -1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_245
timestamp 1486834041
transform 1 0 14056 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_253
timestamp 1486834041
transform 1 0 14504 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_279
timestamp 1486834041
transform 1 0 15960 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_338
timestamp 1486834041
transform 1 0 19264 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_346
timestamp 1486834041
transform 1 0 19712 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_360
timestamp 1486834041
transform 1 0 20496 0 -1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_392
timestamp 1486834041
transform 1 0 22288 0 -1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_408
timestamp 1486834041
transform 1 0 23184 0 -1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_416
timestamp 1486834041
transform 1 0 23632 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_422
timestamp 1486834041
transform 1 0 23968 0 -1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_426
timestamp 1486834041
transform 1 0 24192 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_428
timestamp 1486834041
transform 1 0 24304 0 -1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_2
timestamp 1486834041
transform 1 0 448 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_6
timestamp 1486834041
transform 1 0 672 0 1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_15
timestamp 1486834041
transform 1 0 1176 0 1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_31
timestamp 1486834041
transform 1 0 2072 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_45
timestamp 1486834041
transform 1 0 2856 0 1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_77
timestamp 1486834041
transform 1 0 4648 0 1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_93
timestamp 1486834041
transform 1 0 5544 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_115
timestamp 1486834041
transform 1 0 6776 0 1 2744
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_147
timestamp 1486834041
transform 1 0 8568 0 1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_163
timestamp 1486834041
transform 1 0 9464 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_171
timestamp 1486834041
transform 1 0 9912 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_177
timestamp 1486834041
transform 1 0 10248 0 1 2744
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_241
timestamp 1486834041
transform 1 0 13832 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_247
timestamp 1486834041
transform 1 0 14168 0 1 2744
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_255
timestamp 1486834041
transform 1 0 14616 0 1 2744
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_259
timestamp 1486834041
transform 1 0 14840 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_261
timestamp 1486834041
transform 1 0 14952 0 1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_270
timestamp 1486834041
transform 1 0 15456 0 1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_341
timestamp 1486834041
transform 1 0 19432 0 1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_357
timestamp 1486834041
transform 1 0 20328 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_367
timestamp 1486834041
transform 1 0 20888 0 1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_383
timestamp 1486834041
transform 1 0 21784 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_387
timestamp 1486834041
transform 1 0 22008 0 1 2744
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_403
timestamp 1486834041
transform 1 0 22904 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_405
timestamp 1486834041
transform 1 0 23016 0 1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_422
timestamp 1486834041
transform 1 0 23968 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_424
timestamp 1486834041
transform 1 0 24080 0 1 2744
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_2
timestamp 1486834041
transform 1 0 448 0 -1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_34
timestamp 1486834041
transform 1 0 2240 0 -1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_50
timestamp 1486834041
transform 1 0 3136 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_58
timestamp 1486834041
transform 1 0 3584 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_72
timestamp 1486834041
transform 1 0 4368 0 -1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_104
timestamp 1486834041
transform 1 0 6160 0 -1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_120
timestamp 1486834041
transform 1 0 7056 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_128
timestamp 1486834041
transform 1 0 7504 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_150
timestamp 1486834041
transform 1 0 8736 0 -1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_182
timestamp 1486834041
transform 1 0 10528 0 -1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_198
timestamp 1486834041
transform 1 0 11424 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_206
timestamp 1486834041
transform 1 0 11872 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_212
timestamp 1486834041
transform 1 0 12208 0 -1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_228
timestamp 1486834041
transform 1 0 13104 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_244
timestamp 1486834041
transform 1 0 14000 0 -1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_260
timestamp 1486834041
transform 1 0 14896 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_264
timestamp 1486834041
transform 1 0 15120 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_274
timestamp 1486834041
transform 1 0 15680 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_278
timestamp 1486834041
transform 1 0 15904 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_282
timestamp 1486834041
transform 1 0 16128 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_290
timestamp 1486834041
transform 1 0 16576 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_302
timestamp 1486834041
transform 1 0 17248 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_306
timestamp 1486834041
transform 1 0 17472 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_315
timestamp 1486834041
transform 1 0 17976 0 -1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_347
timestamp 1486834041
transform 1 0 19768 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_349
timestamp 1486834041
transform 1 0 19880 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_352
timestamp 1486834041
transform 1 0 20048 0 -1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_368
timestamp 1486834041
transform 1 0 20944 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_377
timestamp 1486834041
transform 1 0 21448 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_385
timestamp 1486834041
transform 1 0 21896 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_387
timestamp 1486834041
transform 1 0 22008 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_396
timestamp 1486834041
transform 1 0 22512 0 -1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_412
timestamp 1486834041
transform 1 0 23408 0 -1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_422
timestamp 1486834041
transform 1 0 23968 0 -1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_426
timestamp 1486834041
transform 1 0 24192 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_428
timestamp 1486834041
transform 1 0 24304 0 -1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_2
timestamp 1486834041
transform 1 0 448 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_6
timestamp 1486834041
transform 1 0 672 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_15
timestamp 1486834041
transform 1 0 1176 0 1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_31
timestamp 1486834041
transform 1 0 2072 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_37
timestamp 1486834041
transform 1 0 2408 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_41
timestamp 1486834041
transform 1 0 2632 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_43
timestamp 1486834041
transform 1 0 2744 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_52
timestamp 1486834041
transform 1 0 3248 0 1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_76
timestamp 1486834041
transform 1 0 4592 0 1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_92
timestamp 1486834041
transform 1 0 5488 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_100
timestamp 1486834041
transform 1 0 5936 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_104
timestamp 1486834041
transform 1 0 6160 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_107
timestamp 1486834041
transform 1 0 6328 0 1 3528
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_171
timestamp 1486834041
transform 1 0 9912 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_177
timestamp 1486834041
transform 1 0 10248 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_185
timestamp 1486834041
transform 1 0 10696 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_197
timestamp 1486834041
transform 1 0 11368 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_205
timestamp 1486834041
transform 1 0 11816 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_209
timestamp 1486834041
transform 1 0 12040 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_211
timestamp 1486834041
transform 1 0 12152 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_220
timestamp 1486834041
transform 1 0 12656 0 1 3528
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_236
timestamp 1486834041
transform 1 0 13552 0 1 3528
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_244
timestamp 1486834041
transform 1 0 14000 0 1 3528
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_247
timestamp 1486834041
transform 1 0 14168 0 1 3528
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_311
timestamp 1486834041
transform 1 0 17752 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_317
timestamp 1486834041
transform 1 0 18088 0 1 3528
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_381
timestamp 1486834041
transform 1 0 21672 0 1 3528
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_387
timestamp 1486834041
transform 1 0 22008 0 1 3528
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_2
timestamp 1486834041
transform 1 0 448 0 -1 4312
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_66
timestamp 1486834041
transform 1 0 4032 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_72
timestamp 1486834041
transform 1 0 4368 0 -1 4312
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_136
timestamp 1486834041
transform 1 0 7952 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_142
timestamp 1486834041
transform 1 0 8288 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_150
timestamp 1486834041
transform 1 0 8736 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_154
timestamp 1486834041
transform 1 0 8960 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_156
timestamp 1486834041
transform 1 0 9072 0 -1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_165
timestamp 1486834041
transform 1 0 9576 0 -1 4312
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_197
timestamp 1486834041
transform 1 0 11368 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_201
timestamp 1486834041
transform 1 0 11592 0 -1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_212
timestamp 1486834041
transform 1 0 12208 0 -1 4312
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_244
timestamp 1486834041
transform 1 0 14000 0 -1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_260
timestamp 1486834041
transform 1 0 14896 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_262
timestamp 1486834041
transform 1 0 15008 0 -1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_271
timestamp 1486834041
transform 1 0 15512 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_279
timestamp 1486834041
transform 1 0 15960 0 -1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_282
timestamp 1486834041
transform 1 0 16128 0 -1 4312
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_346
timestamp 1486834041
transform 1 0 19712 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_352
timestamp 1486834041
transform 1 0 20048 0 -1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_368
timestamp 1486834041
transform 1 0 20944 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_372
timestamp 1486834041
transform 1 0 21168 0 -1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_381
timestamp 1486834041
transform 1 0 21672 0 -1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_397
timestamp 1486834041
transform 1 0 22568 0 -1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_405
timestamp 1486834041
transform 1 0 23016 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_407
timestamp 1486834041
transform 1 0 23128 0 -1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_416
timestamp 1486834041
transform 1 0 23632 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_422
timestamp 1486834041
transform 1 0 23968 0 -1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_426
timestamp 1486834041
transform 1 0 24192 0 -1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_2
timestamp 1486834041
transform 1 0 448 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_18
timestamp 1486834041
transform 1 0 1344 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_26
timestamp 1486834041
transform 1 0 1792 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_37
timestamp 1486834041
transform 1 0 2408 0 1 4312
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_69
timestamp 1486834041
transform 1 0 4200 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_85
timestamp 1486834041
transform 1 0 5096 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_95
timestamp 1486834041
transform 1 0 5656 0 1 4312
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_103
timestamp 1486834041
transform 1 0 6104 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_107
timestamp 1486834041
transform 1 0 6328 0 1 4312
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_171
timestamp 1486834041
transform 1 0 9912 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_177
timestamp 1486834041
transform 1 0 10248 0 1 4312
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_241
timestamp 1486834041
transform 1 0 13832 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_247
timestamp 1486834041
transform 1 0 14168 0 1 4312
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_311
timestamp 1486834041
transform 1 0 17752 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_317
timestamp 1486834041
transform 1 0 18088 0 1 4312
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_381
timestamp 1486834041
transform 1 0 21672 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_387
timestamp 1486834041
transform 1 0 22008 0 1 4312
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_391
timestamp 1486834041
transform 1 0 22232 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_393
timestamp 1486834041
transform 1 0 22344 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_402
timestamp 1486834041
transform 1 0 22848 0 1 4312
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_418
timestamp 1486834041
transform 1 0 23744 0 1 4312
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_2
timestamp 1486834041
transform 1 0 448 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_6
timestamp 1486834041
transform 1 0 672 0 -1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_15
timestamp 1486834041
transform 1 0 1176 0 -1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_31
timestamp 1486834041
transform 1 0 2072 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_47
timestamp 1486834041
transform 1 0 2968 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_63
timestamp 1486834041
transform 1 0 3864 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_67
timestamp 1486834041
transform 1 0 4088 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_69
timestamp 1486834041
transform 1 0 4200 0 -1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_72
timestamp 1486834041
transform 1 0 4368 0 -1 5096
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_104
timestamp 1486834041
transform 1 0 6160 0 -1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_120
timestamp 1486834041
transform 1 0 7056 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_128
timestamp 1486834041
transform 1 0 7504 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_142
timestamp 1486834041
transform 1 0 8288 0 -1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_158
timestamp 1486834041
transform 1 0 9184 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_162
timestamp 1486834041
transform 1 0 9408 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_164
timestamp 1486834041
transform 1 0 9520 0 -1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_173
timestamp 1486834041
transform 1 0 10024 0 -1 5096
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_205
timestamp 1486834041
transform 1 0 11816 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_209
timestamp 1486834041
transform 1 0 12040 0 -1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_212
timestamp 1486834041
transform 1 0 12208 0 -1 5096
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_276
timestamp 1486834041
transform 1 0 15792 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_290
timestamp 1486834041
transform 1 0 16576 0 -1 5096
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_322
timestamp 1486834041
transform 1 0 18368 0 -1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_338
timestamp 1486834041
transform 1 0 19264 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_346
timestamp 1486834041
transform 1 0 19712 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_352
timestamp 1486834041
transform 1 0 20048 0 -1 5096
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_384
timestamp 1486834041
transform 1 0 21840 0 -1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_400
timestamp 1486834041
transform 1 0 22736 0 -1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_408
timestamp 1486834041
transform 1 0 23184 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_422
timestamp 1486834041
transform 1 0 23968 0 -1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_426
timestamp 1486834041
transform 1 0 24192 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_428
timestamp 1486834041
transform 1 0 24304 0 -1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_2
timestamp 1486834041
transform 1 0 448 0 1 5096
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1486834041
transform 1 0 2240 0 1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_37
timestamp 1486834041
transform 1 0 2408 0 1 5096
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_101
timestamp 1486834041
transform 1 0 5992 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_107
timestamp 1486834041
transform 1 0 6328 0 1 5096
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_171
timestamp 1486834041
transform 1 0 9912 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_177
timestamp 1486834041
transform 1 0 10248 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_185
timestamp 1486834041
transform 1 0 10696 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_189
timestamp 1486834041
transform 1 0 10920 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_191
timestamp 1486834041
transform 1 0 11032 0 1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_200
timestamp 1486834041
transform 1 0 11536 0 1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_216
timestamp 1486834041
transform 1 0 12432 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_224
timestamp 1486834041
transform 1 0 12880 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_228
timestamp 1486834041
transform 1 0 13104 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_230
timestamp 1486834041
transform 1 0 13216 0 1 5096
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_239
timestamp 1486834041
transform 1 0 13720 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_243
timestamp 1486834041
transform 1 0 13944 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_247
timestamp 1486834041
transform 1 0 14168 0 1 5096
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_279
timestamp 1486834041
transform 1 0 15960 0 1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_295
timestamp 1486834041
transform 1 0 16856 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_303
timestamp 1486834041
transform 1 0 17304 0 1 5096
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_317
timestamp 1486834041
transform 1 0 18088 0 1 5096
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_325
timestamp 1486834041
transform 1 0 18536 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_335
timestamp 1486834041
transform 1 0 19096 0 1 5096
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_367
timestamp 1486834041
transform 1 0 20888 0 1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_383
timestamp 1486834041
transform 1 0 21784 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_387
timestamp 1486834041
transform 1 0 22008 0 1 5096
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_403
timestamp 1486834041
transform 1 0 22904 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_2
timestamp 1486834041
transform 1 0 448 0 -1 5880
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_66
timestamp 1486834041
transform 1 0 4032 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_72
timestamp 1486834041
transform 1 0 4368 0 -1 5880
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_104
timestamp 1486834041
transform 1 0 6160 0 -1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_120
timestamp 1486834041
transform 1 0 7056 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_124
timestamp 1486834041
transform 1 0 7280 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_126
timestamp 1486834041
transform 1 0 7392 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_135
timestamp 1486834041
transform 1 0 7896 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_139
timestamp 1486834041
transform 1 0 8120 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_142
timestamp 1486834041
transform 1 0 8288 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_158
timestamp 1486834041
transform 1 0 9184 0 -1 5880
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_190
timestamp 1486834041
transform 1 0 10976 0 -1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_206
timestamp 1486834041
transform 1 0 11872 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_212
timestamp 1486834041
transform 1 0 12208 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_214
timestamp 1486834041
transform 1 0 12320 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_223
timestamp 1486834041
transform 1 0 12824 0 -1 5880
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_255
timestamp 1486834041
transform 1 0 14616 0 -1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_271
timestamp 1486834041
transform 1 0 15512 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_279
timestamp 1486834041
transform 1 0 15960 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_282
timestamp 1486834041
transform 1 0 16128 0 -1 5880
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_314
timestamp 1486834041
transform 1 0 17920 0 -1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_330
timestamp 1486834041
transform 1 0 18816 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_332
timestamp 1486834041
transform 1 0 18928 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_341
timestamp 1486834041
transform 1 0 19432 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_349
timestamp 1486834041
transform 1 0 19880 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_352
timestamp 1486834041
transform 1 0 20048 0 -1 5880
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_384
timestamp 1486834041
transform 1 0 21840 0 -1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_392
timestamp 1486834041
transform 1 0 22288 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_396
timestamp 1486834041
transform 1 0 22512 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_422
timestamp 1486834041
transform 1 0 23968 0 -1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_426
timestamp 1486834041
transform 1 0 24192 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_428
timestamp 1486834041
transform 1 0 24304 0 -1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_2
timestamp 1486834041
transform 1 0 448 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_10
timestamp 1486834041
transform 1 0 896 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_20
timestamp 1486834041
transform 1 0 1456 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_28
timestamp 1486834041
transform 1 0 1904 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_32
timestamp 1486834041
transform 1 0 2128 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1486834041
transform 1 0 2240 0 1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_37
timestamp 1486834041
transform 1 0 2408 0 1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_53
timestamp 1486834041
transform 1 0 3304 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_63
timestamp 1486834041
transform 1 0 3864 0 1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_79
timestamp 1486834041
transform 1 0 4760 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_81
timestamp 1486834041
transform 1 0 4872 0 1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_90
timestamp 1486834041
transform 1 0 5376 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_98
timestamp 1486834041
transform 1 0 5824 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_102
timestamp 1486834041
transform 1 0 6048 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_104
timestamp 1486834041
transform 1 0 6160 0 1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_107
timestamp 1486834041
transform 1 0 6328 0 1 5880
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_171
timestamp 1486834041
transform 1 0 9912 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_177
timestamp 1486834041
transform 1 0 10248 0 1 5880
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_241
timestamp 1486834041
transform 1 0 13832 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_247
timestamp 1486834041
transform 1 0 14168 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_255
timestamp 1486834041
transform 1 0 14616 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_273
timestamp 1486834041
transform 1 0 15624 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_277
timestamp 1486834041
transform 1 0 15848 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_279
timestamp 1486834041
transform 1 0 15960 0 1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_286
timestamp 1486834041
transform 1 0 16352 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_288
timestamp 1486834041
transform 1 0 16464 0 1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_305
timestamp 1486834041
transform 1 0 17416 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_313
timestamp 1486834041
transform 1 0 17864 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_317
timestamp 1486834041
transform 1 0 18088 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_325
timestamp 1486834041
transform 1 0 18536 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_327
timestamp 1486834041
transform 1 0 18648 0 1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_336
timestamp 1486834041
transform 1 0 19152 0 1 5880
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_352
timestamp 1486834041
transform 1 0 20048 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_376
timestamp 1486834041
transform 1 0 21392 0 1 5880
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_384
timestamp 1486834041
transform 1 0 21840 0 1 5880
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_395
timestamp 1486834041
transform 1 0 22456 0 1 5880
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_2
timestamp 1486834041
transform 1 0 448 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_6
timestamp 1486834041
transform 1 0 672 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_8
timestamp 1486834041
transform 1 0 784 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_15
timestamp 1486834041
transform 1 0 1176 0 -1 6664
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_31
timestamp 1486834041
transform 1 0 2072 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_33
timestamp 1486834041
transform 1 0 2184 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_50
timestamp 1486834041
transform 1 0 3136 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_52
timestamp 1486834041
transform 1 0 3248 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_67
timestamp 1486834041
transform 1 0 4088 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_70
timestamp 1486834041
transform 1 0 4256 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_74
timestamp 1486834041
transform 1 0 4480 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_89
timestamp 1486834041
transform 1 0 5320 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_97
timestamp 1486834041
transform 1 0 5768 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_101
timestamp 1486834041
transform 1 0 5992 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_118
timestamp 1486834041
transform 1 0 6944 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_133
timestamp 1486834041
transform 1 0 7784 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_135
timestamp 1486834041
transform 1 0 7896 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_138
timestamp 1486834041
transform 1 0 8064 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_140
timestamp 1486834041
transform 1 0 8176 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_155
timestamp 1486834041
transform 1 0 9016 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_172
timestamp 1486834041
transform 1 0 9968 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_180
timestamp 1486834041
transform 1 0 10416 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_184
timestamp 1486834041
transform 1 0 10640 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_199
timestamp 1486834041
transform 1 0 11480 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_203
timestamp 1486834041
transform 1 0 11704 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_206
timestamp 1486834041
transform 1 0 11872 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_221
timestamp 1486834041
transform 1 0 12712 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_223
timestamp 1486834041
transform 1 0 12824 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_240
timestamp 1486834041
transform 1 0 13776 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_248
timestamp 1486834041
transform 1 0 14224 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_250
timestamp 1486834041
transform 1 0 14336 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_265
timestamp 1486834041
transform 1 0 15176 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_269
timestamp 1486834041
transform 1 0 15400 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_271
timestamp 1486834041
transform 1 0 15512 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_288
timestamp 1486834041
transform 1 0 16464 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_308
timestamp 1486834041
transform 1 0 17584 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_316
timestamp 1486834041
transform 1 0 18032 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_331
timestamp 1486834041
transform 1 0 18872 0 -1 6664
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_339
timestamp 1486834041
transform 1 0 19320 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_356
timestamp 1486834041
transform 1 0 20272 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_376
timestamp 1486834041
transform 1 0 21392 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_380
timestamp 1486834041
transform 1 0 21616 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_382
timestamp 1486834041
transform 1 0 21728 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_397
timestamp 1486834041
transform 1 0 22568 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_399
timestamp 1486834041
transform 1 0 22680 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_424
timestamp 1486834041
transform 1 0 24080 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_426
timestamp 1486834041
transform 1 0 24192 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_441
timestamp 1486834041
transform 1 0 25032 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_452
timestamp 1486834041
transform 1 0 25648 0 -1 6664
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_456
timestamp 1486834041
transform 1 0 25872 0 -1 6664
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output1
timestamp 1486834041
transform 1 0 24248 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output2
timestamp 1486834041
transform 1 0 24360 0 -1 2744
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output3
timestamp 1486834041
transform -1 0 25816 0 1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output4
timestamp 1486834041
transform 1 0 25144 0 -1 2744
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output5
timestamp 1486834041
transform 1 0 24360 0 -1 3528
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output6
timestamp 1486834041
transform 1 0 25032 0 1 2744
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output7
timestamp 1486834041
transform 1 0 24248 0 1 3528
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output8
timestamp 1486834041
transform 1 0 25144 0 -1 3528
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output9
timestamp 1486834041
transform 1 0 25144 0 -1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output10
timestamp 1486834041
transform 1 0 25032 0 1 3528
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output11
timestamp 1486834041
transform 1 0 25032 0 1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output12
timestamp 1486834041
transform 1 0 23464 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output13
timestamp 1486834041
transform 1 0 25144 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output14
timestamp 1486834041
transform 1 0 25032 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output15
timestamp 1486834041
transform 1 0 25144 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output16
timestamp 1486834041
transform 1 0 24248 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output17
timestamp 1486834041
transform 1 0 25032 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output18
timestamp 1486834041
transform 1 0 24360 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output19
timestamp 1486834041
transform 1 0 24248 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output20
timestamp 1486834041
transform 1 0 24360 0 -1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output21
timestamp 1486834041
transform 1 0 24248 0 1 4312
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output22
timestamp 1486834041
transform 1 0 23464 0 1 5096
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output23
timestamp 1486834041
transform 1 0 23520 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output24
timestamp 1486834041
transform 1 0 23072 0 -1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output25
timestamp 1486834041
transform -1 0 23464 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output26
timestamp 1486834041
transform 1 0 24304 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output27
timestamp 1486834041
transform 1 0 24360 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output28
timestamp 1486834041
transform 1 0 25144 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output29
timestamp 1486834041
transform 1 0 24360 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output30
timestamp 1486834041
transform 1 0 25032 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output31
timestamp 1486834041
transform 1 0 24248 0 1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output32
timestamp 1486834041
transform 1 0 25144 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output33
timestamp 1486834041
transform -1 0 3136 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output34
timestamp 1486834041
transform -1 0 15176 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output35
timestamp 1486834041
transform -1 0 16464 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output36
timestamp 1486834041
transform -1 0 17472 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output37
timestamp 1486834041
transform -1 0 18872 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output38
timestamp 1486834041
transform 1 0 19488 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output39
timestamp 1486834041
transform -1 0 21280 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output40
timestamp 1486834041
transform 1 0 21784 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output41
timestamp 1486834041
transform 1 0 23296 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output42
timestamp 1486834041
transform 1 0 24248 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output43
timestamp 1486834041
transform 1 0 23464 0 1 5880
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output44
timestamp 1486834041
transform -1 0 4088 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output45
timestamp 1486834041
transform -1 0 5320 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output46
timestamp 1486834041
transform -1 0 6944 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output47
timestamp 1486834041
transform -1 0 7784 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output48
timestamp 1486834041
transform -1 0 9016 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output49
timestamp 1486834041
transform -1 0 9856 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output50
timestamp 1486834041
transform -1 0 11480 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output51
timestamp 1486834041
transform -1 0 12712 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output52
timestamp 1486834041
transform -1 0 13664 0 -1 6664
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output53
timestamp 1486834041
transform 1 0 11312 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output54
timestamp 1486834041
transform 1 0 10192 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output55
timestamp 1486834041
transform 1 0 11928 0 1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output56
timestamp 1486834041
transform 1 0 11312 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output57
timestamp 1486834041
transform 1 0 11704 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output58
timestamp 1486834041
transform 1 0 10976 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output59
timestamp 1486834041
transform 1 0 12712 0 1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output60
timestamp 1486834041
transform 1 0 12488 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output61
timestamp 1486834041
transform 1 0 12936 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output62
timestamp 1486834041
transform 1 0 12096 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output63
timestamp 1486834041
transform 1 0 12824 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output64
timestamp 1486834041
transform 1 0 13272 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output65
timestamp 1486834041
transform -1 0 13664 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output66
timestamp 1486834041
transform 1 0 13776 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output67
timestamp 1486834041
transform 1 0 13608 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output68
timestamp 1486834041
transform 1 0 14560 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output69
timestamp 1486834041
transform 1 0 14392 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output70
timestamp 1486834041
transform 1 0 14168 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output71
timestamp 1486834041
transform 1 0 14056 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output72
timestamp 1486834041
transform 1 0 15176 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output73
timestamp 1486834041
transform 1 0 15680 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output74
timestamp 1486834041
transform 1 0 16128 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output75
timestamp 1486834041
transform 1 0 16520 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output76
timestamp 1486834041
transform 1 0 17584 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output77
timestamp 1486834041
transform -1 0 16968 0 1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output78
timestamp 1486834041
transform -1 0 18480 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output79
timestamp 1486834041
transform -1 0 17696 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output80
timestamp 1486834041
transform 1 0 14952 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output81
timestamp 1486834041
transform 1 0 14840 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output82
timestamp 1486834041
transform 1 0 14616 0 1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output83
timestamp 1486834041
transform 1 0 16464 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output84
timestamp 1486834041
transform 1 0 15736 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output85
timestamp 1486834041
transform 1 0 16128 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output86
timestamp 1486834041
transform 1 0 15400 0 1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output87
timestamp 1486834041
transform 1 0 15176 0 -1 2744
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output88
timestamp 1486834041
transform 1 0 16912 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output89
timestamp 1486834041
transform 1 0 16128 0 -1 2744
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output90
timestamp 1486834041
transform -1 0 19264 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output91
timestamp 1486834041
transform -1 0 18480 0 -1 2744
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output92
timestamp 1486834041
transform -1 0 19656 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output93
timestamp 1486834041
transform -1 0 18872 0 1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output94
timestamp 1486834041
transform -1 0 21056 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output95
timestamp 1486834041
transform -1 0 19264 0 -1 2744
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output96
timestamp 1486834041
transform 1 0 18368 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output97
timestamp 1486834041
transform 1 0 16968 0 1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output98
timestamp 1486834041
transform 1 0 16408 0 1 2744
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output99
timestamp 1486834041
transform 1 0 18480 0 -1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output100
timestamp 1486834041
transform -1 0 18480 0 -1 1960
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output101
timestamp 1486834041
transform -1 0 18872 0 1 1176
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output102
timestamp 1486834041
transform -1 0 17696 0 -1 2744
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output103
timestamp 1486834041
transform -1 0 20272 0 1 392
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output104
timestamp 1486834041
transform -1 0 17976 0 1 2744
box -43 -43 827 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output105
timestamp 1486834041
transform -1 0 1176 0 -1 6664
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_16
timestamp 1486834041
transform 1 0 336 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1486834041
transform -1 0 26040 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_17
timestamp 1486834041
transform 1 0 336 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1486834041
transform -1 0 26040 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_18
timestamp 1486834041
transform 1 0 336 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1486834041
transform -1 0 26040 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_19
timestamp 1486834041
transform 1 0 336 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1486834041
transform -1 0 26040 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_20
timestamp 1486834041
transform 1 0 336 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1486834041
transform -1 0 26040 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_21
timestamp 1486834041
transform 1 0 336 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1486834041
transform -1 0 26040 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_22
timestamp 1486834041
transform 1 0 336 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1486834041
transform -1 0 26040 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_23
timestamp 1486834041
transform 1 0 336 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1486834041
transform -1 0 26040 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_24
timestamp 1486834041
transform 1 0 336 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1486834041
transform -1 0 26040 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_25
timestamp 1486834041
transform 1 0 336 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1486834041
transform -1 0 26040 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_26
timestamp 1486834041
transform 1 0 336 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1486834041
transform -1 0 26040 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_27
timestamp 1486834041
transform 1 0 336 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1486834041
transform -1 0 26040 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_28
timestamp 1486834041
transform 1 0 336 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1486834041
transform -1 0 26040 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_29
timestamp 1486834041
transform 1 0 336 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1486834041
transform -1 0 26040 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_30
timestamp 1486834041
transform 1 0 336 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1486834041
transform -1 0 26040 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_31
timestamp 1486834041
transform 1 0 336 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1486834041
transform -1 0 26040 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_32
timestamp 1486834041
transform 1 0 2240 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_33
timestamp 1486834041
transform 1 0 4144 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_34
timestamp 1486834041
transform 1 0 6048 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_35
timestamp 1486834041
transform 1 0 7952 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_36
timestamp 1486834041
transform 1 0 9856 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_37
timestamp 1486834041
transform 1 0 11760 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_38
timestamp 1486834041
transform 1 0 13664 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_39
timestamp 1486834041
transform 1 0 15568 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_40
timestamp 1486834041
transform 1 0 17472 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_41
timestamp 1486834041
transform 1 0 19376 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_42
timestamp 1486834041
transform 1 0 21280 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_43
timestamp 1486834041
transform 1 0 23184 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_44
timestamp 1486834041
transform 1 0 25088 0 1 392
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_45
timestamp 1486834041
transform 1 0 4256 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_46
timestamp 1486834041
transform 1 0 8176 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_47
timestamp 1486834041
transform 1 0 12096 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_48
timestamp 1486834041
transform 1 0 16016 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_49
timestamp 1486834041
transform 1 0 19936 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_50
timestamp 1486834041
transform 1 0 23856 0 -1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_51
timestamp 1486834041
transform 1 0 2296 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_52
timestamp 1486834041
transform 1 0 6216 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_53
timestamp 1486834041
transform 1 0 10136 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_54
timestamp 1486834041
transform 1 0 14056 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_55
timestamp 1486834041
transform 1 0 17976 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_56
timestamp 1486834041
transform 1 0 21896 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_57
timestamp 1486834041
transform 1 0 25816 0 1 1176
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_58
timestamp 1486834041
transform 1 0 4256 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_59
timestamp 1486834041
transform 1 0 8176 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_60
timestamp 1486834041
transform 1 0 12096 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_61
timestamp 1486834041
transform 1 0 16016 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_62
timestamp 1486834041
transform 1 0 19936 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_63
timestamp 1486834041
transform 1 0 23856 0 -1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_64
timestamp 1486834041
transform 1 0 2296 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_65
timestamp 1486834041
transform 1 0 6216 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_66
timestamp 1486834041
transform 1 0 10136 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_67
timestamp 1486834041
transform 1 0 14056 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_68
timestamp 1486834041
transform 1 0 17976 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_69
timestamp 1486834041
transform 1 0 21896 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_70
timestamp 1486834041
transform 1 0 25816 0 1 1960
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_71
timestamp 1486834041
transform 1 0 4256 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_72
timestamp 1486834041
transform 1 0 8176 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_73
timestamp 1486834041
transform 1 0 12096 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_74
timestamp 1486834041
transform 1 0 16016 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_75
timestamp 1486834041
transform 1 0 19936 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_76
timestamp 1486834041
transform 1 0 23856 0 -1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_77
timestamp 1486834041
transform 1 0 2296 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_78
timestamp 1486834041
transform 1 0 6216 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_79
timestamp 1486834041
transform 1 0 10136 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_80
timestamp 1486834041
transform 1 0 14056 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_81
timestamp 1486834041
transform 1 0 17976 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_82
timestamp 1486834041
transform 1 0 21896 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_83
timestamp 1486834041
transform 1 0 25816 0 1 2744
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_84
timestamp 1486834041
transform 1 0 4256 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_85
timestamp 1486834041
transform 1 0 8176 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_86
timestamp 1486834041
transform 1 0 12096 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_87
timestamp 1486834041
transform 1 0 16016 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_88
timestamp 1486834041
transform 1 0 19936 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_89
timestamp 1486834041
transform 1 0 23856 0 -1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_90
timestamp 1486834041
transform 1 0 2296 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_91
timestamp 1486834041
transform 1 0 6216 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_92
timestamp 1486834041
transform 1 0 10136 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_93
timestamp 1486834041
transform 1 0 14056 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_94
timestamp 1486834041
transform 1 0 17976 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_95
timestamp 1486834041
transform 1 0 21896 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_96
timestamp 1486834041
transform 1 0 25816 0 1 3528
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_97
timestamp 1486834041
transform 1 0 4256 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_98
timestamp 1486834041
transform 1 0 8176 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_99
timestamp 1486834041
transform 1 0 12096 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_100
timestamp 1486834041
transform 1 0 16016 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_101
timestamp 1486834041
transform 1 0 19936 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_102
timestamp 1486834041
transform 1 0 23856 0 -1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_103
timestamp 1486834041
transform 1 0 2296 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_104
timestamp 1486834041
transform 1 0 6216 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_105
timestamp 1486834041
transform 1 0 10136 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_106
timestamp 1486834041
transform 1 0 14056 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_107
timestamp 1486834041
transform 1 0 17976 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_108
timestamp 1486834041
transform 1 0 21896 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_109
timestamp 1486834041
transform 1 0 25816 0 1 4312
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_110
timestamp 1486834041
transform 1 0 4256 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_111
timestamp 1486834041
transform 1 0 8176 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_112
timestamp 1486834041
transform 1 0 12096 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_113
timestamp 1486834041
transform 1 0 16016 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_114
timestamp 1486834041
transform 1 0 19936 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_115
timestamp 1486834041
transform 1 0 23856 0 -1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_116
timestamp 1486834041
transform 1 0 2296 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_117
timestamp 1486834041
transform 1 0 6216 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_118
timestamp 1486834041
transform 1 0 10136 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_119
timestamp 1486834041
transform 1 0 14056 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_120
timestamp 1486834041
transform 1 0 17976 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_121
timestamp 1486834041
transform 1 0 21896 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_122
timestamp 1486834041
transform 1 0 25816 0 1 5096
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_123
timestamp 1486834041
transform 1 0 4256 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_124
timestamp 1486834041
transform 1 0 8176 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_125
timestamp 1486834041
transform 1 0 12096 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_126
timestamp 1486834041
transform 1 0 16016 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_127
timestamp 1486834041
transform 1 0 19936 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_128
timestamp 1486834041
transform 1 0 23856 0 -1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_129
timestamp 1486834041
transform 1 0 2296 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_130
timestamp 1486834041
transform 1 0 6216 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_131
timestamp 1486834041
transform 1 0 10136 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_132
timestamp 1486834041
transform 1 0 14056 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_133
timestamp 1486834041
transform 1 0 17976 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_134
timestamp 1486834041
transform 1 0 21896 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_135
timestamp 1486834041
transform 1 0 25816 0 1 5880
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_136
timestamp 1486834041
transform 1 0 2240 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_137
timestamp 1486834041
transform 1 0 4144 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_138
timestamp 1486834041
transform 1 0 6048 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_139
timestamp 1486834041
transform 1 0 7952 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_140
timestamp 1486834041
transform 1 0 9856 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_141
timestamp 1486834041
transform 1 0 11760 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_142
timestamp 1486834041
transform 1 0 13664 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_143
timestamp 1486834041
transform 1 0 15568 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_144
timestamp 1486834041
transform 1 0 17472 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_145
timestamp 1486834041
transform 1 0 19376 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_146
timestamp 1486834041
transform 1 0 21280 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_147
timestamp 1486834041
transform 1 0 23184 0 -1 6664
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_148
timestamp 1486834041
transform 1 0 25088 0 -1 6664
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 0 56 56 0 FreeSans 224 0 0 0 FrameData[0]
port 0 nsew signal input
flabel metal3 s 0 2240 56 2296 0 FreeSans 224 0 0 0 FrameData[10]
port 1 nsew signal input
flabel metal3 s 0 2464 56 2520 0 FreeSans 224 0 0 0 FrameData[11]
port 2 nsew signal input
flabel metal3 s 0 2688 56 2744 0 FreeSans 224 0 0 0 FrameData[12]
port 3 nsew signal input
flabel metal3 s 0 2912 56 2968 0 FreeSans 224 0 0 0 FrameData[13]
port 4 nsew signal input
flabel metal3 s 0 3136 56 3192 0 FreeSans 224 0 0 0 FrameData[14]
port 5 nsew signal input
flabel metal3 s 0 3360 56 3416 0 FreeSans 224 0 0 0 FrameData[15]
port 6 nsew signal input
flabel metal3 s 0 3584 56 3640 0 FreeSans 224 0 0 0 FrameData[16]
port 7 nsew signal input
flabel metal3 s 0 3808 56 3864 0 FreeSans 224 0 0 0 FrameData[17]
port 8 nsew signal input
flabel metal3 s 0 4032 56 4088 0 FreeSans 224 0 0 0 FrameData[18]
port 9 nsew signal input
flabel metal3 s 0 4256 56 4312 0 FreeSans 224 0 0 0 FrameData[19]
port 10 nsew signal input
flabel metal3 s 0 224 56 280 0 FreeSans 224 0 0 0 FrameData[1]
port 11 nsew signal input
flabel metal3 s 0 4480 56 4536 0 FreeSans 224 0 0 0 FrameData[20]
port 12 nsew signal input
flabel metal3 s 0 4704 56 4760 0 FreeSans 224 0 0 0 FrameData[21]
port 13 nsew signal input
flabel metal3 s 0 4928 56 4984 0 FreeSans 224 0 0 0 FrameData[22]
port 14 nsew signal input
flabel metal3 s 0 5152 56 5208 0 FreeSans 224 0 0 0 FrameData[23]
port 15 nsew signal input
flabel metal3 s 0 5376 56 5432 0 FreeSans 224 0 0 0 FrameData[24]
port 16 nsew signal input
flabel metal3 s 0 5600 56 5656 0 FreeSans 224 0 0 0 FrameData[25]
port 17 nsew signal input
flabel metal3 s 0 5824 56 5880 0 FreeSans 224 0 0 0 FrameData[26]
port 18 nsew signal input
flabel metal3 s 0 6048 56 6104 0 FreeSans 224 0 0 0 FrameData[27]
port 19 nsew signal input
flabel metal3 s 0 6272 56 6328 0 FreeSans 224 0 0 0 FrameData[28]
port 20 nsew signal input
flabel metal3 s 0 6496 56 6552 0 FreeSans 224 0 0 0 FrameData[29]
port 21 nsew signal input
flabel metal3 s 0 448 56 504 0 FreeSans 224 0 0 0 FrameData[2]
port 22 nsew signal input
flabel metal3 s 0 6720 56 6776 0 FreeSans 224 0 0 0 FrameData[30]
port 23 nsew signal input
flabel metal3 s 0 6944 56 7000 0 FreeSans 224 0 0 0 FrameData[31]
port 24 nsew signal input
flabel metal3 s 0 672 56 728 0 FreeSans 224 0 0 0 FrameData[3]
port 25 nsew signal input
flabel metal3 s 0 896 56 952 0 FreeSans 224 0 0 0 FrameData[4]
port 26 nsew signal input
flabel metal3 s 0 1120 56 1176 0 FreeSans 224 0 0 0 FrameData[5]
port 27 nsew signal input
flabel metal3 s 0 1344 56 1400 0 FreeSans 224 0 0 0 FrameData[6]
port 28 nsew signal input
flabel metal3 s 0 1568 56 1624 0 FreeSans 224 0 0 0 FrameData[7]
port 29 nsew signal input
flabel metal3 s 0 1792 56 1848 0 FreeSans 224 0 0 0 FrameData[8]
port 30 nsew signal input
flabel metal3 s 0 2016 56 2072 0 FreeSans 224 0 0 0 FrameData[9]
port 31 nsew signal input
flabel metal3 s 26320 0 26376 56 0 FreeSans 224 0 0 0 FrameData_O[0]
port 32 nsew signal output
flabel metal3 s 26320 2240 26376 2296 0 FreeSans 224 0 0 0 FrameData_O[10]
port 33 nsew signal output
flabel metal3 s 26320 2464 26376 2520 0 FreeSans 224 0 0 0 FrameData_O[11]
port 34 nsew signal output
flabel metal3 s 26320 2688 26376 2744 0 FreeSans 224 0 0 0 FrameData_O[12]
port 35 nsew signal output
flabel metal3 s 26320 2912 26376 2968 0 FreeSans 224 0 0 0 FrameData_O[13]
port 36 nsew signal output
flabel metal3 s 26320 3136 26376 3192 0 FreeSans 224 0 0 0 FrameData_O[14]
port 37 nsew signal output
flabel metal3 s 26320 3360 26376 3416 0 FreeSans 224 0 0 0 FrameData_O[15]
port 38 nsew signal output
flabel metal3 s 26320 3584 26376 3640 0 FreeSans 224 0 0 0 FrameData_O[16]
port 39 nsew signal output
flabel metal3 s 26320 3808 26376 3864 0 FreeSans 224 0 0 0 FrameData_O[17]
port 40 nsew signal output
flabel metal3 s 26320 4032 26376 4088 0 FreeSans 224 0 0 0 FrameData_O[18]
port 41 nsew signal output
flabel metal3 s 26320 4256 26376 4312 0 FreeSans 224 0 0 0 FrameData_O[19]
port 42 nsew signal output
flabel metal3 s 26320 224 26376 280 0 FreeSans 224 0 0 0 FrameData_O[1]
port 43 nsew signal output
flabel metal3 s 26320 4480 26376 4536 0 FreeSans 224 0 0 0 FrameData_O[20]
port 44 nsew signal output
flabel metal3 s 26320 4704 26376 4760 0 FreeSans 224 0 0 0 FrameData_O[21]
port 45 nsew signal output
flabel metal3 s 26320 4928 26376 4984 0 FreeSans 224 0 0 0 FrameData_O[22]
port 46 nsew signal output
flabel metal3 s 26320 5152 26376 5208 0 FreeSans 224 0 0 0 FrameData_O[23]
port 47 nsew signal output
flabel metal3 s 26320 5376 26376 5432 0 FreeSans 224 0 0 0 FrameData_O[24]
port 48 nsew signal output
flabel metal3 s 26320 5600 26376 5656 0 FreeSans 224 0 0 0 FrameData_O[25]
port 49 nsew signal output
flabel metal3 s 26320 5824 26376 5880 0 FreeSans 224 0 0 0 FrameData_O[26]
port 50 nsew signal output
flabel metal3 s 26320 6048 26376 6104 0 FreeSans 224 0 0 0 FrameData_O[27]
port 51 nsew signal output
flabel metal3 s 26320 6272 26376 6328 0 FreeSans 224 0 0 0 FrameData_O[28]
port 52 nsew signal output
flabel metal3 s 26320 6496 26376 6552 0 FreeSans 224 0 0 0 FrameData_O[29]
port 53 nsew signal output
flabel metal3 s 26320 448 26376 504 0 FreeSans 224 0 0 0 FrameData_O[2]
port 54 nsew signal output
flabel metal3 s 26320 6720 26376 6776 0 FreeSans 224 0 0 0 FrameData_O[30]
port 55 nsew signal output
flabel metal3 s 26320 6944 26376 7000 0 FreeSans 224 0 0 0 FrameData_O[31]
port 56 nsew signal output
flabel metal3 s 26320 672 26376 728 0 FreeSans 224 0 0 0 FrameData_O[3]
port 57 nsew signal output
flabel metal3 s 26320 896 26376 952 0 FreeSans 224 0 0 0 FrameData_O[4]
port 58 nsew signal output
flabel metal3 s 26320 1120 26376 1176 0 FreeSans 224 0 0 0 FrameData_O[5]
port 59 nsew signal output
flabel metal3 s 26320 1344 26376 1400 0 FreeSans 224 0 0 0 FrameData_O[6]
port 60 nsew signal output
flabel metal3 s 26320 1568 26376 1624 0 FreeSans 224 0 0 0 FrameData_O[7]
port 61 nsew signal output
flabel metal3 s 26320 1792 26376 1848 0 FreeSans 224 0 0 0 FrameData_O[8]
port 62 nsew signal output
flabel metal3 s 26320 2016 26376 2072 0 FreeSans 224 0 0 0 FrameData_O[9]
port 63 nsew signal output
flabel metal2 s 17920 0 17976 56 0 FreeSans 224 0 0 0 FrameStrobe[0]
port 64 nsew signal input
flabel metal2 s 19040 0 19096 56 0 FreeSans 224 0 0 0 FrameStrobe[10]
port 65 nsew signal input
flabel metal2 s 19152 0 19208 56 0 FreeSans 224 0 0 0 FrameStrobe[11]
port 66 nsew signal input
flabel metal2 s 19264 0 19320 56 0 FreeSans 224 0 0 0 FrameStrobe[12]
port 67 nsew signal input
flabel metal2 s 19376 0 19432 56 0 FreeSans 224 0 0 0 FrameStrobe[13]
port 68 nsew signal input
flabel metal2 s 19488 0 19544 56 0 FreeSans 224 0 0 0 FrameStrobe[14]
port 69 nsew signal input
flabel metal2 s 19600 0 19656 56 0 FreeSans 224 0 0 0 FrameStrobe[15]
port 70 nsew signal input
flabel metal2 s 19712 0 19768 56 0 FreeSans 224 0 0 0 FrameStrobe[16]
port 71 nsew signal input
flabel metal2 s 19824 0 19880 56 0 FreeSans 224 0 0 0 FrameStrobe[17]
port 72 nsew signal input
flabel metal2 s 19936 0 19992 56 0 FreeSans 224 0 0 0 FrameStrobe[18]
port 73 nsew signal input
flabel metal2 s 20048 0 20104 56 0 FreeSans 224 0 0 0 FrameStrobe[19]
port 74 nsew signal input
flabel metal2 s 18032 0 18088 56 0 FreeSans 224 0 0 0 FrameStrobe[1]
port 75 nsew signal input
flabel metal2 s 18144 0 18200 56 0 FreeSans 224 0 0 0 FrameStrobe[2]
port 76 nsew signal input
flabel metal2 s 18256 0 18312 56 0 FreeSans 224 0 0 0 FrameStrobe[3]
port 77 nsew signal input
flabel metal2 s 18368 0 18424 56 0 FreeSans 224 0 0 0 FrameStrobe[4]
port 78 nsew signal input
flabel metal2 s 18480 0 18536 56 0 FreeSans 224 0 0 0 FrameStrobe[5]
port 79 nsew signal input
flabel metal2 s 18592 0 18648 56 0 FreeSans 224 0 0 0 FrameStrobe[6]
port 80 nsew signal input
flabel metal2 s 18704 0 18760 56 0 FreeSans 224 0 0 0 FrameStrobe[7]
port 81 nsew signal input
flabel metal2 s 18816 0 18872 56 0 FreeSans 224 0 0 0 FrameStrobe[8]
port 82 nsew signal input
flabel metal2 s 18928 0 18984 56 0 FreeSans 224 0 0 0 FrameStrobe[9]
port 83 nsew signal input
flabel metal2 s 2016 7056 2072 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[0]
port 84 nsew signal output
flabel metal2 s 14336 7056 14392 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[10]
port 85 nsew signal output
flabel metal2 s 15568 7056 15624 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[11]
port 86 nsew signal output
flabel metal2 s 16800 7056 16856 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[12]
port 87 nsew signal output
flabel metal2 s 18032 7056 18088 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[13]
port 88 nsew signal output
flabel metal2 s 19264 7056 19320 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[14]
port 89 nsew signal output
flabel metal2 s 20496 7056 20552 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[15]
port 90 nsew signal output
flabel metal2 s 21728 7056 21784 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[16]
port 91 nsew signal output
flabel metal2 s 22960 7056 23016 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[17]
port 92 nsew signal output
flabel metal2 s 24192 7056 24248 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[18]
port 93 nsew signal output
flabel metal2 s 25424 7056 25480 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[19]
port 94 nsew signal output
flabel metal2 s 3248 7056 3304 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[1]
port 95 nsew signal output
flabel metal2 s 4480 7056 4536 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[2]
port 96 nsew signal output
flabel metal2 s 5712 7056 5768 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[3]
port 97 nsew signal output
flabel metal2 s 6944 7056 7000 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[4]
port 98 nsew signal output
flabel metal2 s 8176 7056 8232 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[5]
port 99 nsew signal output
flabel metal2 s 9408 7056 9464 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[6]
port 100 nsew signal output
flabel metal2 s 10640 7056 10696 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[7]
port 101 nsew signal output
flabel metal2 s 11872 7056 11928 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[8]
port 102 nsew signal output
flabel metal2 s 13104 7056 13160 7112 0 FreeSans 224 0 0 0 FrameStrobe_O[9]
port 103 nsew signal output
flabel metal2 s 6160 0 6216 56 0 FreeSans 224 0 0 0 N1END[0]
port 104 nsew signal input
flabel metal2 s 6272 0 6328 56 0 FreeSans 224 0 0 0 N1END[1]
port 105 nsew signal input
flabel metal2 s 6384 0 6440 56 0 FreeSans 224 0 0 0 N1END[2]
port 106 nsew signal input
flabel metal2 s 6496 0 6552 56 0 FreeSans 224 0 0 0 N1END[3]
port 107 nsew signal input
flabel metal2 s 7504 0 7560 56 0 FreeSans 224 0 0 0 N2END[0]
port 108 nsew signal input
flabel metal2 s 7616 0 7672 56 0 FreeSans 224 0 0 0 N2END[1]
port 109 nsew signal input
flabel metal2 s 7728 0 7784 56 0 FreeSans 224 0 0 0 N2END[2]
port 110 nsew signal input
flabel metal2 s 7840 0 7896 56 0 FreeSans 224 0 0 0 N2END[3]
port 111 nsew signal input
flabel metal2 s 7952 0 8008 56 0 FreeSans 224 0 0 0 N2END[4]
port 112 nsew signal input
flabel metal2 s 8064 0 8120 56 0 FreeSans 224 0 0 0 N2END[5]
port 113 nsew signal input
flabel metal2 s 8176 0 8232 56 0 FreeSans 224 0 0 0 N2END[6]
port 114 nsew signal input
flabel metal2 s 8288 0 8344 56 0 FreeSans 224 0 0 0 N2END[7]
port 115 nsew signal input
flabel metal2 s 6608 0 6664 56 0 FreeSans 224 0 0 0 N2MID[0]
port 116 nsew signal input
flabel metal2 s 6720 0 6776 56 0 FreeSans 224 0 0 0 N2MID[1]
port 117 nsew signal input
flabel metal2 s 6832 0 6888 56 0 FreeSans 224 0 0 0 N2MID[2]
port 118 nsew signal input
flabel metal2 s 6944 0 7000 56 0 FreeSans 224 0 0 0 N2MID[3]
port 119 nsew signal input
flabel metal2 s 7056 0 7112 56 0 FreeSans 224 0 0 0 N2MID[4]
port 120 nsew signal input
flabel metal2 s 7168 0 7224 56 0 FreeSans 224 0 0 0 N2MID[5]
port 121 nsew signal input
flabel metal2 s 7280 0 7336 56 0 FreeSans 224 0 0 0 N2MID[6]
port 122 nsew signal input
flabel metal2 s 7392 0 7448 56 0 FreeSans 224 0 0 0 N2MID[7]
port 123 nsew signal input
flabel metal2 s 8400 0 8456 56 0 FreeSans 224 0 0 0 N4END[0]
port 124 nsew signal input
flabel metal2 s 9520 0 9576 56 0 FreeSans 224 0 0 0 N4END[10]
port 125 nsew signal input
flabel metal2 s 9632 0 9688 56 0 FreeSans 224 0 0 0 N4END[11]
port 126 nsew signal input
flabel metal2 s 9744 0 9800 56 0 FreeSans 224 0 0 0 N4END[12]
port 127 nsew signal input
flabel metal2 s 9856 0 9912 56 0 FreeSans 224 0 0 0 N4END[13]
port 128 nsew signal input
flabel metal2 s 9968 0 10024 56 0 FreeSans 224 0 0 0 N4END[14]
port 129 nsew signal input
flabel metal2 s 10080 0 10136 56 0 FreeSans 224 0 0 0 N4END[15]
port 130 nsew signal input
flabel metal2 s 8512 0 8568 56 0 FreeSans 224 0 0 0 N4END[1]
port 131 nsew signal input
flabel metal2 s 8624 0 8680 56 0 FreeSans 224 0 0 0 N4END[2]
port 132 nsew signal input
flabel metal2 s 8736 0 8792 56 0 FreeSans 224 0 0 0 N4END[3]
port 133 nsew signal input
flabel metal2 s 8848 0 8904 56 0 FreeSans 224 0 0 0 N4END[4]
port 134 nsew signal input
flabel metal2 s 8960 0 9016 56 0 FreeSans 224 0 0 0 N4END[5]
port 135 nsew signal input
flabel metal2 s 9072 0 9128 56 0 FreeSans 224 0 0 0 N4END[6]
port 136 nsew signal input
flabel metal2 s 9184 0 9240 56 0 FreeSans 224 0 0 0 N4END[7]
port 137 nsew signal input
flabel metal2 s 9296 0 9352 56 0 FreeSans 224 0 0 0 N4END[8]
port 138 nsew signal input
flabel metal2 s 9408 0 9464 56 0 FreeSans 224 0 0 0 N4END[9]
port 139 nsew signal input
flabel metal2 s 10192 0 10248 56 0 FreeSans 224 0 0 0 NN4END[0]
port 140 nsew signal input
flabel metal2 s 11312 0 11368 56 0 FreeSans 224 0 0 0 NN4END[10]
port 141 nsew signal input
flabel metal2 s 11424 0 11480 56 0 FreeSans 224 0 0 0 NN4END[11]
port 142 nsew signal input
flabel metal2 s 11536 0 11592 56 0 FreeSans 224 0 0 0 NN4END[12]
port 143 nsew signal input
flabel metal2 s 11648 0 11704 56 0 FreeSans 224 0 0 0 NN4END[13]
port 144 nsew signal input
flabel metal2 s 11760 0 11816 56 0 FreeSans 224 0 0 0 NN4END[14]
port 145 nsew signal input
flabel metal2 s 11872 0 11928 56 0 FreeSans 224 0 0 0 NN4END[15]
port 146 nsew signal input
flabel metal2 s 10304 0 10360 56 0 FreeSans 224 0 0 0 NN4END[1]
port 147 nsew signal input
flabel metal2 s 10416 0 10472 56 0 FreeSans 224 0 0 0 NN4END[2]
port 148 nsew signal input
flabel metal2 s 10528 0 10584 56 0 FreeSans 224 0 0 0 NN4END[3]
port 149 nsew signal input
flabel metal2 s 10640 0 10696 56 0 FreeSans 224 0 0 0 NN4END[4]
port 150 nsew signal input
flabel metal2 s 10752 0 10808 56 0 FreeSans 224 0 0 0 NN4END[5]
port 151 nsew signal input
flabel metal2 s 10864 0 10920 56 0 FreeSans 224 0 0 0 NN4END[6]
port 152 nsew signal input
flabel metal2 s 10976 0 11032 56 0 FreeSans 224 0 0 0 NN4END[7]
port 153 nsew signal input
flabel metal2 s 11088 0 11144 56 0 FreeSans 224 0 0 0 NN4END[8]
port 154 nsew signal input
flabel metal2 s 11200 0 11256 56 0 FreeSans 224 0 0 0 NN4END[9]
port 155 nsew signal input
flabel metal2 s 11984 0 12040 56 0 FreeSans 224 0 0 0 S1BEG[0]
port 156 nsew signal output
flabel metal2 s 12096 0 12152 56 0 FreeSans 224 0 0 0 S1BEG[1]
port 157 nsew signal output
flabel metal2 s 12208 0 12264 56 0 FreeSans 224 0 0 0 S1BEG[2]
port 158 nsew signal output
flabel metal2 s 12320 0 12376 56 0 FreeSans 224 0 0 0 S1BEG[3]
port 159 nsew signal output
flabel metal2 s 12432 0 12488 56 0 FreeSans 224 0 0 0 S2BEG[0]
port 160 nsew signal output
flabel metal2 s 12544 0 12600 56 0 FreeSans 224 0 0 0 S2BEG[1]
port 161 nsew signal output
flabel metal2 s 12656 0 12712 56 0 FreeSans 224 0 0 0 S2BEG[2]
port 162 nsew signal output
flabel metal2 s 12768 0 12824 56 0 FreeSans 224 0 0 0 S2BEG[3]
port 163 nsew signal output
flabel metal2 s 12880 0 12936 56 0 FreeSans 224 0 0 0 S2BEG[4]
port 164 nsew signal output
flabel metal2 s 12992 0 13048 56 0 FreeSans 224 0 0 0 S2BEG[5]
port 165 nsew signal output
flabel metal2 s 13104 0 13160 56 0 FreeSans 224 0 0 0 S2BEG[6]
port 166 nsew signal output
flabel metal2 s 13216 0 13272 56 0 FreeSans 224 0 0 0 S2BEG[7]
port 167 nsew signal output
flabel metal2 s 13328 0 13384 56 0 FreeSans 224 0 0 0 S2BEGb[0]
port 168 nsew signal output
flabel metal2 s 13440 0 13496 56 0 FreeSans 224 0 0 0 S2BEGb[1]
port 169 nsew signal output
flabel metal2 s 13552 0 13608 56 0 FreeSans 224 0 0 0 S2BEGb[2]
port 170 nsew signal output
flabel metal2 s 13664 0 13720 56 0 FreeSans 224 0 0 0 S2BEGb[3]
port 171 nsew signal output
flabel metal2 s 13776 0 13832 56 0 FreeSans 224 0 0 0 S2BEGb[4]
port 172 nsew signal output
flabel metal2 s 13888 0 13944 56 0 FreeSans 224 0 0 0 S2BEGb[5]
port 173 nsew signal output
flabel metal2 s 14000 0 14056 56 0 FreeSans 224 0 0 0 S2BEGb[6]
port 174 nsew signal output
flabel metal2 s 14112 0 14168 56 0 FreeSans 224 0 0 0 S2BEGb[7]
port 175 nsew signal output
flabel metal2 s 14224 0 14280 56 0 FreeSans 224 0 0 0 S4BEG[0]
port 176 nsew signal output
flabel metal2 s 15344 0 15400 56 0 FreeSans 224 0 0 0 S4BEG[10]
port 177 nsew signal output
flabel metal2 s 15456 0 15512 56 0 FreeSans 224 0 0 0 S4BEG[11]
port 178 nsew signal output
flabel metal2 s 15568 0 15624 56 0 FreeSans 224 0 0 0 S4BEG[12]
port 179 nsew signal output
flabel metal2 s 15680 0 15736 56 0 FreeSans 224 0 0 0 S4BEG[13]
port 180 nsew signal output
flabel metal2 s 15792 0 15848 56 0 FreeSans 224 0 0 0 S4BEG[14]
port 181 nsew signal output
flabel metal2 s 15904 0 15960 56 0 FreeSans 224 0 0 0 S4BEG[15]
port 182 nsew signal output
flabel metal2 s 14336 0 14392 56 0 FreeSans 224 0 0 0 S4BEG[1]
port 183 nsew signal output
flabel metal2 s 14448 0 14504 56 0 FreeSans 224 0 0 0 S4BEG[2]
port 184 nsew signal output
flabel metal2 s 14560 0 14616 56 0 FreeSans 224 0 0 0 S4BEG[3]
port 185 nsew signal output
flabel metal2 s 14672 0 14728 56 0 FreeSans 224 0 0 0 S4BEG[4]
port 186 nsew signal output
flabel metal2 s 14784 0 14840 56 0 FreeSans 224 0 0 0 S4BEG[5]
port 187 nsew signal output
flabel metal2 s 14896 0 14952 56 0 FreeSans 224 0 0 0 S4BEG[6]
port 188 nsew signal output
flabel metal2 s 15008 0 15064 56 0 FreeSans 224 0 0 0 S4BEG[7]
port 189 nsew signal output
flabel metal2 s 15120 0 15176 56 0 FreeSans 224 0 0 0 S4BEG[8]
port 190 nsew signal output
flabel metal2 s 15232 0 15288 56 0 FreeSans 224 0 0 0 S4BEG[9]
port 191 nsew signal output
flabel metal2 s 16016 0 16072 56 0 FreeSans 224 0 0 0 SS4BEG[0]
port 192 nsew signal output
flabel metal2 s 17136 0 17192 56 0 FreeSans 224 0 0 0 SS4BEG[10]
port 193 nsew signal output
flabel metal2 s 17248 0 17304 56 0 FreeSans 224 0 0 0 SS4BEG[11]
port 194 nsew signal output
flabel metal2 s 17360 0 17416 56 0 FreeSans 224 0 0 0 SS4BEG[12]
port 195 nsew signal output
flabel metal2 s 17472 0 17528 56 0 FreeSans 224 0 0 0 SS4BEG[13]
port 196 nsew signal output
flabel metal2 s 17584 0 17640 56 0 FreeSans 224 0 0 0 SS4BEG[14]
port 197 nsew signal output
flabel metal2 s 17696 0 17752 56 0 FreeSans 224 0 0 0 SS4BEG[15]
port 198 nsew signal output
flabel metal2 s 16128 0 16184 56 0 FreeSans 224 0 0 0 SS4BEG[1]
port 199 nsew signal output
flabel metal2 s 16240 0 16296 56 0 FreeSans 224 0 0 0 SS4BEG[2]
port 200 nsew signal output
flabel metal2 s 16352 0 16408 56 0 FreeSans 224 0 0 0 SS4BEG[3]
port 201 nsew signal output
flabel metal2 s 16464 0 16520 56 0 FreeSans 224 0 0 0 SS4BEG[4]
port 202 nsew signal output
flabel metal2 s 16576 0 16632 56 0 FreeSans 224 0 0 0 SS4BEG[5]
port 203 nsew signal output
flabel metal2 s 16688 0 16744 56 0 FreeSans 224 0 0 0 SS4BEG[6]
port 204 nsew signal output
flabel metal2 s 16800 0 16856 56 0 FreeSans 224 0 0 0 SS4BEG[7]
port 205 nsew signal output
flabel metal2 s 16912 0 16968 56 0 FreeSans 224 0 0 0 SS4BEG[8]
port 206 nsew signal output
flabel metal2 s 17024 0 17080 56 0 FreeSans 224 0 0 0 SS4BEG[9]
port 207 nsew signal output
flabel metal2 s 17808 0 17864 56 0 FreeSans 224 0 0 0 UserCLK
port 208 nsew signal input
flabel metal2 s 784 7056 840 7112 0 FreeSans 224 0 0 0 UserCLKo
port 209 nsew signal output
flabel metal4 s 1888 0 2048 7112 0 FreeSans 736 90 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 1888 0 2048 28 0 FreeSans 184 0 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 1888 7084 2048 7112 0 FreeSans 184 0 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 11888 0 12048 7112 0 FreeSans 736 90 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 11888 0 12048 28 0 FreeSans 184 0 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 11888 7084 12048 7112 0 FreeSans 184 0 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 21888 0 22048 7112 0 FreeSans 736 90 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 21888 0 22048 28 0 FreeSans 184 0 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 21888 7084 22048 7112 0 FreeSans 184 0 0 0 VDD
port 210 nsew power bidirectional
flabel metal4 s 2218 0 2378 7112 0 FreeSans 736 90 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 2218 0 2378 28 0 FreeSans 184 0 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 2218 7084 2378 7112 0 FreeSans 184 0 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 12218 0 12378 7112 0 FreeSans 736 90 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 12218 0 12378 28 0 FreeSans 184 0 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 12218 7084 12378 7112 0 FreeSans 184 0 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 22218 0 22378 7112 0 FreeSans 736 90 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 22218 0 22378 28 0 FreeSans 184 0 0 0 VSS
port 211 nsew ground bidirectional
flabel metal4 s 22218 7084 22378 7112 0 FreeSans 184 0 0 0 VSS
port 211 nsew ground bidirectional
rlabel metal1 13188 6272 13188 6272 0 VDD
rlabel metal1 13188 6664 13188 6664 0 VSS
rlabel metal2 4956 644 4956 644 0 FrameData[0]
rlabel metal3 1575 2268 1575 2268 0 FrameData[10]
rlabel metal3 1491 2492 1491 2492 0 FrameData[11]
rlabel metal3 931 2716 931 2716 0 FrameData[12]
rlabel metal3 1071 2940 1071 2940 0 FrameData[13]
rlabel metal2 2548 2996 2548 2996 0 FrameData[14]
rlabel metal3 931 3388 931 3388 0 FrameData[15]
rlabel metal3 1323 3612 1323 3612 0 FrameData[16]
rlabel metal3 1491 3836 1491 3836 0 FrameData[17]
rlabel metal3 1771 4060 1771 4060 0 FrameData[18]
rlabel metal3 623 4284 623 4284 0 FrameData[19]
rlabel metal2 5292 1008 5292 1008 0 FrameData[1]
rlabel metal3 1547 4508 1547 4508 0 FrameData[20]
rlabel metal3 931 4732 931 4732 0 FrameData[21]
rlabel metal3 1407 4956 1407 4956 0 FrameData[22]
rlabel metal3 1071 5180 1071 5180 0 FrameData[23]
rlabel metal2 24780 4060 24780 4060 0 FrameData[24]
rlabel metal3 1771 5628 1771 5628 0 FrameData[25]
rlabel metal3 259 5852 259 5852 0 FrameData[26]
rlabel metal3 203 6076 203 6076 0 FrameData[27]
rlabel metal3 315 6300 315 6300 0 FrameData[28]
rlabel metal3 847 6524 847 6524 0 FrameData[29]
rlabel metal3 679 476 679 476 0 FrameData[2]
rlabel metal2 1148 6412 1148 6412 0 FrameData[30]
rlabel metal2 23492 6412 23492 6412 0 FrameData[31]
rlabel metal3 1687 700 1687 700 0 FrameData[3]
rlabel metal2 5404 1092 5404 1092 0 FrameData[4]
rlabel metal3 707 1148 707 1148 0 FrameData[5]
rlabel metal2 6524 2240 6524 2240 0 FrameData[6]
rlabel metal3 931 1596 931 1596 0 FrameData[7]
rlabel metal3 875 1820 875 1820 0 FrameData[8]
rlabel metal2 1484 1708 1484 1708 0 FrameData[9]
rlabel metal3 25893 28 25893 28 0 FrameData_O[0]
rlabel metal3 25949 2268 25949 2268 0 FrameData_O[10]
rlabel metal3 25893 2492 25893 2492 0 FrameData_O[11]
rlabel metal2 25620 2660 25620 2660 0 FrameData_O[12]
rlabel metal3 25613 2940 25613 2940 0 FrameData_O[13]
rlabel metal2 25620 3108 25620 3108 0 FrameData_O[14]
rlabel metal3 25585 3388 25585 3388 0 FrameData_O[15]
rlabel metal2 25732 3444 25732 3444 0 FrameData_O[16]
rlabel metal3 26033 3836 26033 3836 0 FrameData_O[17]
rlabel metal2 25620 3948 25620 3948 0 FrameData_O[18]
rlabel metal3 25921 4284 25921 4284 0 FrameData_O[19]
rlabel metal3 25837 252 25837 252 0 FrameData_O[1]
rlabel metal3 26033 4508 26033 4508 0 FrameData_O[20]
rlabel metal3 25921 4732 25921 4732 0 FrameData_O[21]
rlabel metal3 26033 4956 26033 4956 0 FrameData_O[22]
rlabel metal3 25585 5180 25585 5180 0 FrameData_O[23]
rlabel metal3 25977 5404 25977 5404 0 FrameData_O[24]
rlabel metal3 25641 5628 25641 5628 0 FrameData_O[25]
rlabel metal3 25921 5852 25921 5852 0 FrameData_O[26]
rlabel metal3 25312 4844 25312 4844 0 FrameData_O[27]
rlabel metal3 25088 4620 25088 4620 0 FrameData_O[28]
rlabel metal2 24052 5432 24052 5432 0 FrameData_O[29]
rlabel metal3 25221 476 25221 476 0 FrameData_O[2]
rlabel metal3 24388 5740 24388 5740 0 FrameData_O[30]
rlabel metal3 25697 6972 25697 6972 0 FrameData_O[31]
rlabel metal3 25613 700 25613 700 0 FrameData_O[3]
rlabel metal3 25641 924 25641 924 0 FrameData_O[4]
rlabel metal2 25732 1036 25732 1036 0 FrameData_O[5]
rlabel metal3 25921 1372 25921 1372 0 FrameData_O[6]
rlabel metal2 25564 1512 25564 1512 0 FrameData_O[7]
rlabel metal3 25529 1820 25529 1820 0 FrameData_O[8]
rlabel metal2 25732 1876 25732 1876 0 FrameData_O[9]
rlabel metal2 17948 63 17948 63 0 FrameStrobe[0]
rlabel metal2 19040 2660 19040 2660 0 FrameStrobe[10]
rlabel metal2 19180 371 19180 371 0 FrameStrobe[11]
rlabel metal2 19292 595 19292 595 0 FrameStrobe[12]
rlabel metal2 19404 1295 19404 1295 0 FrameStrobe[13]
rlabel metal2 19516 2947 19516 2947 0 FrameStrobe[14]
rlabel metal2 19628 427 19628 427 0 FrameStrobe[15]
rlabel metal2 19740 539 19740 539 0 FrameStrobe[16]
rlabel metal2 19852 399 19852 399 0 FrameStrobe[17]
rlabel metal2 22820 3556 22820 3556 0 FrameStrobe[18]
rlabel metal2 20076 259 20076 259 0 FrameStrobe[19]
rlabel metal3 16744 3388 16744 3388 0 FrameStrobe[1]
rlabel metal2 18172 707 18172 707 0 FrameStrobe[2]
rlabel metal2 18284 343 18284 343 0 FrameStrobe[3]
rlabel metal2 18396 455 18396 455 0 FrameStrobe[4]
rlabel metal2 18508 259 18508 259 0 FrameStrobe[5]
rlabel metal2 18620 287 18620 287 0 FrameStrobe[6]
rlabel metal2 18732 203 18732 203 0 FrameStrobe[7]
rlabel metal2 18844 203 18844 203 0 FrameStrobe[8]
rlabel metal2 18956 315 18956 315 0 FrameStrobe[9]
rlabel metal2 2044 6797 2044 6797 0 FrameStrobe_O[0]
rlabel metal2 14364 7049 14364 7049 0 FrameStrobe_O[10]
rlabel metal2 15596 7049 15596 7049 0 FrameStrobe_O[11]
rlabel metal2 16828 6741 16828 6741 0 FrameStrobe_O[12]
rlabel metal2 18060 7049 18060 7049 0 FrameStrobe_O[13]
rlabel metal2 19292 6825 19292 6825 0 FrameStrobe_O[14]
rlabel metal2 20524 7049 20524 7049 0 FrameStrobe_O[15]
rlabel metal2 21868 6832 21868 6832 0 FrameStrobe_O[16]
rlabel metal2 22988 6825 22988 6825 0 FrameStrobe_O[17]
rlabel metal2 24220 6825 24220 6825 0 FrameStrobe_O[18]
rlabel metal3 24752 6188 24752 6188 0 FrameStrobe_O[19]
rlabel metal2 3276 7049 3276 7049 0 FrameStrobe_O[1]
rlabel metal2 4508 7049 4508 7049 0 FrameStrobe_O[2]
rlabel metal2 5740 6797 5740 6797 0 FrameStrobe_O[3]
rlabel metal2 6972 7049 6972 7049 0 FrameStrobe_O[4]
rlabel metal2 8204 7049 8204 7049 0 FrameStrobe_O[5]
rlabel metal2 9436 6741 9436 6741 0 FrameStrobe_O[6]
rlabel metal2 10668 7049 10668 7049 0 FrameStrobe_O[7]
rlabel metal2 11900 7049 11900 7049 0 FrameStrobe_O[8]
rlabel metal2 13132 6741 13132 6741 0 FrameStrobe_O[9]
rlabel metal2 1260 1064 1260 1064 0 N1END[0]
rlabel metal3 2156 4004 2156 4004 0 N1END[1]
rlabel metal2 1148 1904 1148 1904 0 N1END[2]
rlabel metal2 6524 259 6524 259 0 N1END[3]
rlabel metal2 7532 1435 7532 1435 0 N2END[0]
rlabel metal3 7504 2548 7504 2548 0 N2END[1]
rlabel metal2 7756 861 7756 861 0 N2END[2]
rlabel metal2 7868 1687 7868 1687 0 N2END[3]
rlabel metal3 8820 3500 8820 3500 0 N2END[4]
rlabel metal3 8680 2884 8680 2884 0 N2END[5]
rlabel metal3 10500 2940 10500 2940 0 N2END[6]
rlabel metal2 8316 63 8316 63 0 N2END[7]
rlabel metal3 3318 2548 3318 2548 0 N2MID[0]
rlabel metal2 3164 2240 3164 2240 0 N2MID[1]
rlabel metal2 4172 3304 4172 3304 0 N2MID[2]
rlabel metal2 6972 1827 6972 1827 0 N2MID[3]
rlabel metal2 7084 511 7084 511 0 N2MID[4]
rlabel metal2 7196 1463 7196 1463 0 N2MID[5]
rlabel metal2 7308 427 7308 427 0 N2MID[6]
rlabel metal2 7420 427 7420 427 0 N2MID[7]
rlabel metal2 8428 259 8428 259 0 N4END[0]
rlabel metal3 10836 5628 10836 5628 0 N4END[10]
rlabel metal3 9968 3332 9968 3332 0 N4END[11]
rlabel metal3 10668 1932 10668 1932 0 N4END[12]
rlabel metal3 10444 3612 10444 3612 0 N4END[13]
rlabel metal2 9996 861 9996 861 0 N4END[14]
rlabel metal2 10108 861 10108 861 0 N4END[15]
rlabel metal2 19348 1540 19348 1540 0 N4END[1]
rlabel metal2 8652 427 8652 427 0 N4END[2]
rlabel metal2 8764 371 8764 371 0 N4END[3]
rlabel metal2 8876 455 8876 455 0 N4END[4]
rlabel metal2 8988 483 8988 483 0 N4END[5]
rlabel metal2 9100 861 9100 861 0 N4END[6]
rlabel metal2 9212 511 9212 511 0 N4END[7]
rlabel metal2 9324 175 9324 175 0 N4END[8]
rlabel metal2 9436 651 9436 651 0 N4END[9]
rlabel metal2 24668 2632 24668 2632 0 NN4END[0]
rlabel metal2 11340 203 11340 203 0 NN4END[10]
rlabel metal2 11452 595 11452 595 0 NN4END[11]
rlabel metal3 12152 1820 12152 1820 0 NN4END[12]
rlabel metal2 11676 315 11676 315 0 NN4END[13]
rlabel metal2 11788 119 11788 119 0 NN4END[14]
rlabel metal2 14420 840 14420 840 0 NN4END[15]
rlabel metal3 14532 840 14532 840 0 NN4END[1]
rlabel metal2 14196 476 14196 476 0 NN4END[2]
rlabel metal2 21308 4060 21308 4060 0 NN4END[3]
rlabel metal2 21084 2912 21084 2912 0 NN4END[4]
rlabel metal2 13524 364 13524 364 0 NN4END[5]
rlabel metal2 13524 1064 13524 1064 0 NN4END[6]
rlabel metal2 11004 735 11004 735 0 NN4END[7]
rlabel metal2 11116 1351 11116 1351 0 NN4END[8]
rlabel metal2 11228 1295 11228 1295 0 NN4END[9]
rlabel metal2 12012 371 12012 371 0 S1BEG[0]
rlabel metal2 12124 91 12124 91 0 S1BEG[1]
rlabel metal2 12236 175 12236 175 0 S1BEG[2]
rlabel metal2 12348 175 12348 175 0 S1BEG[3]
rlabel metal2 12460 343 12460 343 0 S2BEG[0]
rlabel metal2 12572 147 12572 147 0 S2BEG[1]
rlabel metal2 12684 861 12684 861 0 S2BEG[2]
rlabel metal2 12796 651 12796 651 0 S2BEG[3]
rlabel metal2 13300 1120 13300 1120 0 S2BEG[4]
rlabel metal2 13020 287 13020 287 0 S2BEG[5]
rlabel metal2 13132 455 13132 455 0 S2BEG[6]
rlabel metal2 13636 980 13636 980 0 S2BEG[7]
rlabel metal2 13356 259 13356 259 0 S2BEGb[0]
rlabel metal2 13468 259 13468 259 0 S2BEGb[1]
rlabel metal2 13580 231 13580 231 0 S2BEGb[2]
rlabel metal2 13692 147 13692 147 0 S2BEGb[3]
rlabel metal2 13804 175 13804 175 0 S2BEGb[4]
rlabel metal2 13916 343 13916 343 0 S2BEGb[5]
rlabel metal2 14028 427 14028 427 0 S2BEGb[6]
rlabel metal2 14140 119 14140 119 0 S2BEGb[7]
rlabel metal2 14252 259 14252 259 0 S4BEG[0]
rlabel metal3 15932 1708 15932 1708 0 S4BEG[10]
rlabel metal2 15484 371 15484 371 0 S4BEG[11]
rlabel metal2 15596 147 15596 147 0 S4BEG[12]
rlabel metal2 15708 427 15708 427 0 S4BEG[13]
rlabel metal2 15820 455 15820 455 0 S4BEG[14]
rlabel metal2 15932 847 15932 847 0 S4BEG[15]
rlabel metal2 14364 315 14364 315 0 S4BEG[1]
rlabel metal2 14476 371 14476 371 0 S4BEG[2]
rlabel metal3 14784 2044 14784 2044 0 S4BEG[3]
rlabel metal2 14700 287 14700 287 0 S4BEG[4]
rlabel metal2 14812 343 14812 343 0 S4BEG[5]
rlabel metal2 14924 203 14924 203 0 S4BEG[6]
rlabel metal2 15036 539 15036 539 0 S4BEG[7]
rlabel metal3 15344 2436 15344 2436 0 S4BEG[8]
rlabel metal2 15260 175 15260 175 0 S4BEG[9]
rlabel metal2 16044 175 16044 175 0 SS4BEG[0]
rlabel metal2 17164 511 17164 511 0 SS4BEG[10]
rlabel metal2 17276 119 17276 119 0 SS4BEG[11]
rlabel metal2 17388 91 17388 91 0 SS4BEG[12]
rlabel metal2 17500 427 17500 427 0 SS4BEG[13]
rlabel metal2 17612 287 17612 287 0 SS4BEG[14]
rlabel metal2 17724 399 17724 399 0 SS4BEG[15]
rlabel metal2 16156 119 16156 119 0 SS4BEG[1]
rlabel metal2 16268 147 16268 147 0 SS4BEG[2]
rlabel metal2 16464 2324 16464 2324 0 SS4BEG[3]
rlabel metal2 16492 175 16492 175 0 SS4BEG[4]
rlabel metal2 16604 427 16604 427 0 SS4BEG[5]
rlabel metal2 16716 679 16716 679 0 SS4BEG[6]
rlabel metal2 16828 203 16828 203 0 SS4BEG[7]
rlabel metal2 16940 91 16940 91 0 SS4BEG[8]
rlabel metal2 17052 735 17052 735 0 SS4BEG[9]
rlabel metal3 17052 3836 17052 3836 0 UserCLK
rlabel metal2 924 6692 924 6692 0 UserCLKo
rlabel metal2 24332 1008 24332 1008 0 net1
rlabel metal2 3780 4564 3780 4564 0 net10
rlabel metal2 18452 2352 18452 2352 0 net100
rlabel metal2 18816 1372 18816 1372 0 net101
rlabel metal2 17612 2744 17612 2744 0 net102
rlabel metal2 20048 588 20048 588 0 net103
rlabel metal2 20412 2660 20412 2660 0 net104
rlabel metal2 2492 5824 2492 5824 0 net105
rlabel metal3 24332 4060 24332 4060 0 net11
rlabel metal2 23548 1428 23548 1428 0 net12
rlabel metal3 23996 4564 23996 4564 0 net13
rlabel metal2 25116 4816 25116 4816 0 net14
rlabel metal3 24724 3780 24724 3780 0 net15
rlabel metal2 24388 5264 24388 5264 0 net16
rlabel metal2 25088 6020 25088 6020 0 net17
rlabel metal2 3780 5768 3780 5768 0 net18
rlabel metal2 24164 4788 24164 4788 0 net19
rlabel metal3 24276 2212 24276 2212 0 net2
rlabel metal3 24108 4900 24108 4900 0 net20
rlabel metal2 24388 4788 24388 4788 0 net21
rlabel metal2 23464 5236 23464 5236 0 net22
rlabel metal2 23716 1148 23716 1148 0 net23
rlabel metal2 1372 6272 1372 6272 0 net24
rlabel metal3 24416 6076 24416 6076 0 net25
rlabel metal2 24388 952 24388 952 0 net26
rlabel metal2 24500 1316 24500 1316 0 net27
rlabel metal3 24500 980 24500 980 0 net28
rlabel metal2 22764 1148 22764 1148 0 net29
rlabel metal2 25592 644 25592 644 0 net3
rlabel metal2 25116 1568 25116 1568 0 net30
rlabel metal2 24388 2352 24388 2352 0 net31
rlabel metal3 2156 1428 2156 1428 0 net32
rlabel metal2 3052 6636 3052 6636 0 net33
rlabel metal2 14868 6300 14868 6300 0 net34
rlabel metal3 16716 6132 16716 6132 0 net35
rlabel metal3 18060 5348 18060 5348 0 net36
rlabel metal2 19040 5740 19040 5740 0 net37
rlabel metal2 19572 6300 19572 6300 0 net38
rlabel metal2 20860 6300 20860 6300 0 net39
rlabel metal3 24864 2604 24864 2604 0 net4
rlabel metal2 21476 4396 21476 4396 0 net40
rlabel metal2 23380 6300 23380 6300 0 net41
rlabel metal3 23744 6468 23744 6468 0 net42
rlabel metal3 22960 6020 22960 6020 0 net43
rlabel metal2 4004 6020 4004 6020 0 net44
rlabel metal2 5236 6048 5236 6048 0 net45
rlabel metal2 8820 6104 8820 6104 0 net46
rlabel metal4 13412 4770 13412 4770 0 net47
rlabel metal2 8932 6440 8932 6440 0 net48
rlabel metal2 12628 5880 12628 5880 0 net49
rlabel metal2 3332 2324 3332 2324 0 net5
rlabel metal2 11256 5348 11256 5348 0 net50
rlabel metal2 12516 6048 12516 6048 0 net51
rlabel metal2 13468 5908 13468 5908 0 net52
rlabel metal2 2660 2408 2660 2408 0 net53
rlabel metal2 3556 1148 3556 1148 0 net54
rlabel metal3 1876 3444 1876 3444 0 net55
rlabel metal2 2604 1568 2604 1568 0 net56
rlabel metal3 10220 1372 10220 1372 0 net57
rlabel metal2 6412 1372 6412 1372 0 net58
rlabel metal2 5908 2576 5908 2576 0 net59
rlabel metal2 2772 2828 2772 2828 0 net6
rlabel metal2 12628 1148 12628 1148 0 net60
rlabel metal2 4228 2800 4228 2800 0 net61
rlabel metal2 3948 2632 3948 2632 0 net62
rlabel metal2 3724 2408 3724 2408 0 net63
rlabel metal2 6356 2044 6356 2044 0 net64
rlabel metal2 13664 588 13664 588 0 net65
rlabel metal3 13636 588 13636 588 0 net66
rlabel metal2 9492 4032 9492 4032 0 net67
rlabel metal2 14644 672 14644 672 0 net68
rlabel metal3 9772 1148 9772 1148 0 net69
rlabel metal2 2156 4144 2156 4144 0 net7
rlabel metal3 12124 4648 12124 4648 0 net70
rlabel metal2 7084 2632 7084 2632 0 net71
rlabel metal2 15260 1344 15260 1344 0 net72
rlabel metal2 15764 336 15764 336 0 net73
rlabel metal2 8988 1260 8988 1260 0 net74
rlabel metal3 16100 2716 16100 2716 0 net75
rlabel metal3 16996 2604 16996 2604 0 net76
rlabel metal3 17248 1428 17248 1428 0 net77
rlabel metal3 19012 980 19012 980 0 net78
rlabel metal2 17920 3276 17920 3276 0 net79
rlabel metal2 25228 3192 25228 3192 0 net8
rlabel metal2 15036 1512 15036 1512 0 net80
rlabel metal2 14924 2744 14924 2744 0 net81
rlabel metal3 13272 2156 13272 2156 0 net82
rlabel metal2 15876 756 15876 756 0 net83
rlabel metal2 15820 1484 15820 1484 0 net84
rlabel metal2 16212 1176 16212 1176 0 net85
rlabel metal3 11144 3892 11144 3892 0 net86
rlabel metal3 10584 3164 10584 3164 0 net87
rlabel metal3 12628 2072 12628 2072 0 net88
rlabel metal3 15652 2548 15652 2548 0 net89
rlabel metal3 24920 4116 24920 4116 0 net9
rlabel metal2 20804 2352 20804 2352 0 net90
rlabel metal2 18396 2940 18396 2940 0 net91
rlabel metal3 20552 1372 20552 1372 0 net92
rlabel metal2 22372 3108 22372 3108 0 net93
rlabel metal2 23884 1708 23884 1708 0 net94
rlabel metal2 24948 2772 24948 2772 0 net95
rlabel metal2 18508 756 18508 756 0 net96
rlabel metal2 17164 2716 17164 2716 0 net97
rlabel metal2 14532 2352 14532 2352 0 net98
rlabel metal2 18536 1036 18536 1036 0 net99
<< properties >>
string FIXED_BBOX 0 0 26376 7112
<< end >>
