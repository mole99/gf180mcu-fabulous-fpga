magic
tech gf180mcuD
magscale 1 10
timestamp 1764324324
<< metal1 >>
rect 672 56474 27888 56508
rect 672 56422 3806 56474
rect 3858 56422 3910 56474
rect 3962 56422 4014 56474
rect 4066 56422 23806 56474
rect 23858 56422 23910 56474
rect 23962 56422 24014 56474
rect 24066 56422 27888 56474
rect 672 56388 27888 56422
rect 3614 56306 3666 56318
rect 3614 56242 3666 56254
rect 5518 56306 5570 56318
rect 5518 56242 5570 56254
rect 8990 56306 9042 56318
rect 8990 56242 9042 56254
rect 10558 56306 10610 56318
rect 10558 56242 10610 56254
rect 13022 56306 13074 56318
rect 13022 56242 13074 56254
rect 14590 56306 14642 56318
rect 14590 56242 14642 56254
rect 16494 56306 16546 56318
rect 16494 56242 16546 56254
rect 18510 56306 18562 56318
rect 18510 56242 18562 56254
rect 20638 56306 20690 56318
rect 20638 56242 20690 56254
rect 21870 56306 21922 56318
rect 21870 56242 21922 56254
rect 24446 56306 24498 56318
rect 24446 56242 24498 56254
rect 26014 56306 26066 56318
rect 26014 56242 26066 56254
rect 7410 56142 7422 56194
rect 7474 56142 7486 56194
rect 5170 56030 5182 56082
rect 5234 56030 5246 56082
rect 20178 56030 20190 56082
rect 20242 56030 20254 56082
rect 25666 56030 25678 56082
rect 25730 56030 25742 56082
rect 1026 55918 1038 55970
rect 1090 55918 1102 55970
rect 3042 55918 3054 55970
rect 3106 55918 3118 55970
rect 8082 55918 8094 55970
rect 8146 55918 8158 55970
rect 9986 55918 9998 55970
rect 10050 55918 10062 55970
rect 11554 55918 11566 55970
rect 11618 55918 11630 55970
rect 14018 55918 14030 55970
rect 14082 55918 14094 55970
rect 15586 55918 15598 55970
rect 15650 55918 15662 55970
rect 17490 55918 17502 55970
rect 17554 55918 17566 55970
rect 19506 55918 19518 55970
rect 19570 55918 19582 55970
rect 22866 55918 22878 55970
rect 22930 55918 22942 55970
rect 23874 55918 23886 55970
rect 23938 55918 23950 55970
rect 1374 55858 1426 55870
rect 1374 55794 1426 55806
rect 672 55690 27888 55724
rect 672 55638 4466 55690
rect 4518 55638 4570 55690
rect 4622 55638 4674 55690
rect 4726 55638 24466 55690
rect 24518 55638 24570 55690
rect 24622 55638 24674 55690
rect 24726 55638 27888 55690
rect 672 55604 27888 55638
rect 18846 55410 18898 55422
rect 21634 55358 21646 55410
rect 21698 55358 21710 55410
rect 18846 55346 18898 55358
rect 19406 55298 19458 55310
rect 20526 55298 20578 55310
rect 3490 55246 3502 55298
rect 3554 55246 3566 55298
rect 7522 55246 7534 55298
rect 7586 55246 7598 55298
rect 12898 55246 12910 55298
rect 12962 55246 12974 55298
rect 18274 55246 18286 55298
rect 18338 55246 18350 55298
rect 20066 55246 20078 55298
rect 20130 55246 20142 55298
rect 20962 55246 20974 55298
rect 21026 55246 21038 55298
rect 23650 55246 23662 55298
rect 23714 55246 23726 55298
rect 24882 55246 24894 55298
rect 24946 55246 24958 55298
rect 26226 55246 26238 55298
rect 26290 55246 26302 55298
rect 19406 55234 19458 55246
rect 20526 55234 20578 55246
rect 2494 55186 2546 55198
rect 2494 55122 2546 55134
rect 6526 55186 6578 55198
rect 6526 55122 6578 55134
rect 11902 55186 11954 55198
rect 11902 55122 11954 55134
rect 17278 55186 17330 55198
rect 17278 55122 17330 55134
rect 22654 55186 22706 55198
rect 25554 55134 25566 55186
rect 25618 55134 25630 55186
rect 22654 55122 22706 55134
rect 27246 55074 27298 55086
rect 27246 55010 27298 55022
rect 672 54906 27888 54940
rect 672 54854 3806 54906
rect 3858 54854 3910 54906
rect 3962 54854 4014 54906
rect 4066 54854 23806 54906
rect 23858 54854 23910 54906
rect 23962 54854 24014 54906
rect 24066 54854 27888 54906
rect 672 54820 27888 54854
rect 22542 54738 22594 54750
rect 22542 54674 22594 54686
rect 24110 54738 24162 54750
rect 24110 54674 24162 54686
rect 19518 54626 19570 54638
rect 21074 54574 21086 54626
rect 21138 54574 21150 54626
rect 25442 54574 25454 54626
rect 25506 54574 25518 54626
rect 19518 54562 19570 54574
rect 21522 54350 21534 54402
rect 21586 54350 21598 54402
rect 23090 54350 23102 54402
rect 23154 54350 23166 54402
rect 24658 54350 24670 54402
rect 24722 54350 24734 54402
rect 26226 54350 26238 54402
rect 26290 54350 26302 54402
rect 27010 54350 27022 54402
rect 27074 54350 27086 54402
rect 18958 54290 19010 54302
rect 18958 54226 19010 54238
rect 20638 54290 20690 54302
rect 20638 54226 20690 54238
rect 672 54122 27888 54156
rect 672 54070 4466 54122
rect 4518 54070 4570 54122
rect 4622 54070 4674 54122
rect 4726 54070 24466 54122
rect 24518 54070 24570 54122
rect 24622 54070 24674 54122
rect 24726 54070 27888 54122
rect 672 54036 27888 54070
rect 1038 53730 1090 53742
rect 1038 53666 1090 53678
rect 20526 53730 20578 53742
rect 20526 53666 20578 53678
rect 20862 53730 20914 53742
rect 21858 53678 21870 53730
rect 21922 53678 21934 53730
rect 22866 53678 22878 53730
rect 22930 53678 22942 53730
rect 24658 53678 24670 53730
rect 24722 53678 24734 53730
rect 26226 53678 26238 53730
rect 26290 53678 26302 53730
rect 20862 53666 20914 53678
rect 19966 53618 20018 53630
rect 23774 53618 23826 53630
rect 1474 53566 1486 53618
rect 1538 53566 1550 53618
rect 21298 53566 21310 53618
rect 21362 53566 21374 53618
rect 22194 53566 22206 53618
rect 22258 53566 22270 53618
rect 25554 53566 25566 53618
rect 25618 53566 25630 53618
rect 19966 53554 20018 53566
rect 23774 53554 23826 53566
rect 27246 53506 27298 53518
rect 27246 53442 27298 53454
rect 672 53338 27888 53372
rect 672 53286 3806 53338
rect 3858 53286 3910 53338
rect 3962 53286 4014 53338
rect 4066 53286 23806 53338
rect 23858 53286 23910 53338
rect 23962 53286 24014 53338
rect 24066 53286 27888 53338
rect 672 53252 27888 53286
rect 24110 53170 24162 53182
rect 24110 53106 24162 53118
rect 21746 53006 21758 53058
rect 21810 53006 21822 53058
rect 22642 53006 22654 53058
rect 22706 53006 22718 53058
rect 27122 53006 27134 53058
rect 27186 53006 27198 53058
rect 1598 52834 1650 52846
rect 1598 52770 1650 52782
rect 21310 52834 21362 52846
rect 23090 52782 23102 52834
rect 23154 52782 23166 52834
rect 24658 52782 24670 52834
rect 24722 52782 24734 52834
rect 25442 52782 25454 52834
rect 25506 52782 25518 52834
rect 26226 52782 26238 52834
rect 26290 52782 26302 52834
rect 21310 52770 21362 52782
rect 1038 52722 1090 52734
rect 1038 52658 1090 52670
rect 22206 52722 22258 52734
rect 22206 52658 22258 52670
rect 672 52554 27888 52588
rect 672 52502 4466 52554
rect 4518 52502 4570 52554
rect 4622 52502 4674 52554
rect 4726 52502 24466 52554
rect 24518 52502 24570 52554
rect 24622 52502 24674 52554
rect 24726 52502 27888 52554
rect 672 52468 27888 52502
rect 21870 52274 21922 52286
rect 22754 52222 22766 52274
rect 22818 52222 22830 52274
rect 23538 52222 23550 52274
rect 23602 52222 23614 52274
rect 24658 52222 24670 52274
rect 24722 52222 24734 52274
rect 21870 52210 21922 52222
rect 22430 52162 22482 52174
rect 26226 52110 26238 52162
rect 26290 52110 26302 52162
rect 22430 52098 22482 52110
rect 25554 51998 25566 52050
rect 25618 51998 25630 52050
rect 27246 51938 27298 51950
rect 27246 51874 27298 51886
rect 672 51770 27888 51804
rect 672 51718 3806 51770
rect 3858 51718 3910 51770
rect 3962 51718 4014 51770
rect 4066 51718 23806 51770
rect 23858 51718 23910 51770
rect 23962 51718 24014 51770
rect 24066 51718 27888 51770
rect 672 51684 27888 51718
rect 24334 51490 24386 51502
rect 1474 51438 1486 51490
rect 1538 51438 1550 51490
rect 23202 51438 23214 51490
rect 23266 51438 23278 51490
rect 25330 51438 25342 51490
rect 25394 51438 25406 51490
rect 24334 51426 24386 51438
rect 24882 51326 24894 51378
rect 24946 51326 24958 51378
rect 26226 51214 26238 51266
rect 26290 51214 26302 51266
rect 27010 51214 27022 51266
rect 27074 51214 27086 51266
rect 1038 51154 1090 51166
rect 1038 51090 1090 51102
rect 22766 51154 22818 51166
rect 22766 51090 22818 51102
rect 23774 51154 23826 51166
rect 23774 51090 23826 51102
rect 672 50986 27888 51020
rect 672 50934 4466 50986
rect 4518 50934 4570 50986
rect 4622 50934 4674 50986
rect 4726 50934 24466 50986
rect 24518 50934 24570 50986
rect 24622 50934 24674 50986
rect 24726 50934 27888 50986
rect 672 50900 27888 50934
rect 23438 50706 23490 50718
rect 26226 50654 26238 50706
rect 26290 50654 26302 50706
rect 23438 50642 23490 50654
rect 23874 50542 23886 50594
rect 23938 50542 23950 50594
rect 24658 50542 24670 50594
rect 24722 50542 24734 50594
rect 25554 50430 25566 50482
rect 25618 50430 25630 50482
rect 27246 50370 27298 50382
rect 27246 50306 27298 50318
rect 672 50202 27888 50236
rect 672 50150 3806 50202
rect 3858 50150 3910 50202
rect 3962 50150 4014 50202
rect 4066 50150 23806 50202
rect 23858 50150 23910 50202
rect 23962 50150 24014 50202
rect 24066 50150 27888 50202
rect 672 50116 27888 50150
rect 24210 49870 24222 49922
rect 24274 49870 24286 49922
rect 27122 49870 27134 49922
rect 27186 49870 27198 49922
rect 24882 49758 24894 49810
rect 24946 49758 24958 49810
rect 26338 49758 26350 49810
rect 26402 49758 26414 49810
rect 1598 49698 1650 49710
rect 25442 49646 25454 49698
rect 25506 49646 25518 49698
rect 1598 49634 1650 49646
rect 1038 49586 1090 49598
rect 1038 49522 1090 49534
rect 23774 49586 23826 49598
rect 23774 49522 23826 49534
rect 672 49418 27888 49452
rect 672 49366 4466 49418
rect 4518 49366 4570 49418
rect 4622 49366 4674 49418
rect 4726 49366 24466 49418
rect 24518 49366 24570 49418
rect 24622 49366 24674 49418
rect 24726 49366 27888 49418
rect 672 49332 27888 49366
rect 1038 49026 1090 49038
rect 24658 48974 24670 49026
rect 24722 48974 24734 49026
rect 26226 48974 26238 49026
rect 26290 48974 26302 49026
rect 1038 48962 1090 48974
rect 1598 48914 1650 48926
rect 25554 48862 25566 48914
rect 25618 48862 25630 48914
rect 1598 48850 1650 48862
rect 27246 48802 27298 48814
rect 27246 48738 27298 48750
rect 672 48634 27888 48668
rect 672 48582 3806 48634
rect 3858 48582 3910 48634
rect 3962 48582 4014 48634
rect 4066 48582 23806 48634
rect 23858 48582 23910 48634
rect 23962 48582 24014 48634
rect 24066 48582 27888 48634
rect 672 48548 27888 48582
rect 25778 48302 25790 48354
rect 25842 48302 25854 48354
rect 25006 48130 25058 48142
rect 26226 48078 26238 48130
rect 26290 48078 26302 48130
rect 27010 48078 27022 48130
rect 27074 48078 27086 48130
rect 25006 48066 25058 48078
rect 24446 48018 24498 48030
rect 24446 47954 24498 47966
rect 25342 48018 25394 48030
rect 25342 47954 25394 47966
rect 672 47850 27888 47884
rect 672 47798 4466 47850
rect 4518 47798 4570 47850
rect 4622 47798 4674 47850
rect 4726 47798 24466 47850
rect 24518 47798 24570 47850
rect 24622 47798 24674 47850
rect 24726 47798 27888 47850
rect 672 47764 27888 47798
rect 1038 47458 1090 47470
rect 24658 47406 24670 47458
rect 24722 47406 24734 47458
rect 26226 47406 26238 47458
rect 26290 47406 26302 47458
rect 1038 47394 1090 47406
rect 1598 47346 1650 47358
rect 1598 47282 1650 47294
rect 25678 47346 25730 47358
rect 25678 47282 25730 47294
rect 27246 47234 27298 47246
rect 27246 47170 27298 47182
rect 672 47066 27888 47100
rect 672 47014 3806 47066
rect 3858 47014 3910 47066
rect 3962 47014 4014 47066
rect 4066 47014 23806 47066
rect 23858 47014 23910 47066
rect 23962 47014 24014 47066
rect 24066 47014 27888 47066
rect 672 46980 27888 47014
rect 25678 46786 25730 46798
rect 27122 46734 27134 46786
rect 27186 46734 27198 46786
rect 25678 46722 25730 46734
rect 24658 46510 24670 46562
rect 24722 46510 24734 46562
rect 26226 46510 26238 46562
rect 26290 46510 26302 46562
rect 672 46282 27888 46316
rect 672 46230 4466 46282
rect 4518 46230 4570 46282
rect 4622 46230 4674 46282
rect 4726 46230 24466 46282
rect 24518 46230 24570 46282
rect 24622 46230 24674 46282
rect 24726 46230 27888 46282
rect 672 46196 27888 46230
rect 1038 45890 1090 45902
rect 24770 45838 24782 45890
rect 24834 45838 24846 45890
rect 26450 45838 26462 45890
rect 26514 45838 26526 45890
rect 1038 45826 1090 45838
rect 1474 45726 1486 45778
rect 1538 45726 1550 45778
rect 25678 45666 25730 45678
rect 25678 45602 25730 45614
rect 27246 45666 27298 45678
rect 27246 45602 27298 45614
rect 672 45498 27888 45532
rect 672 45446 3806 45498
rect 3858 45446 3910 45498
rect 3962 45446 4014 45498
rect 4066 45446 23806 45498
rect 23858 45446 23910 45498
rect 23962 45446 24014 45498
rect 24066 45446 27888 45498
rect 672 45412 27888 45446
rect 26338 45054 26350 45106
rect 26402 45054 26414 45106
rect 27010 44942 27022 44994
rect 27074 44942 27086 44994
rect 672 44714 27888 44748
rect 672 44662 4466 44714
rect 4518 44662 4570 44714
rect 4622 44662 4674 44714
rect 4726 44662 24466 44714
rect 24518 44662 24570 44714
rect 24622 44662 24674 44714
rect 24726 44662 27888 44714
rect 672 44628 27888 44662
rect 1038 44322 1090 44334
rect 24658 44270 24670 44322
rect 24722 44270 24734 44322
rect 26226 44270 26238 44322
rect 26290 44270 26302 44322
rect 1038 44258 1090 44270
rect 25678 44210 25730 44222
rect 1474 44158 1486 44210
rect 1538 44158 1550 44210
rect 25678 44146 25730 44158
rect 27246 44098 27298 44110
rect 27246 44034 27298 44046
rect 672 43930 27888 43964
rect 672 43878 3806 43930
rect 3858 43878 3910 43930
rect 3962 43878 4014 43930
rect 4066 43878 23806 43930
rect 23858 43878 23910 43930
rect 23962 43878 24014 43930
rect 24066 43878 27888 43930
rect 672 43844 27888 43878
rect 25678 43650 25730 43662
rect 27122 43598 27134 43650
rect 27186 43598 27198 43650
rect 25678 43586 25730 43598
rect 24882 43486 24894 43538
rect 24946 43486 24958 43538
rect 1598 43426 1650 43438
rect 26226 43374 26238 43426
rect 26290 43374 26302 43426
rect 1598 43362 1650 43374
rect 1038 43314 1090 43326
rect 1038 43250 1090 43262
rect 672 43146 27888 43180
rect 672 43094 4466 43146
rect 4518 43094 4570 43146
rect 4622 43094 4674 43146
rect 4726 43094 24466 43146
rect 24518 43094 24570 43146
rect 24622 43094 24674 43146
rect 24726 43094 27888 43146
rect 672 43060 27888 43094
rect 1138 42702 1150 42754
rect 1202 42702 1214 42754
rect 24658 42702 24670 42754
rect 24722 42702 24734 42754
rect 26226 42702 26238 42754
rect 26290 42702 26302 42754
rect 1598 42642 1650 42654
rect 1598 42578 1650 42590
rect 25678 42530 25730 42542
rect 25678 42466 25730 42478
rect 27246 42530 27298 42542
rect 27246 42466 27298 42478
rect 672 42362 27888 42396
rect 672 42310 3806 42362
rect 3858 42310 3910 42362
rect 3962 42310 4014 42362
rect 4066 42310 23806 42362
rect 23858 42310 23910 42362
rect 23962 42310 24014 42362
rect 24066 42310 27888 42362
rect 672 42276 27888 42310
rect 3614 41970 3666 41982
rect 16258 41918 16270 41970
rect 16322 41918 16334 41970
rect 3614 41906 3666 41918
rect 1598 41858 1650 41870
rect 1598 41794 1650 41806
rect 4174 41858 4226 41870
rect 18386 41806 18398 41858
rect 18450 41806 18462 41858
rect 26226 41806 26238 41858
rect 26290 41806 26302 41858
rect 27010 41806 27022 41858
rect 27074 41806 27086 41858
rect 4174 41794 4226 41806
rect 1038 41746 1090 41758
rect 1038 41682 1090 41694
rect 672 41578 27888 41612
rect 672 41526 4466 41578
rect 4518 41526 4570 41578
rect 4622 41526 4674 41578
rect 4726 41526 24466 41578
rect 24518 41526 24570 41578
rect 24622 41526 24674 41578
rect 24726 41526 27888 41578
rect 672 41492 27888 41526
rect 6078 41410 6130 41422
rect 6078 41346 6130 41358
rect 2046 41298 2098 41310
rect 2046 41234 2098 41246
rect 2606 41298 2658 41310
rect 6638 41298 6690 41310
rect 4274 41246 4286 41298
rect 4338 41246 4350 41298
rect 10546 41246 10558 41298
rect 10610 41246 10622 41298
rect 2606 41234 2658 41246
rect 6638 41234 6690 41246
rect 1038 41186 1090 41198
rect 8878 41186 8930 41198
rect 3826 41134 3838 41186
rect 3890 41134 3902 41186
rect 10098 41134 10110 41186
rect 10162 41134 10174 41186
rect 24658 41134 24670 41186
rect 24722 41134 24734 41186
rect 26226 41134 26238 41186
rect 26290 41134 26302 41186
rect 1038 41122 1090 41134
rect 8878 41122 8930 41134
rect 25678 41074 25730 41086
rect 1474 41022 1486 41074
rect 1538 41022 1550 41074
rect 9314 41022 9326 41074
rect 9378 41022 9390 41074
rect 25678 41010 25730 41022
rect 5518 40962 5570 40974
rect 5518 40898 5570 40910
rect 11790 40962 11842 40974
rect 11790 40898 11842 40910
rect 27246 40962 27298 40974
rect 27246 40898 27298 40910
rect 672 40794 27888 40828
rect 672 40742 3806 40794
rect 3858 40742 3910 40794
rect 3962 40742 4014 40794
rect 4066 40742 23806 40794
rect 23858 40742 23910 40794
rect 23962 40742 24014 40794
rect 24066 40742 27888 40794
rect 672 40708 27888 40742
rect 2158 40514 2210 40526
rect 2158 40450 2210 40462
rect 6974 40514 7026 40526
rect 25678 40514 25730 40526
rect 13346 40462 13358 40514
rect 13410 40462 13422 40514
rect 15474 40462 15486 40514
rect 15538 40462 15550 40514
rect 27122 40462 27134 40514
rect 27186 40462 27198 40514
rect 6974 40450 7026 40462
rect 25678 40450 25730 40462
rect 4286 40402 4338 40414
rect 8766 40402 8818 40414
rect 1698 40350 1710 40402
rect 1762 40350 1774 40402
rect 2594 40350 2606 40402
rect 2658 40350 2670 40402
rect 7634 40350 7646 40402
rect 7698 40350 7710 40402
rect 8082 40350 8094 40402
rect 8146 40350 8158 40402
rect 9538 40350 9550 40402
rect 9602 40350 9614 40402
rect 10434 40350 10446 40402
rect 10498 40350 10510 40402
rect 17714 40350 17726 40402
rect 17778 40350 17790 40402
rect 18386 40350 18398 40402
rect 18450 40350 18462 40402
rect 24658 40350 24670 40402
rect 24722 40350 24734 40402
rect 26450 40350 26462 40402
rect 26514 40350 26526 40402
rect 4286 40338 4338 40350
rect 8766 40338 8818 40350
rect 7310 40290 7362 40302
rect 3042 40238 3054 40290
rect 3106 40238 3118 40290
rect 8306 40238 8318 40290
rect 8370 40238 8382 40290
rect 7310 40226 7362 40238
rect 6414 40178 6466 40190
rect 6414 40114 6466 40126
rect 12910 40178 12962 40190
rect 12910 40114 12962 40126
rect 672 40010 27888 40044
rect 672 39958 4466 40010
rect 4518 39958 4570 40010
rect 4622 39958 4674 40010
rect 4726 39958 24466 40010
rect 24518 39958 24570 40010
rect 24622 39958 24674 40010
rect 24726 39958 27888 40010
rect 672 39924 27888 39958
rect 6066 39790 6078 39842
rect 6130 39790 6142 39842
rect 9874 39790 9886 39842
rect 9938 39790 9950 39842
rect 12450 39790 12462 39842
rect 12514 39790 12526 39842
rect 2494 39730 2546 39742
rect 2494 39666 2546 39678
rect 5070 39730 5122 39742
rect 5070 39666 5122 39678
rect 12910 39730 12962 39742
rect 12910 39666 12962 39678
rect 6750 39618 6802 39630
rect 11006 39618 11058 39630
rect 1138 39566 1150 39618
rect 1202 39566 1214 39618
rect 2034 39566 2046 39618
rect 2098 39566 2110 39618
rect 5506 39566 5518 39618
rect 5570 39566 5582 39618
rect 5842 39566 5854 39618
rect 5906 39566 5918 39618
rect 7074 39566 7086 39618
rect 7138 39566 7150 39618
rect 7298 39566 7310 39618
rect 7362 39566 7374 39618
rect 8194 39566 8206 39618
rect 8258 39566 8270 39618
rect 9426 39566 9438 39618
rect 9490 39566 9502 39618
rect 11778 39566 11790 39618
rect 11842 39566 11854 39618
rect 12338 39566 12350 39618
rect 12402 39566 12414 39618
rect 13570 39566 13582 39618
rect 13634 39566 13646 39618
rect 14578 39566 14590 39618
rect 14642 39566 14654 39618
rect 16706 39566 16718 39618
rect 16770 39566 16782 39618
rect 24882 39566 24894 39618
rect 24946 39566 24958 39618
rect 26226 39566 26238 39618
rect 26290 39566 26302 39618
rect 6750 39554 6802 39566
rect 11006 39554 11058 39566
rect 11454 39506 11506 39518
rect 1474 39454 1486 39506
rect 1538 39454 1550 39506
rect 18722 39454 18734 39506
rect 18786 39454 18798 39506
rect 11454 39442 11506 39454
rect 25678 39394 25730 39406
rect 25678 39330 25730 39342
rect 27246 39394 27298 39406
rect 27246 39330 27298 39342
rect 672 39226 27888 39260
rect 672 39174 3806 39226
rect 3858 39174 3910 39226
rect 3962 39174 4014 39226
rect 4066 39174 23806 39226
rect 23858 39174 23910 39226
rect 23962 39174 24014 39226
rect 24066 39174 27888 39226
rect 672 39140 27888 39174
rect 7198 39058 7250 39070
rect 7198 38994 7250 39006
rect 13346 38894 13358 38946
rect 13410 38894 13422 38946
rect 12910 38834 12962 38846
rect 2706 38782 2718 38834
rect 2770 38782 2782 38834
rect 5506 38782 5518 38834
rect 5570 38782 5582 38834
rect 10546 38782 10558 38834
rect 10610 38782 10622 38834
rect 15250 38782 15262 38834
rect 15314 38782 15326 38834
rect 12910 38770 12962 38782
rect 1598 38722 1650 38734
rect 4286 38722 4338 38734
rect 3042 38670 3054 38722
rect 3106 38670 3118 38722
rect 5954 38670 5966 38722
rect 6018 38670 6030 38722
rect 18610 38670 18622 38722
rect 18674 38670 18686 38722
rect 26226 38670 26238 38722
rect 26290 38670 26302 38722
rect 27010 38670 27022 38722
rect 27074 38670 27086 38722
rect 1598 38658 1650 38670
rect 4286 38658 4338 38670
rect 1038 38610 1090 38622
rect 12126 38610 12178 38622
rect 10994 38558 11006 38610
rect 11058 38558 11070 38610
rect 1038 38546 1090 38558
rect 12126 38546 12178 38558
rect 672 38442 27888 38476
rect 672 38390 4466 38442
rect 4518 38390 4570 38442
rect 4622 38390 4674 38442
rect 4726 38390 24466 38442
rect 24518 38390 24570 38442
rect 24622 38390 24674 38442
rect 24726 38390 27888 38442
rect 672 38356 27888 38390
rect 6302 38274 6354 38286
rect 12562 38222 12574 38274
rect 12626 38222 12638 38274
rect 15138 38222 15150 38274
rect 15202 38222 15214 38274
rect 6302 38210 6354 38222
rect 3838 38162 3890 38174
rect 7758 38162 7810 38174
rect 2258 38110 2270 38162
rect 2322 38110 2334 38162
rect 5058 38110 5070 38162
rect 5122 38110 5134 38162
rect 9986 38110 9998 38162
rect 10050 38110 10062 38162
rect 3838 38098 3890 38110
rect 7758 38098 7810 38110
rect 6750 38050 6802 38062
rect 3378 37998 3390 38050
rect 3442 37998 3454 38050
rect 4610 37998 4622 38050
rect 4674 37998 4686 38050
rect 6750 37986 6802 37998
rect 8318 38050 8370 38062
rect 11118 38050 11170 38062
rect 15486 38050 15538 38062
rect 9426 37998 9438 38050
rect 9490 37998 9502 38050
rect 11890 37998 11902 38050
rect 11954 37998 11966 38050
rect 12450 37998 12462 38050
rect 12514 37998 12526 38050
rect 13122 37998 13134 38050
rect 13186 37998 13198 38050
rect 13570 37998 13582 38050
rect 13634 37998 13646 38050
rect 14690 37998 14702 38050
rect 14754 37998 14766 38050
rect 16706 37998 16718 38050
rect 16770 37998 16782 38050
rect 17490 37998 17502 38050
rect 17554 37998 17566 38050
rect 24658 37998 24670 38050
rect 24722 37998 24734 38050
rect 26226 37998 26238 38050
rect 26290 37998 26302 38050
rect 8318 37986 8370 37998
rect 11118 37986 11170 37998
rect 15486 37986 15538 37998
rect 11566 37938 11618 37950
rect 25678 37938 25730 37950
rect 2706 37886 2718 37938
rect 2770 37886 2782 37938
rect 7186 37886 7198 37938
rect 7250 37886 7262 37938
rect 19730 37886 19742 37938
rect 19794 37886 19806 37938
rect 11566 37874 11618 37886
rect 25678 37874 25730 37886
rect 1150 37826 1202 37838
rect 1150 37762 1202 37774
rect 27246 37826 27298 37838
rect 27246 37762 27298 37774
rect 672 37658 27888 37692
rect 672 37606 3806 37658
rect 3858 37606 3910 37658
rect 3962 37606 4014 37658
rect 4066 37606 23806 37658
rect 23858 37606 23910 37658
rect 23962 37606 24014 37658
rect 24066 37606 27888 37658
rect 672 37572 27888 37606
rect 6750 37490 6802 37502
rect 6750 37426 6802 37438
rect 2494 37378 2546 37390
rect 3266 37326 3278 37378
rect 3330 37326 3342 37378
rect 16258 37326 16270 37378
rect 16322 37326 16334 37378
rect 27122 37326 27134 37378
rect 27186 37326 27198 37378
rect 2494 37314 2546 37326
rect 8990 37266 9042 37278
rect 1138 37214 1150 37266
rect 1202 37214 1214 37266
rect 5170 37214 5182 37266
rect 5234 37214 5246 37266
rect 7858 37214 7870 37266
rect 7922 37214 7934 37266
rect 8306 37214 8318 37266
rect 8370 37214 8382 37266
rect 9538 37214 9550 37266
rect 9602 37214 9614 37266
rect 10658 37214 10670 37266
rect 10722 37214 10734 37266
rect 18610 37214 18622 37266
rect 18674 37214 18686 37266
rect 24882 37214 24894 37266
rect 24946 37214 24958 37266
rect 8990 37202 9042 37214
rect 1598 37154 1650 37166
rect 7534 37154 7586 37166
rect 5506 37102 5518 37154
rect 5570 37102 5582 37154
rect 8530 37102 8542 37154
rect 8594 37102 8606 37154
rect 16594 37102 16606 37154
rect 16658 37102 16670 37154
rect 25442 37102 25454 37154
rect 25506 37102 25518 37154
rect 26226 37102 26238 37154
rect 26290 37102 26302 37154
rect 1598 37090 1650 37102
rect 7534 37090 7586 37102
rect 1934 37042 1986 37054
rect 1934 36978 1986 36990
rect 2830 37042 2882 37054
rect 2830 36978 2882 36990
rect 672 36874 27888 36908
rect 672 36822 4466 36874
rect 4518 36822 4570 36874
rect 4622 36822 4674 36874
rect 4726 36822 24466 36874
rect 24518 36822 24570 36874
rect 24622 36822 24674 36874
rect 24726 36822 27888 36874
rect 672 36788 27888 36822
rect 1698 36654 1710 36706
rect 1762 36654 1774 36706
rect 3938 36654 3950 36706
rect 4002 36654 4014 36706
rect 18846 36594 18898 36606
rect 10098 36542 10110 36594
rect 10162 36542 10174 36594
rect 12226 36542 12238 36594
rect 12290 36542 12302 36594
rect 15698 36542 15710 36594
rect 15762 36542 15774 36594
rect 18846 36530 18898 36542
rect 6190 36482 6242 36494
rect 1250 36430 1262 36482
rect 1314 36430 1326 36482
rect 6190 36418 6242 36430
rect 8318 36482 8370 36494
rect 8318 36418 8370 36430
rect 14366 36482 14418 36494
rect 14366 36418 14418 36430
rect 14814 36482 14866 36494
rect 18286 36482 18338 36494
rect 15922 36430 15934 36482
rect 15986 36430 15998 36482
rect 17826 36430 17838 36482
rect 17890 36430 17902 36482
rect 24658 36430 24670 36482
rect 24722 36430 24734 36482
rect 26338 36430 26350 36482
rect 26402 36430 26414 36482
rect 14814 36418 14866 36430
rect 18286 36418 18338 36430
rect 7758 36370 7810 36382
rect 3490 36318 3502 36370
rect 3554 36318 3566 36370
rect 6626 36318 6638 36370
rect 6690 36318 6702 36370
rect 10546 36318 10558 36370
rect 10610 36318 10622 36370
rect 11778 36318 11790 36370
rect 11842 36318 11854 36370
rect 13906 36318 13918 36370
rect 13970 36318 13982 36370
rect 17042 36318 17054 36370
rect 17106 36318 17118 36370
rect 7758 36306 7810 36318
rect 2830 36258 2882 36270
rect 2830 36194 2882 36206
rect 5070 36258 5122 36270
rect 5070 36194 5122 36206
rect 8990 36258 9042 36270
rect 8990 36194 9042 36206
rect 13358 36258 13410 36270
rect 13358 36194 13410 36206
rect 15150 36258 15202 36270
rect 15150 36194 15202 36206
rect 25678 36258 25730 36270
rect 25678 36194 25730 36206
rect 27246 36258 27298 36270
rect 27246 36194 27298 36206
rect 672 36090 27888 36124
rect 672 36038 3806 36090
rect 3858 36038 3910 36090
rect 3962 36038 4014 36090
rect 4066 36038 23806 36090
rect 23858 36038 23910 36090
rect 23962 36038 24014 36090
rect 24066 36038 27888 36090
rect 672 36004 27888 36038
rect 11454 35810 11506 35822
rect 5842 35758 5854 35810
rect 5906 35758 5918 35810
rect 12898 35758 12910 35810
rect 12962 35758 12974 35810
rect 15474 35758 15486 35810
rect 15538 35758 15550 35810
rect 11454 35746 11506 35758
rect 9326 35698 9378 35710
rect 2594 35646 2606 35698
rect 2658 35646 2670 35698
rect 8194 35646 8206 35698
rect 8258 35646 8270 35698
rect 8642 35646 8654 35698
rect 8706 35646 8718 35698
rect 9874 35646 9886 35698
rect 9938 35646 9950 35698
rect 10882 35646 10894 35698
rect 10946 35646 10958 35698
rect 11890 35646 11902 35698
rect 11954 35646 11966 35698
rect 18386 35646 18398 35698
rect 18450 35646 18462 35698
rect 26338 35646 26350 35698
rect 26402 35646 26414 35698
rect 9326 35634 9378 35646
rect 1598 35586 1650 35598
rect 1598 35522 1650 35534
rect 7870 35586 7922 35598
rect 13358 35586 13410 35598
rect 8866 35534 8878 35586
rect 8930 35534 8942 35586
rect 27010 35534 27022 35586
rect 27074 35534 27086 35586
rect 7870 35522 7922 35534
rect 13358 35522 13410 35534
rect 1038 35474 1090 35486
rect 4286 35474 4338 35486
rect 7422 35474 7474 35486
rect 3154 35422 3166 35474
rect 3218 35422 3230 35474
rect 6290 35422 6302 35474
rect 6354 35422 6366 35474
rect 1038 35410 1090 35422
rect 4286 35410 4338 35422
rect 7422 35410 7474 35422
rect 672 35306 27888 35340
rect 672 35254 4466 35306
rect 4518 35254 4570 35306
rect 4622 35254 4674 35306
rect 4726 35254 24466 35306
rect 24518 35254 24570 35306
rect 24622 35254 24674 35306
rect 24726 35254 27888 35306
rect 672 35220 27888 35254
rect 16830 35138 16882 35150
rect 19854 35138 19906 35150
rect 6066 35086 6078 35138
rect 6130 35086 6142 35138
rect 10994 35086 11006 35138
rect 11058 35086 11070 35138
rect 13570 35086 13582 35138
rect 13634 35086 13646 35138
rect 17938 35086 17950 35138
rect 18002 35086 18014 35138
rect 16830 35074 16882 35086
rect 19854 35074 19906 35086
rect 1598 35026 1650 35038
rect 14030 35026 14082 35038
rect 20414 35026 20466 35038
rect 3154 34974 3166 35026
rect 3218 34974 3230 35026
rect 18050 34974 18062 35026
rect 18114 34974 18126 35026
rect 1598 34962 1650 34974
rect 14030 34962 14082 34974
rect 20414 34962 20466 34974
rect 1038 34914 1090 34926
rect 4286 34914 4338 34926
rect 6750 34914 6802 34926
rect 18958 34914 19010 34926
rect 2594 34862 2606 34914
rect 2658 34862 2670 34914
rect 5394 34862 5406 34914
rect 5458 34862 5470 34914
rect 5842 34862 5854 34914
rect 5906 34862 5918 34914
rect 7186 34862 7198 34914
rect 7250 34862 7262 34914
rect 8194 34862 8206 34914
rect 8258 34862 8270 34914
rect 12898 34862 12910 34914
rect 12962 34862 12974 34914
rect 13346 34862 13358 34914
rect 13410 34862 13422 34914
rect 14690 34862 14702 34914
rect 14754 34862 14766 34914
rect 15586 34862 15598 34914
rect 15650 34862 15662 34914
rect 24770 34862 24782 34914
rect 24834 34862 24846 34914
rect 26226 34862 26238 34914
rect 26290 34862 26302 34914
rect 1038 34850 1090 34862
rect 4286 34850 4338 34862
rect 6750 34850 6802 34862
rect 18958 34850 19010 34862
rect 5070 34802 5122 34814
rect 12574 34802 12626 34814
rect 19518 34802 19570 34814
rect 10546 34750 10558 34802
rect 10610 34750 10622 34802
rect 18386 34750 18398 34802
rect 18450 34750 18462 34802
rect 5070 34738 5122 34750
rect 12574 34738 12626 34750
rect 19518 34738 19570 34750
rect 25678 34802 25730 34814
rect 25678 34738 25730 34750
rect 12126 34690 12178 34702
rect 12126 34626 12178 34638
rect 27246 34690 27298 34702
rect 27246 34626 27298 34638
rect 672 34522 27888 34556
rect 672 34470 3806 34522
rect 3858 34470 3910 34522
rect 3962 34470 4014 34522
rect 4066 34470 23806 34522
rect 23858 34470 23910 34522
rect 23962 34470 24014 34522
rect 24066 34470 27888 34522
rect 672 34436 27888 34470
rect 6750 34354 6802 34366
rect 6750 34290 6802 34302
rect 25678 34242 25730 34254
rect 9090 34190 9102 34242
rect 9154 34190 9166 34242
rect 16706 34190 16718 34242
rect 16770 34190 16782 34242
rect 27122 34190 27134 34242
rect 27186 34190 27198 34242
rect 25678 34178 25730 34190
rect 2830 34130 2882 34142
rect 1474 34078 1486 34130
rect 1538 34078 1550 34130
rect 1922 34078 1934 34130
rect 1986 34078 1998 34130
rect 3154 34078 3166 34130
rect 3218 34078 3230 34130
rect 4162 34078 4174 34130
rect 4226 34078 4238 34130
rect 5170 34078 5182 34130
rect 5234 34078 5246 34130
rect 18498 34078 18510 34130
rect 18562 34078 18574 34130
rect 2830 34066 2882 34078
rect 1150 34018 1202 34030
rect 8642 33966 8654 34018
rect 8706 33966 8718 34018
rect 24658 33966 24670 34018
rect 24722 33966 24734 34018
rect 26226 33966 26238 34018
rect 26290 33966 26302 34018
rect 1150 33954 1202 33966
rect 7534 33906 7586 33918
rect 2146 33854 2158 33906
rect 2210 33854 2222 33906
rect 5618 33854 5630 33906
rect 5682 33854 5694 33906
rect 7534 33842 7586 33854
rect 672 33738 27888 33772
rect 672 33686 4466 33738
rect 4518 33686 4570 33738
rect 4622 33686 4674 33738
rect 4726 33686 24466 33738
rect 24518 33686 24570 33738
rect 24622 33686 24674 33738
rect 24726 33686 27888 33738
rect 672 33652 27888 33686
rect 3278 33570 3330 33582
rect 6066 33518 6078 33570
rect 6130 33518 6142 33570
rect 3278 33506 3330 33518
rect 3838 33458 3890 33470
rect 1586 33406 1598 33458
rect 1650 33406 1662 33458
rect 3838 33394 3890 33406
rect 8206 33458 8258 33470
rect 14590 33458 14642 33470
rect 9874 33406 9886 33458
rect 9938 33406 9950 33458
rect 12226 33406 12238 33458
rect 12290 33406 12302 33458
rect 8206 33394 8258 33406
rect 14590 33394 14642 33406
rect 15150 33458 15202 33470
rect 15150 33394 15202 33406
rect 16830 33458 16882 33470
rect 18274 33406 18286 33458
rect 18338 33406 18350 33458
rect 16830 33394 16882 33406
rect 7646 33346 7698 33358
rect 17390 33346 17442 33358
rect 9538 33294 9550 33346
rect 9602 33294 9614 33346
rect 11778 33294 11790 33346
rect 11842 33294 11854 33346
rect 24882 33294 24894 33346
rect 24946 33294 24958 33346
rect 26226 33294 26238 33346
rect 26290 33294 26302 33346
rect 7646 33282 7698 33294
rect 17390 33282 17442 33294
rect 1250 33182 1262 33234
rect 1314 33182 1326 33234
rect 5618 33182 5630 33234
rect 5682 33182 5694 33234
rect 17938 33182 17950 33234
rect 18002 33182 18014 33234
rect 2830 33122 2882 33134
rect 2830 33058 2882 33070
rect 7198 33122 7250 33134
rect 7198 33058 7250 33070
rect 11118 33122 11170 33134
rect 11118 33058 11170 33070
rect 13470 33122 13522 33134
rect 13470 33058 13522 33070
rect 19518 33122 19570 33134
rect 19518 33058 19570 33070
rect 25678 33122 25730 33134
rect 25678 33058 25730 33070
rect 27246 33122 27298 33134
rect 27246 33058 27298 33070
rect 672 32954 27888 32988
rect 672 32902 3806 32954
rect 3858 32902 3910 32954
rect 3962 32902 4014 32954
rect 4066 32902 23806 32954
rect 23858 32902 23910 32954
rect 23962 32902 24014 32954
rect 24066 32902 27888 32954
rect 672 32868 27888 32902
rect 18286 32786 18338 32798
rect 18286 32722 18338 32734
rect 14366 32674 14418 32686
rect 1698 32622 1710 32674
rect 1762 32622 1774 32674
rect 13346 32622 13358 32674
rect 13410 32622 13422 32674
rect 17378 32622 17390 32674
rect 17442 32622 17454 32674
rect 14366 32610 14418 32622
rect 7758 32562 7810 32574
rect 6738 32510 6750 32562
rect 6802 32510 6814 32562
rect 7074 32510 7086 32562
rect 7138 32510 7150 32562
rect 8418 32510 8430 32562
rect 8482 32510 8494 32562
rect 9214 32557 9266 32569
rect 18622 32562 18674 32574
rect 7758 32498 7810 32510
rect 10546 32510 10558 32562
rect 10610 32510 10622 32562
rect 13010 32510 13022 32562
rect 13074 32510 13086 32562
rect 15138 32510 15150 32562
rect 15202 32510 15214 32562
rect 19394 32510 19406 32562
rect 19458 32510 19470 32562
rect 9214 32493 9266 32505
rect 18622 32498 18674 32510
rect 4286 32450 4338 32462
rect 2146 32398 2158 32450
rect 2210 32398 2222 32450
rect 4286 32386 4338 32398
rect 6302 32450 6354 32462
rect 7298 32398 7310 32450
rect 7362 32398 7374 32450
rect 15586 32398 15598 32450
rect 15650 32398 15662 32450
rect 19170 32398 19182 32450
rect 19234 32398 19246 32450
rect 26226 32398 26238 32450
rect 26290 32398 26302 32450
rect 27010 32398 27022 32450
rect 27074 32398 27086 32450
rect 6302 32386 6354 32398
rect 3278 32338 3330 32350
rect 3278 32274 3330 32286
rect 3726 32338 3778 32350
rect 12126 32338 12178 32350
rect 10994 32286 11006 32338
rect 11058 32286 11070 32338
rect 3726 32274 3778 32286
rect 12126 32274 12178 32286
rect 13806 32338 13858 32350
rect 13806 32274 13858 32286
rect 16830 32338 16882 32350
rect 16830 32274 16882 32286
rect 17838 32338 17890 32350
rect 17838 32274 17890 32286
rect 672 32170 27888 32204
rect 672 32118 4466 32170
rect 4518 32118 4570 32170
rect 4622 32118 4674 32170
rect 4726 32118 24466 32170
rect 24518 32118 24570 32170
rect 24622 32118 24674 32170
rect 24726 32118 27888 32170
rect 672 32084 27888 32118
rect 13010 31950 13022 32002
rect 13074 31950 13086 32002
rect 17714 31950 17726 32002
rect 17778 31950 17790 32002
rect 3278 31890 3330 31902
rect 2818 31838 2830 31890
rect 2882 31838 2894 31890
rect 3278 31826 3330 31838
rect 9438 31890 9490 31902
rect 9438 31826 9490 31838
rect 13470 31890 13522 31902
rect 13470 31826 13522 31838
rect 18174 31890 18226 31902
rect 18174 31826 18226 31838
rect 8878 31778 8930 31790
rect 16718 31778 16770 31790
rect 2258 31726 2270 31778
rect 2322 31726 2334 31778
rect 2706 31726 2718 31778
rect 2770 31726 2782 31778
rect 4050 31726 4062 31778
rect 4114 31726 4126 31778
rect 4834 31726 4846 31778
rect 4898 31726 4910 31778
rect 7298 31726 7310 31778
rect 7362 31726 7374 31778
rect 12338 31726 12350 31778
rect 12402 31726 12414 31778
rect 12898 31726 12910 31778
rect 12962 31726 12974 31778
rect 14018 31726 14030 31778
rect 14082 31726 14094 31778
rect 15026 31726 15038 31778
rect 15090 31726 15102 31778
rect 17042 31726 17054 31778
rect 17106 31726 17118 31778
rect 17490 31726 17502 31778
rect 17554 31726 17566 31778
rect 18946 31726 18958 31778
rect 19010 31726 19022 31778
rect 19842 31726 19854 31778
rect 19906 31726 19918 31778
rect 24770 31726 24782 31778
rect 24834 31726 24846 31778
rect 26338 31726 26350 31778
rect 26402 31726 26414 31778
rect 8878 31714 8930 31726
rect 16718 31714 16770 31726
rect 1822 31666 1874 31678
rect 1822 31602 1874 31614
rect 12014 31666 12066 31678
rect 12014 31602 12066 31614
rect 25678 31666 25730 31678
rect 25678 31602 25730 31614
rect 7646 31554 7698 31566
rect 7646 31490 7698 31502
rect 27246 31554 27298 31566
rect 27246 31490 27298 31502
rect 672 31386 27888 31420
rect 672 31334 3806 31386
rect 3858 31334 3910 31386
rect 3962 31334 4014 31386
rect 4066 31334 23806 31386
rect 23858 31334 23910 31386
rect 23962 31334 24014 31386
rect 24066 31334 27888 31386
rect 672 31300 27888 31334
rect 15822 31218 15874 31230
rect 15822 31154 15874 31166
rect 4398 31106 4450 31118
rect 11902 31106 11954 31118
rect 6626 31054 6638 31106
rect 6690 31054 6702 31106
rect 7186 31054 7198 31106
rect 7250 31054 7262 31106
rect 10770 31054 10782 31106
rect 10834 31054 10846 31106
rect 4398 31042 4450 31054
rect 11902 31042 11954 31054
rect 11342 30994 11394 31006
rect 18398 30994 18450 31006
rect 1250 30942 1262 30994
rect 1314 30942 1326 30994
rect 2370 30942 2382 30994
rect 2434 30942 2446 30994
rect 3490 30942 3502 30994
rect 3554 30942 3566 30994
rect 3938 30942 3950 30994
rect 4002 30942 4014 30994
rect 8082 30942 8094 30994
rect 8146 30942 8158 30994
rect 10434 30942 10446 30994
rect 10498 30942 10510 30994
rect 14242 30942 14254 30994
rect 14306 30942 14318 30994
rect 17154 30942 17166 30994
rect 17218 30942 17230 30994
rect 17490 30942 17502 30994
rect 17554 30942 17566 30994
rect 18722 30942 18734 30994
rect 18786 30942 18798 30994
rect 19842 30942 19854 30994
rect 19906 30942 19918 30994
rect 24882 30942 24894 30994
rect 24946 30942 24958 30994
rect 26450 30942 26462 30994
rect 26514 30942 26526 30994
rect 11342 30930 11394 30942
rect 18398 30930 18450 30942
rect 2942 30882 2994 30894
rect 16718 30882 16770 30894
rect 8642 30830 8654 30882
rect 8706 30830 8718 30882
rect 14578 30830 14590 30882
rect 14642 30830 14654 30882
rect 17714 30830 17726 30882
rect 17778 30830 17790 30882
rect 25442 30830 25454 30882
rect 25506 30830 25518 30882
rect 27010 30830 27022 30882
rect 27074 30830 27086 30882
rect 2942 30818 2994 30830
rect 16718 30818 16770 30830
rect 6190 30770 6242 30782
rect 3378 30718 3390 30770
rect 3442 30718 3454 30770
rect 6190 30706 6242 30718
rect 7646 30770 7698 30782
rect 7646 30706 7698 30718
rect 9774 30770 9826 30782
rect 9774 30706 9826 30718
rect 672 30602 27888 30636
rect 672 30550 4466 30602
rect 4518 30550 4570 30602
rect 4622 30550 4674 30602
rect 4726 30550 24466 30602
rect 24518 30550 24570 30602
rect 24622 30550 24674 30602
rect 24726 30550 27888 30602
rect 672 30516 27888 30550
rect 3166 30434 3218 30446
rect 3166 30370 3218 30382
rect 3502 30434 3554 30446
rect 6066 30382 6078 30434
rect 6130 30382 6142 30434
rect 10434 30382 10446 30434
rect 10498 30382 10510 30434
rect 3502 30370 3554 30382
rect 4062 30322 4114 30334
rect 17378 30270 17390 30322
rect 17442 30270 17454 30322
rect 4062 30258 4114 30270
rect 6750 30210 6802 30222
rect 9438 30210 9490 30222
rect 14142 30210 14194 30222
rect 18510 30210 18562 30222
rect 2258 30158 2270 30210
rect 2322 30158 2334 30210
rect 5394 30158 5406 30210
rect 5458 30158 5470 30210
rect 5842 30158 5854 30210
rect 5906 30158 5918 30210
rect 7074 30158 7086 30210
rect 7138 30158 7150 30210
rect 8194 30158 8206 30210
rect 8258 30158 8270 30210
rect 9762 30158 9774 30210
rect 9826 30158 9838 30210
rect 10210 30158 10222 30210
rect 10274 30158 10286 30210
rect 10994 30158 11006 30210
rect 11058 30158 11070 30210
rect 11442 30158 11454 30210
rect 11506 30158 11518 30210
rect 12450 30158 12462 30210
rect 12514 30158 12526 30210
rect 15698 30158 15710 30210
rect 15762 30158 15774 30210
rect 16818 30158 16830 30210
rect 16882 30158 16894 30210
rect 26450 30158 26462 30210
rect 26514 30158 26526 30210
rect 6750 30146 6802 30158
rect 9438 30146 9490 30158
rect 14142 30146 14194 30158
rect 18510 30146 18562 30158
rect 1262 30098 1314 30110
rect 5070 30098 5122 30110
rect 2706 30046 2718 30098
rect 2770 30046 2782 30098
rect 1262 30034 1314 30046
rect 5070 30034 5122 30046
rect 14702 30098 14754 30110
rect 16034 30046 16046 30098
rect 16098 30046 16110 30098
rect 27122 30046 27134 30098
rect 27186 30046 27198 30098
rect 14702 30034 14754 30046
rect 672 29818 27888 29852
rect 672 29766 3806 29818
rect 3858 29766 3910 29818
rect 3962 29766 4014 29818
rect 4066 29766 23806 29818
rect 23858 29766 23910 29818
rect 23962 29766 24014 29818
rect 24066 29766 27888 29818
rect 672 29732 27888 29766
rect 2830 29650 2882 29662
rect 2830 29586 2882 29598
rect 6750 29650 6802 29662
rect 6750 29586 6802 29598
rect 17502 29650 17554 29662
rect 17502 29586 17554 29598
rect 27246 29538 27298 29550
rect 3714 29486 3726 29538
rect 3778 29486 3790 29538
rect 5170 29486 5182 29538
rect 5234 29486 5246 29538
rect 12114 29486 12126 29538
rect 12178 29486 12190 29538
rect 27246 29474 27298 29486
rect 1138 29374 1150 29426
rect 1202 29374 1214 29426
rect 3378 29374 3390 29426
rect 3442 29374 3454 29426
rect 8530 29374 8542 29426
rect 8594 29374 8606 29426
rect 11778 29374 11790 29426
rect 11842 29374 11854 29426
rect 13570 29374 13582 29426
rect 13634 29374 13646 29426
rect 15810 29374 15822 29426
rect 15874 29374 15886 29426
rect 18050 29374 18062 29426
rect 18114 29374 18126 29426
rect 1698 29262 1710 29314
rect 1762 29262 1774 29314
rect 8866 29262 8878 29314
rect 8930 29262 8942 29314
rect 16258 29262 16270 29314
rect 16322 29262 16334 29314
rect 18498 29262 18510 29314
rect 18562 29262 18574 29314
rect 26226 29262 26238 29314
rect 26290 29262 26302 29314
rect 10110 29202 10162 29214
rect 15262 29202 15314 29214
rect 5618 29150 5630 29202
rect 5682 29150 5694 29202
rect 14130 29150 14142 29202
rect 14194 29150 14206 29202
rect 10110 29138 10162 29150
rect 15262 29138 15314 29150
rect 19742 29202 19794 29214
rect 19742 29138 19794 29150
rect 672 29034 27888 29068
rect 672 28982 4466 29034
rect 4518 28982 4570 29034
rect 4622 28982 4674 29034
rect 4726 28982 24466 29034
rect 24518 28982 24570 29034
rect 24622 28982 24674 29034
rect 24726 28982 27888 29034
rect 672 28948 27888 28982
rect 2830 28866 2882 28878
rect 2830 28802 2882 28814
rect 5070 28866 5122 28878
rect 11330 28814 11342 28866
rect 11394 28814 11406 28866
rect 13906 28814 13918 28866
rect 13970 28814 13982 28866
rect 5070 28802 5122 28814
rect 12910 28754 12962 28766
rect 1586 28702 1598 28754
rect 1650 28702 1662 28754
rect 3826 28702 3838 28754
rect 3890 28702 3902 28754
rect 6962 28702 6974 28754
rect 7026 28702 7038 28754
rect 12910 28690 12962 28702
rect 18398 28754 18450 28766
rect 19854 28754 19906 28766
rect 19394 28702 19406 28754
rect 19458 28702 19470 28754
rect 26226 28702 26238 28754
rect 26290 28702 26302 28754
rect 18398 28690 18450 28702
rect 19854 28690 19906 28702
rect 5518 28642 5570 28654
rect 12462 28642 12514 28654
rect 14366 28642 14418 28654
rect 1138 28590 1150 28642
rect 1202 28590 1214 28642
rect 5954 28590 5966 28642
rect 6018 28590 6030 28642
rect 13234 28590 13246 28642
rect 13298 28590 13310 28642
rect 13682 28590 13694 28642
rect 13746 28590 13758 28642
rect 14914 28590 14926 28642
rect 14978 28590 14990 28642
rect 16034 28590 16046 28642
rect 16098 28590 16110 28642
rect 18834 28590 18846 28642
rect 18898 28590 18910 28642
rect 19170 28590 19182 28642
rect 19234 28590 19246 28642
rect 20402 28590 20414 28642
rect 20466 28590 20478 28642
rect 21410 28590 21422 28642
rect 21474 28590 21486 28642
rect 5518 28578 5570 28590
rect 12462 28578 12514 28590
rect 14366 28578 14418 28590
rect 27246 28530 27298 28542
rect 3490 28478 3502 28530
rect 3554 28478 3566 28530
rect 6626 28478 6638 28530
rect 6690 28478 6702 28530
rect 10882 28478 10894 28530
rect 10946 28478 10958 28530
rect 27246 28466 27298 28478
rect 8206 28418 8258 28430
rect 8206 28354 8258 28366
rect 672 28250 27888 28284
rect 672 28198 3806 28250
rect 3858 28198 3910 28250
rect 3962 28198 4014 28250
rect 4066 28198 23806 28250
rect 23858 28198 23910 28250
rect 23962 28198 24014 28250
rect 24066 28198 27888 28250
rect 672 28164 27888 28198
rect 19070 28082 19122 28094
rect 19070 28018 19122 28030
rect 27246 28082 27298 28094
rect 27246 28018 27298 28030
rect 1598 27970 1650 27982
rect 8990 27970 9042 27982
rect 2706 27918 2718 27970
rect 2770 27918 2782 27970
rect 1598 27906 1650 27918
rect 8990 27906 9042 27918
rect 13582 27970 13634 27982
rect 20078 27970 20130 27982
rect 17490 27918 17502 27970
rect 17554 27918 17566 27970
rect 13582 27906 13634 27918
rect 20078 27906 20130 27918
rect 25678 27970 25730 27982
rect 25678 27906 25730 27918
rect 1038 27858 1090 27870
rect 1038 27794 1090 27806
rect 4286 27858 4338 27870
rect 10446 27858 10498 27870
rect 15262 27858 15314 27870
rect 19518 27858 19570 27870
rect 5282 27806 5294 27858
rect 5346 27806 5358 27858
rect 5730 27806 5742 27858
rect 5794 27806 5806 27858
rect 6514 27806 6526 27858
rect 6578 27806 6590 27858
rect 7074 27806 7086 27858
rect 7138 27806 7150 27858
rect 8082 27806 8094 27858
rect 8146 27806 8158 27858
rect 9314 27806 9326 27858
rect 9378 27806 9390 27858
rect 9762 27806 9774 27858
rect 9826 27806 9838 27858
rect 10994 27806 11006 27858
rect 11058 27806 11070 27858
rect 12114 27806 12126 27858
rect 12178 27806 12190 27858
rect 14018 27806 14030 27858
rect 14082 27806 14094 27858
rect 14354 27806 14366 27858
rect 14418 27806 14430 27858
rect 15810 27806 15822 27858
rect 15874 27806 15886 27858
rect 16594 27806 16606 27858
rect 16658 27806 16670 27858
rect 24658 27806 24670 27858
rect 24722 27806 24734 27858
rect 26338 27806 26350 27858
rect 26402 27806 26414 27858
rect 4286 27794 4338 27806
rect 10446 27794 10498 27806
rect 15262 27794 15314 27806
rect 19518 27794 19570 27806
rect 4958 27746 5010 27758
rect 3154 27694 3166 27746
rect 3218 27694 3230 27746
rect 5954 27694 5966 27746
rect 6018 27694 6030 27746
rect 17938 27694 17950 27746
rect 18002 27694 18014 27746
rect 4958 27682 5010 27694
rect 9986 27582 9998 27634
rect 10050 27582 10062 27634
rect 14578 27582 14590 27634
rect 14642 27582 14654 27634
rect 672 27466 27888 27500
rect 672 27414 4466 27466
rect 4518 27414 4570 27466
rect 4622 27414 4674 27466
rect 4726 27414 24466 27466
rect 24518 27414 24570 27466
rect 24622 27414 24674 27466
rect 24726 27414 27888 27466
rect 672 27380 27888 27414
rect 6526 27298 6578 27310
rect 5394 27246 5406 27298
rect 5458 27246 5470 27298
rect 6526 27234 6578 27246
rect 10222 27298 10274 27310
rect 10222 27234 10274 27246
rect 12910 27298 12962 27310
rect 15150 27298 15202 27310
rect 14018 27246 14030 27298
rect 14082 27246 14094 27298
rect 12910 27234 12962 27246
rect 15150 27234 15202 27246
rect 15598 27298 15650 27310
rect 15598 27234 15650 27246
rect 16158 27186 16210 27198
rect 1586 27134 1598 27186
rect 1650 27134 1662 27186
rect 11666 27134 11678 27186
rect 11730 27134 11742 27186
rect 18274 27134 18286 27186
rect 18338 27134 18350 27186
rect 24658 27134 24670 27186
rect 24722 27134 24734 27186
rect 26226 27134 26238 27186
rect 26290 27134 26302 27186
rect 16158 27122 16210 27134
rect 1138 27022 1150 27074
rect 1202 27022 1214 27074
rect 3378 27022 3390 27074
rect 3442 27022 3454 27074
rect 4834 27022 4846 27074
rect 4898 27022 4910 27074
rect 13458 27022 13470 27074
rect 13522 27022 13534 27074
rect 17826 27022 17838 27074
rect 17890 27022 17902 27074
rect 10782 26962 10834 26974
rect 27246 26962 27298 26974
rect 3714 26910 3726 26962
rect 3778 26910 3790 26962
rect 11330 26910 11342 26962
rect 11394 26910 11406 26962
rect 10782 26898 10834 26910
rect 27246 26898 27298 26910
rect 2830 26850 2882 26862
rect 2830 26786 2882 26798
rect 19406 26850 19458 26862
rect 19406 26786 19458 26798
rect 25678 26850 25730 26862
rect 25678 26786 25730 26798
rect 672 26682 27888 26716
rect 672 26630 3806 26682
rect 3858 26630 3910 26682
rect 3962 26630 4014 26682
rect 4066 26630 23806 26682
rect 23858 26630 23910 26682
rect 23962 26630 24014 26682
rect 24066 26630 27888 26682
rect 672 26596 27888 26630
rect 27246 26514 27298 26526
rect 27246 26450 27298 26462
rect 4286 26402 4338 26414
rect 1698 26350 1710 26402
rect 1762 26350 1774 26402
rect 4286 26338 4338 26350
rect 13358 26402 13410 26414
rect 14466 26350 14478 26402
rect 14530 26350 14542 26402
rect 13358 26338 13410 26350
rect 19182 26290 19234 26302
rect 7634 26238 7646 26290
rect 7698 26238 7710 26290
rect 16370 26238 16382 26290
rect 16434 26238 16446 26290
rect 19182 26226 19234 26238
rect 19742 26178 19794 26190
rect 7970 26126 7982 26178
rect 8034 26126 8046 26178
rect 16930 26126 16942 26178
rect 16994 26126 17006 26178
rect 26226 26126 26238 26178
rect 26290 26126 26302 26178
rect 19742 26114 19794 26126
rect 3278 26066 3330 26078
rect 2146 26014 2158 26066
rect 2210 26014 2222 26066
rect 3278 26002 3330 26014
rect 3726 26066 3778 26078
rect 3726 26002 3778 26014
rect 9214 26066 9266 26078
rect 9214 26002 9266 26014
rect 12798 26066 12850 26078
rect 12798 26002 12850 26014
rect 14030 26066 14082 26078
rect 14030 26002 14082 26014
rect 18062 26066 18114 26078
rect 18062 26002 18114 26014
rect 672 25898 27888 25932
rect 672 25846 4466 25898
rect 4518 25846 4570 25898
rect 4622 25846 4674 25898
rect 4726 25846 24466 25898
rect 24518 25846 24570 25898
rect 24622 25846 24674 25898
rect 24726 25846 27888 25898
rect 672 25812 27888 25846
rect 1038 25730 1090 25742
rect 3042 25678 3054 25730
rect 3106 25678 3118 25730
rect 13122 25678 13134 25730
rect 13186 25678 13198 25730
rect 1038 25666 1090 25678
rect 2046 25618 2098 25630
rect 2046 25554 2098 25566
rect 3502 25618 3554 25630
rect 9438 25618 9490 25630
rect 15262 25618 15314 25630
rect 6626 25566 6638 25618
rect 6690 25566 6702 25618
rect 10882 25566 10894 25618
rect 10946 25566 10958 25618
rect 18498 25566 18510 25618
rect 18562 25566 18574 25618
rect 24658 25566 24670 25618
rect 24722 25566 24734 25618
rect 3502 25554 3554 25566
rect 9438 25554 9490 25566
rect 15262 25554 15314 25566
rect 8878 25506 8930 25518
rect 14702 25506 14754 25518
rect 19182 25506 19234 25518
rect 2482 25454 2494 25506
rect 2546 25454 2558 25506
rect 2930 25454 2942 25506
rect 2994 25454 3006 25506
rect 4050 25454 4062 25506
rect 4114 25454 4126 25506
rect 5058 25454 5070 25506
rect 5122 25454 5134 25506
rect 6290 25454 6302 25506
rect 6354 25454 6366 25506
rect 12562 25454 12574 25506
rect 12626 25454 12638 25506
rect 17938 25454 17950 25506
rect 18002 25454 18014 25506
rect 18274 25454 18286 25506
rect 18338 25454 18350 25506
rect 19730 25454 19742 25506
rect 19794 25454 19806 25506
rect 20626 25454 20638 25506
rect 20690 25454 20702 25506
rect 26226 25454 26238 25506
rect 26290 25454 26302 25506
rect 8878 25442 8930 25454
rect 14702 25442 14754 25454
rect 19182 25442 19234 25454
rect 1598 25394 1650 25406
rect 17502 25394 17554 25406
rect 10434 25342 10446 25394
rect 10498 25342 10510 25394
rect 1598 25330 1650 25342
rect 17502 25330 17554 25342
rect 27246 25394 27298 25406
rect 27246 25330 27298 25342
rect 7870 25282 7922 25294
rect 7870 25218 7922 25230
rect 12014 25282 12066 25294
rect 12014 25218 12066 25230
rect 14254 25282 14306 25294
rect 14254 25218 14306 25230
rect 25678 25282 25730 25294
rect 25678 25218 25730 25230
rect 672 25114 27888 25148
rect 672 25062 3806 25114
rect 3858 25062 3910 25114
rect 3962 25062 4014 25114
rect 4066 25062 23806 25114
rect 23858 25062 23910 25114
rect 23962 25062 24014 25114
rect 24066 25062 27888 25114
rect 672 25028 27888 25062
rect 6190 24834 6242 24846
rect 19518 24834 19570 24846
rect 18162 24782 18174 24834
rect 18226 24782 18238 24834
rect 27122 24782 27134 24834
rect 27186 24782 27198 24834
rect 6190 24770 6242 24782
rect 19518 24770 19570 24782
rect 2718 24722 2770 24734
rect 9214 24722 9266 24734
rect 14366 24722 14418 24734
rect 16606 24722 16658 24734
rect 1362 24670 1374 24722
rect 1426 24670 1438 24722
rect 2370 24670 2382 24722
rect 2434 24670 2446 24722
rect 3490 24670 3502 24722
rect 3554 24670 3566 24722
rect 4050 24670 4062 24722
rect 4114 24670 4126 24722
rect 7858 24670 7870 24722
rect 7922 24670 7934 24722
rect 8306 24670 8318 24722
rect 8370 24670 8382 24722
rect 9538 24670 9550 24722
rect 9602 24670 9614 24722
rect 10658 24670 10670 24722
rect 10722 24670 10734 24722
rect 13346 24670 13358 24722
rect 13410 24670 13422 24722
rect 13682 24670 13694 24722
rect 13746 24670 13758 24722
rect 14914 24670 14926 24722
rect 14978 24670 14990 24722
rect 15922 24670 15934 24722
rect 15986 24670 15998 24722
rect 2718 24658 2770 24670
rect 9214 24658 9266 24670
rect 14366 24658 14418 24670
rect 16606 24658 16658 24670
rect 18958 24722 19010 24734
rect 18958 24658 19010 24670
rect 4398 24610 4450 24622
rect 4398 24546 4450 24558
rect 7534 24610 7586 24622
rect 12238 24610 12290 24622
rect 8530 24558 8542 24610
rect 8594 24558 8606 24610
rect 7534 24546 7586 24558
rect 12238 24546 12290 24558
rect 12910 24610 12962 24622
rect 13906 24558 13918 24610
rect 13970 24558 13982 24610
rect 17714 24558 17726 24610
rect 17778 24558 17790 24610
rect 24658 24558 24670 24610
rect 24722 24558 24734 24610
rect 25442 24558 25454 24610
rect 25506 24558 25518 24610
rect 26226 24558 26238 24610
rect 26290 24558 26302 24610
rect 12910 24546 12962 24558
rect 5630 24498 5682 24510
rect 3378 24446 3390 24498
rect 3442 24446 3454 24498
rect 5630 24434 5682 24446
rect 12014 24498 12066 24510
rect 12014 24434 12066 24446
rect 12126 24498 12178 24510
rect 12126 24434 12178 24446
rect 672 24330 27888 24364
rect 672 24278 4466 24330
rect 4518 24278 4570 24330
rect 4622 24278 4674 24330
rect 4726 24278 24466 24330
rect 24518 24278 24570 24330
rect 24622 24278 24674 24330
rect 24726 24278 27888 24330
rect 672 24244 27888 24278
rect 1038 24162 1090 24174
rect 1038 24098 1090 24110
rect 2494 24162 2546 24174
rect 5618 24110 5630 24162
rect 5682 24110 5694 24162
rect 11218 24110 11230 24162
rect 11282 24110 11294 24162
rect 13794 24110 13806 24162
rect 13858 24110 13870 24162
rect 17938 24110 17950 24162
rect 18002 24110 18014 24162
rect 2494 24098 2546 24110
rect 6078 24050 6130 24062
rect 3602 23998 3614 24050
rect 3666 23998 3678 24050
rect 6078 23986 6130 23998
rect 9326 24050 9378 24062
rect 9326 23986 9378 23998
rect 19966 24050 20018 24062
rect 19966 23986 20018 23998
rect 9886 23938 9938 23950
rect 14254 23938 14306 23950
rect 4050 23886 4062 23938
rect 4114 23886 4126 23938
rect 5058 23886 5070 23938
rect 5122 23886 5134 23938
rect 5394 23886 5406 23938
rect 5458 23886 5470 23938
rect 6850 23886 6862 23938
rect 6914 23886 6926 23938
rect 7634 23886 7646 23938
rect 7698 23886 7710 23938
rect 13122 23886 13134 23938
rect 13186 23886 13198 23938
rect 13682 23886 13694 23938
rect 13746 23886 13758 23938
rect 15026 23886 15038 23938
rect 15090 23886 15102 23938
rect 15922 23886 15934 23938
rect 15986 23886 15998 23938
rect 18386 23886 18398 23938
rect 18450 23886 18462 23938
rect 19506 23886 19518 23938
rect 19570 23886 19582 23938
rect 24882 23886 24894 23938
rect 24946 23886 24958 23938
rect 26226 23886 26238 23938
rect 26290 23886 26302 23938
rect 9886 23874 9938 23886
rect 14254 23874 14306 23886
rect 1598 23826 1650 23838
rect 1598 23762 1650 23774
rect 4622 23826 4674 23838
rect 12350 23826 12402 23838
rect 10770 23774 10782 23826
rect 10834 23774 10846 23826
rect 4622 23762 4674 23774
rect 12350 23762 12402 23774
rect 12798 23826 12850 23838
rect 12798 23762 12850 23774
rect 27246 23826 27298 23838
rect 27246 23762 27298 23774
rect 16830 23714 16882 23726
rect 16830 23650 16882 23662
rect 25678 23714 25730 23726
rect 25678 23650 25730 23662
rect 672 23546 27888 23580
rect 672 23494 3806 23546
rect 3858 23494 3910 23546
rect 3962 23494 4014 23546
rect 4066 23494 23806 23546
rect 23858 23494 23910 23546
rect 23962 23494 24014 23546
rect 24066 23494 27888 23546
rect 672 23460 27888 23494
rect 3838 23378 3890 23390
rect 11666 23326 11678 23378
rect 11730 23326 11742 23378
rect 3838 23314 3890 23326
rect 16942 23266 16994 23278
rect 1586 23214 1598 23266
rect 1650 23214 1662 23266
rect 2258 23214 2270 23266
rect 2322 23214 2334 23266
rect 18946 23214 18958 23266
rect 19010 23214 19022 23266
rect 27122 23214 27134 23266
rect 27186 23214 27198 23266
rect 16942 23202 16994 23214
rect 6190 23154 6242 23166
rect 1250 23102 1262 23154
rect 1314 23102 1326 23154
rect 5730 23102 5742 23154
rect 5794 23102 5806 23154
rect 6738 23102 6750 23154
rect 6802 23102 6814 23154
rect 8978 23102 8990 23154
rect 9042 23102 9054 23154
rect 11442 23102 11454 23154
rect 11506 23102 11518 23154
rect 13122 23102 13134 23154
rect 13186 23102 13198 23154
rect 13682 23102 13694 23154
rect 13746 23102 13758 23154
rect 14354 23102 14366 23154
rect 14418 23102 14430 23154
rect 14802 23102 14814 23154
rect 14866 23102 14878 23154
rect 15922 23102 15934 23154
rect 15986 23102 15998 23154
rect 26338 23102 26350 23154
rect 26402 23102 26414 23154
rect 6190 23090 6242 23102
rect 10558 23042 10610 23054
rect 12238 23042 12290 23054
rect 2594 22990 2606 23042
rect 2658 22990 2670 23042
rect 9426 22990 9438 23042
rect 9490 22990 9502 23042
rect 12002 22990 12014 23042
rect 12066 22990 12078 23042
rect 10558 22978 10610 22990
rect 12238 22978 12290 22990
rect 12798 23042 12850 23054
rect 13794 22990 13806 23042
rect 13858 22990 13870 23042
rect 12798 22978 12850 22990
rect 8318 22930 8370 22942
rect 16382 22930 16434 22942
rect 7186 22878 7198 22930
rect 7250 22878 7262 22930
rect 11778 22878 11790 22930
rect 11842 22878 11854 22930
rect 8318 22866 8370 22878
rect 16382 22866 16434 22878
rect 17390 22930 17442 22942
rect 18498 22878 18510 22930
rect 18562 22878 18574 22930
rect 17390 22866 17442 22878
rect 672 22762 27888 22796
rect 672 22710 4466 22762
rect 4518 22710 4570 22762
rect 4622 22710 4674 22762
rect 4726 22710 24466 22762
rect 24518 22710 24570 22762
rect 24622 22710 24674 22762
rect 24726 22710 27888 22762
rect 672 22676 27888 22710
rect 1710 22594 1762 22606
rect 2706 22542 2718 22594
rect 2770 22542 2782 22594
rect 5954 22542 5966 22594
rect 6018 22542 6030 22594
rect 9874 22542 9886 22594
rect 9938 22542 9950 22594
rect 15138 22542 15150 22594
rect 15202 22542 15214 22594
rect 1710 22530 1762 22542
rect 1150 22482 1202 22494
rect 1150 22418 1202 22430
rect 10334 22482 10386 22494
rect 10334 22418 10386 22430
rect 14702 22482 14754 22494
rect 18610 22430 18622 22482
rect 18674 22430 18686 22482
rect 26226 22430 26238 22482
rect 26290 22430 26302 22482
rect 14702 22418 14754 22430
rect 16830 22370 16882 22382
rect 2146 22318 2158 22370
rect 2210 22318 2222 22370
rect 5282 22318 5294 22370
rect 5346 22318 5358 22370
rect 5730 22318 5742 22370
rect 5794 22318 5806 22370
rect 6514 22318 6526 22370
rect 6578 22318 6590 22370
rect 6962 22318 6974 22370
rect 7026 22318 7038 22370
rect 8082 22318 8094 22370
rect 8146 22318 8158 22370
rect 9202 22318 9214 22370
rect 9266 22318 9278 22370
rect 9762 22318 9774 22370
rect 9826 22318 9838 22370
rect 10882 22318 10894 22370
rect 10946 22318 10958 22370
rect 11890 22318 11902 22370
rect 11954 22318 11966 22370
rect 13010 22318 13022 22370
rect 13074 22318 13086 22370
rect 13906 22318 13918 22370
rect 13970 22318 13982 22370
rect 15362 22318 15374 22370
rect 15426 22318 15438 22370
rect 15810 22318 15822 22370
rect 15874 22318 15886 22370
rect 19058 22318 19070 22370
rect 19122 22318 19134 22370
rect 24882 22318 24894 22370
rect 24946 22318 24958 22370
rect 16830 22306 16882 22318
rect 4958 22258 5010 22270
rect 4958 22194 5010 22206
rect 8878 22258 8930 22270
rect 8878 22194 8930 22206
rect 16158 22258 16210 22270
rect 16158 22194 16210 22206
rect 27246 22258 27298 22270
rect 27246 22194 27298 22206
rect 3838 22146 3890 22158
rect 3838 22082 3890 22094
rect 16718 22146 16770 22158
rect 16718 22082 16770 22094
rect 17390 22146 17442 22158
rect 17390 22082 17442 22094
rect 25678 22146 25730 22158
rect 25678 22082 25730 22094
rect 672 21978 27888 22012
rect 672 21926 3806 21978
rect 3858 21926 3910 21978
rect 3962 21926 4014 21978
rect 4066 21926 23806 21978
rect 23858 21926 23910 21978
rect 23962 21926 24014 21978
rect 24066 21926 27888 21978
rect 672 21892 27888 21926
rect 4286 21810 4338 21822
rect 4286 21746 4338 21758
rect 11678 21810 11730 21822
rect 11678 21746 11730 21758
rect 12798 21810 12850 21822
rect 12798 21746 12850 21758
rect 13134 21810 13186 21822
rect 13134 21746 13186 21758
rect 6302 21698 6354 21710
rect 5506 21646 5518 21698
rect 5570 21646 5582 21698
rect 6302 21634 6354 21646
rect 16718 21698 16770 21710
rect 18722 21646 18734 21698
rect 18786 21646 18798 21698
rect 27122 21646 27134 21698
rect 27186 21646 27198 21698
rect 16718 21634 16770 21646
rect 1038 21586 1090 21598
rect 2594 21534 2606 21586
rect 2658 21534 2670 21586
rect 6738 21534 6750 21586
rect 6802 21534 6814 21586
rect 7074 21534 7086 21586
rect 7138 21534 7150 21586
rect 7858 21534 7870 21586
rect 7922 21534 7934 21586
rect 8306 21534 8318 21586
rect 8370 21534 8382 21586
rect 9426 21534 9438 21586
rect 9490 21534 9502 21586
rect 10098 21534 10110 21586
rect 10162 21534 10174 21586
rect 13570 21534 13582 21586
rect 13634 21534 13646 21586
rect 14466 21534 14478 21586
rect 14530 21534 14542 21586
rect 15810 21534 15822 21586
rect 15874 21534 15886 21586
rect 16370 21534 16382 21586
rect 16434 21534 16446 21586
rect 1038 21522 1090 21534
rect 1598 21474 1650 21486
rect 12238 21474 12290 21486
rect 3154 21422 3166 21474
rect 3218 21422 3230 21474
rect 10434 21422 10446 21474
rect 10498 21422 10510 21474
rect 1598 21410 1650 21422
rect 12238 21410 12290 21422
rect 15262 21474 15314 21486
rect 15262 21410 15314 21422
rect 17166 21474 17218 21486
rect 19294 21474 19346 21486
rect 18274 21422 18286 21474
rect 18338 21422 18350 21474
rect 17166 21410 17218 21422
rect 19294 21410 19346 21422
rect 25342 21474 25394 21486
rect 26226 21422 26238 21474
rect 26290 21422 26302 21474
rect 25342 21410 25394 21422
rect 5966 21362 6018 21374
rect 12126 21362 12178 21374
rect 7298 21310 7310 21362
rect 7362 21310 7374 21362
rect 5966 21298 6018 21310
rect 12126 21298 12178 21310
rect 12910 21362 12962 21374
rect 19854 21362 19906 21374
rect 15698 21310 15710 21362
rect 15762 21310 15774 21362
rect 12910 21298 12962 21310
rect 19854 21298 19906 21310
rect 25902 21362 25954 21374
rect 25902 21298 25954 21310
rect 672 21194 27888 21228
rect 672 21142 4466 21194
rect 4518 21142 4570 21194
rect 4622 21142 4674 21194
rect 4726 21142 24466 21194
rect 24518 21142 24570 21194
rect 24622 21142 24674 21194
rect 24726 21142 27888 21194
rect 672 21108 27888 21142
rect 7870 21026 7922 21038
rect 7870 20962 7922 20974
rect 9774 21026 9826 21038
rect 9774 20962 9826 20974
rect 17614 21026 17666 21038
rect 19854 21026 19906 21038
rect 18722 20974 18734 21026
rect 18786 20974 18798 21026
rect 17614 20962 17666 20974
rect 19854 20962 19906 20974
rect 27470 21026 27522 21038
rect 27470 20962 27522 20974
rect 1374 20914 1426 20926
rect 1374 20850 1426 20862
rect 1934 20914 1986 20926
rect 1934 20850 1986 20862
rect 2270 20914 2322 20926
rect 3726 20914 3778 20926
rect 9886 20914 9938 20926
rect 17054 20914 17106 20926
rect 26014 20914 26066 20926
rect 3266 20862 3278 20914
rect 3330 20862 3342 20914
rect 6626 20862 6638 20914
rect 6690 20862 6702 20914
rect 13906 20862 13918 20914
rect 13970 20862 13982 20914
rect 20402 20862 20414 20914
rect 20466 20862 20478 20914
rect 20738 20862 20750 20914
rect 20802 20862 20814 20914
rect 2270 20850 2322 20862
rect 3726 20850 3778 20862
rect 9886 20850 9938 20862
rect 17054 20850 17106 20862
rect 26014 20850 26066 20862
rect 26910 20914 26962 20926
rect 26910 20850 26962 20862
rect 9998 20802 10050 20814
rect 2594 20750 2606 20802
rect 2658 20750 2670 20802
rect 3042 20750 3054 20802
rect 3106 20750 3118 20802
rect 4498 20750 4510 20802
rect 4562 20750 4574 20802
rect 5282 20750 5294 20802
rect 5346 20750 5358 20802
rect 6178 20750 6190 20802
rect 6242 20750 6254 20802
rect 9426 20750 9438 20802
rect 9490 20750 9502 20802
rect 9998 20738 10050 20750
rect 10446 20802 10498 20814
rect 14590 20802 14642 20814
rect 20190 20802 20242 20814
rect 10994 20750 11006 20802
rect 11058 20750 11070 20802
rect 11554 20750 11566 20802
rect 11618 20750 11630 20802
rect 11890 20750 11902 20802
rect 11954 20750 11966 20802
rect 13346 20750 13358 20802
rect 13410 20750 13422 20802
rect 13794 20750 13806 20802
rect 13858 20750 13870 20802
rect 14914 20750 14926 20802
rect 14978 20750 14990 20802
rect 15922 20750 15934 20802
rect 15986 20750 15998 20802
rect 16706 20750 16718 20802
rect 16770 20750 16782 20802
rect 10446 20738 10498 20750
rect 14590 20738 14642 20750
rect 20190 20738 20242 20750
rect 26574 20802 26626 20814
rect 26574 20738 26626 20750
rect 12910 20690 12962 20702
rect 11778 20638 11790 20690
rect 11842 20638 11854 20690
rect 19170 20638 19182 20690
rect 19234 20638 19246 20690
rect 12910 20626 12962 20638
rect 16718 20578 16770 20590
rect 10770 20526 10782 20578
rect 10834 20526 10846 20578
rect 16718 20514 16770 20526
rect 672 20410 27888 20444
rect 672 20358 3806 20410
rect 3858 20358 3910 20410
rect 3962 20358 4014 20410
rect 4066 20358 23806 20410
rect 23858 20358 23910 20410
rect 23962 20358 24014 20410
rect 24066 20358 27888 20410
rect 672 20324 27888 20358
rect 12002 20190 12014 20242
rect 12066 20190 12078 20242
rect 16034 20190 16046 20242
rect 16098 20190 16110 20242
rect 2046 20130 2098 20142
rect 2046 20066 2098 20078
rect 2830 20130 2882 20142
rect 2830 20066 2882 20078
rect 6190 20130 6242 20142
rect 10558 20130 10610 20142
rect 6738 20078 6750 20130
rect 6802 20078 6814 20130
rect 6190 20066 6242 20078
rect 10558 20066 10610 20078
rect 12910 20130 12962 20142
rect 19742 20130 19794 20142
rect 15026 20078 15038 20130
rect 15090 20078 15102 20130
rect 18162 20078 18174 20130
rect 18226 20078 18238 20130
rect 27010 20078 27022 20130
rect 27074 20078 27086 20130
rect 12910 20066 12962 20078
rect 19742 20066 19794 20078
rect 8318 20018 8370 20030
rect 11454 20018 11506 20030
rect 13246 20018 13298 20030
rect 15822 20018 15874 20030
rect 27470 20018 27522 20030
rect 1026 19966 1038 20018
rect 1090 19966 1102 20018
rect 1250 19966 1262 20018
rect 1314 19966 1326 20018
rect 3602 19966 3614 20018
rect 3666 19966 3678 20018
rect 6626 19966 6638 20018
rect 6690 19966 6702 20018
rect 8978 19966 8990 20018
rect 9042 19966 9054 20018
rect 12226 19966 12238 20018
rect 12290 19966 12302 20018
rect 14690 19966 14702 20018
rect 14754 19966 14766 20018
rect 16034 19966 16046 20018
rect 16098 19966 16110 20018
rect 8318 19954 8370 19966
rect 11454 19954 11506 19966
rect 13246 19954 13298 19966
rect 15822 19954 15874 19966
rect 27470 19954 27522 19966
rect 15486 19906 15538 19918
rect 7186 19854 7198 19906
rect 7250 19854 7262 19906
rect 9314 19854 9326 19906
rect 9378 19854 9390 19906
rect 11666 19854 11678 19906
rect 11730 19854 11742 19906
rect 13458 19854 13470 19906
rect 13522 19854 13534 19906
rect 13794 19854 13806 19906
rect 13858 19854 13870 19906
rect 14018 19854 14030 19906
rect 14082 19854 14094 19906
rect 15698 19854 15710 19906
rect 15762 19854 15774 19906
rect 15486 19842 15538 19854
rect 5630 19794 5682 19806
rect 15598 19794 15650 19806
rect 11778 19742 11790 19794
rect 11842 19742 11854 19794
rect 18610 19742 18622 19794
rect 18674 19742 18686 19794
rect 5630 19730 5682 19742
rect 15598 19730 15650 19742
rect 672 19626 27888 19660
rect 672 19574 4466 19626
rect 4518 19574 4570 19626
rect 4622 19574 4674 19626
rect 4726 19574 24466 19626
rect 24518 19574 24570 19626
rect 24622 19574 24674 19626
rect 24726 19574 27888 19626
rect 672 19540 27888 19574
rect 1598 19458 1650 19470
rect 5742 19458 5794 19470
rect 2706 19406 2718 19458
rect 2770 19406 2782 19458
rect 1598 19394 1650 19406
rect 5742 19394 5794 19406
rect 8206 19458 8258 19470
rect 27470 19458 27522 19470
rect 11554 19406 11566 19458
rect 11618 19406 11630 19458
rect 8206 19394 8258 19406
rect 27470 19394 27522 19406
rect 11118 19346 11170 19358
rect 4498 19294 4510 19346
rect 4562 19294 4574 19346
rect 7074 19294 7086 19346
rect 7138 19294 7150 19346
rect 11118 19282 11170 19294
rect 12574 19346 12626 19358
rect 14366 19346 14418 19358
rect 13906 19294 13918 19346
rect 13970 19294 13982 19346
rect 12574 19282 12626 19294
rect 14366 19282 14418 19294
rect 16718 19346 16770 19358
rect 16718 19282 16770 19294
rect 16942 19346 16994 19358
rect 16942 19282 16994 19294
rect 26014 19346 26066 19358
rect 26014 19282 26066 19294
rect 26574 19234 26626 19246
rect 9538 19182 9550 19234
rect 9602 19182 9614 19234
rect 10322 19182 10334 19234
rect 10386 19182 10398 19234
rect 11778 19182 11790 19234
rect 11842 19182 11854 19234
rect 12226 19182 12238 19234
rect 12290 19182 12302 19234
rect 13346 19182 13358 19234
rect 13410 19182 13422 19234
rect 13682 19182 13694 19234
rect 13746 19182 13758 19234
rect 15026 19182 15038 19234
rect 15090 19182 15102 19234
rect 15922 19182 15934 19234
rect 15986 19182 15998 19234
rect 26574 19170 26626 19182
rect 12910 19122 12962 19134
rect 3154 19070 3166 19122
rect 3218 19070 3230 19122
rect 4162 19070 4174 19122
rect 4226 19070 4238 19122
rect 6626 19070 6638 19122
rect 6690 19070 6702 19122
rect 12910 19058 12962 19070
rect 16830 19122 16882 19134
rect 27010 19070 27022 19122
rect 27074 19070 27086 19122
rect 16830 19058 16882 19070
rect 672 18842 27888 18876
rect 672 18790 3806 18842
rect 3858 18790 3910 18842
rect 3962 18790 4014 18842
rect 4066 18790 23806 18842
rect 23858 18790 23910 18842
rect 23962 18790 24014 18842
rect 24066 18790 27888 18842
rect 672 18756 27888 18790
rect 13806 18674 13858 18686
rect 13806 18610 13858 18622
rect 15822 18674 15874 18686
rect 15822 18610 15874 18622
rect 16046 18562 16098 18574
rect 8082 18510 8094 18562
rect 8146 18510 8158 18562
rect 10322 18510 10334 18562
rect 10386 18510 10398 18562
rect 16046 18498 16098 18510
rect 17054 18562 17106 18574
rect 26114 18510 26126 18562
rect 26178 18510 26190 18562
rect 17054 18498 17106 18510
rect 3166 18450 3218 18462
rect 2706 18398 2718 18450
rect 2770 18398 2782 18450
rect 3166 18386 3218 18398
rect 4398 18450 4450 18462
rect 7198 18450 7250 18462
rect 15598 18450 15650 18462
rect 5618 18398 5630 18450
rect 5682 18398 5694 18450
rect 14578 18398 14590 18450
rect 14642 18398 14654 18450
rect 4398 18386 4450 18398
rect 7198 18386 7250 18398
rect 15598 18386 15650 18398
rect 16494 18450 16546 18462
rect 16494 18386 16546 18398
rect 19518 18450 19570 18462
rect 19518 18386 19570 18398
rect 26910 18450 26962 18462
rect 26910 18386 26962 18398
rect 27470 18450 27522 18462
rect 27470 18386 27522 18398
rect 11902 18338 11954 18350
rect 15262 18338 15314 18350
rect 2258 18286 2270 18338
rect 2322 18286 2334 18338
rect 8530 18286 8542 18338
rect 8594 18286 8606 18338
rect 10658 18286 10670 18338
rect 10722 18286 10734 18338
rect 14466 18286 14478 18338
rect 14530 18286 14542 18338
rect 11902 18274 11954 18286
rect 15262 18274 15314 18286
rect 17390 18338 17442 18350
rect 17390 18274 17442 18286
rect 1710 18226 1762 18238
rect 1710 18162 1762 18174
rect 3838 18226 3890 18238
rect 9662 18226 9714 18238
rect 6066 18174 6078 18226
rect 6130 18174 6142 18226
rect 3838 18162 3890 18174
rect 9662 18162 9714 18174
rect 13470 18226 13522 18238
rect 13470 18162 13522 18174
rect 15150 18226 15202 18238
rect 15150 18162 15202 18174
rect 16270 18226 16322 18238
rect 16270 18162 16322 18174
rect 16382 18226 16434 18238
rect 16382 18162 16434 18174
rect 16942 18226 16994 18238
rect 16942 18162 16994 18174
rect 17166 18226 17218 18238
rect 17166 18162 17218 18174
rect 18958 18226 19010 18238
rect 18958 18162 19010 18174
rect 26574 18226 26626 18238
rect 26574 18162 26626 18174
rect 672 18058 27888 18092
rect 672 18006 4466 18058
rect 4518 18006 4570 18058
rect 4622 18006 4674 18058
rect 4726 18006 24466 18058
rect 24518 18006 24570 18058
rect 24622 18006 24674 18058
rect 24726 18006 27888 18058
rect 672 17972 27888 18006
rect 1038 17890 1090 17902
rect 1038 17826 1090 17838
rect 3726 17890 3778 17902
rect 27470 17890 27522 17902
rect 4834 17838 4846 17890
rect 4898 17838 4910 17890
rect 3726 17826 3778 17838
rect 27470 17826 27522 17838
rect 1598 17778 1650 17790
rect 14030 17778 14082 17790
rect 16046 17778 16098 17790
rect 2594 17726 2606 17778
rect 2658 17726 2670 17778
rect 6962 17726 6974 17778
rect 7026 17726 7038 17778
rect 9986 17726 9998 17778
rect 10050 17726 10062 17778
rect 14466 17726 14478 17778
rect 14530 17726 14542 17778
rect 1598 17714 1650 17726
rect 14030 17714 14082 17726
rect 16046 17714 16098 17726
rect 26014 17778 26066 17790
rect 26014 17714 26066 17726
rect 26910 17778 26962 17790
rect 26910 17714 26962 17726
rect 26574 17666 26626 17678
rect 2146 17614 2158 17666
rect 2210 17614 2222 17666
rect 4274 17614 4286 17666
rect 4338 17614 4350 17666
rect 6626 17614 6638 17666
rect 6690 17614 6702 17666
rect 12338 17614 12350 17666
rect 12402 17614 12414 17666
rect 13234 17614 13246 17666
rect 13298 17614 13310 17666
rect 14578 17602 14590 17654
rect 14642 17602 14654 17654
rect 15026 17614 15038 17666
rect 15090 17614 15102 17666
rect 26574 17602 26626 17614
rect 11230 17554 11282 17566
rect 9650 17502 9662 17554
rect 9714 17502 9726 17554
rect 11230 17490 11282 17502
rect 15486 17554 15538 17566
rect 16146 17502 16158 17554
rect 16210 17502 16222 17554
rect 15486 17490 15538 17502
rect 5966 17442 6018 17454
rect 5966 17378 6018 17390
rect 8206 17442 8258 17454
rect 8206 17378 8258 17390
rect 15822 17442 15874 17454
rect 15822 17378 15874 17390
rect 672 17274 27888 17308
rect 672 17222 3806 17274
rect 3858 17222 3910 17274
rect 3962 17222 4014 17274
rect 4066 17222 23806 17274
rect 23858 17222 23910 17274
rect 23962 17222 24014 17274
rect 24066 17222 27888 17274
rect 672 17188 27888 17222
rect 8318 17106 8370 17118
rect 8318 17042 8370 17054
rect 13134 17106 13186 17118
rect 13134 17042 13186 17054
rect 14254 17106 14306 17118
rect 14254 17042 14306 17054
rect 2494 16994 2546 17006
rect 12238 16994 12290 17006
rect 1474 16942 1486 16994
rect 1538 16942 1550 16994
rect 3266 16942 3278 16994
rect 3330 16942 3342 16994
rect 5842 16942 5854 16994
rect 5906 16942 5918 16994
rect 10210 16942 10222 16994
rect 10274 16942 10286 16994
rect 12898 16942 12910 16994
rect 12962 16942 12974 16994
rect 27010 16942 27022 16994
rect 27074 16942 27086 16994
rect 2494 16930 2546 16942
rect 12238 16930 12290 16942
rect 1934 16882 1986 16894
rect 1138 16830 1150 16882
rect 1202 16830 1214 16882
rect 1934 16818 1986 16830
rect 2830 16882 2882 16894
rect 2830 16818 2882 16830
rect 3838 16882 3890 16894
rect 10894 16882 10946 16894
rect 4274 16830 4286 16882
rect 4338 16830 4350 16882
rect 4946 16830 4958 16882
rect 5010 16830 5022 16882
rect 6626 16830 6638 16882
rect 6690 16830 6702 16882
rect 10546 16830 10558 16882
rect 10610 16830 10622 16882
rect 3838 16818 3890 16830
rect 10894 16818 10946 16830
rect 11006 16882 11058 16894
rect 13806 16882 13858 16894
rect 27470 16882 27522 16894
rect 11778 16830 11790 16882
rect 11842 16830 11854 16882
rect 14018 16830 14030 16882
rect 14082 16830 14094 16882
rect 14354 16830 14366 16882
rect 14418 16830 14430 16882
rect 15250 16830 15262 16882
rect 15314 16830 15326 16882
rect 15810 16830 15822 16882
rect 15874 16830 15886 16882
rect 16482 16830 16494 16882
rect 16546 16830 16558 16882
rect 16930 16830 16942 16882
rect 16994 16830 17006 16882
rect 17938 16830 17950 16882
rect 18002 16830 18014 16882
rect 11006 16818 11058 16830
rect 13806 16818 13858 16830
rect 27470 16818 27522 16830
rect 9886 16770 9938 16782
rect 7074 16718 7086 16770
rect 7138 16718 7150 16770
rect 9886 16706 9938 16718
rect 10110 16770 10162 16782
rect 10110 16706 10162 16718
rect 11342 16770 11394 16782
rect 11342 16706 11394 16718
rect 12910 16770 12962 16782
rect 12910 16706 12962 16718
rect 14926 16770 14978 16782
rect 15922 16718 15934 16770
rect 15986 16718 15998 16770
rect 14926 16706 14978 16718
rect 11230 16658 11282 16670
rect 11230 16594 11282 16606
rect 14590 16658 14642 16670
rect 14590 16594 14642 16606
rect 672 16490 27888 16524
rect 672 16438 4466 16490
rect 4518 16438 4570 16490
rect 4622 16438 4674 16490
rect 4726 16438 24466 16490
rect 24518 16438 24570 16490
rect 24622 16438 24674 16490
rect 24726 16438 27888 16490
rect 672 16404 27888 16438
rect 27470 16322 27522 16334
rect 11778 16270 11790 16322
rect 11842 16270 11854 16322
rect 17938 16270 17950 16322
rect 18002 16270 18014 16322
rect 27470 16258 27522 16270
rect 9550 16210 9602 16222
rect 3154 16158 3166 16210
rect 3218 16158 3230 16210
rect 4722 16158 4734 16210
rect 4786 16158 4798 16210
rect 6850 16158 6862 16210
rect 6914 16158 6926 16210
rect 9550 16146 9602 16158
rect 10110 16210 10162 16222
rect 10110 16146 10162 16158
rect 10334 16210 10386 16222
rect 10334 16146 10386 16158
rect 10782 16210 10834 16222
rect 10782 16146 10834 16158
rect 12238 16210 12290 16222
rect 12238 16146 12290 16158
rect 15262 16210 15314 16222
rect 15262 16146 15314 16158
rect 15710 16210 15762 16222
rect 15710 16146 15762 16158
rect 9886 16098 9938 16110
rect 3490 16046 3502 16098
rect 3554 16046 3566 16098
rect 4274 16046 4286 16098
rect 4338 16046 4350 16098
rect 6514 16046 6526 16098
rect 6578 16046 6590 16098
rect 9090 16046 9102 16098
rect 9154 16046 9166 16098
rect 9314 16046 9326 16098
rect 9378 16046 9390 16098
rect 9886 16034 9938 16046
rect 9998 16098 10050 16110
rect 16270 16098 16322 16110
rect 11106 16046 11118 16098
rect 11170 16046 11182 16098
rect 11666 16046 11678 16098
rect 11730 16046 11742 16098
rect 12786 16046 12798 16098
rect 12850 16046 12862 16098
rect 13010 16046 13022 16098
rect 13074 16046 13086 16098
rect 13906 16046 13918 16098
rect 13970 16046 13982 16098
rect 15922 16046 15934 16098
rect 15986 16046 15998 16098
rect 9998 16034 10050 16046
rect 16270 16034 16322 16046
rect 26574 16098 26626 16110
rect 26574 16034 26626 16046
rect 8094 15986 8146 15998
rect 8094 15922 8146 15934
rect 15374 15986 15426 15998
rect 26014 15986 26066 15998
rect 18386 15934 18398 15986
rect 18450 15934 18462 15986
rect 27010 15934 27022 15986
rect 27074 15934 27086 15986
rect 15374 15922 15426 15934
rect 26014 15922 26066 15934
rect 1934 15874 1986 15886
rect 1934 15810 1986 15822
rect 5854 15874 5906 15886
rect 5854 15810 5906 15822
rect 9662 15874 9714 15886
rect 9662 15810 9714 15822
rect 16046 15874 16098 15886
rect 16046 15810 16098 15822
rect 16830 15874 16882 15886
rect 16830 15810 16882 15822
rect 672 15706 27888 15740
rect 672 15654 3806 15706
rect 3858 15654 3910 15706
rect 3962 15654 4014 15706
rect 4066 15654 23806 15706
rect 23858 15654 23910 15706
rect 23962 15654 24014 15706
rect 24066 15654 27888 15706
rect 672 15620 27888 15654
rect 7310 15538 7362 15550
rect 7310 15474 7362 15486
rect 11230 15538 11282 15550
rect 11230 15474 11282 15486
rect 11902 15538 11954 15550
rect 11902 15474 11954 15486
rect 9550 15426 9602 15438
rect 5730 15374 5742 15426
rect 5794 15374 5806 15426
rect 9550 15362 9602 15374
rect 11006 15426 11058 15438
rect 11006 15362 11058 15374
rect 15262 15426 15314 15438
rect 26114 15374 26126 15426
rect 26178 15374 26190 15426
rect 27010 15374 27022 15426
rect 27074 15374 27086 15426
rect 15262 15362 15314 15374
rect 10558 15314 10610 15326
rect 3602 15262 3614 15314
rect 3666 15262 3678 15314
rect 7858 15262 7870 15314
rect 7922 15262 7934 15314
rect 10558 15250 10610 15262
rect 11454 15314 11506 15326
rect 15374 15314 15426 15326
rect 27470 15314 27522 15326
rect 13570 15262 13582 15314
rect 13634 15262 13646 15314
rect 18610 15262 18622 15314
rect 18674 15262 18686 15314
rect 11454 15250 11506 15262
rect 15374 15250 15426 15262
rect 27470 15250 27522 15262
rect 10110 15202 10162 15214
rect 3042 15150 3054 15202
rect 3106 15150 3118 15202
rect 6178 15150 6190 15202
rect 6242 15150 6254 15202
rect 8306 15150 8318 15202
rect 8370 15150 8382 15202
rect 10110 15138 10162 15150
rect 11790 15202 11842 15214
rect 11790 15138 11842 15150
rect 11902 15202 11954 15214
rect 11902 15138 11954 15150
rect 13358 15202 13410 15214
rect 13358 15138 13410 15150
rect 14926 15202 14978 15214
rect 14926 15138 14978 15150
rect 15150 15202 15202 15214
rect 15150 15138 15202 15150
rect 15822 15202 15874 15214
rect 15822 15138 15874 15150
rect 15934 15202 15986 15214
rect 15934 15138 15986 15150
rect 16046 15202 16098 15214
rect 16046 15138 16098 15150
rect 16942 15202 16994 15214
rect 18050 15150 18062 15202
rect 18114 15150 18126 15202
rect 16942 15138 16994 15150
rect 1934 15090 1986 15102
rect 1934 15026 1986 15038
rect 9998 15090 10050 15102
rect 9998 15026 10050 15038
rect 10670 15090 10722 15102
rect 10670 15026 10722 15038
rect 10782 15090 10834 15102
rect 26574 15090 26626 15102
rect 16482 15038 16494 15090
rect 16546 15038 16558 15090
rect 10782 15026 10834 15038
rect 26574 15026 26626 15038
rect 672 14922 27888 14956
rect 672 14870 4466 14922
rect 4518 14870 4570 14922
rect 4622 14870 4674 14922
rect 4726 14870 24466 14922
rect 24518 14870 24570 14922
rect 24622 14870 24674 14922
rect 24726 14870 27888 14922
rect 672 14836 27888 14870
rect 1038 14754 1090 14766
rect 1038 14690 1090 14702
rect 2830 14754 2882 14766
rect 2830 14690 2882 14702
rect 11118 14754 11170 14766
rect 11118 14690 11170 14702
rect 11230 14754 11282 14766
rect 11230 14690 11282 14702
rect 15486 14754 15538 14766
rect 15486 14690 15538 14702
rect 16270 14754 16322 14766
rect 16270 14690 16322 14702
rect 17614 14754 17666 14766
rect 17614 14690 17666 14702
rect 27470 14754 27522 14766
rect 27470 14690 27522 14702
rect 2494 14642 2546 14654
rect 5966 14642 6018 14654
rect 5506 14590 5518 14642
rect 5570 14590 5582 14642
rect 2494 14578 2546 14590
rect 5966 14578 6018 14590
rect 9438 14642 9490 14654
rect 9438 14578 9490 14590
rect 9550 14642 9602 14654
rect 9550 14578 9602 14590
rect 10110 14642 10162 14654
rect 10110 14578 10162 14590
rect 10222 14642 10274 14654
rect 16046 14642 16098 14654
rect 14242 14590 14254 14642
rect 14306 14590 14318 14642
rect 10222 14578 10274 14590
rect 16046 14578 16098 14590
rect 1934 14530 1986 14542
rect 9998 14530 10050 14542
rect 15934 14530 15986 14542
rect 4834 14478 4846 14530
rect 4898 14478 4910 14530
rect 5282 14478 5294 14530
rect 5346 14478 5358 14530
rect 6514 14478 6526 14530
rect 6578 14478 6590 14530
rect 7634 14478 7646 14530
rect 7698 14478 7710 14530
rect 10658 14478 10670 14530
rect 10722 14478 10734 14530
rect 1934 14466 1986 14478
rect 9998 14466 10050 14478
rect 15934 14466 15986 14478
rect 16718 14530 16770 14542
rect 16718 14466 16770 14478
rect 17166 14530 17218 14542
rect 17166 14466 17218 14478
rect 17390 14530 17442 14542
rect 17390 14466 17442 14478
rect 26574 14530 26626 14542
rect 26574 14466 26626 14478
rect 1598 14418 1650 14430
rect 4510 14418 4562 14430
rect 26910 14418 26962 14430
rect 3266 14366 3278 14418
rect 3330 14366 3342 14418
rect 13906 14366 13918 14418
rect 13970 14366 13982 14418
rect 17490 14366 17502 14418
rect 17554 14366 17566 14418
rect 26114 14366 26126 14418
rect 26178 14366 26190 14418
rect 1598 14354 1650 14366
rect 4510 14354 4562 14366
rect 26910 14354 26962 14366
rect 9438 14306 9490 14318
rect 9438 14242 9490 14254
rect 11006 14306 11058 14318
rect 11006 14242 11058 14254
rect 16942 14306 16994 14318
rect 16942 14242 16994 14254
rect 672 14138 27888 14172
rect 672 14086 3806 14138
rect 3858 14086 3910 14138
rect 3962 14086 4014 14138
rect 4066 14086 23806 14138
rect 23858 14086 23910 14138
rect 23962 14086 24014 14138
rect 24066 14086 27888 14138
rect 672 14052 27888 14086
rect 7422 13970 7474 13982
rect 7422 13906 7474 13918
rect 15374 13970 15426 13982
rect 15374 13906 15426 13918
rect 17390 13970 17442 13982
rect 17390 13906 17442 13918
rect 16382 13858 16434 13870
rect 16382 13794 16434 13806
rect 2606 13746 2658 13758
rect 16046 13746 16098 13758
rect 1474 13694 1486 13746
rect 1538 13694 1550 13746
rect 1922 13694 1934 13746
rect 1986 13694 1998 13746
rect 3378 13694 3390 13746
rect 3442 13694 3454 13746
rect 4274 13694 4286 13746
rect 4338 13694 4350 13746
rect 5170 13694 5182 13746
rect 5234 13694 5246 13746
rect 8194 13694 8206 13746
rect 8258 13694 8270 13746
rect 9314 13694 9326 13746
rect 9378 13694 9390 13746
rect 13122 13694 13134 13746
rect 13186 13694 13198 13746
rect 15698 13694 15710 13746
rect 15762 13694 15774 13746
rect 2606 13682 2658 13694
rect 16046 13682 16098 13694
rect 16158 13746 16210 13758
rect 16158 13682 16210 13694
rect 16494 13746 16546 13758
rect 17054 13746 17106 13758
rect 16818 13694 16830 13746
rect 16882 13694 16894 13746
rect 16494 13682 16546 13694
rect 17054 13682 17106 13694
rect 17278 13746 17330 13758
rect 17278 13682 17330 13694
rect 27470 13746 27522 13758
rect 27470 13682 27522 13694
rect 1150 13634 1202 13646
rect 15262 13634 15314 13646
rect 5618 13582 5630 13634
rect 5682 13582 5694 13634
rect 9762 13582 9774 13634
rect 9826 13582 9838 13634
rect 13682 13582 13694 13634
rect 13746 13582 13758 13634
rect 1150 13570 1202 13582
rect 15262 13570 15314 13582
rect 26910 13634 26962 13646
rect 26910 13570 26962 13582
rect 6750 13522 6802 13534
rect 2146 13470 2158 13522
rect 2210 13470 2222 13522
rect 6750 13458 6802 13470
rect 11006 13522 11058 13534
rect 11006 13458 11058 13470
rect 14814 13522 14866 13534
rect 14814 13458 14866 13470
rect 672 13354 27888 13388
rect 672 13302 4466 13354
rect 4518 13302 4570 13354
rect 4622 13302 4674 13354
rect 4726 13302 24466 13354
rect 24518 13302 24570 13354
rect 24622 13302 24674 13354
rect 24726 13302 27888 13354
rect 672 13268 27888 13302
rect 7758 13186 7810 13198
rect 7758 13122 7810 13134
rect 15374 13186 15426 13198
rect 15374 13122 15426 13134
rect 16046 13186 16098 13198
rect 16046 13122 16098 13134
rect 27470 13186 27522 13198
rect 27470 13122 27522 13134
rect 12798 13074 12850 13086
rect 2594 13022 2606 13074
rect 2658 13022 2670 13074
rect 5170 13022 5182 13074
rect 5234 13022 5246 13074
rect 9426 13022 9438 13074
rect 9490 13022 9502 13074
rect 12798 13010 12850 13022
rect 14478 13074 14530 13086
rect 14478 13010 14530 13022
rect 14814 13074 14866 13086
rect 14814 13010 14866 13022
rect 15262 13074 15314 13086
rect 15262 13010 15314 13022
rect 26014 13074 26066 13086
rect 26014 13010 26066 13022
rect 1038 12962 1090 12974
rect 3726 12962 3778 12974
rect 5854 12962 5906 12974
rect 11342 12962 11394 12974
rect 2146 12910 2158 12962
rect 2210 12910 2222 12962
rect 4498 12910 4510 12962
rect 4562 12910 4574 12962
rect 4946 12910 4958 12962
rect 5010 12910 5022 12962
rect 6402 12910 6414 12962
rect 6466 12910 6478 12962
rect 7298 12910 7310 12962
rect 7362 12910 7374 12962
rect 1038 12898 1090 12910
rect 3726 12898 3778 12910
rect 5854 12898 5906 12910
rect 11342 12898 11394 12910
rect 12238 12962 12290 12974
rect 12238 12898 12290 12910
rect 15486 12962 15538 12974
rect 15486 12898 15538 12910
rect 16158 12962 16210 12974
rect 16158 12898 16210 12910
rect 26574 12962 26626 12974
rect 26574 12898 26626 12910
rect 1598 12850 1650 12862
rect 1598 12786 1650 12798
rect 4174 12850 4226 12862
rect 11902 12850 11954 12862
rect 8194 12798 8206 12850
rect 8258 12798 8270 12850
rect 9090 12798 9102 12850
rect 9154 12798 9166 12850
rect 27010 12798 27022 12850
rect 27074 12798 27086 12850
rect 4174 12786 4226 12798
rect 11902 12786 11954 12798
rect 10670 12738 10722 12750
rect 10670 12674 10722 12686
rect 672 12570 27888 12604
rect 672 12518 3806 12570
rect 3858 12518 3910 12570
rect 3962 12518 4014 12570
rect 4066 12518 23806 12570
rect 23858 12518 23910 12570
rect 23962 12518 24014 12570
rect 24066 12518 27888 12570
rect 672 12484 27888 12518
rect 1038 12290 1090 12302
rect 4286 12290 4338 12302
rect 3266 12238 3278 12290
rect 3330 12238 3342 12290
rect 1038 12226 1090 12238
rect 4286 12226 4338 12238
rect 5966 12290 6018 12302
rect 5966 12226 6018 12238
rect 26014 12290 26066 12302
rect 26014 12226 26066 12238
rect 26910 12290 26962 12302
rect 26910 12226 26962 12238
rect 1934 12178 1986 12190
rect 3726 12178 3778 12190
rect 8542 12178 8594 12190
rect 10670 12178 10722 12190
rect 27470 12178 27522 12190
rect 1474 12126 1486 12178
rect 1538 12126 1550 12178
rect 2930 12126 2942 12178
rect 2994 12126 3006 12178
rect 5506 12126 5518 12178
rect 5570 12126 5582 12178
rect 6962 12126 6974 12178
rect 7026 12126 7038 12178
rect 9314 12126 9326 12178
rect 9378 12126 9390 12178
rect 9762 12126 9774 12178
rect 9826 12126 9838 12178
rect 11218 12126 11230 12178
rect 11282 12126 11294 12178
rect 12002 12126 12014 12178
rect 12066 12126 12078 12178
rect 13122 12126 13134 12178
rect 13186 12126 13198 12178
rect 13570 12126 13582 12178
rect 13634 12126 13646 12178
rect 15026 12126 15038 12178
rect 15090 12126 15102 12178
rect 15810 12126 15822 12178
rect 15874 12126 15886 12178
rect 1934 12114 1986 12126
rect 3726 12114 3778 12126
rect 8542 12114 8594 12126
rect 10670 12114 10722 12126
rect 27470 12114 27522 12126
rect 2494 12066 2546 12078
rect 8990 12066 9042 12078
rect 12798 12066 12850 12078
rect 7298 12014 7310 12066
rect 7362 12014 7374 12066
rect 9986 12014 9998 12066
rect 10050 12014 10062 12066
rect 2494 12002 2546 12014
rect 8990 12002 9042 12014
rect 12798 12002 12850 12014
rect 14254 12066 14306 12078
rect 14254 12002 14306 12014
rect 26574 11954 26626 11966
rect 13794 11902 13806 11954
rect 13858 11902 13870 11954
rect 26574 11890 26626 11902
rect 672 11786 27888 11820
rect 672 11734 4466 11786
rect 4518 11734 4570 11786
rect 4622 11734 4674 11786
rect 4726 11734 24466 11786
rect 24518 11734 24570 11786
rect 24622 11734 24674 11786
rect 24726 11734 27888 11786
rect 672 11700 27888 11734
rect 2606 11618 2658 11630
rect 27470 11618 27522 11630
rect 4834 11566 4846 11618
rect 4898 11566 4910 11618
rect 7074 11566 7086 11618
rect 7138 11566 7150 11618
rect 10882 11566 10894 11618
rect 10946 11566 10958 11618
rect 2606 11554 2658 11566
rect 27470 11554 27522 11566
rect 9886 11506 9938 11518
rect 26014 11506 26066 11518
rect 2258 11454 2270 11506
rect 2322 11454 2334 11506
rect 14690 11454 14702 11506
rect 14754 11454 14766 11506
rect 15138 11454 15150 11506
rect 15202 11454 15214 11506
rect 9886 11442 9938 11454
rect 26014 11442 26066 11454
rect 8206 11394 8258 11406
rect 26574 11394 26626 11406
rect 6626 11342 6638 11394
rect 6690 11342 6702 11394
rect 10210 11342 10222 11394
rect 10274 11342 10286 11394
rect 10770 11342 10782 11394
rect 10834 11342 10846 11394
rect 11442 11342 11454 11394
rect 11506 11342 11518 11394
rect 12002 11342 12014 11394
rect 12066 11342 12078 11394
rect 12898 11342 12910 11394
rect 12962 11342 12974 11394
rect 8206 11330 8258 11342
rect 26574 11330 26626 11342
rect 3166 11282 3218 11294
rect 26910 11282 26962 11294
rect 4386 11230 4398 11282
rect 4450 11230 4462 11282
rect 3166 11218 3218 11230
rect 26910 11218 26962 11230
rect 1262 11170 1314 11182
rect 1262 11106 1314 11118
rect 5966 11170 6018 11182
rect 5966 11106 6018 11118
rect 14142 11170 14194 11182
rect 14142 11106 14194 11118
rect 14478 11170 14530 11182
rect 14478 11106 14530 11118
rect 672 11002 27888 11036
rect 672 10950 3806 11002
rect 3858 10950 3910 11002
rect 3962 10950 4014 11002
rect 4066 10950 23806 11002
rect 23858 10950 23910 11002
rect 23962 10950 24014 11002
rect 24066 10950 27888 11002
rect 672 10916 27888 10950
rect 12126 10834 12178 10846
rect 12126 10770 12178 10782
rect 1598 10722 1650 10734
rect 5854 10722 5906 10734
rect 2370 10670 2382 10722
rect 2434 10670 2446 10722
rect 3266 10670 3278 10722
rect 3330 10670 3342 10722
rect 1598 10658 1650 10670
rect 5854 10658 5906 10670
rect 6750 10722 6802 10734
rect 6750 10658 6802 10670
rect 14030 10722 14082 10734
rect 14030 10658 14082 10670
rect 14926 10722 14978 10734
rect 14926 10658 14978 10670
rect 26910 10722 26962 10734
rect 26910 10658 26962 10670
rect 1038 10610 1090 10622
rect 1038 10546 1090 10558
rect 1934 10610 1986 10622
rect 5294 10610 5346 10622
rect 8206 10610 8258 10622
rect 14366 10610 14418 10622
rect 2930 10558 2942 10610
rect 2994 10558 3006 10610
rect 7074 10558 7086 10610
rect 7138 10558 7150 10610
rect 7634 10558 7646 10610
rect 7698 10558 7710 10610
rect 8754 10558 8766 10610
rect 8818 10558 8830 10610
rect 9874 10558 9886 10610
rect 9938 10558 9950 10610
rect 10434 10558 10446 10610
rect 10498 10558 10510 10610
rect 13570 10558 13582 10610
rect 13634 10558 13646 10610
rect 1934 10546 1986 10558
rect 5294 10546 5346 10558
rect 8206 10546 8258 10558
rect 14366 10546 14418 10558
rect 27470 10610 27522 10622
rect 27470 10546 27522 10558
rect 10882 10446 10894 10498
rect 10946 10446 10958 10498
rect 7746 10334 7758 10386
rect 7810 10334 7822 10386
rect 672 10218 27888 10252
rect 672 10166 4466 10218
rect 4518 10166 4570 10218
rect 4622 10166 4674 10218
rect 4726 10166 24466 10218
rect 24518 10166 24570 10218
rect 24622 10166 24674 10218
rect 24726 10166 27888 10218
rect 672 10132 27888 10166
rect 7534 10050 7586 10062
rect 7534 9986 7586 9998
rect 27470 10050 27522 10062
rect 27470 9986 27522 9998
rect 3166 9938 3218 9950
rect 3166 9874 3218 9886
rect 4734 9938 4786 9950
rect 4734 9874 4786 9886
rect 10110 9938 10162 9950
rect 26014 9938 26066 9950
rect 11106 9886 11118 9938
rect 11170 9886 11182 9938
rect 10110 9874 10162 9886
rect 26014 9874 26066 9886
rect 26910 9938 26962 9950
rect 26910 9874 26962 9886
rect 11566 9826 11618 9838
rect 26574 9826 26626 9838
rect 2034 9774 2046 9826
rect 2098 9774 2110 9826
rect 2706 9774 2718 9826
rect 2770 9774 2782 9826
rect 5170 9774 5182 9826
rect 5234 9774 5246 9826
rect 10434 9774 10446 9826
rect 10498 9774 10510 9826
rect 10882 9774 10894 9826
rect 10946 9774 10958 9826
rect 12338 9774 12350 9826
rect 12402 9774 12414 9826
rect 13234 9774 13246 9826
rect 13298 9774 13310 9826
rect 11566 9762 11618 9774
rect 26574 9762 26626 9774
rect 7074 9662 7086 9714
rect 7138 9662 7150 9714
rect 1262 9602 1314 9614
rect 1262 9538 1314 9550
rect 672 9434 27888 9468
rect 672 9382 3806 9434
rect 3858 9382 3910 9434
rect 3962 9382 4014 9434
rect 4066 9382 23806 9434
rect 23858 9382 23910 9434
rect 23962 9382 24014 9434
rect 24066 9382 27888 9434
rect 672 9348 27888 9382
rect 8878 9266 8930 9278
rect 8878 9202 8930 9214
rect 11118 9266 11170 9278
rect 11118 9202 11170 9214
rect 26014 9154 26066 9166
rect 1474 9102 1486 9154
rect 1538 9102 1550 9154
rect 9538 9102 9550 9154
rect 9602 9102 9614 9154
rect 27010 9102 27022 9154
rect 27074 9102 27086 9154
rect 26014 9090 26066 9102
rect 27470 9042 27522 9054
rect 1138 8990 1150 9042
rect 1202 8990 1214 9042
rect 2034 8990 2046 9042
rect 2098 8990 2110 9042
rect 7298 8990 7310 9042
rect 7362 8990 7374 9042
rect 27470 8978 27522 8990
rect 2494 8930 2546 8942
rect 7634 8878 7646 8930
rect 7698 8878 7710 8930
rect 9874 8878 9886 8930
rect 9938 8878 9950 8930
rect 2494 8866 2546 8878
rect 26574 8818 26626 8830
rect 26574 8754 26626 8766
rect 672 8650 27888 8684
rect 672 8598 4466 8650
rect 4518 8598 4570 8650
rect 4622 8598 4674 8650
rect 4726 8598 24466 8650
rect 24518 8598 24570 8650
rect 24622 8598 24674 8650
rect 24726 8598 27888 8650
rect 672 8564 27888 8598
rect 1038 8482 1090 8494
rect 1038 8418 1090 8430
rect 7758 8482 7810 8494
rect 7758 8418 7810 8430
rect 11342 8482 11394 8494
rect 11342 8418 11394 8430
rect 27470 8482 27522 8494
rect 27470 8418 27522 8430
rect 26014 8370 26066 8382
rect 10098 8318 10110 8370
rect 10162 8318 10174 8370
rect 26014 8306 26066 8318
rect 1598 8258 1650 8270
rect 26574 8258 26626 8270
rect 9650 8206 9662 8258
rect 9714 8206 9726 8258
rect 1598 8194 1650 8206
rect 26574 8194 26626 8206
rect 8318 8146 8370 8158
rect 8318 8082 8370 8094
rect 26910 8146 26962 8158
rect 26910 8082 26962 8094
rect 672 7866 27888 7900
rect 672 7814 3806 7866
rect 3858 7814 3910 7866
rect 3962 7814 4014 7866
rect 4066 7814 23806 7866
rect 23858 7814 23910 7866
rect 23962 7814 24014 7866
rect 24066 7814 27888 7866
rect 672 7780 27888 7814
rect 10670 7586 10722 7598
rect 1474 7534 1486 7586
rect 1538 7534 1550 7586
rect 10670 7522 10722 7534
rect 11566 7586 11618 7598
rect 11566 7522 11618 7534
rect 1038 7474 1090 7486
rect 1038 7410 1090 7422
rect 10110 7474 10162 7486
rect 10110 7410 10162 7422
rect 11006 7474 11058 7486
rect 11006 7410 11058 7422
rect 26910 7474 26962 7486
rect 26910 7410 26962 7422
rect 27470 7474 27522 7486
rect 27470 7410 27522 7422
rect 672 7082 27888 7116
rect 672 7030 4466 7082
rect 4518 7030 4570 7082
rect 4622 7030 4674 7082
rect 4726 7030 24466 7082
rect 24518 7030 24570 7082
rect 24622 7030 24674 7082
rect 24726 7030 27888 7082
rect 672 6996 27888 7030
rect 27470 6914 27522 6926
rect 27470 6850 27522 6862
rect 26574 6690 26626 6702
rect 2146 6638 2158 6690
rect 2210 6638 2222 6690
rect 26574 6626 26626 6638
rect 26910 6690 26962 6702
rect 26910 6626 26962 6638
rect 1262 6578 1314 6590
rect 1262 6514 1314 6526
rect 26014 6578 26066 6590
rect 26014 6514 26066 6526
rect 672 6298 27888 6332
rect 672 6246 3806 6298
rect 3858 6246 3910 6298
rect 3962 6246 4014 6298
rect 4066 6246 23806 6298
rect 23858 6246 23910 6298
rect 23962 6246 24014 6298
rect 24066 6246 27888 6298
rect 672 6212 27888 6246
rect 1262 6018 1314 6030
rect 1262 5954 1314 5966
rect 26910 6018 26962 6030
rect 26910 5954 26962 5966
rect 27470 5906 27522 5918
rect 2258 5854 2270 5906
rect 2322 5854 2334 5906
rect 27470 5842 27522 5854
rect 26014 5794 26066 5806
rect 26014 5730 26066 5742
rect 26574 5682 26626 5694
rect 26574 5618 26626 5630
rect 672 5514 27888 5548
rect 672 5462 4466 5514
rect 4518 5462 4570 5514
rect 4622 5462 4674 5514
rect 4726 5462 24466 5514
rect 24518 5462 24570 5514
rect 24622 5462 24674 5514
rect 24726 5462 27888 5514
rect 672 5428 27888 5462
rect 27470 5346 27522 5358
rect 27470 5282 27522 5294
rect 26014 5234 26066 5246
rect 26014 5170 26066 5182
rect 26910 5234 26962 5246
rect 26910 5170 26962 5182
rect 26574 5122 26626 5134
rect 26574 5058 26626 5070
rect 672 4730 27888 4764
rect 672 4678 3806 4730
rect 3858 4678 3910 4730
rect 3962 4678 4014 4730
rect 4066 4678 23806 4730
rect 23858 4678 23910 4730
rect 23962 4678 24014 4730
rect 24066 4678 27888 4730
rect 672 4644 27888 4678
rect 1474 4398 1486 4450
rect 1538 4398 1550 4450
rect 27010 4398 27022 4450
rect 27074 4398 27086 4450
rect 27470 4338 27522 4350
rect 27470 4274 27522 4286
rect 1038 4114 1090 4126
rect 1038 4050 1090 4062
rect 672 3946 27888 3980
rect 672 3894 4466 3946
rect 4518 3894 4570 3946
rect 4622 3894 4674 3946
rect 4726 3894 24466 3946
rect 24518 3894 24570 3946
rect 24622 3894 24674 3946
rect 24726 3894 27888 3946
rect 672 3860 27888 3894
rect 27470 3778 27522 3790
rect 27470 3714 27522 3726
rect 26574 3554 26626 3566
rect 26574 3490 26626 3502
rect 26014 3442 26066 3454
rect 26014 3378 26066 3390
rect 26910 3442 26962 3454
rect 26910 3378 26962 3390
rect 672 3162 27888 3196
rect 672 3110 3806 3162
rect 3858 3110 3910 3162
rect 3962 3110 4014 3162
rect 4066 3110 23806 3162
rect 23858 3110 23910 3162
rect 23962 3110 24014 3162
rect 24066 3110 27888 3162
rect 672 3076 27888 3110
rect 26014 2882 26066 2894
rect 26014 2818 26066 2830
rect 26910 2882 26962 2894
rect 26910 2818 26962 2830
rect 27470 2770 27522 2782
rect 27470 2706 27522 2718
rect 26574 2546 26626 2558
rect 26574 2482 26626 2494
rect 672 2378 27888 2412
rect 672 2326 4466 2378
rect 4518 2326 4570 2378
rect 4622 2326 4674 2378
rect 4726 2326 24466 2378
rect 24518 2326 24570 2378
rect 24622 2326 24674 2378
rect 24726 2326 27888 2378
rect 672 2292 27888 2326
rect 27470 2210 27522 2222
rect 27470 2146 27522 2158
rect 26014 2098 26066 2110
rect 26014 2034 26066 2046
rect 26574 1986 26626 1998
rect 26574 1922 26626 1934
rect 27010 1822 27022 1874
rect 27074 1822 27086 1874
rect 672 1594 27888 1628
rect 672 1542 3806 1594
rect 3858 1542 3910 1594
rect 3962 1542 4014 1594
rect 4066 1542 23806 1594
rect 23858 1542 23910 1594
rect 23962 1542 24014 1594
rect 24066 1542 27888 1594
rect 672 1508 27888 1542
rect 5518 1314 5570 1326
rect 5518 1250 5570 1262
rect 26574 1314 26626 1326
rect 26574 1250 26626 1262
rect 24782 1202 24834 1214
rect 27134 1202 27186 1214
rect 26114 1150 26126 1202
rect 26178 1150 26190 1202
rect 24782 1138 24834 1150
rect 27134 1138 27186 1150
rect 6862 1090 6914 1102
rect 6862 1026 6914 1038
rect 25678 1090 25730 1102
rect 25678 1026 25730 1038
rect 4958 978 5010 990
rect 4958 914 5010 926
rect 6302 978 6354 990
rect 6302 914 6354 926
rect 25342 978 25394 990
rect 25342 914 25394 926
rect 672 810 27888 844
rect 672 758 4466 810
rect 4518 758 4570 810
rect 4622 758 4674 810
rect 4726 758 24466 810
rect 24518 758 24570 810
rect 24622 758 24674 810
rect 24726 758 27888 810
rect 672 724 27888 758
<< via1 >>
rect 3806 56422 3858 56474
rect 3910 56422 3962 56474
rect 4014 56422 4066 56474
rect 23806 56422 23858 56474
rect 23910 56422 23962 56474
rect 24014 56422 24066 56474
rect 3614 56254 3666 56306
rect 5518 56254 5570 56306
rect 8990 56254 9042 56306
rect 10558 56254 10610 56306
rect 13022 56254 13074 56306
rect 14590 56254 14642 56306
rect 16494 56254 16546 56306
rect 18510 56254 18562 56306
rect 20638 56254 20690 56306
rect 21870 56254 21922 56306
rect 24446 56254 24498 56306
rect 26014 56254 26066 56306
rect 7422 56142 7474 56194
rect 5182 56030 5234 56082
rect 20190 56030 20242 56082
rect 25678 56030 25730 56082
rect 1038 55918 1090 55970
rect 3054 55918 3106 55970
rect 8094 55918 8146 55970
rect 9998 55918 10050 55970
rect 11566 55918 11618 55970
rect 14030 55918 14082 55970
rect 15598 55918 15650 55970
rect 17502 55918 17554 55970
rect 19518 55918 19570 55970
rect 22878 55918 22930 55970
rect 23886 55918 23938 55970
rect 1374 55806 1426 55858
rect 4466 55638 4518 55690
rect 4570 55638 4622 55690
rect 4674 55638 4726 55690
rect 24466 55638 24518 55690
rect 24570 55638 24622 55690
rect 24674 55638 24726 55690
rect 18846 55358 18898 55410
rect 21646 55358 21698 55410
rect 3502 55246 3554 55298
rect 7534 55246 7586 55298
rect 12910 55246 12962 55298
rect 18286 55246 18338 55298
rect 19406 55246 19458 55298
rect 20078 55246 20130 55298
rect 20526 55246 20578 55298
rect 20974 55246 21026 55298
rect 23662 55246 23714 55298
rect 24894 55246 24946 55298
rect 26238 55246 26290 55298
rect 2494 55134 2546 55186
rect 6526 55134 6578 55186
rect 11902 55134 11954 55186
rect 17278 55134 17330 55186
rect 22654 55134 22706 55186
rect 25566 55134 25618 55186
rect 27246 55022 27298 55074
rect 3806 54854 3858 54906
rect 3910 54854 3962 54906
rect 4014 54854 4066 54906
rect 23806 54854 23858 54906
rect 23910 54854 23962 54906
rect 24014 54854 24066 54906
rect 22542 54686 22594 54738
rect 24110 54686 24162 54738
rect 19518 54574 19570 54626
rect 21086 54574 21138 54626
rect 25454 54574 25506 54626
rect 21534 54350 21586 54402
rect 23102 54350 23154 54402
rect 24670 54350 24722 54402
rect 26238 54350 26290 54402
rect 27022 54350 27074 54402
rect 18958 54238 19010 54290
rect 20638 54238 20690 54290
rect 4466 54070 4518 54122
rect 4570 54070 4622 54122
rect 4674 54070 4726 54122
rect 24466 54070 24518 54122
rect 24570 54070 24622 54122
rect 24674 54070 24726 54122
rect 1038 53678 1090 53730
rect 20526 53678 20578 53730
rect 20862 53678 20914 53730
rect 21870 53678 21922 53730
rect 22878 53678 22930 53730
rect 24670 53678 24722 53730
rect 26238 53678 26290 53730
rect 1486 53566 1538 53618
rect 19966 53566 20018 53618
rect 21310 53566 21362 53618
rect 22206 53566 22258 53618
rect 23774 53566 23826 53618
rect 25566 53566 25618 53618
rect 27246 53454 27298 53506
rect 3806 53286 3858 53338
rect 3910 53286 3962 53338
rect 4014 53286 4066 53338
rect 23806 53286 23858 53338
rect 23910 53286 23962 53338
rect 24014 53286 24066 53338
rect 24110 53118 24162 53170
rect 21758 53006 21810 53058
rect 22654 53006 22706 53058
rect 27134 53006 27186 53058
rect 1598 52782 1650 52834
rect 21310 52782 21362 52834
rect 23102 52782 23154 52834
rect 24670 52782 24722 52834
rect 25454 52782 25506 52834
rect 26238 52782 26290 52834
rect 1038 52670 1090 52722
rect 22206 52670 22258 52722
rect 4466 52502 4518 52554
rect 4570 52502 4622 52554
rect 4674 52502 4726 52554
rect 24466 52502 24518 52554
rect 24570 52502 24622 52554
rect 24674 52502 24726 52554
rect 21870 52222 21922 52274
rect 22766 52222 22818 52274
rect 23550 52222 23602 52274
rect 24670 52222 24722 52274
rect 22430 52110 22482 52162
rect 26238 52110 26290 52162
rect 25566 51998 25618 52050
rect 27246 51886 27298 51938
rect 3806 51718 3858 51770
rect 3910 51718 3962 51770
rect 4014 51718 4066 51770
rect 23806 51718 23858 51770
rect 23910 51718 23962 51770
rect 24014 51718 24066 51770
rect 1486 51438 1538 51490
rect 23214 51438 23266 51490
rect 24334 51438 24386 51490
rect 25342 51438 25394 51490
rect 24894 51326 24946 51378
rect 26238 51214 26290 51266
rect 27022 51214 27074 51266
rect 1038 51102 1090 51154
rect 22766 51102 22818 51154
rect 23774 51102 23826 51154
rect 4466 50934 4518 50986
rect 4570 50934 4622 50986
rect 4674 50934 4726 50986
rect 24466 50934 24518 50986
rect 24570 50934 24622 50986
rect 24674 50934 24726 50986
rect 23438 50654 23490 50706
rect 26238 50654 26290 50706
rect 23886 50542 23938 50594
rect 24670 50542 24722 50594
rect 25566 50430 25618 50482
rect 27246 50318 27298 50370
rect 3806 50150 3858 50202
rect 3910 50150 3962 50202
rect 4014 50150 4066 50202
rect 23806 50150 23858 50202
rect 23910 50150 23962 50202
rect 24014 50150 24066 50202
rect 24222 49870 24274 49922
rect 27134 49870 27186 49922
rect 24894 49758 24946 49810
rect 26350 49758 26402 49810
rect 1598 49646 1650 49698
rect 25454 49646 25506 49698
rect 1038 49534 1090 49586
rect 23774 49534 23826 49586
rect 4466 49366 4518 49418
rect 4570 49366 4622 49418
rect 4674 49366 4726 49418
rect 24466 49366 24518 49418
rect 24570 49366 24622 49418
rect 24674 49366 24726 49418
rect 1038 48974 1090 49026
rect 24670 48974 24722 49026
rect 26238 48974 26290 49026
rect 1598 48862 1650 48914
rect 25566 48862 25618 48914
rect 27246 48750 27298 48802
rect 3806 48582 3858 48634
rect 3910 48582 3962 48634
rect 4014 48582 4066 48634
rect 23806 48582 23858 48634
rect 23910 48582 23962 48634
rect 24014 48582 24066 48634
rect 25790 48302 25842 48354
rect 25006 48078 25058 48130
rect 26238 48078 26290 48130
rect 27022 48078 27074 48130
rect 24446 47966 24498 48018
rect 25342 47966 25394 48018
rect 4466 47798 4518 47850
rect 4570 47798 4622 47850
rect 4674 47798 4726 47850
rect 24466 47798 24518 47850
rect 24570 47798 24622 47850
rect 24674 47798 24726 47850
rect 1038 47406 1090 47458
rect 24670 47406 24722 47458
rect 26238 47406 26290 47458
rect 1598 47294 1650 47346
rect 25678 47294 25730 47346
rect 27246 47182 27298 47234
rect 3806 47014 3858 47066
rect 3910 47014 3962 47066
rect 4014 47014 4066 47066
rect 23806 47014 23858 47066
rect 23910 47014 23962 47066
rect 24014 47014 24066 47066
rect 25678 46734 25730 46786
rect 27134 46734 27186 46786
rect 24670 46510 24722 46562
rect 26238 46510 26290 46562
rect 4466 46230 4518 46282
rect 4570 46230 4622 46282
rect 4674 46230 4726 46282
rect 24466 46230 24518 46282
rect 24570 46230 24622 46282
rect 24674 46230 24726 46282
rect 1038 45838 1090 45890
rect 24782 45838 24834 45890
rect 26462 45838 26514 45890
rect 1486 45726 1538 45778
rect 25678 45614 25730 45666
rect 27246 45614 27298 45666
rect 3806 45446 3858 45498
rect 3910 45446 3962 45498
rect 4014 45446 4066 45498
rect 23806 45446 23858 45498
rect 23910 45446 23962 45498
rect 24014 45446 24066 45498
rect 26350 45054 26402 45106
rect 27022 44942 27074 44994
rect 4466 44662 4518 44714
rect 4570 44662 4622 44714
rect 4674 44662 4726 44714
rect 24466 44662 24518 44714
rect 24570 44662 24622 44714
rect 24674 44662 24726 44714
rect 1038 44270 1090 44322
rect 24670 44270 24722 44322
rect 26238 44270 26290 44322
rect 1486 44158 1538 44210
rect 25678 44158 25730 44210
rect 27246 44046 27298 44098
rect 3806 43878 3858 43930
rect 3910 43878 3962 43930
rect 4014 43878 4066 43930
rect 23806 43878 23858 43930
rect 23910 43878 23962 43930
rect 24014 43878 24066 43930
rect 25678 43598 25730 43650
rect 27134 43598 27186 43650
rect 24894 43486 24946 43538
rect 1598 43374 1650 43426
rect 26238 43374 26290 43426
rect 1038 43262 1090 43314
rect 4466 43094 4518 43146
rect 4570 43094 4622 43146
rect 4674 43094 4726 43146
rect 24466 43094 24518 43146
rect 24570 43094 24622 43146
rect 24674 43094 24726 43146
rect 1150 42702 1202 42754
rect 24670 42702 24722 42754
rect 26238 42702 26290 42754
rect 1598 42590 1650 42642
rect 25678 42478 25730 42530
rect 27246 42478 27298 42530
rect 3806 42310 3858 42362
rect 3910 42310 3962 42362
rect 4014 42310 4066 42362
rect 23806 42310 23858 42362
rect 23910 42310 23962 42362
rect 24014 42310 24066 42362
rect 3614 41918 3666 41970
rect 16270 41918 16322 41970
rect 1598 41806 1650 41858
rect 4174 41806 4226 41858
rect 18398 41806 18450 41858
rect 26238 41806 26290 41858
rect 27022 41806 27074 41858
rect 1038 41694 1090 41746
rect 4466 41526 4518 41578
rect 4570 41526 4622 41578
rect 4674 41526 4726 41578
rect 24466 41526 24518 41578
rect 24570 41526 24622 41578
rect 24674 41526 24726 41578
rect 6078 41358 6130 41410
rect 2046 41246 2098 41298
rect 2606 41246 2658 41298
rect 4286 41246 4338 41298
rect 6638 41246 6690 41298
rect 10558 41246 10610 41298
rect 1038 41134 1090 41186
rect 3838 41134 3890 41186
rect 8878 41134 8930 41186
rect 10110 41134 10162 41186
rect 24670 41134 24722 41186
rect 26238 41134 26290 41186
rect 1486 41022 1538 41074
rect 9326 41022 9378 41074
rect 25678 41022 25730 41074
rect 5518 40910 5570 40962
rect 11790 40910 11842 40962
rect 27246 40910 27298 40962
rect 3806 40742 3858 40794
rect 3910 40742 3962 40794
rect 4014 40742 4066 40794
rect 23806 40742 23858 40794
rect 23910 40742 23962 40794
rect 24014 40742 24066 40794
rect 2158 40462 2210 40514
rect 6974 40462 7026 40514
rect 13358 40462 13410 40514
rect 15486 40462 15538 40514
rect 25678 40462 25730 40514
rect 27134 40462 27186 40514
rect 1710 40350 1762 40402
rect 2606 40350 2658 40402
rect 4286 40350 4338 40402
rect 7646 40350 7698 40402
rect 8094 40350 8146 40402
rect 8766 40350 8818 40402
rect 9550 40350 9602 40402
rect 10446 40350 10498 40402
rect 17726 40350 17778 40402
rect 18398 40350 18450 40402
rect 24670 40350 24722 40402
rect 26462 40350 26514 40402
rect 3054 40238 3106 40290
rect 7310 40238 7362 40290
rect 8318 40238 8370 40290
rect 6414 40126 6466 40178
rect 12910 40126 12962 40178
rect 4466 39958 4518 40010
rect 4570 39958 4622 40010
rect 4674 39958 4726 40010
rect 24466 39958 24518 40010
rect 24570 39958 24622 40010
rect 24674 39958 24726 40010
rect 6078 39790 6130 39842
rect 9886 39790 9938 39842
rect 12462 39790 12514 39842
rect 2494 39678 2546 39730
rect 5070 39678 5122 39730
rect 12910 39678 12962 39730
rect 1150 39566 1202 39618
rect 2046 39566 2098 39618
rect 5518 39566 5570 39618
rect 5854 39566 5906 39618
rect 6750 39566 6802 39618
rect 7086 39566 7138 39618
rect 7310 39566 7362 39618
rect 8206 39566 8258 39618
rect 9438 39566 9490 39618
rect 11006 39566 11058 39618
rect 11790 39566 11842 39618
rect 12350 39566 12402 39618
rect 13582 39566 13634 39618
rect 14590 39566 14642 39618
rect 16718 39566 16770 39618
rect 24894 39566 24946 39618
rect 26238 39566 26290 39618
rect 1486 39454 1538 39506
rect 11454 39454 11506 39506
rect 18734 39454 18786 39506
rect 25678 39342 25730 39394
rect 27246 39342 27298 39394
rect 3806 39174 3858 39226
rect 3910 39174 3962 39226
rect 4014 39174 4066 39226
rect 23806 39174 23858 39226
rect 23910 39174 23962 39226
rect 24014 39174 24066 39226
rect 7198 39006 7250 39058
rect 13358 38894 13410 38946
rect 2718 38782 2770 38834
rect 5518 38782 5570 38834
rect 10558 38782 10610 38834
rect 12910 38782 12962 38834
rect 15262 38782 15314 38834
rect 1598 38670 1650 38722
rect 3054 38670 3106 38722
rect 4286 38670 4338 38722
rect 5966 38670 6018 38722
rect 18622 38670 18674 38722
rect 26238 38670 26290 38722
rect 27022 38670 27074 38722
rect 1038 38558 1090 38610
rect 11006 38558 11058 38610
rect 12126 38558 12178 38610
rect 4466 38390 4518 38442
rect 4570 38390 4622 38442
rect 4674 38390 4726 38442
rect 24466 38390 24518 38442
rect 24570 38390 24622 38442
rect 24674 38390 24726 38442
rect 6302 38222 6354 38274
rect 12574 38222 12626 38274
rect 15150 38222 15202 38274
rect 2270 38110 2322 38162
rect 3838 38110 3890 38162
rect 5070 38110 5122 38162
rect 7758 38110 7810 38162
rect 9998 38110 10050 38162
rect 3390 37998 3442 38050
rect 4622 37998 4674 38050
rect 6750 37998 6802 38050
rect 8318 37998 8370 38050
rect 9438 37998 9490 38050
rect 11118 37998 11170 38050
rect 11902 37998 11954 38050
rect 12462 37998 12514 38050
rect 13134 37998 13186 38050
rect 13582 37998 13634 38050
rect 14702 37998 14754 38050
rect 15486 37998 15538 38050
rect 16718 37998 16770 38050
rect 17502 37998 17554 38050
rect 24670 37998 24722 38050
rect 26238 37998 26290 38050
rect 2718 37886 2770 37938
rect 7198 37886 7250 37938
rect 11566 37886 11618 37938
rect 19742 37886 19794 37938
rect 25678 37886 25730 37938
rect 1150 37774 1202 37826
rect 27246 37774 27298 37826
rect 3806 37606 3858 37658
rect 3910 37606 3962 37658
rect 4014 37606 4066 37658
rect 23806 37606 23858 37658
rect 23910 37606 23962 37658
rect 24014 37606 24066 37658
rect 6750 37438 6802 37490
rect 2494 37326 2546 37378
rect 3278 37326 3330 37378
rect 16270 37326 16322 37378
rect 27134 37326 27186 37378
rect 1150 37214 1202 37266
rect 5182 37214 5234 37266
rect 7870 37214 7922 37266
rect 8318 37214 8370 37266
rect 8990 37214 9042 37266
rect 9550 37214 9602 37266
rect 10670 37214 10722 37266
rect 18622 37214 18674 37266
rect 24894 37214 24946 37266
rect 1598 37102 1650 37154
rect 5518 37102 5570 37154
rect 7534 37102 7586 37154
rect 8542 37102 8594 37154
rect 16606 37102 16658 37154
rect 25454 37102 25506 37154
rect 26238 37102 26290 37154
rect 1934 36990 1986 37042
rect 2830 36990 2882 37042
rect 4466 36822 4518 36874
rect 4570 36822 4622 36874
rect 4674 36822 4726 36874
rect 24466 36822 24518 36874
rect 24570 36822 24622 36874
rect 24674 36822 24726 36874
rect 1710 36654 1762 36706
rect 3950 36654 4002 36706
rect 10110 36542 10162 36594
rect 12238 36542 12290 36594
rect 15710 36542 15762 36594
rect 18846 36542 18898 36594
rect 1262 36430 1314 36482
rect 6190 36430 6242 36482
rect 8318 36430 8370 36482
rect 14366 36430 14418 36482
rect 14814 36430 14866 36482
rect 15934 36430 15986 36482
rect 17838 36430 17890 36482
rect 18286 36430 18338 36482
rect 24670 36430 24722 36482
rect 26350 36430 26402 36482
rect 3502 36318 3554 36370
rect 6638 36318 6690 36370
rect 7758 36318 7810 36370
rect 10558 36318 10610 36370
rect 11790 36318 11842 36370
rect 13918 36318 13970 36370
rect 17054 36318 17106 36370
rect 2830 36206 2882 36258
rect 5070 36206 5122 36258
rect 8990 36206 9042 36258
rect 13358 36206 13410 36258
rect 15150 36206 15202 36258
rect 25678 36206 25730 36258
rect 27246 36206 27298 36258
rect 3806 36038 3858 36090
rect 3910 36038 3962 36090
rect 4014 36038 4066 36090
rect 23806 36038 23858 36090
rect 23910 36038 23962 36090
rect 24014 36038 24066 36090
rect 5854 35758 5906 35810
rect 11454 35758 11506 35810
rect 12910 35758 12962 35810
rect 15486 35758 15538 35810
rect 2606 35646 2658 35698
rect 8206 35646 8258 35698
rect 8654 35646 8706 35698
rect 9326 35646 9378 35698
rect 9886 35646 9938 35698
rect 10894 35646 10946 35698
rect 11902 35646 11954 35698
rect 18398 35646 18450 35698
rect 26350 35646 26402 35698
rect 1598 35534 1650 35586
rect 7870 35534 7922 35586
rect 8878 35534 8930 35586
rect 13358 35534 13410 35586
rect 27022 35534 27074 35586
rect 1038 35422 1090 35474
rect 3166 35422 3218 35474
rect 4286 35422 4338 35474
rect 6302 35422 6354 35474
rect 7422 35422 7474 35474
rect 4466 35254 4518 35306
rect 4570 35254 4622 35306
rect 4674 35254 4726 35306
rect 24466 35254 24518 35306
rect 24570 35254 24622 35306
rect 24674 35254 24726 35306
rect 6078 35086 6130 35138
rect 11006 35086 11058 35138
rect 13582 35086 13634 35138
rect 16830 35086 16882 35138
rect 17950 35086 18002 35138
rect 19854 35086 19906 35138
rect 1598 34974 1650 35026
rect 3166 34974 3218 35026
rect 14030 34974 14082 35026
rect 18062 34974 18114 35026
rect 20414 34974 20466 35026
rect 1038 34862 1090 34914
rect 2606 34862 2658 34914
rect 4286 34862 4338 34914
rect 5406 34862 5458 34914
rect 5854 34862 5906 34914
rect 6750 34862 6802 34914
rect 7198 34862 7250 34914
rect 8206 34862 8258 34914
rect 12910 34862 12962 34914
rect 13358 34862 13410 34914
rect 14702 34862 14754 34914
rect 15598 34862 15650 34914
rect 18958 34862 19010 34914
rect 24782 34862 24834 34914
rect 26238 34862 26290 34914
rect 5070 34750 5122 34802
rect 10558 34750 10610 34802
rect 12574 34750 12626 34802
rect 18398 34750 18450 34802
rect 19518 34750 19570 34802
rect 25678 34750 25730 34802
rect 12126 34638 12178 34690
rect 27246 34638 27298 34690
rect 3806 34470 3858 34522
rect 3910 34470 3962 34522
rect 4014 34470 4066 34522
rect 23806 34470 23858 34522
rect 23910 34470 23962 34522
rect 24014 34470 24066 34522
rect 6750 34302 6802 34354
rect 9102 34190 9154 34242
rect 16718 34190 16770 34242
rect 25678 34190 25730 34242
rect 27134 34190 27186 34242
rect 1486 34078 1538 34130
rect 1934 34078 1986 34130
rect 2830 34078 2882 34130
rect 3166 34078 3218 34130
rect 4174 34078 4226 34130
rect 5182 34078 5234 34130
rect 18510 34078 18562 34130
rect 1150 33966 1202 34018
rect 8654 33966 8706 34018
rect 24670 33966 24722 34018
rect 26238 33966 26290 34018
rect 2158 33854 2210 33906
rect 5630 33854 5682 33906
rect 7534 33854 7586 33906
rect 4466 33686 4518 33738
rect 4570 33686 4622 33738
rect 4674 33686 4726 33738
rect 24466 33686 24518 33738
rect 24570 33686 24622 33738
rect 24674 33686 24726 33738
rect 3278 33518 3330 33570
rect 6078 33518 6130 33570
rect 1598 33406 1650 33458
rect 3838 33406 3890 33458
rect 8206 33406 8258 33458
rect 9886 33406 9938 33458
rect 12238 33406 12290 33458
rect 14590 33406 14642 33458
rect 15150 33406 15202 33458
rect 16830 33406 16882 33458
rect 18286 33406 18338 33458
rect 7646 33294 7698 33346
rect 9550 33294 9602 33346
rect 11790 33294 11842 33346
rect 17390 33294 17442 33346
rect 24894 33294 24946 33346
rect 26238 33294 26290 33346
rect 1262 33182 1314 33234
rect 5630 33182 5682 33234
rect 17950 33182 18002 33234
rect 2830 33070 2882 33122
rect 7198 33070 7250 33122
rect 11118 33070 11170 33122
rect 13470 33070 13522 33122
rect 19518 33070 19570 33122
rect 25678 33070 25730 33122
rect 27246 33070 27298 33122
rect 3806 32902 3858 32954
rect 3910 32902 3962 32954
rect 4014 32902 4066 32954
rect 23806 32902 23858 32954
rect 23910 32902 23962 32954
rect 24014 32902 24066 32954
rect 18286 32734 18338 32786
rect 1710 32622 1762 32674
rect 13358 32622 13410 32674
rect 14366 32622 14418 32674
rect 17390 32622 17442 32674
rect 6750 32510 6802 32562
rect 7086 32510 7138 32562
rect 7758 32510 7810 32562
rect 8430 32510 8482 32562
rect 9214 32505 9266 32557
rect 10558 32510 10610 32562
rect 13022 32510 13074 32562
rect 15150 32510 15202 32562
rect 18622 32510 18674 32562
rect 19406 32510 19458 32562
rect 2158 32398 2210 32450
rect 4286 32398 4338 32450
rect 6302 32398 6354 32450
rect 7310 32398 7362 32450
rect 15598 32398 15650 32450
rect 19182 32398 19234 32450
rect 26238 32398 26290 32450
rect 27022 32398 27074 32450
rect 3278 32286 3330 32338
rect 3726 32286 3778 32338
rect 11006 32286 11058 32338
rect 12126 32286 12178 32338
rect 13806 32286 13858 32338
rect 16830 32286 16882 32338
rect 17838 32286 17890 32338
rect 4466 32118 4518 32170
rect 4570 32118 4622 32170
rect 4674 32118 4726 32170
rect 24466 32118 24518 32170
rect 24570 32118 24622 32170
rect 24674 32118 24726 32170
rect 13022 31950 13074 32002
rect 17726 31950 17778 32002
rect 2830 31838 2882 31890
rect 3278 31838 3330 31890
rect 9438 31838 9490 31890
rect 13470 31838 13522 31890
rect 18174 31838 18226 31890
rect 2270 31726 2322 31778
rect 2718 31726 2770 31778
rect 4062 31726 4114 31778
rect 4846 31726 4898 31778
rect 7310 31726 7362 31778
rect 8878 31726 8930 31778
rect 12350 31726 12402 31778
rect 12910 31726 12962 31778
rect 14030 31726 14082 31778
rect 15038 31726 15090 31778
rect 16718 31726 16770 31778
rect 17054 31726 17106 31778
rect 17502 31726 17554 31778
rect 18958 31726 19010 31778
rect 19854 31726 19906 31778
rect 24782 31726 24834 31778
rect 26350 31726 26402 31778
rect 1822 31614 1874 31666
rect 12014 31614 12066 31666
rect 25678 31614 25730 31666
rect 7646 31502 7698 31554
rect 27246 31502 27298 31554
rect 3806 31334 3858 31386
rect 3910 31334 3962 31386
rect 4014 31334 4066 31386
rect 23806 31334 23858 31386
rect 23910 31334 23962 31386
rect 24014 31334 24066 31386
rect 15822 31166 15874 31218
rect 4398 31054 4450 31106
rect 6638 31054 6690 31106
rect 7198 31054 7250 31106
rect 10782 31054 10834 31106
rect 11902 31054 11954 31106
rect 1262 30942 1314 30994
rect 2382 30942 2434 30994
rect 3502 30942 3554 30994
rect 3950 30942 4002 30994
rect 8094 30942 8146 30994
rect 10446 30942 10498 30994
rect 11342 30942 11394 30994
rect 14254 30942 14306 30994
rect 17166 30942 17218 30994
rect 17502 30942 17554 30994
rect 18398 30942 18450 30994
rect 18734 30942 18786 30994
rect 19854 30942 19906 30994
rect 24894 30942 24946 30994
rect 26462 30942 26514 30994
rect 2942 30830 2994 30882
rect 8654 30830 8706 30882
rect 14590 30830 14642 30882
rect 16718 30830 16770 30882
rect 17726 30830 17778 30882
rect 25454 30830 25506 30882
rect 27022 30830 27074 30882
rect 3390 30718 3442 30770
rect 6190 30718 6242 30770
rect 7646 30718 7698 30770
rect 9774 30718 9826 30770
rect 4466 30550 4518 30602
rect 4570 30550 4622 30602
rect 4674 30550 4726 30602
rect 24466 30550 24518 30602
rect 24570 30550 24622 30602
rect 24674 30550 24726 30602
rect 3166 30382 3218 30434
rect 3502 30382 3554 30434
rect 6078 30382 6130 30434
rect 10446 30382 10498 30434
rect 4062 30270 4114 30322
rect 17390 30270 17442 30322
rect 2270 30158 2322 30210
rect 5406 30158 5458 30210
rect 5854 30158 5906 30210
rect 6750 30158 6802 30210
rect 7086 30158 7138 30210
rect 8206 30158 8258 30210
rect 9438 30158 9490 30210
rect 9774 30158 9826 30210
rect 10222 30158 10274 30210
rect 11006 30158 11058 30210
rect 11454 30158 11506 30210
rect 12462 30158 12514 30210
rect 14142 30158 14194 30210
rect 15710 30158 15762 30210
rect 16830 30158 16882 30210
rect 18510 30158 18562 30210
rect 26462 30158 26514 30210
rect 1262 30046 1314 30098
rect 2718 30046 2770 30098
rect 5070 30046 5122 30098
rect 14702 30046 14754 30098
rect 16046 30046 16098 30098
rect 27134 30046 27186 30098
rect 3806 29766 3858 29818
rect 3910 29766 3962 29818
rect 4014 29766 4066 29818
rect 23806 29766 23858 29818
rect 23910 29766 23962 29818
rect 24014 29766 24066 29818
rect 2830 29598 2882 29650
rect 6750 29598 6802 29650
rect 17502 29598 17554 29650
rect 3726 29486 3778 29538
rect 5182 29486 5234 29538
rect 12126 29486 12178 29538
rect 27246 29486 27298 29538
rect 1150 29374 1202 29426
rect 3390 29374 3442 29426
rect 8542 29374 8594 29426
rect 11790 29374 11842 29426
rect 13582 29374 13634 29426
rect 15822 29374 15874 29426
rect 18062 29374 18114 29426
rect 1710 29262 1762 29314
rect 8878 29262 8930 29314
rect 16270 29262 16322 29314
rect 18510 29262 18562 29314
rect 26238 29262 26290 29314
rect 5630 29150 5682 29202
rect 10110 29150 10162 29202
rect 14142 29150 14194 29202
rect 15262 29150 15314 29202
rect 19742 29150 19794 29202
rect 4466 28982 4518 29034
rect 4570 28982 4622 29034
rect 4674 28982 4726 29034
rect 24466 28982 24518 29034
rect 24570 28982 24622 29034
rect 24674 28982 24726 29034
rect 2830 28814 2882 28866
rect 5070 28814 5122 28866
rect 11342 28814 11394 28866
rect 13918 28814 13970 28866
rect 1598 28702 1650 28754
rect 3838 28702 3890 28754
rect 6974 28702 7026 28754
rect 12910 28702 12962 28754
rect 18398 28702 18450 28754
rect 19406 28702 19458 28754
rect 19854 28702 19906 28754
rect 26238 28702 26290 28754
rect 1150 28590 1202 28642
rect 5518 28590 5570 28642
rect 5966 28590 6018 28642
rect 12462 28590 12514 28642
rect 13246 28590 13298 28642
rect 13694 28590 13746 28642
rect 14366 28590 14418 28642
rect 14926 28590 14978 28642
rect 16046 28590 16098 28642
rect 18846 28590 18898 28642
rect 19182 28590 19234 28642
rect 20414 28590 20466 28642
rect 21422 28590 21474 28642
rect 3502 28478 3554 28530
rect 6638 28478 6690 28530
rect 10894 28478 10946 28530
rect 27246 28478 27298 28530
rect 8206 28366 8258 28418
rect 3806 28198 3858 28250
rect 3910 28198 3962 28250
rect 4014 28198 4066 28250
rect 23806 28198 23858 28250
rect 23910 28198 23962 28250
rect 24014 28198 24066 28250
rect 19070 28030 19122 28082
rect 27246 28030 27298 28082
rect 1598 27918 1650 27970
rect 2718 27918 2770 27970
rect 8990 27918 9042 27970
rect 13582 27918 13634 27970
rect 17502 27918 17554 27970
rect 20078 27918 20130 27970
rect 25678 27918 25730 27970
rect 1038 27806 1090 27858
rect 4286 27806 4338 27858
rect 5294 27806 5346 27858
rect 5742 27806 5794 27858
rect 6526 27806 6578 27858
rect 7086 27806 7138 27858
rect 8094 27806 8146 27858
rect 9326 27806 9378 27858
rect 9774 27806 9826 27858
rect 10446 27806 10498 27858
rect 11006 27806 11058 27858
rect 12126 27806 12178 27858
rect 14030 27806 14082 27858
rect 14366 27806 14418 27858
rect 15262 27806 15314 27858
rect 15822 27806 15874 27858
rect 16606 27806 16658 27858
rect 19518 27806 19570 27858
rect 24670 27806 24722 27858
rect 26350 27806 26402 27858
rect 3166 27694 3218 27746
rect 4958 27694 5010 27746
rect 5966 27694 6018 27746
rect 17950 27694 18002 27746
rect 9998 27582 10050 27634
rect 14590 27582 14642 27634
rect 4466 27414 4518 27466
rect 4570 27414 4622 27466
rect 4674 27414 4726 27466
rect 24466 27414 24518 27466
rect 24570 27414 24622 27466
rect 24674 27414 24726 27466
rect 5406 27246 5458 27298
rect 6526 27246 6578 27298
rect 10222 27246 10274 27298
rect 12910 27246 12962 27298
rect 14030 27246 14082 27298
rect 15150 27246 15202 27298
rect 15598 27246 15650 27298
rect 1598 27134 1650 27186
rect 11678 27134 11730 27186
rect 16158 27134 16210 27186
rect 18286 27134 18338 27186
rect 24670 27134 24722 27186
rect 26238 27134 26290 27186
rect 1150 27022 1202 27074
rect 3390 27022 3442 27074
rect 4846 27022 4898 27074
rect 13470 27022 13522 27074
rect 17838 27022 17890 27074
rect 3726 26910 3778 26962
rect 10782 26910 10834 26962
rect 11342 26910 11394 26962
rect 27246 26910 27298 26962
rect 2830 26798 2882 26850
rect 19406 26798 19458 26850
rect 25678 26798 25730 26850
rect 3806 26630 3858 26682
rect 3910 26630 3962 26682
rect 4014 26630 4066 26682
rect 23806 26630 23858 26682
rect 23910 26630 23962 26682
rect 24014 26630 24066 26682
rect 27246 26462 27298 26514
rect 1710 26350 1762 26402
rect 4286 26350 4338 26402
rect 13358 26350 13410 26402
rect 14478 26350 14530 26402
rect 7646 26238 7698 26290
rect 16382 26238 16434 26290
rect 19182 26238 19234 26290
rect 7982 26126 8034 26178
rect 16942 26126 16994 26178
rect 19742 26126 19794 26178
rect 26238 26126 26290 26178
rect 2158 26014 2210 26066
rect 3278 26014 3330 26066
rect 3726 26014 3778 26066
rect 9214 26014 9266 26066
rect 12798 26014 12850 26066
rect 14030 26014 14082 26066
rect 18062 26014 18114 26066
rect 4466 25846 4518 25898
rect 4570 25846 4622 25898
rect 4674 25846 4726 25898
rect 24466 25846 24518 25898
rect 24570 25846 24622 25898
rect 24674 25846 24726 25898
rect 1038 25678 1090 25730
rect 3054 25678 3106 25730
rect 13134 25678 13186 25730
rect 2046 25566 2098 25618
rect 3502 25566 3554 25618
rect 6638 25566 6690 25618
rect 9438 25566 9490 25618
rect 10894 25566 10946 25618
rect 15262 25566 15314 25618
rect 18510 25566 18562 25618
rect 24670 25566 24722 25618
rect 2494 25454 2546 25506
rect 2942 25454 2994 25506
rect 4062 25454 4114 25506
rect 5070 25454 5122 25506
rect 6302 25454 6354 25506
rect 8878 25454 8930 25506
rect 12574 25454 12626 25506
rect 14702 25454 14754 25506
rect 17950 25454 18002 25506
rect 18286 25454 18338 25506
rect 19182 25454 19234 25506
rect 19742 25454 19794 25506
rect 20638 25454 20690 25506
rect 26238 25454 26290 25506
rect 1598 25342 1650 25394
rect 10446 25342 10498 25394
rect 17502 25342 17554 25394
rect 27246 25342 27298 25394
rect 7870 25230 7922 25282
rect 12014 25230 12066 25282
rect 14254 25230 14306 25282
rect 25678 25230 25730 25282
rect 3806 25062 3858 25114
rect 3910 25062 3962 25114
rect 4014 25062 4066 25114
rect 23806 25062 23858 25114
rect 23910 25062 23962 25114
rect 24014 25062 24066 25114
rect 6190 24782 6242 24834
rect 18174 24782 18226 24834
rect 19518 24782 19570 24834
rect 27134 24782 27186 24834
rect 1374 24670 1426 24722
rect 2382 24670 2434 24722
rect 2718 24670 2770 24722
rect 3502 24670 3554 24722
rect 4062 24670 4114 24722
rect 7870 24670 7922 24722
rect 8318 24670 8370 24722
rect 9214 24670 9266 24722
rect 9550 24670 9602 24722
rect 10670 24670 10722 24722
rect 13358 24670 13410 24722
rect 13694 24670 13746 24722
rect 14366 24670 14418 24722
rect 14926 24670 14978 24722
rect 15934 24670 15986 24722
rect 16606 24670 16658 24722
rect 18958 24670 19010 24722
rect 4398 24558 4450 24610
rect 7534 24558 7586 24610
rect 8542 24558 8594 24610
rect 12238 24558 12290 24610
rect 12910 24558 12962 24610
rect 13918 24558 13970 24610
rect 17726 24558 17778 24610
rect 24670 24558 24722 24610
rect 25454 24558 25506 24610
rect 26238 24558 26290 24610
rect 3390 24446 3442 24498
rect 5630 24446 5682 24498
rect 12014 24446 12066 24498
rect 12126 24446 12178 24498
rect 4466 24278 4518 24330
rect 4570 24278 4622 24330
rect 4674 24278 4726 24330
rect 24466 24278 24518 24330
rect 24570 24278 24622 24330
rect 24674 24278 24726 24330
rect 1038 24110 1090 24162
rect 2494 24110 2546 24162
rect 5630 24110 5682 24162
rect 11230 24110 11282 24162
rect 13806 24110 13858 24162
rect 17950 24110 18002 24162
rect 3614 23998 3666 24050
rect 6078 23998 6130 24050
rect 9326 23998 9378 24050
rect 19966 23998 20018 24050
rect 4062 23886 4114 23938
rect 5070 23886 5122 23938
rect 5406 23886 5458 23938
rect 6862 23886 6914 23938
rect 7646 23886 7698 23938
rect 9886 23886 9938 23938
rect 13134 23886 13186 23938
rect 13694 23886 13746 23938
rect 14254 23886 14306 23938
rect 15038 23886 15090 23938
rect 15934 23886 15986 23938
rect 18398 23886 18450 23938
rect 19518 23886 19570 23938
rect 24894 23886 24946 23938
rect 26238 23886 26290 23938
rect 1598 23774 1650 23826
rect 4622 23774 4674 23826
rect 10782 23774 10834 23826
rect 12350 23774 12402 23826
rect 12798 23774 12850 23826
rect 27246 23774 27298 23826
rect 16830 23662 16882 23714
rect 25678 23662 25730 23714
rect 3806 23494 3858 23546
rect 3910 23494 3962 23546
rect 4014 23494 4066 23546
rect 23806 23494 23858 23546
rect 23910 23494 23962 23546
rect 24014 23494 24066 23546
rect 3838 23326 3890 23378
rect 11678 23326 11730 23378
rect 1598 23214 1650 23266
rect 2270 23214 2322 23266
rect 16942 23214 16994 23266
rect 18958 23214 19010 23266
rect 27134 23214 27186 23266
rect 1262 23102 1314 23154
rect 5742 23102 5794 23154
rect 6190 23102 6242 23154
rect 6750 23102 6802 23154
rect 8990 23102 9042 23154
rect 11454 23102 11506 23154
rect 13134 23102 13186 23154
rect 13694 23102 13746 23154
rect 14366 23102 14418 23154
rect 14814 23102 14866 23154
rect 15934 23102 15986 23154
rect 26350 23102 26402 23154
rect 2606 22990 2658 23042
rect 9438 22990 9490 23042
rect 10558 22990 10610 23042
rect 12014 22990 12066 23042
rect 12238 22990 12290 23042
rect 12798 22990 12850 23042
rect 13806 22990 13858 23042
rect 7198 22878 7250 22930
rect 8318 22878 8370 22930
rect 11790 22878 11842 22930
rect 16382 22878 16434 22930
rect 17390 22878 17442 22930
rect 18510 22878 18562 22930
rect 4466 22710 4518 22762
rect 4570 22710 4622 22762
rect 4674 22710 4726 22762
rect 24466 22710 24518 22762
rect 24570 22710 24622 22762
rect 24674 22710 24726 22762
rect 1710 22542 1762 22594
rect 2718 22542 2770 22594
rect 5966 22542 6018 22594
rect 9886 22542 9938 22594
rect 15150 22542 15202 22594
rect 1150 22430 1202 22482
rect 10334 22430 10386 22482
rect 14702 22430 14754 22482
rect 18622 22430 18674 22482
rect 26238 22430 26290 22482
rect 2158 22318 2210 22370
rect 5294 22318 5346 22370
rect 5742 22318 5794 22370
rect 6526 22318 6578 22370
rect 6974 22318 7026 22370
rect 8094 22318 8146 22370
rect 9214 22318 9266 22370
rect 9774 22318 9826 22370
rect 10894 22318 10946 22370
rect 11902 22318 11954 22370
rect 13022 22318 13074 22370
rect 13918 22318 13970 22370
rect 15374 22318 15426 22370
rect 15822 22318 15874 22370
rect 16830 22318 16882 22370
rect 19070 22318 19122 22370
rect 24894 22318 24946 22370
rect 4958 22206 5010 22258
rect 8878 22206 8930 22258
rect 16158 22206 16210 22258
rect 27246 22206 27298 22258
rect 3838 22094 3890 22146
rect 16718 22094 16770 22146
rect 17390 22094 17442 22146
rect 25678 22094 25730 22146
rect 3806 21926 3858 21978
rect 3910 21926 3962 21978
rect 4014 21926 4066 21978
rect 23806 21926 23858 21978
rect 23910 21926 23962 21978
rect 24014 21926 24066 21978
rect 4286 21758 4338 21810
rect 11678 21758 11730 21810
rect 12798 21758 12850 21810
rect 13134 21758 13186 21810
rect 5518 21646 5570 21698
rect 6302 21646 6354 21698
rect 16718 21646 16770 21698
rect 18734 21646 18786 21698
rect 27134 21646 27186 21698
rect 1038 21534 1090 21586
rect 2606 21534 2658 21586
rect 6750 21534 6802 21586
rect 7086 21534 7138 21586
rect 7870 21534 7922 21586
rect 8318 21534 8370 21586
rect 9438 21534 9490 21586
rect 10110 21534 10162 21586
rect 13582 21534 13634 21586
rect 14478 21534 14530 21586
rect 15822 21534 15874 21586
rect 16382 21534 16434 21586
rect 1598 21422 1650 21474
rect 3166 21422 3218 21474
rect 10446 21422 10498 21474
rect 12238 21422 12290 21474
rect 15262 21422 15314 21474
rect 17166 21422 17218 21474
rect 18286 21422 18338 21474
rect 19294 21422 19346 21474
rect 25342 21422 25394 21474
rect 26238 21422 26290 21474
rect 5966 21310 6018 21362
rect 7310 21310 7362 21362
rect 12126 21310 12178 21362
rect 12910 21310 12962 21362
rect 15710 21310 15762 21362
rect 19854 21310 19906 21362
rect 25902 21310 25954 21362
rect 4466 21142 4518 21194
rect 4570 21142 4622 21194
rect 4674 21142 4726 21194
rect 24466 21142 24518 21194
rect 24570 21142 24622 21194
rect 24674 21142 24726 21194
rect 7870 20974 7922 21026
rect 9774 20974 9826 21026
rect 17614 20974 17666 21026
rect 18734 20974 18786 21026
rect 19854 20974 19906 21026
rect 27470 20974 27522 21026
rect 1374 20862 1426 20914
rect 1934 20862 1986 20914
rect 2270 20862 2322 20914
rect 3278 20862 3330 20914
rect 3726 20862 3778 20914
rect 6638 20862 6690 20914
rect 9886 20862 9938 20914
rect 13918 20862 13970 20914
rect 17054 20862 17106 20914
rect 20414 20862 20466 20914
rect 20750 20862 20802 20914
rect 26014 20862 26066 20914
rect 26910 20862 26962 20914
rect 2606 20750 2658 20802
rect 3054 20750 3106 20802
rect 4510 20750 4562 20802
rect 5294 20750 5346 20802
rect 6190 20750 6242 20802
rect 9438 20750 9490 20802
rect 9998 20750 10050 20802
rect 10446 20750 10498 20802
rect 11006 20750 11058 20802
rect 11566 20750 11618 20802
rect 11902 20750 11954 20802
rect 13358 20750 13410 20802
rect 13806 20750 13858 20802
rect 14590 20750 14642 20802
rect 14926 20750 14978 20802
rect 15934 20750 15986 20802
rect 16718 20750 16770 20802
rect 20190 20750 20242 20802
rect 26574 20750 26626 20802
rect 11790 20638 11842 20690
rect 12910 20638 12962 20690
rect 19182 20638 19234 20690
rect 10782 20526 10834 20578
rect 16718 20526 16770 20578
rect 3806 20358 3858 20410
rect 3910 20358 3962 20410
rect 4014 20358 4066 20410
rect 23806 20358 23858 20410
rect 23910 20358 23962 20410
rect 24014 20358 24066 20410
rect 12014 20190 12066 20242
rect 16046 20190 16098 20242
rect 2046 20078 2098 20130
rect 2830 20078 2882 20130
rect 6190 20078 6242 20130
rect 6750 20078 6802 20130
rect 10558 20078 10610 20130
rect 12910 20078 12962 20130
rect 15038 20078 15090 20130
rect 18174 20078 18226 20130
rect 19742 20078 19794 20130
rect 27022 20078 27074 20130
rect 1038 19966 1090 20018
rect 1262 19966 1314 20018
rect 3614 19966 3666 20018
rect 6638 19966 6690 20018
rect 8318 19966 8370 20018
rect 8990 19966 9042 20018
rect 11454 19966 11506 20018
rect 12238 19966 12290 20018
rect 13246 19966 13298 20018
rect 14702 19966 14754 20018
rect 15822 19966 15874 20018
rect 16046 19966 16098 20018
rect 27470 19966 27522 20018
rect 7198 19854 7250 19906
rect 9326 19854 9378 19906
rect 11678 19854 11730 19906
rect 13470 19854 13522 19906
rect 13806 19854 13858 19906
rect 14030 19854 14082 19906
rect 15486 19854 15538 19906
rect 15710 19854 15762 19906
rect 5630 19742 5682 19794
rect 11790 19742 11842 19794
rect 15598 19742 15650 19794
rect 18622 19742 18674 19794
rect 4466 19574 4518 19626
rect 4570 19574 4622 19626
rect 4674 19574 4726 19626
rect 24466 19574 24518 19626
rect 24570 19574 24622 19626
rect 24674 19574 24726 19626
rect 1598 19406 1650 19458
rect 2718 19406 2770 19458
rect 5742 19406 5794 19458
rect 8206 19406 8258 19458
rect 11566 19406 11618 19458
rect 27470 19406 27522 19458
rect 4510 19294 4562 19346
rect 7086 19294 7138 19346
rect 11118 19294 11170 19346
rect 12574 19294 12626 19346
rect 13918 19294 13970 19346
rect 14366 19294 14418 19346
rect 16718 19294 16770 19346
rect 16942 19294 16994 19346
rect 26014 19294 26066 19346
rect 9550 19182 9602 19234
rect 10334 19182 10386 19234
rect 11790 19182 11842 19234
rect 12238 19182 12290 19234
rect 13358 19182 13410 19234
rect 13694 19182 13746 19234
rect 15038 19182 15090 19234
rect 15934 19182 15986 19234
rect 26574 19182 26626 19234
rect 3166 19070 3218 19122
rect 4174 19070 4226 19122
rect 6638 19070 6690 19122
rect 12910 19070 12962 19122
rect 16830 19070 16882 19122
rect 27022 19070 27074 19122
rect 3806 18790 3858 18842
rect 3910 18790 3962 18842
rect 4014 18790 4066 18842
rect 23806 18790 23858 18842
rect 23910 18790 23962 18842
rect 24014 18790 24066 18842
rect 13806 18622 13858 18674
rect 15822 18622 15874 18674
rect 8094 18510 8146 18562
rect 10334 18510 10386 18562
rect 16046 18510 16098 18562
rect 17054 18510 17106 18562
rect 26126 18510 26178 18562
rect 2718 18398 2770 18450
rect 3166 18398 3218 18450
rect 4398 18398 4450 18450
rect 5630 18398 5682 18450
rect 7198 18398 7250 18450
rect 14590 18398 14642 18450
rect 15598 18398 15650 18450
rect 16494 18398 16546 18450
rect 19518 18398 19570 18450
rect 26910 18398 26962 18450
rect 27470 18398 27522 18450
rect 2270 18286 2322 18338
rect 8542 18286 8594 18338
rect 10670 18286 10722 18338
rect 11902 18286 11954 18338
rect 14478 18286 14530 18338
rect 15262 18286 15314 18338
rect 17390 18286 17442 18338
rect 1710 18174 1762 18226
rect 3838 18174 3890 18226
rect 6078 18174 6130 18226
rect 9662 18174 9714 18226
rect 13470 18174 13522 18226
rect 15150 18174 15202 18226
rect 16270 18174 16322 18226
rect 16382 18174 16434 18226
rect 16942 18174 16994 18226
rect 17166 18174 17218 18226
rect 18958 18174 19010 18226
rect 26574 18174 26626 18226
rect 4466 18006 4518 18058
rect 4570 18006 4622 18058
rect 4674 18006 4726 18058
rect 24466 18006 24518 18058
rect 24570 18006 24622 18058
rect 24674 18006 24726 18058
rect 1038 17838 1090 17890
rect 3726 17838 3778 17890
rect 4846 17838 4898 17890
rect 27470 17838 27522 17890
rect 1598 17726 1650 17778
rect 2606 17726 2658 17778
rect 6974 17726 7026 17778
rect 9998 17726 10050 17778
rect 14030 17726 14082 17778
rect 14478 17726 14530 17778
rect 16046 17726 16098 17778
rect 26014 17726 26066 17778
rect 26910 17726 26962 17778
rect 2158 17614 2210 17666
rect 4286 17614 4338 17666
rect 6638 17614 6690 17666
rect 12350 17614 12402 17666
rect 13246 17614 13298 17666
rect 14590 17602 14642 17654
rect 15038 17614 15090 17666
rect 26574 17614 26626 17666
rect 9662 17502 9714 17554
rect 11230 17502 11282 17554
rect 15486 17502 15538 17554
rect 16158 17502 16210 17554
rect 5966 17390 6018 17442
rect 8206 17390 8258 17442
rect 15822 17390 15874 17442
rect 3806 17222 3858 17274
rect 3910 17222 3962 17274
rect 4014 17222 4066 17274
rect 23806 17222 23858 17274
rect 23910 17222 23962 17274
rect 24014 17222 24066 17274
rect 8318 17054 8370 17106
rect 13134 17054 13186 17106
rect 14254 17054 14306 17106
rect 1486 16942 1538 16994
rect 2494 16942 2546 16994
rect 3278 16942 3330 16994
rect 5854 16942 5906 16994
rect 10222 16942 10274 16994
rect 12238 16942 12290 16994
rect 12910 16942 12962 16994
rect 27022 16942 27074 16994
rect 1150 16830 1202 16882
rect 1934 16830 1986 16882
rect 2830 16830 2882 16882
rect 3838 16830 3890 16882
rect 4286 16830 4338 16882
rect 4958 16830 5010 16882
rect 6638 16830 6690 16882
rect 10558 16830 10610 16882
rect 10894 16830 10946 16882
rect 11006 16830 11058 16882
rect 11790 16830 11842 16882
rect 13806 16830 13858 16882
rect 14030 16830 14082 16882
rect 14366 16830 14418 16882
rect 15262 16830 15314 16882
rect 15822 16830 15874 16882
rect 16494 16830 16546 16882
rect 16942 16830 16994 16882
rect 17950 16830 18002 16882
rect 27470 16830 27522 16882
rect 7086 16718 7138 16770
rect 9886 16718 9938 16770
rect 10110 16718 10162 16770
rect 11342 16718 11394 16770
rect 12910 16718 12962 16770
rect 14926 16718 14978 16770
rect 15934 16718 15986 16770
rect 11230 16606 11282 16658
rect 14590 16606 14642 16658
rect 4466 16438 4518 16490
rect 4570 16438 4622 16490
rect 4674 16438 4726 16490
rect 24466 16438 24518 16490
rect 24570 16438 24622 16490
rect 24674 16438 24726 16490
rect 11790 16270 11842 16322
rect 17950 16270 18002 16322
rect 27470 16270 27522 16322
rect 3166 16158 3218 16210
rect 4734 16158 4786 16210
rect 6862 16158 6914 16210
rect 9550 16158 9602 16210
rect 10110 16158 10162 16210
rect 10334 16158 10386 16210
rect 10782 16158 10834 16210
rect 12238 16158 12290 16210
rect 15262 16158 15314 16210
rect 15710 16158 15762 16210
rect 3502 16046 3554 16098
rect 4286 16046 4338 16098
rect 6526 16046 6578 16098
rect 9102 16046 9154 16098
rect 9326 16046 9378 16098
rect 9886 16046 9938 16098
rect 9998 16046 10050 16098
rect 11118 16046 11170 16098
rect 11678 16046 11730 16098
rect 12798 16046 12850 16098
rect 13022 16046 13074 16098
rect 13918 16046 13970 16098
rect 15934 16046 15986 16098
rect 16270 16046 16322 16098
rect 26574 16046 26626 16098
rect 8094 15934 8146 15986
rect 15374 15934 15426 15986
rect 18398 15934 18450 15986
rect 26014 15934 26066 15986
rect 27022 15934 27074 15986
rect 1934 15822 1986 15874
rect 5854 15822 5906 15874
rect 9662 15822 9714 15874
rect 16046 15822 16098 15874
rect 16830 15822 16882 15874
rect 3806 15654 3858 15706
rect 3910 15654 3962 15706
rect 4014 15654 4066 15706
rect 23806 15654 23858 15706
rect 23910 15654 23962 15706
rect 24014 15654 24066 15706
rect 7310 15486 7362 15538
rect 11230 15486 11282 15538
rect 11902 15486 11954 15538
rect 5742 15374 5794 15426
rect 9550 15374 9602 15426
rect 11006 15374 11058 15426
rect 15262 15374 15314 15426
rect 26126 15374 26178 15426
rect 27022 15374 27074 15426
rect 3614 15262 3666 15314
rect 7870 15262 7922 15314
rect 10558 15262 10610 15314
rect 11454 15262 11506 15314
rect 13582 15262 13634 15314
rect 15374 15262 15426 15314
rect 18622 15262 18674 15314
rect 27470 15262 27522 15314
rect 3054 15150 3106 15202
rect 6190 15150 6242 15202
rect 8318 15150 8370 15202
rect 10110 15150 10162 15202
rect 11790 15150 11842 15202
rect 11902 15150 11954 15202
rect 13358 15150 13410 15202
rect 14926 15150 14978 15202
rect 15150 15150 15202 15202
rect 15822 15150 15874 15202
rect 15934 15150 15986 15202
rect 16046 15150 16098 15202
rect 16942 15150 16994 15202
rect 18062 15150 18114 15202
rect 1934 15038 1986 15090
rect 9998 15038 10050 15090
rect 10670 15038 10722 15090
rect 10782 15038 10834 15090
rect 16494 15038 16546 15090
rect 26574 15038 26626 15090
rect 4466 14870 4518 14922
rect 4570 14870 4622 14922
rect 4674 14870 4726 14922
rect 24466 14870 24518 14922
rect 24570 14870 24622 14922
rect 24674 14870 24726 14922
rect 1038 14702 1090 14754
rect 2830 14702 2882 14754
rect 11118 14702 11170 14754
rect 11230 14702 11282 14754
rect 15486 14702 15538 14754
rect 16270 14702 16322 14754
rect 17614 14702 17666 14754
rect 27470 14702 27522 14754
rect 2494 14590 2546 14642
rect 5518 14590 5570 14642
rect 5966 14590 6018 14642
rect 9438 14590 9490 14642
rect 9550 14590 9602 14642
rect 10110 14590 10162 14642
rect 10222 14590 10274 14642
rect 14254 14590 14306 14642
rect 16046 14590 16098 14642
rect 1934 14478 1986 14530
rect 4846 14478 4898 14530
rect 5294 14478 5346 14530
rect 6526 14478 6578 14530
rect 7646 14478 7698 14530
rect 9998 14478 10050 14530
rect 10670 14478 10722 14530
rect 15934 14478 15986 14530
rect 16718 14478 16770 14530
rect 17166 14478 17218 14530
rect 17390 14478 17442 14530
rect 26574 14478 26626 14530
rect 1598 14366 1650 14418
rect 3278 14366 3330 14418
rect 4510 14366 4562 14418
rect 13918 14366 13970 14418
rect 17502 14366 17554 14418
rect 26126 14366 26178 14418
rect 26910 14366 26962 14418
rect 9438 14254 9490 14306
rect 11006 14254 11058 14306
rect 16942 14254 16994 14306
rect 3806 14086 3858 14138
rect 3910 14086 3962 14138
rect 4014 14086 4066 14138
rect 23806 14086 23858 14138
rect 23910 14086 23962 14138
rect 24014 14086 24066 14138
rect 7422 13918 7474 13970
rect 15374 13918 15426 13970
rect 17390 13918 17442 13970
rect 16382 13806 16434 13858
rect 1486 13694 1538 13746
rect 1934 13694 1986 13746
rect 2606 13694 2658 13746
rect 3390 13694 3442 13746
rect 4286 13694 4338 13746
rect 5182 13694 5234 13746
rect 8206 13694 8258 13746
rect 9326 13694 9378 13746
rect 13134 13694 13186 13746
rect 15710 13694 15762 13746
rect 16046 13694 16098 13746
rect 16158 13694 16210 13746
rect 16494 13694 16546 13746
rect 16830 13694 16882 13746
rect 17054 13694 17106 13746
rect 17278 13694 17330 13746
rect 27470 13694 27522 13746
rect 1150 13582 1202 13634
rect 5630 13582 5682 13634
rect 9774 13582 9826 13634
rect 13694 13582 13746 13634
rect 15262 13582 15314 13634
rect 26910 13582 26962 13634
rect 2158 13470 2210 13522
rect 6750 13470 6802 13522
rect 11006 13470 11058 13522
rect 14814 13470 14866 13522
rect 4466 13302 4518 13354
rect 4570 13302 4622 13354
rect 4674 13302 4726 13354
rect 24466 13302 24518 13354
rect 24570 13302 24622 13354
rect 24674 13302 24726 13354
rect 7758 13134 7810 13186
rect 15374 13134 15426 13186
rect 16046 13134 16098 13186
rect 27470 13134 27522 13186
rect 2606 13022 2658 13074
rect 5182 13022 5234 13074
rect 9438 13022 9490 13074
rect 12798 13022 12850 13074
rect 14478 13022 14530 13074
rect 14814 13022 14866 13074
rect 15262 13022 15314 13074
rect 26014 13022 26066 13074
rect 1038 12910 1090 12962
rect 2158 12910 2210 12962
rect 3726 12910 3778 12962
rect 4510 12910 4562 12962
rect 4958 12910 5010 12962
rect 5854 12910 5906 12962
rect 6414 12910 6466 12962
rect 7310 12910 7362 12962
rect 11342 12910 11394 12962
rect 12238 12910 12290 12962
rect 15486 12910 15538 12962
rect 16158 12910 16210 12962
rect 26574 12910 26626 12962
rect 1598 12798 1650 12850
rect 4174 12798 4226 12850
rect 8206 12798 8258 12850
rect 9102 12798 9154 12850
rect 11902 12798 11954 12850
rect 27022 12798 27074 12850
rect 10670 12686 10722 12738
rect 3806 12518 3858 12570
rect 3910 12518 3962 12570
rect 4014 12518 4066 12570
rect 23806 12518 23858 12570
rect 23910 12518 23962 12570
rect 24014 12518 24066 12570
rect 1038 12238 1090 12290
rect 3278 12238 3330 12290
rect 4286 12238 4338 12290
rect 5966 12238 6018 12290
rect 26014 12238 26066 12290
rect 26910 12238 26962 12290
rect 1486 12126 1538 12178
rect 1934 12126 1986 12178
rect 2942 12126 2994 12178
rect 3726 12126 3778 12178
rect 5518 12126 5570 12178
rect 6974 12126 7026 12178
rect 8542 12126 8594 12178
rect 9326 12126 9378 12178
rect 9774 12126 9826 12178
rect 10670 12126 10722 12178
rect 11230 12126 11282 12178
rect 12014 12126 12066 12178
rect 13134 12126 13186 12178
rect 13582 12126 13634 12178
rect 15038 12126 15090 12178
rect 15822 12126 15874 12178
rect 27470 12126 27522 12178
rect 2494 12014 2546 12066
rect 7310 12014 7362 12066
rect 8990 12014 9042 12066
rect 9998 12014 10050 12066
rect 12798 12014 12850 12066
rect 14254 12014 14306 12066
rect 13806 11902 13858 11954
rect 26574 11902 26626 11954
rect 4466 11734 4518 11786
rect 4570 11734 4622 11786
rect 4674 11734 4726 11786
rect 24466 11734 24518 11786
rect 24570 11734 24622 11786
rect 24674 11734 24726 11786
rect 2606 11566 2658 11618
rect 4846 11566 4898 11618
rect 7086 11566 7138 11618
rect 10894 11566 10946 11618
rect 27470 11566 27522 11618
rect 2270 11454 2322 11506
rect 9886 11454 9938 11506
rect 14702 11454 14754 11506
rect 15150 11454 15202 11506
rect 26014 11454 26066 11506
rect 6638 11342 6690 11394
rect 8206 11342 8258 11394
rect 10222 11342 10274 11394
rect 10782 11342 10834 11394
rect 11454 11342 11506 11394
rect 12014 11342 12066 11394
rect 12910 11342 12962 11394
rect 26574 11342 26626 11394
rect 3166 11230 3218 11282
rect 4398 11230 4450 11282
rect 26910 11230 26962 11282
rect 1262 11118 1314 11170
rect 5966 11118 6018 11170
rect 14142 11118 14194 11170
rect 14478 11118 14530 11170
rect 3806 10950 3858 11002
rect 3910 10950 3962 11002
rect 4014 10950 4066 11002
rect 23806 10950 23858 11002
rect 23910 10950 23962 11002
rect 24014 10950 24066 11002
rect 12126 10782 12178 10834
rect 1598 10670 1650 10722
rect 2382 10670 2434 10722
rect 3278 10670 3330 10722
rect 5854 10670 5906 10722
rect 6750 10670 6802 10722
rect 14030 10670 14082 10722
rect 14926 10670 14978 10722
rect 26910 10670 26962 10722
rect 1038 10558 1090 10610
rect 1934 10558 1986 10610
rect 2942 10558 2994 10610
rect 5294 10558 5346 10610
rect 7086 10558 7138 10610
rect 7646 10558 7698 10610
rect 8206 10558 8258 10610
rect 8766 10558 8818 10610
rect 9886 10558 9938 10610
rect 10446 10558 10498 10610
rect 13582 10558 13634 10610
rect 14366 10558 14418 10610
rect 27470 10558 27522 10610
rect 10894 10446 10946 10498
rect 7758 10334 7810 10386
rect 4466 10166 4518 10218
rect 4570 10166 4622 10218
rect 4674 10166 4726 10218
rect 24466 10166 24518 10218
rect 24570 10166 24622 10218
rect 24674 10166 24726 10218
rect 7534 9998 7586 10050
rect 27470 9998 27522 10050
rect 3166 9886 3218 9938
rect 4734 9886 4786 9938
rect 10110 9886 10162 9938
rect 11118 9886 11170 9938
rect 26014 9886 26066 9938
rect 26910 9886 26962 9938
rect 2046 9774 2098 9826
rect 2718 9774 2770 9826
rect 5182 9774 5234 9826
rect 10446 9774 10498 9826
rect 10894 9774 10946 9826
rect 11566 9774 11618 9826
rect 12350 9774 12402 9826
rect 13246 9774 13298 9826
rect 26574 9774 26626 9826
rect 7086 9662 7138 9714
rect 1262 9550 1314 9602
rect 3806 9382 3858 9434
rect 3910 9382 3962 9434
rect 4014 9382 4066 9434
rect 23806 9382 23858 9434
rect 23910 9382 23962 9434
rect 24014 9382 24066 9434
rect 8878 9214 8930 9266
rect 11118 9214 11170 9266
rect 1486 9102 1538 9154
rect 9550 9102 9602 9154
rect 26014 9102 26066 9154
rect 27022 9102 27074 9154
rect 1150 8990 1202 9042
rect 2046 8990 2098 9042
rect 7310 8990 7362 9042
rect 27470 8990 27522 9042
rect 2494 8878 2546 8930
rect 7646 8878 7698 8930
rect 9886 8878 9938 8930
rect 26574 8766 26626 8818
rect 4466 8598 4518 8650
rect 4570 8598 4622 8650
rect 4674 8598 4726 8650
rect 24466 8598 24518 8650
rect 24570 8598 24622 8650
rect 24674 8598 24726 8650
rect 1038 8430 1090 8482
rect 7758 8430 7810 8482
rect 11342 8430 11394 8482
rect 27470 8430 27522 8482
rect 10110 8318 10162 8370
rect 26014 8318 26066 8370
rect 1598 8206 1650 8258
rect 9662 8206 9714 8258
rect 26574 8206 26626 8258
rect 8318 8094 8370 8146
rect 26910 8094 26962 8146
rect 3806 7814 3858 7866
rect 3910 7814 3962 7866
rect 4014 7814 4066 7866
rect 23806 7814 23858 7866
rect 23910 7814 23962 7866
rect 24014 7814 24066 7866
rect 1486 7534 1538 7586
rect 10670 7534 10722 7586
rect 11566 7534 11618 7586
rect 1038 7422 1090 7474
rect 10110 7422 10162 7474
rect 11006 7422 11058 7474
rect 26910 7422 26962 7474
rect 27470 7422 27522 7474
rect 4466 7030 4518 7082
rect 4570 7030 4622 7082
rect 4674 7030 4726 7082
rect 24466 7030 24518 7082
rect 24570 7030 24622 7082
rect 24674 7030 24726 7082
rect 27470 6862 27522 6914
rect 2158 6638 2210 6690
rect 26574 6638 26626 6690
rect 26910 6638 26962 6690
rect 1262 6526 1314 6578
rect 26014 6526 26066 6578
rect 3806 6246 3858 6298
rect 3910 6246 3962 6298
rect 4014 6246 4066 6298
rect 23806 6246 23858 6298
rect 23910 6246 23962 6298
rect 24014 6246 24066 6298
rect 1262 5966 1314 6018
rect 26910 5966 26962 6018
rect 2270 5854 2322 5906
rect 27470 5854 27522 5906
rect 26014 5742 26066 5794
rect 26574 5630 26626 5682
rect 4466 5462 4518 5514
rect 4570 5462 4622 5514
rect 4674 5462 4726 5514
rect 24466 5462 24518 5514
rect 24570 5462 24622 5514
rect 24674 5462 24726 5514
rect 27470 5294 27522 5346
rect 26014 5182 26066 5234
rect 26910 5182 26962 5234
rect 26574 5070 26626 5122
rect 3806 4678 3858 4730
rect 3910 4678 3962 4730
rect 4014 4678 4066 4730
rect 23806 4678 23858 4730
rect 23910 4678 23962 4730
rect 24014 4678 24066 4730
rect 1486 4398 1538 4450
rect 27022 4398 27074 4450
rect 27470 4286 27522 4338
rect 1038 4062 1090 4114
rect 4466 3894 4518 3946
rect 4570 3894 4622 3946
rect 4674 3894 4726 3946
rect 24466 3894 24518 3946
rect 24570 3894 24622 3946
rect 24674 3894 24726 3946
rect 27470 3726 27522 3778
rect 26574 3502 26626 3554
rect 26014 3390 26066 3442
rect 26910 3390 26962 3442
rect 3806 3110 3858 3162
rect 3910 3110 3962 3162
rect 4014 3110 4066 3162
rect 23806 3110 23858 3162
rect 23910 3110 23962 3162
rect 24014 3110 24066 3162
rect 26014 2830 26066 2882
rect 26910 2830 26962 2882
rect 27470 2718 27522 2770
rect 26574 2494 26626 2546
rect 4466 2326 4518 2378
rect 4570 2326 4622 2378
rect 4674 2326 4726 2378
rect 24466 2326 24518 2378
rect 24570 2326 24622 2378
rect 24674 2326 24726 2378
rect 27470 2158 27522 2210
rect 26014 2046 26066 2098
rect 26574 1934 26626 1986
rect 27022 1822 27074 1874
rect 3806 1542 3858 1594
rect 3910 1542 3962 1594
rect 4014 1542 4066 1594
rect 23806 1542 23858 1594
rect 23910 1542 23962 1594
rect 24014 1542 24066 1594
rect 5518 1262 5570 1314
rect 26574 1262 26626 1314
rect 24782 1150 24834 1202
rect 26126 1150 26178 1202
rect 27134 1150 27186 1202
rect 6862 1038 6914 1090
rect 25678 1038 25730 1090
rect 4958 926 5010 978
rect 6302 926 6354 978
rect 25342 926 25394 978
rect 4466 758 4518 810
rect 4570 758 4622 810
rect 4674 758 4726 810
rect 24466 758 24518 810
rect 24570 758 24622 810
rect 24674 758 24726 810
<< metal2 >>
rect 672 57344 784 57456
rect 2016 57344 2128 57456
rect 3360 57344 3472 57456
rect 4704 57344 4816 57456
rect 6048 57344 6160 57456
rect 7392 57344 7504 57456
rect 8736 57344 8848 57456
rect 10080 57344 10192 57456
rect 11424 57344 11536 57456
rect 12768 57344 12880 57456
rect 14112 57344 14224 57456
rect 15456 57344 15568 57456
rect 16800 57344 16912 57456
rect 18144 57344 18256 57456
rect 19488 57344 19600 57456
rect 20832 57344 20944 57456
rect 22176 57344 22288 57456
rect 23520 57344 23632 57456
rect 24864 57344 24976 57456
rect 26208 57344 26320 57456
rect 27552 57344 27664 57456
rect 700 55972 756 57344
rect 1036 55972 1092 55982
rect 700 55970 1092 55972
rect 700 55918 1038 55970
rect 1090 55918 1092 55970
rect 700 55916 1092 55918
rect 1036 55906 1092 55916
rect 1372 55858 1428 55870
rect 1372 55806 1374 55858
rect 1426 55806 1428 55858
rect 1036 53730 1092 53742
rect 1036 53678 1038 53730
rect 1090 53678 1092 53730
rect 1036 53620 1092 53678
rect 1036 53554 1092 53564
rect 1372 52948 1428 55806
rect 2044 55468 2100 57344
rect 3388 56308 3444 57344
rect 4732 57316 4788 57344
rect 4732 57250 4788 57260
rect 5516 57316 5572 57326
rect 3804 56476 4068 56486
rect 3860 56420 3908 56476
rect 3964 56420 4012 56476
rect 3804 56410 4068 56420
rect 3612 56308 3668 56318
rect 3388 56306 3668 56308
rect 3388 56254 3614 56306
rect 3666 56254 3668 56306
rect 3388 56252 3668 56254
rect 3612 56242 3668 56252
rect 5516 56306 5572 57260
rect 5516 56254 5518 56306
rect 5570 56254 5572 56306
rect 5516 56242 5572 56254
rect 5180 56082 5236 56094
rect 5180 56030 5182 56082
rect 5234 56030 5236 56082
rect 3052 55972 3108 55982
rect 3052 55878 3108 55916
rect 4464 55692 4728 55702
rect 4520 55636 4568 55692
rect 4624 55636 4672 55692
rect 4464 55626 4728 55636
rect 5180 55468 5236 56030
rect 6076 55468 6132 57344
rect 7420 56194 7476 57344
rect 8764 56644 8820 57344
rect 10108 56756 10164 57344
rect 10108 56700 10612 56756
rect 8764 56588 9044 56644
rect 8988 56306 9044 56588
rect 8988 56254 8990 56306
rect 9042 56254 9044 56306
rect 8988 56242 9044 56254
rect 10556 56306 10612 56700
rect 10556 56254 10558 56306
rect 10610 56254 10612 56306
rect 10556 56242 10612 56254
rect 7420 56142 7422 56194
rect 7474 56142 7476 56194
rect 7420 56130 7476 56142
rect 8092 55972 8148 55982
rect 8092 55878 8148 55916
rect 9996 55970 10052 55982
rect 9996 55918 9998 55970
rect 10050 55918 10052 55970
rect 2044 55412 2548 55468
rect 5180 55412 5348 55468
rect 6076 55412 6580 55468
rect 2492 55186 2548 55412
rect 2492 55134 2494 55186
rect 2546 55134 2548 55186
rect 2492 55122 2548 55134
rect 3500 55298 3556 55310
rect 3500 55246 3502 55298
rect 3554 55246 3556 55298
rect 1372 52882 1428 52892
rect 1484 53618 1540 53630
rect 1484 53566 1486 53618
rect 1538 53566 1540 53618
rect 252 52836 308 52846
rect 140 28756 196 28766
rect 140 19796 196 28700
rect 252 26628 308 52780
rect 1036 52722 1092 52734
rect 1036 52670 1038 52722
rect 1090 52670 1092 52722
rect 1036 52276 1092 52670
rect 1036 52210 1092 52220
rect 1484 51716 1540 53566
rect 1596 52836 1652 52846
rect 1596 52742 1652 52780
rect 1484 51660 1652 51716
rect 1484 51492 1540 51502
rect 812 51490 1540 51492
rect 812 51438 1486 51490
rect 1538 51438 1540 51490
rect 812 51436 1540 51438
rect 476 49924 532 49934
rect 476 38668 532 49868
rect 364 38612 532 38668
rect 588 41860 644 41870
rect 364 27636 420 38612
rect 364 27570 420 27580
rect 476 30996 532 31006
rect 252 26562 308 26572
rect 364 27076 420 27086
rect 140 19730 196 19740
rect 252 26404 308 26414
rect 252 17780 308 26348
rect 364 20692 420 27020
rect 364 20626 420 20636
rect 252 17714 308 17724
rect 364 17108 420 17118
rect 364 10836 420 17052
rect 476 14420 532 30940
rect 588 29316 644 41804
rect 700 41076 756 41086
rect 700 33012 756 41020
rect 812 40068 868 51436
rect 1484 51426 1540 51436
rect 1036 51154 1092 51166
rect 1036 51102 1038 51154
rect 1090 51102 1092 51154
rect 1036 50932 1092 51102
rect 1036 50866 1092 50876
rect 1596 49924 1652 51660
rect 1596 49858 1652 49868
rect 1596 49700 1652 49710
rect 1596 49606 1652 49644
rect 1036 49588 1092 49598
rect 1036 49494 1092 49532
rect 1036 49026 1092 49038
rect 1036 48974 1038 49026
rect 1090 48974 1092 49026
rect 1036 48244 1092 48974
rect 1596 48916 1652 48926
rect 1596 48822 1652 48860
rect 1036 48178 1092 48188
rect 1036 47458 1092 47470
rect 1036 47406 1038 47458
rect 1090 47406 1092 47458
rect 1036 46900 1092 47406
rect 1036 46834 1092 46844
rect 1596 47346 1652 47358
rect 1596 47294 1598 47346
rect 1650 47294 1652 47346
rect 1036 45890 1092 45902
rect 1036 45838 1038 45890
rect 1090 45838 1092 45890
rect 1036 45556 1092 45838
rect 1484 45780 1540 45790
rect 1484 45686 1540 45724
rect 1036 45490 1092 45500
rect 1036 44322 1092 44334
rect 1036 44270 1038 44322
rect 1090 44270 1092 44322
rect 1036 44212 1092 44270
rect 1036 44146 1092 44156
rect 1484 44210 1540 44222
rect 1484 44158 1486 44210
rect 1538 44158 1540 44210
rect 1484 43652 1540 44158
rect 1596 43764 1652 47294
rect 1596 43698 1652 43708
rect 1484 43586 1540 43596
rect 3500 43652 3556 55246
rect 3804 54908 4068 54918
rect 3860 54852 3908 54908
rect 3964 54852 4012 54908
rect 3804 54842 4068 54852
rect 4464 54124 4728 54134
rect 4520 54068 4568 54124
rect 4624 54068 4672 54124
rect 4464 54058 4728 54068
rect 3804 53340 4068 53350
rect 3860 53284 3908 53340
rect 3964 53284 4012 53340
rect 3804 53274 4068 53284
rect 4464 52556 4728 52566
rect 4520 52500 4568 52556
rect 4624 52500 4672 52556
rect 4464 52490 4728 52500
rect 3804 51772 4068 51782
rect 3860 51716 3908 51772
rect 3964 51716 4012 51772
rect 3804 51706 4068 51716
rect 4464 50988 4728 50998
rect 4520 50932 4568 50988
rect 4624 50932 4672 50988
rect 4464 50922 4728 50932
rect 3804 50204 4068 50214
rect 3860 50148 3908 50204
rect 3964 50148 4012 50204
rect 3804 50138 4068 50148
rect 4464 49420 4728 49430
rect 4520 49364 4568 49420
rect 4624 49364 4672 49420
rect 4464 49354 4728 49364
rect 3804 48636 4068 48646
rect 3860 48580 3908 48636
rect 3964 48580 4012 48636
rect 3804 48570 4068 48580
rect 4464 47852 4728 47862
rect 4520 47796 4568 47852
rect 4624 47796 4672 47852
rect 4464 47786 4728 47796
rect 3804 47068 4068 47078
rect 3860 47012 3908 47068
rect 3964 47012 4012 47068
rect 3804 47002 4068 47012
rect 4464 46284 4728 46294
rect 4520 46228 4568 46284
rect 4624 46228 4672 46284
rect 4464 46218 4728 46228
rect 3804 45500 4068 45510
rect 3860 45444 3908 45500
rect 3964 45444 4012 45500
rect 3804 45434 4068 45444
rect 4464 44716 4728 44726
rect 4520 44660 4568 44716
rect 4624 44660 4672 44716
rect 4464 44650 4728 44660
rect 3804 43932 4068 43942
rect 3860 43876 3908 43932
rect 3964 43876 4012 43932
rect 3804 43866 4068 43876
rect 3500 43586 3556 43596
rect 3612 43764 3668 43774
rect 1596 43428 1652 43438
rect 1596 43334 1652 43372
rect 1036 43316 1092 43326
rect 924 43314 1092 43316
rect 924 43262 1038 43314
rect 1090 43262 1092 43314
rect 924 43260 1092 43262
rect 924 42868 980 43260
rect 1036 43250 1092 43260
rect 924 42802 980 42812
rect 1148 42754 1204 42766
rect 1148 42702 1150 42754
rect 1202 42702 1204 42754
rect 1036 41748 1092 41758
rect 924 41746 1092 41748
rect 924 41694 1038 41746
rect 1090 41694 1092 41746
rect 924 41692 1092 41694
rect 924 40180 980 41692
rect 1036 41682 1092 41692
rect 1148 41524 1204 42702
rect 1596 42644 1652 42654
rect 1596 42642 1876 42644
rect 1596 42590 1598 42642
rect 1650 42590 1876 42642
rect 1596 42588 1876 42590
rect 1596 42578 1652 42588
rect 1820 42532 1876 42588
rect 1820 42466 1876 42476
rect 2156 42084 2212 42094
rect 1596 41860 1652 41870
rect 1596 41766 1652 41804
rect 1148 41458 1204 41468
rect 2044 41300 2100 41310
rect 2044 41206 2100 41244
rect 924 40114 980 40124
rect 1036 41186 1092 41198
rect 1036 41134 1038 41186
rect 1090 41134 1092 41186
rect 812 40002 868 40012
rect 1036 38836 1092 41134
rect 1484 41076 1540 41086
rect 1484 40982 1540 41020
rect 2156 40514 2212 42028
rect 3612 41972 3668 43708
rect 4464 43148 4728 43158
rect 4520 43092 4568 43148
rect 4624 43092 4672 43148
rect 4464 43082 4728 43092
rect 3804 42364 4068 42374
rect 3860 42308 3908 42364
rect 3964 42308 4012 42364
rect 3804 42298 4068 42308
rect 3500 41970 3668 41972
rect 3500 41918 3614 41970
rect 3666 41918 3668 41970
rect 3500 41916 3668 41918
rect 2604 41860 2660 41870
rect 2492 41412 2548 41422
rect 2156 40462 2158 40514
rect 2210 40462 2212 40514
rect 2156 40450 2212 40462
rect 2380 41300 2436 41310
rect 1708 40402 1764 40414
rect 1708 40350 1710 40402
rect 1762 40350 1764 40402
rect 1708 40292 1764 40350
rect 1708 40226 1764 40236
rect 2268 40292 2324 40302
rect 1932 40068 1988 40078
rect 1036 38770 1092 38780
rect 1148 39618 1204 39630
rect 1148 39566 1150 39618
rect 1202 39566 1204 39618
rect 1036 38612 1092 38622
rect 924 38610 1092 38612
rect 924 38558 1038 38610
rect 1090 38558 1092 38610
rect 924 38556 1092 38558
rect 700 32946 756 32956
rect 812 36820 868 36830
rect 812 30100 868 36764
rect 924 36148 980 38556
rect 1036 38546 1092 38556
rect 1148 38052 1204 39566
rect 1036 37996 1204 38052
rect 1484 39506 1540 39518
rect 1484 39454 1486 39506
rect 1538 39454 1540 39506
rect 1036 37492 1092 37996
rect 1148 37828 1204 37838
rect 1148 37826 1316 37828
rect 1148 37774 1150 37826
rect 1202 37774 1316 37826
rect 1148 37772 1316 37774
rect 1148 37762 1204 37772
rect 1036 37426 1092 37436
rect 924 36082 980 36092
rect 1036 37268 1092 37278
rect 1036 35700 1092 37212
rect 1148 37266 1204 37278
rect 1148 37214 1150 37266
rect 1202 37214 1204 37266
rect 1148 35812 1204 37214
rect 1260 37044 1316 37772
rect 1484 37380 1540 39454
rect 1596 38722 1652 38734
rect 1596 38670 1598 38722
rect 1650 38670 1652 38722
rect 1596 38052 1652 38670
rect 1596 37996 1764 38052
rect 1484 37314 1540 37324
rect 1596 37156 1652 37166
rect 1596 37062 1652 37100
rect 1260 36988 1540 37044
rect 1260 36820 1316 36830
rect 1260 36482 1316 36764
rect 1260 36430 1262 36482
rect 1314 36430 1316 36482
rect 1260 36418 1316 36430
rect 1148 35756 1428 35812
rect 1036 35644 1316 35700
rect 1036 35476 1092 35486
rect 924 35474 1092 35476
rect 924 35422 1038 35474
rect 1090 35422 1092 35474
rect 924 35420 1092 35422
rect 924 33460 980 35420
rect 1036 35410 1092 35420
rect 924 33394 980 33404
rect 1036 34914 1092 34926
rect 1036 34862 1038 34914
rect 1090 34862 1092 34914
rect 1036 32116 1092 34862
rect 1148 34018 1204 34030
rect 1148 33966 1150 34018
rect 1202 33966 1204 34018
rect 1148 33460 1204 33966
rect 1260 33572 1316 35644
rect 1372 34804 1428 35756
rect 1372 34738 1428 34748
rect 1484 34130 1540 36988
rect 1708 36932 1764 37996
rect 1932 37042 1988 40012
rect 2044 39620 2100 39630
rect 2044 39526 2100 39564
rect 1932 36990 1934 37042
rect 1986 36990 1988 37042
rect 1708 36876 1876 36932
rect 1708 36708 1764 36718
rect 1708 36614 1764 36652
rect 1708 36260 1764 36270
rect 1596 35588 1652 35598
rect 1596 35494 1652 35532
rect 1708 35364 1764 36204
rect 1596 35308 1764 35364
rect 1596 35026 1652 35308
rect 1820 35252 1876 36876
rect 1932 36372 1988 36990
rect 1932 36306 1988 36316
rect 2268 38162 2324 40236
rect 2268 38110 2270 38162
rect 2322 38110 2324 38162
rect 1596 34974 1598 35026
rect 1650 34974 1652 35026
rect 1596 34962 1652 34974
rect 1708 35196 1876 35252
rect 1484 34078 1486 34130
rect 1538 34078 1540 34130
rect 1484 34066 1540 34078
rect 1260 33516 1540 33572
rect 1148 33404 1428 33460
rect 1260 33234 1316 33246
rect 1260 33182 1262 33234
rect 1314 33182 1316 33234
rect 1260 32676 1316 33182
rect 1036 32050 1092 32060
rect 1148 32620 1260 32676
rect 812 30034 868 30044
rect 588 29250 644 29260
rect 1036 29428 1092 29438
rect 588 29092 644 29102
rect 588 20468 644 29036
rect 1036 27858 1092 29372
rect 1036 27806 1038 27858
rect 1090 27806 1092 27858
rect 1036 27794 1092 27806
rect 1148 29426 1204 32620
rect 1260 32610 1316 32620
rect 1260 31668 1316 31678
rect 1260 30996 1316 31612
rect 1260 30902 1316 30940
rect 1148 29374 1150 29426
rect 1202 29374 1204 29426
rect 1148 28642 1204 29374
rect 1148 28590 1150 28642
rect 1202 28590 1204 28642
rect 1036 27636 1092 27646
rect 1036 26908 1092 27580
rect 1148 27188 1204 28590
rect 1260 30100 1316 30110
rect 1260 28532 1316 30044
rect 1260 28466 1316 28476
rect 1148 27074 1204 27132
rect 1148 27022 1150 27074
rect 1202 27022 1204 27074
rect 1148 27010 1204 27022
rect 1036 26852 1204 26908
rect 1036 26740 1092 26750
rect 700 26628 756 26638
rect 700 23156 756 26572
rect 1036 25730 1092 26684
rect 1036 25678 1038 25730
rect 1090 25678 1092 25730
rect 1036 25666 1092 25678
rect 1036 25396 1092 25406
rect 1036 24162 1092 25340
rect 1036 24110 1038 24162
rect 1090 24110 1092 24162
rect 1036 24098 1092 24110
rect 700 23090 756 23100
rect 924 24052 980 24062
rect 588 20402 644 20412
rect 700 22932 756 22942
rect 700 17892 756 22876
rect 812 22708 868 22718
rect 812 19796 868 22652
rect 924 21588 980 23996
rect 1148 22708 1204 26852
rect 1372 25620 1428 33404
rect 1372 25554 1428 25564
rect 1484 27188 1540 33516
rect 1596 33460 1652 33470
rect 1596 33366 1652 33404
rect 1596 33012 1652 33022
rect 1596 28756 1652 32956
rect 1708 32900 1764 35196
rect 1932 34132 1988 34142
rect 1708 32834 1764 32844
rect 1820 34130 1988 34132
rect 1820 34078 1934 34130
rect 1986 34078 1988 34130
rect 1820 34076 1988 34078
rect 1708 32676 1764 32686
rect 1708 32582 1764 32620
rect 1820 32452 1876 34076
rect 1932 34066 1988 34076
rect 2156 33906 2212 33918
rect 2156 33854 2158 33906
rect 2210 33854 2212 33906
rect 2156 33572 2212 33854
rect 2156 33506 2212 33516
rect 2268 33348 2324 38110
rect 1708 32396 1876 32452
rect 1932 33292 2324 33348
rect 1708 31668 1764 32396
rect 1708 31602 1764 31612
rect 1820 31666 1876 31678
rect 1820 31614 1822 31666
rect 1874 31614 1876 31666
rect 1820 30884 1876 31614
rect 1820 30818 1876 30828
rect 1708 29316 1764 29326
rect 1708 29222 1764 29260
rect 1596 28662 1652 28700
rect 1596 27972 1652 27982
rect 1932 27972 1988 33292
rect 2380 33236 2436 41244
rect 2492 39730 2548 41356
rect 2604 41298 2660 41804
rect 2604 41246 2606 41298
rect 2658 41246 2660 41298
rect 2604 41234 2660 41246
rect 3500 41076 3556 41916
rect 3612 41906 3668 41916
rect 4172 41860 4228 41870
rect 4172 41766 4228 41804
rect 4464 41580 4728 41590
rect 4520 41524 4568 41580
rect 4624 41524 4672 41580
rect 4464 41514 4728 41524
rect 4284 41300 4340 41310
rect 4284 41206 4340 41244
rect 3836 41188 3892 41198
rect 2492 39678 2494 39730
rect 2546 39678 2548 39730
rect 2492 39666 2548 39678
rect 2604 40402 2660 40414
rect 2604 40350 2606 40402
rect 2658 40350 2660 40402
rect 2492 37380 2548 37390
rect 2492 37286 2548 37324
rect 2604 35698 2660 40350
rect 3052 40292 3108 40302
rect 2940 39620 2996 39630
rect 2940 38948 2996 39564
rect 2716 38836 2772 38846
rect 2716 38742 2772 38780
rect 2716 37938 2772 37950
rect 2716 37886 2718 37938
rect 2770 37886 2772 37938
rect 2716 36820 2772 37886
rect 2940 37380 2996 38892
rect 3052 38722 3108 40236
rect 3052 38670 3054 38722
rect 3106 38670 3108 38722
rect 3052 38658 3108 38670
rect 3388 38050 3444 38062
rect 3388 37998 3390 38050
rect 3442 37998 3444 38050
rect 3276 37828 3332 37838
rect 2940 37324 3108 37380
rect 2716 36754 2772 36764
rect 2828 37042 2884 37054
rect 2828 36990 2830 37042
rect 2882 36990 2884 37042
rect 2828 36932 2884 36990
rect 2828 36708 2884 36876
rect 2828 36642 2884 36652
rect 2940 36820 2996 36830
rect 2604 35646 2606 35698
rect 2658 35646 2660 35698
rect 2604 35252 2660 35646
rect 2604 34916 2660 35196
rect 2156 33180 2436 33236
rect 2492 34914 2660 34916
rect 2492 34862 2606 34914
rect 2658 34862 2660 34914
rect 2492 34860 2660 34862
rect 1596 27970 1988 27972
rect 1596 27918 1598 27970
rect 1650 27918 1988 27970
rect 1596 27916 1988 27918
rect 2044 32900 2100 32910
rect 1596 27906 1652 27916
rect 1820 27636 1876 27646
rect 1596 27188 1652 27198
rect 1484 27186 1652 27188
rect 1484 27134 1598 27186
rect 1650 27134 1652 27186
rect 1484 27132 1652 27134
rect 1484 26180 1540 27132
rect 1596 27122 1652 27132
rect 1708 27188 1764 27198
rect 1708 26964 1764 27132
rect 1708 26402 1764 26908
rect 1708 26350 1710 26402
rect 1762 26350 1764 26402
rect 1708 26338 1764 26350
rect 1484 25396 1540 26124
rect 1260 25340 1540 25396
rect 1596 25396 1652 25406
rect 1260 23154 1316 25340
rect 1596 25302 1652 25340
rect 1820 25172 1876 27580
rect 2044 26068 2100 32844
rect 2156 32450 2212 33180
rect 2156 32398 2158 32450
rect 2210 32398 2212 32450
rect 2156 28756 2212 32398
rect 2268 32116 2324 32126
rect 2268 31778 2324 32060
rect 2268 31726 2270 31778
rect 2322 31726 2324 31778
rect 2268 31714 2324 31726
rect 2380 31108 2436 31118
rect 2380 30994 2436 31052
rect 2380 30942 2382 30994
rect 2434 30942 2436 30994
rect 2380 30930 2436 30942
rect 2492 30772 2548 34860
rect 2604 34850 2660 34860
rect 2716 36596 2772 36606
rect 2716 33460 2772 36540
rect 2828 36258 2884 36270
rect 2828 36206 2830 36258
rect 2882 36206 2884 36258
rect 2828 34130 2884 36206
rect 2828 34078 2830 34130
rect 2882 34078 2884 34130
rect 2828 34066 2884 34078
rect 2380 30716 2548 30772
rect 2604 33404 2716 33460
rect 2156 26908 2212 28700
rect 2268 30210 2324 30222
rect 2268 30158 2270 30210
rect 2322 30158 2324 30210
rect 2268 27076 2324 30158
rect 2268 27010 2324 27020
rect 2156 26852 2324 26908
rect 2156 26068 2212 26078
rect 2044 26012 2156 26068
rect 2156 25974 2212 26012
rect 2268 25844 2324 26852
rect 1708 25116 1876 25172
rect 1932 25788 2324 25844
rect 1372 24948 1428 24958
rect 1372 24722 1428 24892
rect 1372 24670 1374 24722
rect 1426 24670 1428 24722
rect 1372 24658 1428 24670
rect 1260 23102 1262 23154
rect 1314 23102 1316 23154
rect 1260 23090 1316 23102
rect 1372 24164 1428 24174
rect 1148 22652 1316 22708
rect 1148 22484 1204 22494
rect 1148 22390 1204 22428
rect 1036 21588 1092 21598
rect 924 21586 1092 21588
rect 924 21534 1038 21586
rect 1090 21534 1092 21586
rect 924 21532 1092 21534
rect 1036 21522 1092 21532
rect 1148 21364 1204 21374
rect 1036 20692 1092 20702
rect 1036 20018 1092 20636
rect 1036 19966 1038 20018
rect 1090 19966 1092 20018
rect 1036 19954 1092 19966
rect 812 19740 1092 19796
rect 700 17826 756 17836
rect 924 18676 980 18686
rect 700 17444 756 17454
rect 476 14354 532 14364
rect 588 15988 644 15998
rect 364 10770 420 10780
rect 476 13748 532 13758
rect 476 4452 532 13692
rect 588 10724 644 15932
rect 588 10658 644 10668
rect 476 4386 532 4396
rect 700 112 756 17388
rect 924 15148 980 18620
rect 1036 17890 1092 19740
rect 1036 17838 1038 17890
rect 1090 17838 1092 17890
rect 1036 17826 1092 17838
rect 1148 16882 1204 21308
rect 1260 20244 1316 22652
rect 1372 21140 1428 24108
rect 1596 23828 1652 23838
rect 1596 23734 1652 23772
rect 1596 23380 1652 23390
rect 1596 23266 1652 23324
rect 1596 23214 1598 23266
rect 1650 23214 1652 23266
rect 1596 23202 1652 23214
rect 1708 22820 1764 25116
rect 1596 22764 1764 22820
rect 1596 22372 1652 22764
rect 1708 22596 1764 22606
rect 1708 22502 1764 22540
rect 1596 22316 1764 22372
rect 1596 21474 1652 21486
rect 1596 21422 1598 21474
rect 1650 21422 1652 21474
rect 1372 21084 1540 21140
rect 1372 20916 1428 20926
rect 1372 20822 1428 20860
rect 1260 20178 1316 20188
rect 1372 20468 1428 20478
rect 1148 16830 1150 16882
rect 1202 16830 1204 16882
rect 1148 16818 1204 16830
rect 1260 20018 1316 20030
rect 1260 19966 1262 20018
rect 1314 19966 1316 20018
rect 1148 16660 1204 16670
rect 924 15092 1092 15148
rect 1036 14754 1092 15092
rect 1036 14702 1038 14754
rect 1090 14702 1092 14754
rect 1036 14690 1092 14702
rect 1148 14084 1204 16604
rect 812 14028 1204 14084
rect 1260 14532 1316 19966
rect 812 8260 868 14028
rect 1148 13636 1204 13646
rect 1148 13542 1204 13580
rect 1036 13524 1092 13534
rect 1036 12962 1092 13468
rect 1260 13524 1316 14476
rect 1260 13458 1316 13468
rect 1036 12910 1038 12962
rect 1090 12910 1092 12962
rect 1036 12290 1092 12910
rect 1036 12238 1038 12290
rect 1090 12238 1092 12290
rect 1036 12226 1092 12238
rect 1148 13300 1204 13310
rect 924 11956 980 11966
rect 924 8484 980 11900
rect 1036 10724 1092 10734
rect 1036 10610 1092 10668
rect 1036 10558 1038 10610
rect 1090 10558 1092 10610
rect 1036 10546 1092 10558
rect 1036 9380 1092 9390
rect 1036 8708 1092 9324
rect 1148 9042 1204 13244
rect 1260 11170 1316 11182
rect 1260 11118 1262 11170
rect 1314 11118 1316 11170
rect 1260 10612 1316 11118
rect 1260 10546 1316 10556
rect 1260 9602 1316 9614
rect 1260 9550 1262 9602
rect 1314 9550 1316 9602
rect 1260 9268 1316 9550
rect 1260 9202 1316 9212
rect 1372 9156 1428 20412
rect 1484 16994 1540 21084
rect 1596 20580 1652 21422
rect 1596 20514 1652 20524
rect 1596 20132 1652 20142
rect 1596 19684 1652 20076
rect 1596 19618 1652 19628
rect 1596 19460 1652 19470
rect 1596 19366 1652 19404
rect 1708 18452 1764 22316
rect 1932 21140 1988 25788
rect 1708 18386 1764 18396
rect 1820 21084 1988 21140
rect 2044 25620 2100 25630
rect 2044 21700 2100 25564
rect 2380 24948 2436 30716
rect 2604 29316 2660 33404
rect 2716 33394 2772 33404
rect 2828 33122 2884 33134
rect 2828 33070 2830 33122
rect 2882 33070 2884 33122
rect 2828 32116 2884 33070
rect 2828 32050 2884 32060
rect 2828 31892 2884 31902
rect 2828 31798 2884 31836
rect 2716 31778 2772 31790
rect 2716 31726 2718 31778
rect 2770 31726 2772 31778
rect 2716 30996 2772 31726
rect 2940 31108 2996 36764
rect 3052 36596 3108 37324
rect 3276 37378 3332 37772
rect 3276 37326 3278 37378
rect 3330 37326 3332 37378
rect 3276 37314 3332 37326
rect 3052 36530 3108 36540
rect 3388 37044 3444 37998
rect 3276 36372 3332 36382
rect 3164 35474 3220 35486
rect 3164 35422 3166 35474
rect 3218 35422 3220 35474
rect 3164 35364 3220 35422
rect 3164 35298 3220 35308
rect 3164 35028 3220 35038
rect 3276 35028 3332 36316
rect 3388 36260 3444 36988
rect 3500 36820 3556 41020
rect 3612 41186 3892 41188
rect 3612 41134 3838 41186
rect 3890 41134 3892 41186
rect 3612 41132 3892 41134
rect 3612 38836 3668 41132
rect 3836 41122 3892 41132
rect 3804 40796 4068 40806
rect 3860 40740 3908 40796
rect 3964 40740 4012 40796
rect 3804 40730 4068 40740
rect 4284 40404 4340 40414
rect 4284 40310 4340 40348
rect 4464 40012 4728 40022
rect 4520 39956 4568 40012
rect 4624 39956 4672 40012
rect 4464 39946 4728 39956
rect 5068 39732 5124 39742
rect 5068 39638 5124 39676
rect 3804 39228 4068 39238
rect 3860 39172 3908 39228
rect 3964 39172 4012 39228
rect 3804 39162 4068 39172
rect 3612 38770 3668 38780
rect 4284 38724 4340 38762
rect 4284 38658 4340 38668
rect 3836 38612 3892 38622
rect 3836 38162 3892 38556
rect 4464 38444 4728 38454
rect 4520 38388 4568 38444
rect 4624 38388 4672 38444
rect 4464 38378 4728 38388
rect 3836 38110 3838 38162
rect 3890 38110 3892 38162
rect 3836 38098 3892 38110
rect 5068 38162 5124 38174
rect 5068 38110 5070 38162
rect 5122 38110 5124 38162
rect 4620 38052 4676 38062
rect 4172 38050 4676 38052
rect 4172 37998 4622 38050
rect 4674 37998 4676 38050
rect 4172 37996 4676 37998
rect 3804 37660 4068 37670
rect 3860 37604 3908 37660
rect 3964 37604 4012 37660
rect 3804 37594 4068 37604
rect 3948 37044 4004 37054
rect 3500 36754 3556 36764
rect 3612 36932 3668 36942
rect 3612 36708 3668 36876
rect 3388 36194 3444 36204
rect 3500 36370 3556 36382
rect 3500 36318 3502 36370
rect 3554 36318 3556 36370
rect 3164 35026 3332 35028
rect 3164 34974 3166 35026
rect 3218 34974 3332 35026
rect 3164 34972 3332 34974
rect 3164 34962 3220 34972
rect 3164 34132 3220 34142
rect 2716 30930 2772 30940
rect 2828 31052 2996 31108
rect 3052 34130 3220 34132
rect 3052 34078 3166 34130
rect 3218 34078 3220 34130
rect 3052 34076 3220 34078
rect 2828 30324 2884 31052
rect 2828 30258 2884 30268
rect 2940 30882 2996 30894
rect 2940 30830 2942 30882
rect 2994 30830 2996 30882
rect 2716 30098 2772 30110
rect 2716 30046 2718 30098
rect 2770 30046 2772 30098
rect 2716 29988 2772 30046
rect 2716 29922 2772 29932
rect 2828 30100 2884 30110
rect 2828 29650 2884 30044
rect 2828 29598 2830 29650
rect 2882 29598 2884 29650
rect 2828 29586 2884 29598
rect 2604 29092 2660 29260
rect 2604 29026 2660 29036
rect 2828 28868 2884 28878
rect 2940 28868 2996 30830
rect 2828 28866 2996 28868
rect 2828 28814 2830 28866
rect 2882 28814 2996 28866
rect 2828 28812 2996 28814
rect 2828 28802 2884 28812
rect 2716 28532 2772 28542
rect 2716 27970 2772 28476
rect 2716 27918 2718 27970
rect 2770 27918 2772 27970
rect 2716 27906 2772 27918
rect 3052 27188 3108 34076
rect 3164 34066 3220 34076
rect 3276 33796 3332 34972
rect 3164 33740 3332 33796
rect 3388 35924 3444 35934
rect 3388 35364 3444 35868
rect 3164 30660 3220 33740
rect 3276 33572 3332 33582
rect 3276 33478 3332 33516
rect 3276 32338 3332 32350
rect 3276 32286 3278 32338
rect 3330 32286 3332 32338
rect 3276 31890 3332 32286
rect 3276 31838 3278 31890
rect 3330 31838 3332 31890
rect 3276 31826 3332 31838
rect 3388 31220 3444 35308
rect 3500 35252 3556 36318
rect 3500 34132 3556 35196
rect 3500 34066 3556 34076
rect 3612 31556 3668 36652
rect 3948 36706 4004 36988
rect 3948 36654 3950 36706
rect 4002 36654 4004 36706
rect 3948 36642 4004 36654
rect 3804 36092 4068 36102
rect 3860 36036 3908 36092
rect 3964 36036 4012 36092
rect 3804 36026 4068 36036
rect 3804 34524 4068 34534
rect 3860 34468 3908 34524
rect 3964 34468 4012 34524
rect 3804 34458 4068 34468
rect 4172 34356 4228 37996
rect 4620 37986 4676 37996
rect 4844 37492 4900 37502
rect 4464 36876 4728 36886
rect 4520 36820 4568 36876
rect 4624 36820 4672 36876
rect 4464 36810 4728 36820
rect 4284 35474 4340 35486
rect 4284 35422 4286 35474
rect 4338 35422 4340 35474
rect 4284 35140 4340 35422
rect 4464 35308 4728 35318
rect 4520 35252 4568 35308
rect 4624 35252 4672 35308
rect 4464 35242 4728 35252
rect 4284 35074 4340 35084
rect 4284 34916 4340 34926
rect 4284 34822 4340 34860
rect 4172 34300 4340 34356
rect 4060 34244 4116 34254
rect 4060 34132 4116 34188
rect 4172 34132 4228 34142
rect 4060 34130 4228 34132
rect 4060 34078 4174 34130
rect 4226 34078 4228 34130
rect 4060 34076 4228 34078
rect 4172 34066 4228 34076
rect 3836 33908 3892 33918
rect 3836 33458 3892 33852
rect 3836 33406 3838 33458
rect 3890 33406 3892 33458
rect 3836 33394 3892 33406
rect 3804 32956 4068 32966
rect 3860 32900 3908 32956
rect 3964 32900 4012 32956
rect 3804 32890 4068 32900
rect 4284 32676 4340 34300
rect 4464 33740 4728 33750
rect 4520 33684 4568 33740
rect 4624 33684 4672 33740
rect 4464 33674 4728 33684
rect 4172 32620 4340 32676
rect 4396 32676 4452 32686
rect 3724 32338 3780 32350
rect 3724 32286 3726 32338
rect 3778 32286 3780 32338
rect 3724 31892 3780 32286
rect 3724 31826 3780 31836
rect 4060 31780 4116 31790
rect 4060 31686 4116 31724
rect 3612 31490 3668 31500
rect 3804 31388 4068 31398
rect 3860 31332 3908 31388
rect 3964 31332 4012 31388
rect 3804 31322 4068 31332
rect 3388 31164 4116 31220
rect 3500 30996 3556 31006
rect 3500 30902 3556 30940
rect 3948 30994 4004 31006
rect 3948 30942 3950 30994
rect 4002 30942 4004 30994
rect 3388 30770 3444 30782
rect 3388 30718 3390 30770
rect 3442 30718 3444 30770
rect 3164 30604 3332 30660
rect 3164 30436 3220 30446
rect 3164 30342 3220 30380
rect 3164 30212 3220 30222
rect 3164 27746 3220 30156
rect 3164 27694 3166 27746
rect 3218 27694 3220 27746
rect 3164 27636 3220 27694
rect 3164 27570 3220 27580
rect 3276 27412 3332 30604
rect 3388 30436 3444 30718
rect 3388 30370 3444 30380
rect 3500 30772 3556 30782
rect 3500 30434 3556 30716
rect 3500 30382 3502 30434
rect 3554 30382 3556 30434
rect 3500 30370 3556 30382
rect 3948 30100 4004 30942
rect 4060 30322 4116 31164
rect 4060 30270 4062 30322
rect 4114 30270 4116 30322
rect 4060 30258 4116 30270
rect 3948 30034 4004 30044
rect 3804 29820 4068 29830
rect 3860 29764 3908 29820
rect 3964 29764 4012 29820
rect 3804 29754 4068 29764
rect 3724 29540 3780 29550
rect 3724 29446 3780 29484
rect 3388 29426 3444 29438
rect 3388 29374 3390 29426
rect 3442 29374 3444 29426
rect 3388 28084 3444 29374
rect 3836 28756 3892 28766
rect 3612 28754 3892 28756
rect 3612 28702 3838 28754
rect 3890 28702 3892 28754
rect 3612 28700 3892 28702
rect 3500 28532 3556 28542
rect 3500 28438 3556 28476
rect 3388 28018 3444 28028
rect 3052 27122 3108 27132
rect 3164 27356 3332 27412
rect 2828 26852 2884 26862
rect 2492 26850 2884 26852
rect 2492 26798 2830 26850
rect 2882 26798 2884 26850
rect 2492 26796 2884 26798
rect 2492 25506 2548 26796
rect 2828 26786 2884 26796
rect 2940 26516 2996 26526
rect 2492 25454 2494 25506
rect 2546 25454 2548 25506
rect 2492 25442 2548 25454
rect 2828 26292 2884 26302
rect 2828 26068 2884 26236
rect 2156 24892 2436 24948
rect 2156 22370 2212 24892
rect 2268 24724 2324 24734
rect 2268 23828 2324 24668
rect 2380 24722 2436 24734
rect 2716 24724 2772 24734
rect 2380 24670 2382 24722
rect 2434 24670 2436 24722
rect 2380 24052 2436 24670
rect 2492 24722 2772 24724
rect 2492 24670 2718 24722
rect 2770 24670 2772 24722
rect 2492 24668 2772 24670
rect 2492 24162 2548 24668
rect 2716 24658 2772 24668
rect 2492 24110 2494 24162
rect 2546 24110 2548 24162
rect 2492 24098 2548 24110
rect 2380 23986 2436 23996
rect 2380 23828 2436 23838
rect 2268 23772 2380 23828
rect 2268 23492 2324 23502
rect 2268 23266 2324 23436
rect 2268 23214 2270 23266
rect 2322 23214 2324 23266
rect 2268 23202 2324 23214
rect 2156 22318 2158 22370
rect 2210 22318 2212 22370
rect 2156 21812 2212 22318
rect 2156 21746 2212 21756
rect 2380 23044 2436 23772
rect 2716 23156 2772 23166
rect 2604 23044 2660 23054
rect 2380 23042 2660 23044
rect 2380 22990 2606 23042
rect 2658 22990 2660 23042
rect 2380 22988 2660 22990
rect 1708 18226 1764 18238
rect 1708 18174 1710 18226
rect 1762 18174 1764 18226
rect 1708 18116 1764 18174
rect 1596 17780 1652 17790
rect 1596 17686 1652 17724
rect 1708 17444 1764 18060
rect 1484 16942 1486 16994
rect 1538 16942 1540 16994
rect 1484 16930 1540 16942
rect 1596 17388 1764 17444
rect 1596 16436 1652 17388
rect 1820 17332 1876 21084
rect 2044 21028 2100 21644
rect 2044 20962 2100 20972
rect 2156 21588 2212 21598
rect 1932 20916 1988 20926
rect 1932 20822 1988 20860
rect 2044 20132 2100 20142
rect 2044 20038 2100 20076
rect 1708 17276 1876 17332
rect 1932 20020 1988 20030
rect 1708 16660 1764 17276
rect 1932 16882 1988 19964
rect 1932 16830 1934 16882
rect 1986 16830 1988 16882
rect 1932 16818 1988 16830
rect 2044 18228 2100 18238
rect 1708 16594 1764 16604
rect 1596 16380 1764 16436
rect 1708 15764 1764 16380
rect 2044 16324 2100 18172
rect 2156 17780 2212 21532
rect 2268 21028 2324 21038
rect 2268 20914 2324 20972
rect 2268 20862 2270 20914
rect 2322 20862 2324 20914
rect 2268 20850 2324 20862
rect 2156 17666 2212 17724
rect 2156 17614 2158 17666
rect 2210 17614 2212 17666
rect 2156 17602 2212 17614
rect 2268 19124 2324 19134
rect 2268 18338 2324 19068
rect 2268 18286 2270 18338
rect 2322 18286 2324 18338
rect 2268 16660 2324 18286
rect 2380 16772 2436 22988
rect 2604 22978 2660 22988
rect 2716 22596 2772 23100
rect 2492 22594 2772 22596
rect 2492 22542 2718 22594
rect 2770 22542 2772 22594
rect 2492 22540 2772 22542
rect 2492 21924 2548 22540
rect 2716 22530 2772 22540
rect 2828 22260 2884 26012
rect 2940 25508 2996 26460
rect 3052 25732 3108 25742
rect 3052 25638 3108 25676
rect 2940 25506 3108 25508
rect 2940 25454 2942 25506
rect 2994 25454 3108 25506
rect 2940 25452 3108 25454
rect 2940 25442 2996 25452
rect 3052 25284 3108 25452
rect 2492 21858 2548 21868
rect 2716 22204 2884 22260
rect 2940 25060 2996 25070
rect 2604 21588 2660 21598
rect 2604 21494 2660 21532
rect 2492 20804 2548 20814
rect 2492 18116 2548 20748
rect 2604 20802 2660 20814
rect 2604 20750 2606 20802
rect 2658 20750 2660 20802
rect 2604 19460 2660 20750
rect 2716 19908 2772 22204
rect 2828 21812 2884 21822
rect 2828 20130 2884 21756
rect 2940 20804 2996 25004
rect 2940 20738 2996 20748
rect 3052 20802 3108 25228
rect 3164 22372 3220 27356
rect 3388 27076 3444 27086
rect 3388 26982 3444 27020
rect 3276 26068 3332 26078
rect 3276 26066 3556 26068
rect 3276 26014 3278 26066
rect 3330 26014 3556 26066
rect 3276 26012 3556 26014
rect 3276 26002 3332 26012
rect 3500 25618 3556 26012
rect 3500 25566 3502 25618
rect 3554 25566 3556 25618
rect 3500 25554 3556 25566
rect 3276 25508 3332 25518
rect 3276 25060 3332 25452
rect 3612 25396 3668 28700
rect 3836 28690 3892 28700
rect 3804 28252 4068 28262
rect 3860 28196 3908 28252
rect 3964 28196 4012 28252
rect 3804 28186 4068 28196
rect 4172 27636 4228 32620
rect 4284 32452 4340 32462
rect 4396 32452 4452 32620
rect 4284 32450 4452 32452
rect 4284 32398 4286 32450
rect 4338 32398 4452 32450
rect 4284 32396 4452 32398
rect 4284 32386 4340 32396
rect 4464 32172 4728 32182
rect 4520 32116 4568 32172
rect 4624 32116 4672 32172
rect 4464 32106 4728 32116
rect 4844 32004 4900 37436
rect 5068 36708 5124 38110
rect 5068 36642 5124 36652
rect 5180 37604 5236 37614
rect 5180 37266 5236 37548
rect 5180 37214 5182 37266
rect 5234 37214 5236 37266
rect 5068 36260 5124 36270
rect 5068 36166 5124 36204
rect 4620 31948 4900 32004
rect 4956 35140 5012 35150
rect 4396 31108 4452 31118
rect 4396 30884 4452 31052
rect 4620 30996 4676 31948
rect 4732 31780 4788 31790
rect 4732 31444 4788 31724
rect 4844 31778 4900 31790
rect 4844 31726 4846 31778
rect 4898 31726 4900 31778
rect 4844 31668 4900 31726
rect 4844 31602 4900 31612
rect 4732 31388 4900 31444
rect 4620 30930 4676 30940
rect 4844 31220 4900 31388
rect 4396 30818 4452 30828
rect 4464 30604 4728 30614
rect 4520 30548 4568 30604
rect 4624 30548 4672 30604
rect 4464 30538 4728 30548
rect 4464 29036 4728 29046
rect 4520 28980 4568 29036
rect 4624 28980 4672 29036
rect 4464 28970 4728 28980
rect 4732 28532 4788 28542
rect 4284 27860 4340 27870
rect 4284 27766 4340 27804
rect 4732 27636 4788 28476
rect 4844 27748 4900 31164
rect 4956 28644 5012 35084
rect 5068 34804 5124 34814
rect 5068 34710 5124 34748
rect 5180 34356 5236 37214
rect 5068 34300 5236 34356
rect 5068 31556 5124 34300
rect 5180 34132 5236 34142
rect 5180 33684 5236 34076
rect 5180 33618 5236 33628
rect 5068 31490 5124 31500
rect 5180 33012 5236 33022
rect 5068 30098 5124 30110
rect 5068 30046 5070 30098
rect 5122 30046 5124 30098
rect 5068 29540 5124 30046
rect 5068 29474 5124 29484
rect 5180 29538 5236 32956
rect 5180 29486 5182 29538
rect 5234 29486 5236 29538
rect 5068 29092 5124 29102
rect 5068 28866 5124 29036
rect 5068 28814 5070 28866
rect 5122 28814 5124 28866
rect 5068 28802 5124 28814
rect 4956 28588 5124 28644
rect 4956 27748 5012 27758
rect 4844 27746 5012 27748
rect 4844 27694 4958 27746
rect 5010 27694 5012 27746
rect 4844 27692 5012 27694
rect 4172 27580 4340 27636
rect 4732 27580 4900 27636
rect 4172 27188 4228 27198
rect 3724 26964 3780 27002
rect 3724 26898 3780 26908
rect 3804 26684 4068 26694
rect 3860 26628 3908 26684
rect 3964 26628 4012 26684
rect 3804 26618 4068 26628
rect 4172 26516 4228 27132
rect 4284 26628 4340 27580
rect 4464 27468 4728 27478
rect 4520 27412 4568 27468
rect 4624 27412 4672 27468
rect 4464 27402 4728 27412
rect 4844 27074 4900 27580
rect 4956 27412 5012 27692
rect 4956 27346 5012 27356
rect 4844 27022 4846 27074
rect 4898 27022 4900 27074
rect 4844 27010 4900 27022
rect 4956 26964 5012 26974
rect 4284 26562 4340 26572
rect 4396 26852 4452 26862
rect 4060 26460 4228 26516
rect 3724 26066 3780 26078
rect 3724 26014 3726 26066
rect 3778 26014 3780 26066
rect 3724 25732 3780 26014
rect 3724 25666 3780 25676
rect 3276 24994 3332 25004
rect 3500 25284 3556 25294
rect 3500 24722 3556 25228
rect 3500 24670 3502 24722
rect 3554 24670 3556 24722
rect 3500 24658 3556 24670
rect 3388 24500 3444 24510
rect 3276 24498 3444 24500
rect 3276 24446 3390 24498
rect 3442 24446 3444 24498
rect 3276 24444 3444 24446
rect 3276 22596 3332 24444
rect 3388 24434 3444 24444
rect 3612 24052 3668 25340
rect 4060 25506 4116 26460
rect 4284 26404 4340 26414
rect 4396 26404 4452 26796
rect 4284 26402 4452 26404
rect 4284 26350 4286 26402
rect 4338 26350 4452 26402
rect 4284 26348 4452 26350
rect 4284 26338 4340 26348
rect 4464 25900 4728 25910
rect 4520 25844 4568 25900
rect 4624 25844 4672 25900
rect 4464 25834 4728 25844
rect 4060 25454 4062 25506
rect 4114 25454 4116 25506
rect 4060 25284 4116 25454
rect 4060 25228 4340 25284
rect 3804 25116 4068 25126
rect 3860 25060 3908 25116
rect 3964 25060 4012 25116
rect 3804 25050 4068 25060
rect 4060 24724 4116 24734
rect 4060 24722 4228 24724
rect 4060 24670 4062 24722
rect 4114 24670 4228 24722
rect 4060 24668 4228 24670
rect 4060 24658 4116 24668
rect 3276 22530 3332 22540
rect 3500 24050 3668 24052
rect 3500 23998 3614 24050
rect 3666 23998 3668 24050
rect 3500 23996 3668 23998
rect 3164 22316 3332 22372
rect 3164 21924 3220 21934
rect 3164 21474 3220 21868
rect 3164 21422 3166 21474
rect 3218 21422 3220 21474
rect 3164 21410 3220 21422
rect 3276 21140 3332 22316
rect 3052 20750 3054 20802
rect 3106 20750 3108 20802
rect 3052 20738 3108 20750
rect 3164 21084 3332 21140
rect 3164 20580 3220 21084
rect 3276 20916 3332 20926
rect 3276 20822 3332 20860
rect 2828 20078 2830 20130
rect 2882 20078 2884 20130
rect 2828 20066 2884 20078
rect 2940 20524 3220 20580
rect 2716 19852 2884 19908
rect 2604 19394 2660 19404
rect 2716 19684 2772 19694
rect 2716 19458 2772 19628
rect 2716 19406 2718 19458
rect 2770 19406 2772 19458
rect 2716 19348 2772 19406
rect 2716 19282 2772 19292
rect 2492 18050 2548 18060
rect 2604 18452 2660 18462
rect 2604 17778 2660 18396
rect 2716 18452 2772 18462
rect 2828 18452 2884 19852
rect 2716 18450 2884 18452
rect 2716 18398 2718 18450
rect 2770 18398 2884 18450
rect 2716 18396 2884 18398
rect 2716 18386 2772 18396
rect 2940 17892 2996 20524
rect 3388 19348 3444 19358
rect 3164 19124 3220 19134
rect 3164 19030 3220 19068
rect 3164 18452 3220 18462
rect 3164 18358 3220 18396
rect 3388 18004 3444 19292
rect 3500 18676 3556 23996
rect 3612 23986 3668 23996
rect 4060 24500 4116 24510
rect 4060 23940 4116 24444
rect 3724 23938 4116 23940
rect 3724 23886 4062 23938
rect 4114 23886 4116 23938
rect 3724 23884 4116 23886
rect 3724 23716 3780 23884
rect 4060 23874 4116 23884
rect 3612 23660 3780 23716
rect 3612 23492 3668 23660
rect 3804 23548 4068 23558
rect 3860 23492 3908 23548
rect 3964 23492 4012 23548
rect 3804 23482 4068 23492
rect 3612 23426 3668 23436
rect 3836 23380 3892 23390
rect 4172 23380 4228 24668
rect 4284 24612 4340 25228
rect 4396 24612 4452 24622
rect 4284 24610 4452 24612
rect 4284 24558 4398 24610
rect 4450 24558 4452 24610
rect 4284 24556 4452 24558
rect 4284 23940 4340 24556
rect 4396 24546 4452 24556
rect 4956 24500 5012 26908
rect 5068 26908 5124 28588
rect 5180 28532 5236 29486
rect 5180 28466 5236 28476
rect 5292 28084 5348 55412
rect 6524 55186 6580 55412
rect 6524 55134 6526 55186
rect 6578 55134 6580 55186
rect 6524 55122 6580 55134
rect 7532 55298 7588 55310
rect 7532 55246 7534 55298
rect 7586 55246 7588 55298
rect 6524 52276 6580 52286
rect 5740 49700 5796 49710
rect 5516 40962 5572 40974
rect 5516 40910 5518 40962
rect 5570 40910 5572 40962
rect 5516 39618 5572 40910
rect 5516 39566 5518 39618
rect 5570 39566 5572 39618
rect 5516 39554 5572 39566
rect 5516 38836 5572 38846
rect 5516 37604 5572 38780
rect 5516 37538 5572 37548
rect 5516 37154 5572 37166
rect 5516 37102 5518 37154
rect 5570 37102 5572 37154
rect 5516 36708 5572 37102
rect 5516 36642 5572 36652
rect 5516 36260 5572 36270
rect 5404 34916 5460 34926
rect 5404 34822 5460 34860
rect 5404 30210 5460 30222
rect 5404 30158 5406 30210
rect 5458 30158 5460 30210
rect 5404 29092 5460 30158
rect 5404 29026 5460 29036
rect 5516 28868 5572 36204
rect 5740 35364 5796 49644
rect 6076 48916 6132 48926
rect 6076 41412 6132 48860
rect 5852 41410 6132 41412
rect 5852 41358 6078 41410
rect 6130 41358 6132 41410
rect 5852 41356 6132 41358
rect 5852 39956 5908 41356
rect 6076 41346 6132 41356
rect 6412 40180 6468 40190
rect 5852 39890 5908 39900
rect 6076 40178 6468 40180
rect 6076 40126 6414 40178
rect 6466 40126 6468 40178
rect 6076 40124 6468 40126
rect 6076 39842 6132 40124
rect 6412 40114 6468 40124
rect 6076 39790 6078 39842
rect 6130 39790 6132 39842
rect 6076 39778 6132 39790
rect 6188 39956 6244 39966
rect 5852 39618 5908 39630
rect 5852 39566 5854 39618
rect 5906 39566 5908 39618
rect 5852 36036 5908 39566
rect 5964 38948 6020 38958
rect 5964 38722 6020 38892
rect 5964 38670 5966 38722
rect 6018 38670 6020 38722
rect 5964 38658 6020 38670
rect 6188 38668 6244 39900
rect 6076 38612 6244 38668
rect 6300 39508 6356 39518
rect 5852 35980 6020 36036
rect 5852 35812 5908 35822
rect 5852 35718 5908 35756
rect 5964 35588 6020 35980
rect 5628 33908 5684 33918
rect 5740 33908 5796 35308
rect 5852 35532 6020 35588
rect 5852 34914 5908 35532
rect 6076 35364 6132 38612
rect 6300 38274 6356 39452
rect 6524 39284 6580 52220
rect 6636 51380 6692 51390
rect 6636 41298 6692 51324
rect 7420 48916 7476 48926
rect 6636 41246 6638 41298
rect 6690 41246 6692 41298
rect 6636 41234 6692 41246
rect 7084 48244 7140 48254
rect 6636 40628 6692 40638
rect 6636 39508 6692 40572
rect 6972 40516 7028 40526
rect 6972 40422 7028 40460
rect 7084 40292 7140 48188
rect 6972 40236 7140 40292
rect 7308 40290 7364 40302
rect 7308 40238 7310 40290
rect 7362 40238 7364 40290
rect 6636 39442 6692 39452
rect 6748 39618 6804 39630
rect 6748 39566 6750 39618
rect 6802 39566 6804 39618
rect 6524 39228 6692 39284
rect 6636 38668 6692 39228
rect 6748 39060 6804 39566
rect 6748 38994 6804 39004
rect 6300 38222 6302 38274
rect 6354 38222 6356 38274
rect 6300 38210 6356 38222
rect 6412 38612 6692 38668
rect 5852 34862 5854 34914
rect 5906 34862 5908 34914
rect 5852 34468 5908 34862
rect 5852 34402 5908 34412
rect 5964 35308 6132 35364
rect 6188 36482 6244 36494
rect 6188 36430 6190 36482
rect 6242 36430 6244 36482
rect 5628 33906 5796 33908
rect 5628 33854 5630 33906
rect 5682 33854 5796 33906
rect 5628 33852 5796 33854
rect 5628 33842 5684 33852
rect 5628 33234 5684 33246
rect 5628 33182 5630 33234
rect 5682 33182 5684 33234
rect 5628 33012 5684 33182
rect 5628 32946 5684 32956
rect 5740 29988 5796 33852
rect 5852 30212 5908 30222
rect 5852 30118 5908 30156
rect 5740 29932 5908 29988
rect 5180 28028 5348 28084
rect 5404 28812 5572 28868
rect 5628 29202 5684 29214
rect 5628 29150 5630 29202
rect 5682 29150 5684 29202
rect 5180 27636 5236 28028
rect 5292 27860 5348 27870
rect 5292 27766 5348 27804
rect 5180 27580 5348 27636
rect 5068 26852 5236 26908
rect 4956 24434 5012 24444
rect 5068 25506 5124 25518
rect 5068 25454 5070 25506
rect 5122 25454 5124 25506
rect 4464 24332 4728 24342
rect 4520 24276 4568 24332
rect 4624 24276 4672 24332
rect 4464 24266 4728 24276
rect 5068 24164 5124 25454
rect 4956 24108 5124 24164
rect 4284 23874 4340 23884
rect 4620 24052 4676 24062
rect 4620 23826 4676 23996
rect 4620 23774 4622 23826
rect 4674 23774 4676 23826
rect 3836 23378 4228 23380
rect 3836 23326 3838 23378
rect 3890 23326 4228 23378
rect 3836 23324 4228 23326
rect 4284 23604 4340 23614
rect 3836 23314 3892 23324
rect 4284 23268 4340 23548
rect 4172 23212 4340 23268
rect 3836 22148 3892 22158
rect 3612 22146 3892 22148
rect 3612 22094 3838 22146
rect 3890 22094 3892 22146
rect 3612 22092 3892 22094
rect 3612 20916 3668 22092
rect 3836 22082 3892 22092
rect 3804 21980 4068 21990
rect 3860 21924 3908 21980
rect 3964 21924 4012 21980
rect 3804 21914 4068 21924
rect 3724 20916 3780 20926
rect 3612 20914 3780 20916
rect 3612 20862 3726 20914
rect 3778 20862 3780 20914
rect 3612 20860 3780 20862
rect 3724 20850 3780 20860
rect 3804 20412 4068 20422
rect 3860 20356 3908 20412
rect 3964 20356 4012 20412
rect 3804 20346 4068 20356
rect 3836 20132 3892 20142
rect 3612 20018 3668 20030
rect 3612 19966 3614 20018
rect 3666 19966 3668 20018
rect 3612 19124 3668 19966
rect 3612 19058 3668 19068
rect 3836 19012 3892 20076
rect 4172 20132 4228 23212
rect 4620 22932 4676 23774
rect 4956 23716 5012 24108
rect 5068 23940 5124 23950
rect 5180 23940 5236 26852
rect 5068 23938 5236 23940
rect 5068 23886 5070 23938
rect 5122 23886 5236 23938
rect 5068 23884 5236 23886
rect 5068 23874 5124 23884
rect 4956 23660 5124 23716
rect 4620 22876 4900 22932
rect 4464 22764 4728 22774
rect 4520 22708 4568 22764
rect 4624 22708 4672 22764
rect 4464 22698 4728 22708
rect 4844 22260 4900 22876
rect 4956 22260 5012 22270
rect 4844 22258 5012 22260
rect 4844 22206 4958 22258
rect 5010 22206 5012 22258
rect 4844 22204 5012 22206
rect 4284 21812 4340 21822
rect 4284 21718 4340 21756
rect 4464 21196 4728 21206
rect 4520 21140 4568 21196
rect 4624 21140 4672 21196
rect 4464 21130 4728 21140
rect 4172 20066 4228 20076
rect 4508 20802 4564 20814
rect 4508 20750 4510 20802
rect 4562 20750 4564 20802
rect 4508 20020 4564 20750
rect 4508 19954 4564 19964
rect 4464 19628 4728 19638
rect 4520 19572 4568 19628
rect 4624 19572 4672 19628
rect 4464 19562 4728 19572
rect 4508 19348 4564 19358
rect 4508 19254 4564 19292
rect 4172 19124 4228 19134
rect 4172 19122 4340 19124
rect 4172 19070 4174 19122
rect 4226 19070 4340 19122
rect 4172 19068 4340 19070
rect 4172 19058 4228 19068
rect 3836 18946 3892 18956
rect 3500 18610 3556 18620
rect 3612 18900 3668 18910
rect 4284 18900 4340 19068
rect 3612 18452 3668 18844
rect 3804 18844 4068 18854
rect 3860 18788 3908 18844
rect 3964 18788 4012 18844
rect 3804 18778 4068 18788
rect 3164 17948 3444 18004
rect 3500 18396 3668 18452
rect 4172 18676 4228 18686
rect 2940 17836 3108 17892
rect 2604 17726 2606 17778
rect 2658 17726 2660 17778
rect 2604 17714 2660 17726
rect 2492 17668 2548 17678
rect 2492 16994 2548 17612
rect 2492 16942 2494 16994
rect 2546 16942 2548 16994
rect 2492 16930 2548 16942
rect 2828 16882 2884 16894
rect 2828 16830 2830 16882
rect 2882 16830 2884 16882
rect 2380 16716 2772 16772
rect 2268 16594 2324 16604
rect 2044 16268 2436 16324
rect 1932 15876 1988 15886
rect 1932 15782 1988 15820
rect 1708 15698 1764 15708
rect 2156 15764 2212 15774
rect 1484 15092 1540 15102
rect 1484 13746 1540 15036
rect 1932 15092 1988 15102
rect 1932 14998 1988 15036
rect 2044 14980 2100 14990
rect 1820 14868 1876 14878
rect 1708 14644 1764 14654
rect 1596 14418 1652 14430
rect 1596 14366 1598 14418
rect 1650 14366 1652 14418
rect 1596 13860 1652 14366
rect 1596 13794 1652 13804
rect 1484 13694 1486 13746
rect 1538 13694 1540 13746
rect 1484 13682 1540 13694
rect 1596 12850 1652 12862
rect 1596 12798 1598 12850
rect 1650 12798 1652 12850
rect 1484 12178 1540 12190
rect 1484 12126 1486 12178
rect 1538 12126 1540 12178
rect 1484 9380 1540 12126
rect 1596 11396 1652 12798
rect 1708 11956 1764 14588
rect 1820 13748 1876 14812
rect 1932 14532 1988 14570
rect 1932 14466 1988 14476
rect 1932 13748 1988 13758
rect 1820 13692 1932 13748
rect 1932 13654 1988 13692
rect 1932 12180 1988 12190
rect 1932 12086 1988 12124
rect 1708 11900 1988 11956
rect 1596 11330 1652 11340
rect 1596 10836 1652 10846
rect 1596 10722 1652 10780
rect 1596 10670 1598 10722
rect 1650 10670 1652 10722
rect 1596 10658 1652 10670
rect 1932 10610 1988 11900
rect 1932 10558 1934 10610
rect 1986 10558 1988 10610
rect 1932 10546 1988 10558
rect 2044 9826 2100 14924
rect 2156 13748 2212 15708
rect 2156 13682 2212 13692
rect 2156 13524 2212 13534
rect 2156 13522 2324 13524
rect 2156 13470 2158 13522
rect 2210 13470 2324 13522
rect 2156 13468 2324 13470
rect 2156 13458 2212 13468
rect 2156 13300 2212 13310
rect 2156 12962 2212 13244
rect 2156 12910 2158 12962
rect 2210 12910 2212 12962
rect 2156 12898 2212 12910
rect 2268 12180 2324 13468
rect 2268 12114 2324 12124
rect 2268 11620 2324 11630
rect 2268 11506 2324 11564
rect 2268 11454 2270 11506
rect 2322 11454 2324 11506
rect 2268 11442 2324 11454
rect 2380 10722 2436 16268
rect 2604 15876 2660 15886
rect 2492 14644 2548 14654
rect 2492 14550 2548 14588
rect 2492 13972 2548 13982
rect 2492 12628 2548 13916
rect 2604 13746 2660 15820
rect 2604 13694 2606 13746
rect 2658 13694 2660 13746
rect 2604 13682 2660 13694
rect 2604 13076 2660 13086
rect 2716 13076 2772 16716
rect 2828 16660 2884 16830
rect 2828 16594 2884 16604
rect 2940 16884 2996 16894
rect 2828 15204 2884 15214
rect 2828 14754 2884 15148
rect 2828 14702 2830 14754
rect 2882 14702 2884 14754
rect 2828 14690 2884 14702
rect 2604 13074 2772 13076
rect 2604 13022 2606 13074
rect 2658 13022 2772 13074
rect 2604 13020 2772 13022
rect 2604 13010 2660 13020
rect 2492 12572 2660 12628
rect 2492 12068 2548 12078
rect 2492 11974 2548 12012
rect 2604 11618 2660 12572
rect 2604 11566 2606 11618
rect 2658 11566 2660 11618
rect 2604 11554 2660 11566
rect 2380 10670 2382 10722
rect 2434 10670 2436 10722
rect 2380 10658 2436 10670
rect 2044 9774 2046 9826
rect 2098 9774 2100 9826
rect 2044 9762 2100 9774
rect 2156 10500 2212 10510
rect 1484 9314 1540 9324
rect 1596 9604 1652 9614
rect 1484 9156 1540 9166
rect 1372 9154 1540 9156
rect 1372 9102 1486 9154
rect 1538 9102 1540 9154
rect 1372 9100 1540 9102
rect 1484 9090 1540 9100
rect 1148 8990 1150 9042
rect 1202 8990 1204 9042
rect 1148 8978 1204 8990
rect 1036 8652 1204 8708
rect 1036 8484 1092 8494
rect 924 8482 1092 8484
rect 924 8430 1038 8482
rect 1090 8430 1092 8482
rect 924 8428 1092 8430
rect 1036 8418 1092 8428
rect 812 8194 868 8204
rect 1036 7924 1092 7934
rect 1036 7474 1092 7868
rect 1036 7422 1038 7474
rect 1090 7422 1092 7474
rect 1036 7410 1092 7422
rect 1036 4114 1092 4126
rect 1036 4062 1038 4114
rect 1090 4062 1092 4114
rect 1036 3892 1092 4062
rect 1036 3826 1092 3836
rect 1148 2772 1204 8652
rect 1596 8484 1652 9548
rect 2044 9156 2100 9166
rect 2044 9042 2100 9100
rect 2044 8990 2046 9042
rect 2098 8990 2100 9042
rect 2044 8978 2100 8990
rect 1484 8428 1652 8484
rect 1484 7586 1540 8428
rect 1596 8260 1652 8270
rect 1596 8166 1652 8204
rect 1484 7534 1486 7586
rect 1538 7534 1540 7586
rect 1484 7522 1540 7534
rect 2156 6690 2212 10444
rect 2716 9826 2772 13020
rect 2940 12404 2996 16828
rect 3052 16324 3108 17836
rect 3052 16258 3108 16268
rect 3164 16210 3220 17948
rect 3276 16996 3332 17006
rect 3276 16902 3332 16940
rect 3164 16158 3166 16210
rect 3218 16158 3220 16210
rect 3052 16100 3108 16110
rect 3052 15204 3108 16044
rect 3052 15138 3108 15148
rect 3164 15148 3220 16158
rect 3500 16100 3556 18396
rect 3836 18228 3892 18238
rect 3836 18134 3892 18172
rect 3724 17892 3780 17902
rect 3724 17798 3780 17836
rect 3500 16006 3556 16044
rect 3612 17668 3668 17678
rect 3612 15314 3668 17612
rect 3804 17276 4068 17286
rect 3860 17220 3908 17276
rect 3964 17220 4012 17276
rect 3804 17210 4068 17220
rect 3836 16884 3892 16894
rect 3836 16790 3892 16828
rect 3804 15708 4068 15718
rect 3860 15652 3908 15708
rect 3964 15652 4012 15708
rect 3804 15642 4068 15652
rect 3612 15262 3614 15314
rect 3666 15262 3668 15314
rect 3276 15204 3332 15214
rect 2716 9774 2718 9826
rect 2770 9774 2772 9826
rect 2716 9762 2772 9774
rect 2828 12348 2996 12404
rect 3164 15092 3332 15148
rect 2492 8932 2548 8942
rect 2492 8838 2548 8876
rect 2156 6638 2158 6690
rect 2210 6638 2212 6690
rect 2156 6626 2212 6638
rect 1260 6580 1316 6590
rect 1260 6486 1316 6524
rect 1260 6018 1316 6030
rect 1260 5966 1262 6018
rect 1314 5966 1316 6018
rect 1260 5236 1316 5966
rect 2268 5908 2324 5918
rect 2828 5908 2884 12348
rect 2940 12180 2996 12190
rect 3164 12180 3220 15092
rect 3276 14756 3332 14766
rect 3276 14418 3332 14700
rect 3276 14366 3278 14418
rect 3330 14366 3332 14418
rect 3276 14354 3332 14366
rect 3388 13746 3444 13758
rect 3388 13694 3390 13746
rect 3442 13694 3444 13746
rect 3388 13636 3444 13694
rect 3388 13570 3444 13580
rect 3276 12404 3332 12414
rect 3276 12290 3332 12348
rect 3276 12238 3278 12290
rect 3330 12238 3332 12290
rect 3276 12226 3332 12238
rect 2940 12178 3220 12180
rect 2940 12126 2942 12178
rect 2994 12126 3220 12178
rect 2940 12124 3220 12126
rect 2940 12114 2996 12124
rect 3276 11508 3332 11518
rect 2940 11284 2996 11294
rect 2940 10610 2996 11228
rect 3164 11282 3220 11294
rect 3164 11230 3166 11282
rect 3218 11230 3220 11282
rect 3164 11172 3220 11230
rect 3164 11106 3220 11116
rect 3276 10722 3332 11452
rect 3612 11396 3668 15262
rect 4172 15148 4228 18620
rect 4284 17780 4340 18844
rect 4396 18452 4452 18462
rect 4396 18358 4452 18396
rect 4464 18060 4728 18070
rect 4520 18004 4568 18060
rect 4624 18004 4672 18060
rect 4464 17994 4728 18004
rect 4284 17666 4340 17724
rect 4284 17614 4286 17666
rect 4338 17614 4340 17666
rect 4284 17602 4340 17614
rect 4620 17892 4676 17902
rect 4284 16882 4340 16894
rect 4284 16830 4286 16882
rect 4338 16830 4340 16882
rect 4284 16324 4340 16830
rect 4620 16660 4676 17836
rect 4844 17892 4900 17902
rect 4844 17798 4900 17836
rect 4956 17108 5012 22204
rect 5068 21140 5124 23660
rect 5292 22596 5348 27580
rect 5404 27524 5460 28812
rect 5516 28644 5572 28654
rect 5516 28550 5572 28588
rect 5404 27468 5572 27524
rect 5404 27300 5460 27310
rect 5404 27206 5460 27244
rect 5516 27188 5572 27468
rect 5516 27122 5572 27132
rect 5628 26908 5684 29150
rect 5740 27860 5796 27870
rect 5740 27766 5796 27804
rect 5516 26852 5684 26908
rect 5404 24948 5460 24958
rect 5404 24164 5460 24892
rect 5516 24724 5572 26852
rect 5516 24658 5572 24668
rect 5740 26740 5796 26750
rect 5628 24498 5684 24510
rect 5628 24446 5630 24498
rect 5682 24446 5684 24498
rect 5404 24108 5572 24164
rect 5068 21074 5124 21084
rect 5180 22540 5348 22596
rect 5404 23940 5460 23950
rect 5180 18564 5236 22540
rect 5292 22370 5348 22382
rect 5292 22318 5294 22370
rect 5346 22318 5348 22370
rect 5292 21812 5348 22318
rect 5404 22372 5460 23884
rect 5404 22306 5460 22316
rect 5292 21746 5348 21756
rect 5516 21698 5572 24108
rect 5628 24162 5684 24446
rect 5628 24110 5630 24162
rect 5682 24110 5684 24162
rect 5628 24098 5684 24110
rect 5740 23380 5796 26684
rect 5516 21646 5518 21698
rect 5570 21646 5572 21698
rect 5516 21634 5572 21646
rect 5628 23324 5796 23380
rect 5292 21140 5348 21150
rect 5628 21140 5684 23324
rect 5852 23268 5908 29932
rect 5964 28868 6020 35308
rect 6076 35140 6132 35150
rect 6188 35140 6244 36430
rect 6300 35474 6356 35486
rect 6300 35422 6302 35474
rect 6354 35422 6356 35474
rect 6300 35364 6356 35422
rect 6300 35298 6356 35308
rect 6076 35138 6244 35140
rect 6076 35086 6078 35138
rect 6130 35086 6244 35138
rect 6076 35084 6244 35086
rect 6076 35074 6132 35084
rect 6300 34804 6356 34814
rect 6076 33572 6132 33582
rect 6076 33478 6132 33516
rect 6300 32450 6356 34748
rect 6300 32398 6302 32450
rect 6354 32398 6356 32450
rect 6300 30884 6356 32398
rect 6300 30818 6356 30828
rect 6188 30770 6244 30782
rect 6188 30718 6190 30770
rect 6242 30718 6244 30770
rect 6076 30436 6132 30446
rect 6188 30436 6244 30718
rect 6076 30434 6244 30436
rect 6076 30382 6078 30434
rect 6130 30382 6244 30434
rect 6076 30380 6244 30382
rect 6076 30370 6132 30380
rect 6412 30212 6468 38612
rect 6748 38050 6804 38062
rect 6748 37998 6750 38050
rect 6802 37998 6804 38050
rect 6748 37716 6804 37998
rect 6972 37940 7028 40236
rect 7084 39618 7140 39630
rect 7084 39566 7086 39618
rect 7138 39566 7140 39618
rect 7084 38668 7140 39566
rect 7308 39618 7364 40238
rect 7308 39566 7310 39618
rect 7362 39566 7364 39618
rect 7308 39554 7364 39566
rect 7196 39060 7252 39070
rect 7196 38966 7252 39004
rect 7084 38612 7364 38668
rect 7196 37940 7252 37950
rect 6972 37938 7252 37940
rect 6972 37886 7198 37938
rect 7250 37886 7252 37938
rect 6972 37884 7252 37886
rect 7196 37874 7252 37884
rect 6636 37660 6804 37716
rect 6636 37268 6692 37660
rect 7308 37604 7364 38612
rect 7420 37828 7476 48860
rect 7532 39956 7588 55246
rect 9996 54628 10052 55918
rect 11452 55188 11508 57344
rect 12796 56644 12852 57344
rect 14140 56756 14196 57344
rect 14140 56700 14644 56756
rect 12796 56588 13076 56644
rect 13020 56306 13076 56588
rect 13020 56254 13022 56306
rect 13074 56254 13076 56306
rect 13020 56242 13076 56254
rect 14588 56306 14644 56700
rect 14588 56254 14590 56306
rect 14642 56254 14644 56306
rect 14588 56242 14644 56254
rect 15484 56308 15540 57344
rect 16828 57204 16884 57344
rect 16828 57148 16996 57204
rect 15484 56242 15540 56252
rect 16492 56308 16548 56318
rect 16492 56214 16548 56252
rect 11564 55970 11620 55982
rect 11564 55918 11566 55970
rect 11618 55918 11620 55970
rect 11564 55412 11620 55918
rect 11564 55346 11620 55356
rect 14028 55970 14084 55982
rect 14028 55918 14030 55970
rect 14082 55918 14084 55970
rect 12908 55298 12964 55310
rect 12908 55246 12910 55298
rect 12962 55246 12964 55298
rect 11900 55188 11956 55198
rect 11452 55186 11956 55188
rect 11452 55134 11902 55186
rect 11954 55134 11956 55186
rect 11452 55132 11956 55134
rect 11900 55122 11956 55132
rect 9996 54562 10052 54572
rect 10892 54404 10948 54414
rect 9212 54068 9268 54078
rect 8876 41188 8932 41198
rect 8428 41186 8932 41188
rect 8428 41134 8878 41186
rect 8930 41134 8932 41186
rect 8428 41132 8932 41134
rect 7644 40628 7700 40638
rect 7644 40402 7700 40572
rect 7644 40350 7646 40402
rect 7698 40350 7700 40402
rect 7644 40338 7700 40350
rect 8092 40402 8148 40414
rect 8092 40350 8094 40402
rect 8146 40350 8148 40402
rect 7532 39890 7588 39900
rect 8092 39732 8148 40350
rect 8316 40292 8372 40302
rect 8428 40292 8484 41132
rect 8876 41122 8932 41132
rect 8988 41188 9044 41198
rect 8316 40290 8484 40292
rect 8316 40238 8318 40290
rect 8370 40238 8484 40290
rect 8316 40236 8484 40238
rect 8652 40628 8708 40638
rect 8316 40226 8372 40236
rect 7756 38500 7812 38510
rect 7756 38162 7812 38444
rect 7756 38110 7758 38162
rect 7810 38110 7812 38162
rect 7756 38098 7812 38110
rect 7420 37762 7476 37772
rect 7308 37548 8036 37604
rect 6748 37492 6804 37502
rect 6748 37490 7924 37492
rect 6748 37438 6750 37490
rect 6802 37438 7924 37490
rect 6748 37436 7924 37438
rect 6748 37426 6804 37436
rect 6636 37212 6804 37268
rect 6524 37156 6580 37166
rect 6524 33572 6580 37100
rect 6636 36370 6692 36382
rect 6636 36318 6638 36370
rect 6690 36318 6692 36370
rect 6636 35028 6692 36318
rect 6748 35924 6804 37212
rect 7868 37266 7924 37436
rect 7868 37214 7870 37266
rect 7922 37214 7924 37266
rect 7868 37202 7924 37214
rect 6748 35858 6804 35868
rect 6972 37156 7028 37166
rect 6972 35700 7028 37100
rect 7532 37156 7588 37166
rect 7532 37062 7588 37100
rect 6636 34962 6692 34972
rect 6860 35644 7028 35700
rect 7756 36370 7812 36382
rect 7756 36318 7758 36370
rect 7810 36318 7812 36370
rect 6748 34914 6804 34926
rect 6748 34862 6750 34914
rect 6802 34862 6804 34914
rect 6524 33506 6580 33516
rect 6636 34356 6692 34366
rect 6188 30156 6468 30212
rect 6524 31556 6580 31566
rect 5964 28812 6132 28868
rect 5964 28642 6020 28654
rect 5964 28590 5966 28642
rect 6018 28590 6020 28642
rect 5964 27746 6020 28590
rect 5964 27694 5966 27746
rect 6018 27694 6020 27746
rect 5964 27682 6020 27694
rect 6076 27524 6132 28812
rect 5964 27468 6132 27524
rect 5964 27300 6020 27468
rect 5964 26740 6020 27244
rect 5964 26674 6020 26684
rect 6076 27188 6132 27198
rect 5964 26292 6020 26302
rect 5964 25620 6020 26236
rect 5964 25554 6020 25564
rect 6076 24050 6132 27132
rect 6188 25060 6244 30156
rect 6524 30100 6580 31500
rect 6636 31106 6692 34300
rect 6748 34354 6804 34862
rect 6748 34302 6750 34354
rect 6802 34302 6804 34354
rect 6748 34290 6804 34302
rect 6748 32564 6804 32574
rect 6748 32470 6804 32508
rect 6636 31054 6638 31106
rect 6690 31054 6692 31106
rect 6636 31042 6692 31054
rect 6300 30044 6580 30100
rect 6636 30884 6692 30894
rect 6636 30100 6692 30828
rect 6300 26964 6356 30044
rect 6636 30034 6692 30044
rect 6748 30210 6804 30222
rect 6748 30158 6750 30210
rect 6802 30158 6804 30210
rect 6748 29650 6804 30158
rect 6748 29598 6750 29650
rect 6802 29598 6804 29650
rect 6748 29586 6804 29598
rect 6636 28532 6692 28542
rect 6636 28438 6692 28476
rect 6300 26898 6356 26908
rect 6412 28420 6468 28430
rect 6300 26628 6356 26638
rect 6300 26292 6356 26572
rect 6300 25508 6356 26236
rect 6300 25414 6356 25452
rect 6188 25004 6356 25060
rect 6188 24836 6244 24846
rect 6188 24742 6244 24780
rect 6076 23998 6078 24050
rect 6130 23998 6132 24050
rect 6076 23986 6132 23998
rect 6300 23380 6356 25004
rect 6300 23314 6356 23324
rect 5852 23212 6132 23268
rect 5740 23156 5796 23166
rect 5740 23154 6020 23156
rect 5740 23102 5742 23154
rect 5794 23102 6020 23154
rect 5740 23100 6020 23102
rect 5740 23090 5796 23100
rect 5964 22594 6020 23100
rect 5964 22542 5966 22594
rect 6018 22542 6020 22594
rect 5964 22530 6020 22542
rect 5292 20802 5348 21084
rect 5292 20750 5294 20802
rect 5346 20750 5348 20802
rect 5292 20738 5348 20750
rect 5404 21084 5684 21140
rect 5740 22372 5796 22382
rect 5180 18498 5236 18508
rect 5404 17892 5460 21084
rect 5628 20916 5684 20926
rect 5628 19796 5684 20860
rect 5740 20020 5796 22316
rect 5964 21364 6020 21374
rect 5964 21270 6020 21308
rect 6076 20916 6132 23212
rect 6188 23156 6244 23166
rect 6188 23062 6244 23100
rect 6300 21700 6356 21710
rect 6300 21606 6356 21644
rect 5964 20860 6132 20916
rect 6300 21028 6356 21038
rect 5740 19954 5796 19964
rect 5852 20804 5908 20814
rect 5404 17826 5460 17836
rect 5516 19794 5684 19796
rect 5516 19742 5630 19794
rect 5682 19742 5684 19794
rect 5516 19740 5684 19742
rect 5516 18452 5572 19740
rect 5628 19730 5684 19740
rect 5740 19460 5796 19470
rect 5740 19366 5796 19404
rect 5852 19236 5908 20748
rect 5964 19572 6020 20860
rect 6188 20804 6244 20814
rect 6188 20710 6244 20748
rect 6188 20132 6244 20142
rect 6188 20038 6244 20076
rect 5964 19516 6244 19572
rect 5740 19180 5908 19236
rect 5964 19348 6020 19358
rect 5516 17444 5572 18396
rect 5516 17378 5572 17388
rect 5628 18452 5684 18462
rect 5740 18452 5796 19180
rect 5964 18676 6020 19292
rect 5628 18450 5796 18452
rect 5628 18398 5630 18450
rect 5682 18398 5796 18450
rect 5628 18396 5796 18398
rect 5852 18620 6020 18676
rect 4956 17052 5124 17108
rect 4956 16884 5012 16894
rect 4956 16790 5012 16828
rect 5068 16660 5124 17052
rect 4620 16604 4900 16660
rect 4464 16492 4728 16502
rect 4520 16436 4568 16492
rect 4624 16436 4672 16492
rect 4464 16426 4728 16436
rect 4284 16258 4340 16268
rect 4732 16212 4788 16222
rect 4732 16118 4788 16156
rect 4284 16100 4340 16110
rect 4284 16006 4340 16044
rect 4172 15092 4340 15148
rect 4172 14196 4228 14206
rect 3804 14140 4068 14150
rect 3860 14084 3908 14140
rect 3964 14084 4012 14140
rect 3804 14074 4068 14084
rect 4172 13636 4228 14140
rect 4284 13972 4340 15092
rect 4464 14924 4728 14934
rect 4520 14868 4568 14924
rect 4624 14868 4672 14924
rect 4464 14858 4728 14868
rect 4844 14530 4900 16604
rect 4844 14478 4846 14530
rect 4898 14478 4900 14530
rect 4844 14466 4900 14478
rect 4956 16604 5124 16660
rect 5180 16772 5236 16782
rect 4508 14418 4564 14430
rect 4508 14366 4510 14418
rect 4562 14366 4564 14418
rect 4508 14196 4564 14366
rect 4508 14130 4564 14140
rect 4844 14308 4900 14318
rect 4284 13906 4340 13916
rect 4284 13748 4340 13758
rect 4284 13654 4340 13692
rect 3724 12964 3780 12974
rect 3724 12870 3780 12908
rect 4172 12850 4228 13580
rect 4464 13356 4728 13366
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4464 13290 4728 13300
rect 4508 12964 4564 12974
rect 4844 12964 4900 14252
rect 4956 14084 5012 16604
rect 5180 15148 5236 16716
rect 4956 14018 5012 14028
rect 5068 15092 5236 15148
rect 5404 16660 5460 16670
rect 4956 12964 5012 12974
rect 4844 12962 5012 12964
rect 4844 12910 4958 12962
rect 5010 12910 5012 12962
rect 4844 12908 5012 12910
rect 4508 12870 4564 12908
rect 4956 12898 5012 12908
rect 4172 12798 4174 12850
rect 4226 12798 4228 12850
rect 4172 12786 4228 12798
rect 3804 12572 4068 12582
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 3804 12506 4068 12516
rect 4284 12516 4340 12526
rect 4284 12290 4340 12460
rect 4284 12238 4286 12290
rect 4338 12238 4340 12290
rect 4284 12226 4340 12238
rect 3724 12180 3780 12190
rect 3724 12086 3780 12124
rect 4464 11788 4728 11798
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4464 11722 4728 11732
rect 4844 11620 4900 11630
rect 5068 11620 5124 15092
rect 5292 14980 5348 14990
rect 5292 14530 5348 14924
rect 5292 14478 5294 14530
rect 5346 14478 5348 14530
rect 5292 14420 5348 14478
rect 5292 14354 5348 14364
rect 5180 13746 5236 13758
rect 5180 13694 5182 13746
rect 5234 13694 5236 13746
rect 5180 13300 5236 13694
rect 5180 13234 5236 13244
rect 4844 11618 5124 11620
rect 4844 11566 4846 11618
rect 4898 11566 5124 11618
rect 4844 11564 5124 11566
rect 4844 11554 4900 11564
rect 3612 11330 3668 11340
rect 4396 11396 4452 11406
rect 4396 11282 4452 11340
rect 4396 11230 4398 11282
rect 4450 11230 4452 11282
rect 3804 11004 4068 11014
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 3804 10938 4068 10948
rect 3276 10670 3278 10722
rect 3330 10670 3332 10722
rect 3276 10658 3332 10670
rect 2940 10558 2942 10610
rect 2994 10558 2996 10610
rect 2940 10546 2996 10558
rect 4396 10388 4452 11230
rect 5068 10612 5124 11564
rect 5068 10546 5124 10556
rect 5180 13074 5236 13086
rect 5180 13022 5182 13074
rect 5234 13022 5236 13074
rect 4396 10322 4452 10332
rect 4464 10220 4728 10230
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4464 10154 4728 10164
rect 3164 10052 3220 10062
rect 3164 9938 3220 9996
rect 3164 9886 3166 9938
rect 3218 9886 3220 9938
rect 3164 9874 3220 9886
rect 4732 9940 4788 9950
rect 4732 9846 4788 9884
rect 5180 9826 5236 13022
rect 5292 10612 5348 10622
rect 5292 10518 5348 10556
rect 5180 9774 5182 9826
rect 5234 9774 5236 9826
rect 5180 9762 5236 9774
rect 3804 9436 4068 9446
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 3804 9370 4068 9380
rect 4464 8652 4728 8662
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4464 8586 4728 8596
rect 5404 8428 5460 16604
rect 5628 16324 5684 18396
rect 5852 16994 5908 18620
rect 6076 18228 6132 18238
rect 6076 18134 6132 18172
rect 5852 16942 5854 16994
rect 5906 16942 5908 16994
rect 5852 16930 5908 16942
rect 5964 17442 6020 17454
rect 5964 17390 5966 17442
rect 6018 17390 6020 17442
rect 5628 16258 5684 16268
rect 5740 16884 5796 16894
rect 5740 15426 5796 16828
rect 5740 15374 5742 15426
rect 5794 15374 5796 15426
rect 5740 15362 5796 15374
rect 5852 15874 5908 15886
rect 5852 15822 5854 15874
rect 5906 15822 5908 15874
rect 5516 14642 5572 14654
rect 5516 14590 5518 14642
rect 5570 14590 5572 14642
rect 5516 12178 5572 14590
rect 5628 13972 5684 13982
rect 5628 13634 5684 13916
rect 5852 13748 5908 15822
rect 5964 14642 6020 17390
rect 6188 16772 6244 19516
rect 6188 16706 6244 16716
rect 6300 16548 6356 20972
rect 5964 14590 5966 14642
rect 6018 14590 6020 14642
rect 5964 14578 6020 14590
rect 6076 16492 6356 16548
rect 5628 13582 5630 13634
rect 5682 13582 5684 13634
rect 5628 13570 5684 13582
rect 5740 13692 5908 13748
rect 5516 12126 5518 12178
rect 5570 12126 5572 12178
rect 5516 12114 5572 12126
rect 5740 10724 5796 13692
rect 5852 13524 5908 13534
rect 5852 12962 5908 13468
rect 5852 12910 5854 12962
rect 5906 12910 5908 12962
rect 5852 12898 5908 12910
rect 5964 12292 6020 12302
rect 6076 12292 6132 16492
rect 6188 15204 6244 15242
rect 6188 15138 6244 15148
rect 6412 14644 6468 28364
rect 6524 27858 6580 27870
rect 6524 27806 6526 27858
rect 6578 27806 6580 27858
rect 6524 27298 6580 27806
rect 6860 27860 6916 35644
rect 7420 35474 7476 35486
rect 7420 35422 7422 35474
rect 7474 35422 7476 35474
rect 7420 35364 7476 35422
rect 7420 35298 7476 35308
rect 7196 34914 7252 34926
rect 7196 34862 7198 34914
rect 7250 34862 7252 34914
rect 7084 34468 7140 34478
rect 7084 32562 7140 34412
rect 7196 33348 7252 34862
rect 7756 34020 7812 36318
rect 7868 35588 7924 35598
rect 7980 35588 8036 37548
rect 7868 35586 8036 35588
rect 7868 35534 7870 35586
rect 7922 35534 8036 35586
rect 7868 35532 8036 35534
rect 7868 35522 7924 35532
rect 7756 33964 7924 34020
rect 7532 33908 7588 33918
rect 7532 33906 7812 33908
rect 7532 33854 7534 33906
rect 7586 33854 7812 33906
rect 7532 33852 7812 33854
rect 7532 33842 7588 33852
rect 7644 33348 7700 33358
rect 7196 33282 7252 33292
rect 7308 33346 7700 33348
rect 7308 33294 7646 33346
rect 7698 33294 7700 33346
rect 7308 33292 7700 33294
rect 7084 32510 7086 32562
rect 7138 32510 7140 32562
rect 7084 32340 7140 32510
rect 7196 33122 7252 33134
rect 7196 33070 7198 33122
rect 7250 33070 7252 33122
rect 7196 32564 7252 33070
rect 7196 32498 7252 32508
rect 7308 32450 7364 33292
rect 7644 33282 7700 33292
rect 7308 32398 7310 32450
rect 7362 32398 7364 32450
rect 7308 32386 7364 32398
rect 7420 33124 7476 33134
rect 7420 32564 7476 33068
rect 7084 32274 7140 32284
rect 7308 31780 7364 31790
rect 7196 31106 7252 31118
rect 7196 31054 7198 31106
rect 7250 31054 7252 31106
rect 7084 30210 7140 30222
rect 7084 30158 7086 30210
rect 7138 30158 7140 30210
rect 7084 30100 7140 30158
rect 7084 30034 7140 30044
rect 6972 28756 7028 28766
rect 6972 28662 7028 28700
rect 6972 27860 7028 27870
rect 6860 27804 6972 27860
rect 6524 27246 6526 27298
rect 6578 27246 6580 27298
rect 6524 27234 6580 27246
rect 6636 25620 6692 25630
rect 6636 25526 6692 25564
rect 6748 25172 6804 25182
rect 6748 23154 6804 25116
rect 6860 25060 6916 25070
rect 6860 23938 6916 25004
rect 6860 23886 6862 23938
rect 6914 23886 6916 23938
rect 6860 23716 6916 23886
rect 6860 23650 6916 23660
rect 6748 23102 6750 23154
rect 6802 23102 6804 23154
rect 6524 22370 6580 22382
rect 6524 22318 6526 22370
rect 6578 22318 6580 22370
rect 6524 19460 6580 22318
rect 6748 21812 6804 23102
rect 6972 22596 7028 27804
rect 7084 27858 7140 27870
rect 7084 27806 7086 27858
rect 7138 27806 7140 27858
rect 7084 25060 7140 27806
rect 7084 24994 7140 25004
rect 7196 23268 7252 31054
rect 7308 30772 7364 31724
rect 7308 30706 7364 30716
rect 7308 30212 7364 30222
rect 7420 30212 7476 32508
rect 7756 32562 7812 33852
rect 7756 32510 7758 32562
rect 7810 32510 7812 32562
rect 7756 32498 7812 32510
rect 7756 32340 7812 32350
rect 7644 31556 7700 31566
rect 7644 30996 7700 31500
rect 7644 30930 7700 30940
rect 7644 30772 7700 30782
rect 7644 30678 7700 30716
rect 7364 30156 7476 30212
rect 7308 23268 7364 30156
rect 7420 28532 7476 28542
rect 7420 25172 7476 28476
rect 7644 26292 7700 26302
rect 7644 26198 7700 26236
rect 7420 25106 7476 25116
rect 7532 25060 7588 25070
rect 7532 24610 7588 25004
rect 7532 24558 7534 24610
rect 7586 24558 7588 24610
rect 7308 23212 7476 23268
rect 7196 23202 7252 23212
rect 7196 22930 7252 22942
rect 7196 22878 7198 22930
rect 7250 22878 7252 22930
rect 6972 22540 7140 22596
rect 6972 22372 7028 22382
rect 6972 22278 7028 22316
rect 6636 21756 6804 21812
rect 6636 21364 6692 21756
rect 6748 21586 6804 21598
rect 6748 21534 6750 21586
rect 6802 21534 6804 21586
rect 6748 21476 6804 21534
rect 7084 21588 7140 22540
rect 7084 21494 7140 21532
rect 6748 21420 7028 21476
rect 6636 21308 6804 21364
rect 6748 21140 6804 21308
rect 6748 21084 6916 21140
rect 6636 20916 6692 20926
rect 6636 20822 6692 20860
rect 6748 20132 6804 20142
rect 6748 20038 6804 20076
rect 6524 19394 6580 19404
rect 6636 20018 6692 20030
rect 6636 19966 6638 20018
rect 6690 19966 6692 20018
rect 6636 19348 6692 19966
rect 6636 19282 6692 19292
rect 6636 19124 6692 19134
rect 6636 19030 6692 19068
rect 6860 19124 6916 21084
rect 6972 19572 7028 21420
rect 7196 20916 7252 22878
rect 7308 21364 7364 21374
rect 7308 21270 7364 21308
rect 7196 20850 7252 20860
rect 7420 20468 7476 23212
rect 7532 23044 7588 24558
rect 7644 23940 7700 23978
rect 7644 23874 7700 23884
rect 7532 22978 7588 22988
rect 7644 23716 7700 23726
rect 7196 19908 7252 19918
rect 7252 19852 7364 19908
rect 7196 19814 7252 19852
rect 6972 19516 7252 19572
rect 6860 19058 6916 19068
rect 6972 19348 7028 19358
rect 6972 18900 7028 19292
rect 6860 18844 7028 18900
rect 7084 19346 7140 19358
rect 7084 19294 7086 19346
rect 7138 19294 7140 19346
rect 6636 18564 6692 18574
rect 6636 17668 6692 18508
rect 6636 17574 6692 17612
rect 6636 16884 6692 16894
rect 6524 16100 6580 16110
rect 6636 16100 6692 16828
rect 6860 16436 6916 18844
rect 7084 18340 7140 19294
rect 7196 18450 7252 19516
rect 7196 18398 7198 18450
rect 7250 18398 7252 18450
rect 7196 18386 7252 18398
rect 6972 18284 7140 18340
rect 6972 18228 7028 18284
rect 6972 17778 7028 18172
rect 6972 17726 6974 17778
rect 7026 17726 7028 17778
rect 6972 17714 7028 17726
rect 7084 16772 7140 16782
rect 7084 16678 7140 16716
rect 7308 16436 7364 19852
rect 7420 19348 7476 20412
rect 7420 19282 7476 19292
rect 7532 22372 7588 22382
rect 7644 22372 7700 23660
rect 7588 22316 7700 22372
rect 6860 16380 7028 16436
rect 6524 16098 6692 16100
rect 6524 16046 6526 16098
rect 6578 16046 6692 16098
rect 6524 16044 6692 16046
rect 6860 16210 6916 16222
rect 6860 16158 6862 16210
rect 6914 16158 6916 16210
rect 6524 16034 6580 16044
rect 6860 15316 6916 16158
rect 6860 15250 6916 15260
rect 6972 15148 7028 16380
rect 5964 12290 6132 12292
rect 5964 12238 5966 12290
rect 6018 12238 6132 12290
rect 5964 12236 6132 12238
rect 6300 14588 6468 14644
rect 6860 15092 7028 15148
rect 7196 16380 7364 16436
rect 7420 19124 7476 19134
rect 5964 12226 6020 12236
rect 5740 10658 5796 10668
rect 5852 11732 5908 11742
rect 5852 10722 5908 11676
rect 5852 10670 5854 10722
rect 5906 10670 5908 10722
rect 5852 10658 5908 10670
rect 5964 11170 6020 11182
rect 5964 11118 5966 11170
rect 6018 11118 6020 11170
rect 5964 10612 6020 11118
rect 5964 10546 6020 10556
rect 6300 9940 6356 14588
rect 6524 14532 6580 14542
rect 6412 14530 6580 14532
rect 6412 14478 6526 14530
rect 6578 14478 6580 14530
rect 6412 14476 6580 14478
rect 6412 13748 6468 14476
rect 6524 14466 6580 14476
rect 6412 13188 6468 13692
rect 6748 13524 6804 13534
rect 6748 13430 6804 13468
rect 6412 12962 6468 13132
rect 6412 12910 6414 12962
rect 6466 12910 6468 12962
rect 6412 12898 6468 12910
rect 6636 12180 6692 12190
rect 6636 11394 6692 12124
rect 6636 11342 6638 11394
rect 6690 11342 6692 11394
rect 6636 11330 6692 11342
rect 6748 10724 6804 10734
rect 6860 10724 6916 15092
rect 6972 12180 7028 12190
rect 6972 12086 7028 12124
rect 7084 12068 7140 12078
rect 7084 11618 7140 12012
rect 7084 11566 7086 11618
rect 7138 11566 7140 11618
rect 7084 11554 7140 11566
rect 7196 12068 7252 16380
rect 7308 15764 7364 15774
rect 7308 15538 7364 15708
rect 7308 15486 7310 15538
rect 7362 15486 7364 15538
rect 7308 15474 7364 15486
rect 7420 13970 7476 19068
rect 7420 13918 7422 13970
rect 7474 13918 7476 13970
rect 7420 13906 7476 13918
rect 7308 12964 7364 12974
rect 7308 12870 7364 12908
rect 7532 12292 7588 22316
rect 7644 14756 7700 14766
rect 7644 14530 7700 14700
rect 7644 14478 7646 14530
rect 7698 14478 7700 14530
rect 7644 14466 7700 14478
rect 7756 13524 7812 32284
rect 7868 25620 7924 33964
rect 7980 29988 8036 35532
rect 8092 35700 8148 39676
rect 8204 39620 8260 39630
rect 8204 39526 8260 39564
rect 8316 38052 8372 38062
rect 8316 38050 8596 38052
rect 8316 37998 8318 38050
rect 8370 37998 8596 38050
rect 8316 37996 8596 37998
rect 8316 37986 8372 37996
rect 8316 37492 8372 37502
rect 8316 37266 8372 37436
rect 8316 37214 8318 37266
rect 8370 37214 8372 37266
rect 8316 37202 8372 37214
rect 8204 37156 8260 37166
rect 8204 36708 8260 37100
rect 8540 37154 8596 37996
rect 8540 37102 8542 37154
rect 8594 37102 8596 37154
rect 8540 37090 8596 37102
rect 8204 36652 8484 36708
rect 8316 36482 8372 36494
rect 8316 36430 8318 36482
rect 8370 36430 8372 36482
rect 8092 34916 8148 35644
rect 8204 35698 8260 35710
rect 8204 35646 8206 35698
rect 8258 35646 8260 35698
rect 8204 35364 8260 35646
rect 8316 35588 8372 36430
rect 8316 35522 8372 35532
rect 8428 35364 8484 36652
rect 8652 35924 8708 40572
rect 8764 40404 8820 40414
rect 8764 40310 8820 40348
rect 8988 39956 9044 41132
rect 8204 35298 8260 35308
rect 8316 35308 8484 35364
rect 8540 35868 8708 35924
rect 8764 39900 9044 39956
rect 8204 34916 8260 34926
rect 8092 34914 8260 34916
rect 8092 34862 8206 34914
rect 8258 34862 8260 34914
rect 8092 34860 8260 34862
rect 8204 33796 8260 34860
rect 8204 33730 8260 33740
rect 8092 33684 8148 33694
rect 8092 30994 8148 33628
rect 8204 33572 8260 33582
rect 8204 33458 8260 33516
rect 8204 33406 8206 33458
rect 8258 33406 8260 33458
rect 8204 33394 8260 33406
rect 8092 30942 8094 30994
rect 8146 30942 8148 30994
rect 8092 30930 8148 30942
rect 8204 30212 8260 30222
rect 8316 30212 8372 35308
rect 8428 32564 8484 32574
rect 8428 32470 8484 32508
rect 8540 30660 8596 35868
rect 8652 35700 8708 35738
rect 8652 35634 8708 35644
rect 8652 35476 8708 35486
rect 8652 34018 8708 35420
rect 8652 33966 8654 34018
rect 8706 33966 8708 34018
rect 8652 31892 8708 33966
rect 8764 32788 8820 39900
rect 8988 38724 9044 38734
rect 8988 37266 9044 38668
rect 8988 37214 8990 37266
rect 9042 37214 9044 37266
rect 8988 37202 9044 37214
rect 8988 36258 9044 36270
rect 8988 36206 8990 36258
rect 9042 36206 9044 36258
rect 8988 35700 9044 36206
rect 9212 36148 9268 54012
rect 9996 49028 10052 49038
rect 9324 41074 9380 41086
rect 9324 41022 9326 41074
rect 9378 41022 9380 41074
rect 9324 40628 9380 41022
rect 9324 40562 9380 40572
rect 9436 40404 9492 40414
rect 9436 39620 9492 40348
rect 9548 40404 9604 40414
rect 9548 40402 9828 40404
rect 9548 40350 9550 40402
rect 9602 40350 9828 40402
rect 9548 40348 9828 40350
rect 9548 40338 9604 40348
rect 9772 39620 9828 40348
rect 9884 39844 9940 39854
rect 9884 39750 9940 39788
rect 9436 39618 9716 39620
rect 9436 39566 9438 39618
rect 9490 39566 9716 39618
rect 9436 39564 9716 39566
rect 9436 39554 9492 39564
rect 9436 38052 9492 38062
rect 9436 37958 9492 37996
rect 9548 37268 9604 37278
rect 9212 36082 9268 36092
rect 9436 37266 9604 37268
rect 9436 37214 9550 37266
rect 9602 37214 9604 37266
rect 9436 37212 9604 37214
rect 8988 35634 9044 35644
rect 9324 35700 9380 35710
rect 9324 35606 9380 35644
rect 8876 35588 8932 35598
rect 8876 35494 8932 35532
rect 9212 35588 9268 35598
rect 9100 35476 9156 35486
rect 9100 34242 9156 35420
rect 9100 34190 9102 34242
rect 9154 34190 9156 34242
rect 9100 33012 9156 34190
rect 9100 32946 9156 32956
rect 9212 32788 9268 35532
rect 9436 32788 9492 37212
rect 9548 37202 9604 37212
rect 9660 36148 9716 39564
rect 9548 36092 9716 36148
rect 9548 33684 9604 36092
rect 9772 36036 9828 39564
rect 9996 38668 10052 48972
rect 10892 41860 10948 54348
rect 12908 53396 12964 55246
rect 13580 54292 13636 54302
rect 12908 53330 12964 53340
rect 13020 53956 13076 53966
rect 12796 52388 12852 52398
rect 11004 50708 11060 50718
rect 11004 42084 11060 50652
rect 12796 44548 12852 52332
rect 13020 50428 13076 53900
rect 13580 50428 13636 54236
rect 14028 53844 14084 55918
rect 15596 55970 15652 55982
rect 15596 55918 15598 55970
rect 15650 55918 15652 55970
rect 15596 55524 15652 55918
rect 15596 55458 15652 55468
rect 16940 55468 16996 57148
rect 18172 56308 18228 57344
rect 18508 56308 18564 56318
rect 18172 56306 18564 56308
rect 18172 56254 18510 56306
rect 18562 56254 18564 56306
rect 18172 56252 18564 56254
rect 18508 56242 18564 56252
rect 19516 56308 19572 57344
rect 19516 56242 19572 56252
rect 20636 56308 20692 56318
rect 20636 56214 20692 56252
rect 20860 56308 20916 57344
rect 22204 57204 22260 57344
rect 22204 57148 22708 57204
rect 20860 56242 20916 56252
rect 21868 56308 21924 56318
rect 21868 56214 21924 56252
rect 22540 56196 22596 56206
rect 20188 56082 20244 56094
rect 20188 56030 20190 56082
rect 20242 56030 20244 56082
rect 17500 55970 17556 55982
rect 17500 55918 17502 55970
rect 17554 55918 17556 55970
rect 16940 55412 17332 55468
rect 17276 55186 17332 55412
rect 17276 55134 17278 55186
rect 17330 55134 17332 55186
rect 17276 55122 17332 55134
rect 14028 53778 14084 53788
rect 17500 53620 17556 55918
rect 19516 55970 19572 55982
rect 19516 55918 19518 55970
rect 19570 55918 19572 55970
rect 19516 55468 19572 55918
rect 18844 55412 18900 55422
rect 19516 55412 19684 55468
rect 18844 55318 18900 55356
rect 18284 55298 18340 55310
rect 18284 55246 18286 55298
rect 18338 55246 18340 55298
rect 17500 53554 17556 53564
rect 17612 54180 17668 54190
rect 15148 52948 15204 52958
rect 14252 50484 14308 50494
rect 13020 50372 13300 50428
rect 13580 50372 13748 50428
rect 12796 44492 13188 44548
rect 11004 42018 11060 42028
rect 11340 43652 11396 43662
rect 10892 41794 10948 41804
rect 10556 41298 10612 41310
rect 10556 41246 10558 41298
rect 10610 41246 10612 41298
rect 10108 41186 10164 41198
rect 10108 41134 10110 41186
rect 10162 41134 10164 41186
rect 10108 40404 10164 41134
rect 10556 41076 10612 41246
rect 10556 41010 10612 41020
rect 10108 40338 10164 40348
rect 10444 40402 10500 40414
rect 10444 40350 10446 40402
rect 10498 40350 10500 40402
rect 9548 33346 9604 33628
rect 9548 33294 9550 33346
rect 9602 33294 9604 33346
rect 9548 33282 9604 33294
rect 9660 35980 9828 36036
rect 9884 38612 10052 38668
rect 9660 35700 9716 35980
rect 9884 35924 9940 38612
rect 9996 38162 10052 38174
rect 9996 38110 9998 38162
rect 10050 38110 10052 38162
rect 9996 37828 10052 38110
rect 9996 37044 10052 37772
rect 9996 36978 10052 36988
rect 10108 36594 10164 36606
rect 10108 36542 10110 36594
rect 10162 36542 10164 36594
rect 10108 36372 10164 36542
rect 10108 36306 10164 36316
rect 8764 32722 8820 32732
rect 9100 32732 9268 32788
rect 9324 32732 9492 32788
rect 9548 32788 9604 32798
rect 8652 30882 8708 31836
rect 8876 31780 8932 31790
rect 8876 31686 8932 31724
rect 8652 30830 8654 30882
rect 8706 30830 8708 30882
rect 8652 30818 8708 30830
rect 8540 30604 8708 30660
rect 8204 30210 8316 30212
rect 8204 30158 8206 30210
rect 8258 30158 8316 30210
rect 8204 30156 8316 30158
rect 8204 30146 8260 30156
rect 8316 30118 8372 30156
rect 7980 29932 8372 29988
rect 8204 28418 8260 28430
rect 8204 28366 8206 28418
rect 8258 28366 8260 28418
rect 8092 27858 8148 27870
rect 8092 27806 8094 27858
rect 8146 27806 8148 27858
rect 7980 26180 8036 26190
rect 7980 26086 8036 26124
rect 7868 25564 8036 25620
rect 7868 25282 7924 25294
rect 7868 25230 7870 25282
rect 7922 25230 7924 25282
rect 7868 24722 7924 25230
rect 7868 24670 7870 24722
rect 7922 24670 7924 24722
rect 7868 24658 7924 24670
rect 7980 24500 8036 25564
rect 7980 24434 8036 24444
rect 7868 23940 7924 23950
rect 7868 21812 7924 23884
rect 8092 23492 8148 27806
rect 8204 27860 8260 28366
rect 8204 27794 8260 27804
rect 8316 26908 8372 29932
rect 8540 29426 8596 29438
rect 8540 29374 8542 29426
rect 8594 29374 8596 29426
rect 8204 26852 8372 26908
rect 8428 29204 8484 29214
rect 8204 24388 8260 26852
rect 8204 24322 8260 24332
rect 8316 24722 8372 24734
rect 8316 24670 8318 24722
rect 8370 24670 8372 24722
rect 8092 23426 8148 23436
rect 8316 23156 8372 24670
rect 7868 21746 7924 21756
rect 7980 23100 8372 23156
rect 7980 21700 8036 23100
rect 8316 22930 8372 22942
rect 8316 22878 8318 22930
rect 8370 22878 8372 22930
rect 8316 22484 8372 22878
rect 8316 22418 8372 22428
rect 8092 22370 8148 22382
rect 8092 22318 8094 22370
rect 8146 22318 8148 22370
rect 8092 22260 8148 22318
rect 8092 22194 8148 22204
rect 8204 22372 8260 22382
rect 7980 21634 8036 21644
rect 8092 21812 8148 21822
rect 7868 21586 7924 21598
rect 7868 21534 7870 21586
rect 7922 21534 7924 21586
rect 7868 21026 7924 21534
rect 7868 20974 7870 21026
rect 7922 20974 7924 21026
rect 7868 20962 7924 20974
rect 8092 19236 8148 21756
rect 8204 19458 8260 22316
rect 8316 21924 8372 21934
rect 8316 21586 8372 21868
rect 8316 21534 8318 21586
rect 8370 21534 8372 21586
rect 8316 21522 8372 21534
rect 8316 20020 8372 20030
rect 8316 19926 8372 19964
rect 8428 19908 8484 29148
rect 8540 28532 8596 29374
rect 8540 28466 8596 28476
rect 8652 27412 8708 30604
rect 8876 29316 8932 29326
rect 8876 29222 8932 29260
rect 9100 28532 9156 32732
rect 9212 32557 9268 32569
rect 9212 32505 9214 32557
rect 9266 32505 9268 32557
rect 9212 32452 9268 32505
rect 9212 29540 9268 32396
rect 9212 29474 9268 29484
rect 9324 30212 9380 32732
rect 9436 32564 9492 32574
rect 9436 31890 9492 32508
rect 9436 31838 9438 31890
rect 9490 31838 9492 31890
rect 9436 31826 9492 31838
rect 9436 30212 9492 30222
rect 9324 30210 9492 30212
rect 9324 30158 9438 30210
rect 9490 30158 9492 30210
rect 9324 30156 9492 30158
rect 9100 28476 9268 28532
rect 9100 28308 9156 28318
rect 8988 28084 9044 28094
rect 8988 27970 9044 28028
rect 8988 27918 8990 27970
rect 9042 27918 9044 27970
rect 8988 27906 9044 27918
rect 9100 27636 9156 28252
rect 8652 27346 8708 27356
rect 8988 27580 9156 27636
rect 8876 25508 8932 25518
rect 8540 25506 8932 25508
rect 8540 25454 8878 25506
rect 8930 25454 8932 25506
rect 8540 25452 8932 25454
rect 8540 24610 8596 25452
rect 8876 25442 8932 25452
rect 8540 24558 8542 24610
rect 8594 24558 8596 24610
rect 8540 24546 8596 24558
rect 8428 19842 8484 19852
rect 8540 24276 8596 24286
rect 8540 19684 8596 24220
rect 8988 23380 9044 27580
rect 9212 26908 9268 28476
rect 9324 28084 9380 30156
rect 9436 30146 9492 30156
rect 9324 28018 9380 28028
rect 9436 29316 9492 29326
rect 9324 27860 9380 27870
rect 9324 27766 9380 27804
rect 8204 19406 8206 19458
rect 8258 19406 8260 19458
rect 8204 19394 8260 19406
rect 8428 19628 8596 19684
rect 8652 23324 9044 23380
rect 9100 26852 9268 26908
rect 8092 19170 8148 19180
rect 8092 18564 8148 18574
rect 8092 18470 8148 18508
rect 8204 17442 8260 17454
rect 8204 17390 8206 17442
rect 8258 17390 8260 17442
rect 7868 16884 7924 16894
rect 7868 15314 7924 16828
rect 7868 15262 7870 15314
rect 7922 15262 7924 15314
rect 7868 15250 7924 15262
rect 7980 16324 8036 16334
rect 7532 12226 7588 12236
rect 7644 13468 7812 13524
rect 7308 12068 7364 12078
rect 7196 12066 7364 12068
rect 7196 12014 7310 12066
rect 7362 12014 7364 12066
rect 7196 12012 7364 12014
rect 6748 10722 6916 10724
rect 6748 10670 6750 10722
rect 6802 10670 6916 10722
rect 6748 10668 6916 10670
rect 6748 10658 6804 10668
rect 7084 10612 7140 10622
rect 7084 10518 7140 10556
rect 6300 9874 6356 9884
rect 7084 9716 7140 9726
rect 7084 9622 7140 9660
rect 7196 9156 7252 12012
rect 7308 12002 7364 12012
rect 7420 12068 7476 12078
rect 7196 9090 7252 9100
rect 7420 9380 7476 12012
rect 7644 10612 7700 13468
rect 7756 13300 7812 13310
rect 7756 13186 7812 13244
rect 7756 13134 7758 13186
rect 7810 13134 7812 13186
rect 7756 13122 7812 13134
rect 7980 11788 8036 16268
rect 8204 16324 8260 17390
rect 8316 17332 8372 17342
rect 8316 17106 8372 17276
rect 8316 17054 8318 17106
rect 8370 17054 8372 17106
rect 8316 17042 8372 17054
rect 8204 16258 8260 16268
rect 8316 16212 8372 16222
rect 8092 15988 8148 15998
rect 8092 15894 8148 15932
rect 8316 15202 8372 16156
rect 8316 15150 8318 15202
rect 8370 15150 8372 15202
rect 8316 15138 8372 15150
rect 8204 13746 8260 13758
rect 8204 13694 8206 13746
rect 8258 13694 8260 13746
rect 8204 12852 8260 13694
rect 8204 12180 8260 12796
rect 8204 12114 8260 12124
rect 7980 11732 8148 11788
rect 7644 10610 8036 10612
rect 7644 10558 7646 10610
rect 7698 10558 8036 10610
rect 7644 10556 8036 10558
rect 7644 10546 7700 10556
rect 7756 10386 7812 10398
rect 7756 10334 7758 10386
rect 7810 10334 7812 10386
rect 7532 10052 7588 10062
rect 7756 10052 7812 10334
rect 7532 10050 7812 10052
rect 7532 9998 7534 10050
rect 7586 9998 7812 10050
rect 7532 9996 7812 9998
rect 7532 9986 7588 9996
rect 7980 9604 8036 10556
rect 7980 9538 8036 9548
rect 7308 9044 7364 9054
rect 7308 8950 7364 8988
rect 7420 8932 7476 9324
rect 8092 9044 8148 11732
rect 8204 11396 8260 11406
rect 8204 11302 8260 11340
rect 8204 10724 8260 10734
rect 8204 10610 8260 10668
rect 8204 10558 8206 10610
rect 8258 10558 8260 10610
rect 8204 10546 8260 10558
rect 8428 10052 8484 19628
rect 8540 18452 8596 18462
rect 8540 18338 8596 18396
rect 8540 18286 8542 18338
rect 8594 18286 8596 18338
rect 8540 18274 8596 18286
rect 8540 12180 8596 12190
rect 8540 12086 8596 12124
rect 8428 9986 8484 9996
rect 8092 8978 8148 8988
rect 7644 8932 7700 8942
rect 7420 8930 7700 8932
rect 7420 8878 7646 8930
rect 7698 8878 7700 8930
rect 7420 8876 7700 8878
rect 7644 8484 7700 8876
rect 7756 8484 7812 8494
rect 7644 8482 7812 8484
rect 7644 8430 7758 8482
rect 7810 8430 7812 8482
rect 7644 8428 7812 8430
rect 5404 8372 5572 8428
rect 7756 8418 7812 8428
rect 8652 8428 8708 23324
rect 8988 23154 9044 23166
rect 8988 23102 8990 23154
rect 9042 23102 9044 23154
rect 8764 23044 8820 23054
rect 8764 22260 8820 22988
rect 8876 22260 8932 22270
rect 8764 22258 8932 22260
rect 8764 22206 8878 22258
rect 8930 22206 8932 22258
rect 8764 22204 8932 22206
rect 8764 13636 8820 22204
rect 8876 22194 8932 22204
rect 8988 21588 9044 23102
rect 8988 20132 9044 21532
rect 9100 21028 9156 26852
rect 9324 26180 9380 26190
rect 9212 26066 9268 26078
rect 9212 26014 9214 26066
rect 9266 26014 9268 26066
rect 9212 24722 9268 26014
rect 9324 25060 9380 26124
rect 9436 25618 9492 29260
rect 9436 25566 9438 25618
rect 9490 25566 9492 25618
rect 9436 25554 9492 25566
rect 9324 25004 9492 25060
rect 9212 24670 9214 24722
rect 9266 24670 9268 24722
rect 9212 24658 9268 24670
rect 9324 24164 9380 24174
rect 9324 24050 9380 24108
rect 9324 23998 9326 24050
rect 9378 23998 9380 24050
rect 9324 23986 9380 23998
rect 9324 23492 9380 23502
rect 9212 22372 9268 22382
rect 9212 22278 9268 22316
rect 9324 22036 9380 23436
rect 9436 23042 9492 25004
rect 9548 24948 9604 32732
rect 9548 24882 9604 24892
rect 9436 22990 9438 23042
rect 9490 22990 9492 23042
rect 9436 22978 9492 22990
rect 9548 24722 9604 24734
rect 9548 24670 9550 24722
rect 9602 24670 9604 24722
rect 9548 22708 9604 24670
rect 9436 22652 9604 22708
rect 9436 22372 9492 22652
rect 9660 22596 9716 35644
rect 9772 35868 9940 35924
rect 9772 32788 9828 35868
rect 9884 35700 9940 35710
rect 9884 35606 9940 35644
rect 9884 33460 9940 33470
rect 9884 33366 9940 33404
rect 9772 32732 9940 32788
rect 9772 30770 9828 30782
rect 9772 30718 9774 30770
rect 9826 30718 9828 30770
rect 9772 30210 9828 30718
rect 9772 30158 9774 30210
rect 9826 30158 9828 30210
rect 9772 30146 9828 30158
rect 9772 29428 9828 29438
rect 9772 27858 9828 29372
rect 9772 27806 9774 27858
rect 9826 27806 9828 27858
rect 9772 27794 9828 27806
rect 9884 24276 9940 32732
rect 10444 32340 10500 40350
rect 11004 39620 11060 39630
rect 11004 39526 11060 39564
rect 10556 38834 10612 38846
rect 10556 38782 10558 38834
rect 10610 38782 10612 38834
rect 10556 38052 10612 38782
rect 10556 37986 10612 37996
rect 11004 38610 11060 38622
rect 11004 38558 11006 38610
rect 11058 38558 11060 38610
rect 10668 37266 10724 37278
rect 10668 37214 10670 37266
rect 10722 37214 10724 37266
rect 10556 36370 10612 36382
rect 10556 36318 10558 36370
rect 10610 36318 10612 36370
rect 10556 35812 10612 36318
rect 10668 36036 10724 37214
rect 10668 35970 10724 35980
rect 10556 35746 10612 35756
rect 11004 35924 11060 38558
rect 11116 38052 11172 38062
rect 11116 37958 11172 37996
rect 10892 35700 10948 35710
rect 10668 35698 10948 35700
rect 10668 35646 10894 35698
rect 10946 35646 10948 35698
rect 10668 35644 10948 35646
rect 10556 34802 10612 34814
rect 10556 34750 10558 34802
rect 10610 34750 10612 34802
rect 10556 32564 10612 34750
rect 10556 32470 10612 32508
rect 10444 32284 10612 32340
rect 10444 30994 10500 31006
rect 10444 30942 10446 30994
rect 10498 30942 10500 30994
rect 10444 30434 10500 30942
rect 10444 30382 10446 30434
rect 10498 30382 10500 30434
rect 10444 30370 10500 30382
rect 10220 30212 10276 30222
rect 10220 29428 10276 30156
rect 10220 29362 10276 29372
rect 10108 29204 10164 29214
rect 10108 29202 10500 29204
rect 10108 29150 10110 29202
rect 10162 29150 10500 29202
rect 10108 29148 10500 29150
rect 10108 29138 10164 29148
rect 10444 27858 10500 29148
rect 10444 27806 10446 27858
rect 10498 27806 10500 27858
rect 10444 27794 10500 27806
rect 9996 27636 10052 27646
rect 9996 27634 10164 27636
rect 9996 27582 9998 27634
rect 10050 27582 10164 27634
rect 9996 27580 10164 27582
rect 9996 27570 10052 27580
rect 10108 27300 10164 27580
rect 10220 27300 10276 27310
rect 10108 27298 10276 27300
rect 10108 27246 10222 27298
rect 10274 27246 10276 27298
rect 10108 27244 10276 27246
rect 10220 27234 10276 27244
rect 10556 26908 10612 32284
rect 9884 24210 9940 24220
rect 10220 26852 10612 26908
rect 9436 22306 9492 22316
rect 9548 22540 9716 22596
rect 9884 23938 9940 23950
rect 9884 23886 9886 23938
rect 9938 23886 9940 23938
rect 9884 22594 9940 23886
rect 9884 22542 9886 22594
rect 9938 22542 9940 22594
rect 9436 22036 9492 22046
rect 9324 21980 9436 22036
rect 9436 21586 9492 21980
rect 9436 21534 9438 21586
rect 9490 21534 9492 21586
rect 9436 21522 9492 21534
rect 9100 20972 9268 21028
rect 8988 20018 9044 20076
rect 8988 19966 8990 20018
rect 9042 19966 9044 20018
rect 8988 18564 9044 19966
rect 8988 18498 9044 18508
rect 9100 16098 9156 16110
rect 9100 16046 9102 16098
rect 9154 16046 9156 16098
rect 9100 15540 9156 16046
rect 9100 15474 9156 15484
rect 9212 14308 9268 20972
rect 9436 20802 9492 20814
rect 9436 20750 9438 20802
rect 9490 20750 9492 20802
rect 9436 20244 9492 20750
rect 9548 20580 9604 22540
rect 9884 22530 9940 22542
rect 9660 22372 9716 22382
rect 9660 21924 9716 22316
rect 9660 20692 9716 21868
rect 9772 22370 9828 22382
rect 9772 22318 9774 22370
rect 9826 22318 9828 22370
rect 9772 21700 9828 22318
rect 9772 21634 9828 21644
rect 10108 21588 10164 21598
rect 10108 21494 10164 21532
rect 9772 21364 9828 21374
rect 9772 21026 9828 21308
rect 9772 20974 9774 21026
rect 9826 20974 9828 21026
rect 9772 20962 9828 20974
rect 9884 20916 9940 20926
rect 9884 20822 9940 20860
rect 9996 20802 10052 20814
rect 9996 20750 9998 20802
rect 10050 20750 10052 20802
rect 9660 20636 9940 20692
rect 9548 20524 9828 20580
rect 9436 20178 9492 20188
rect 9324 19908 9380 19918
rect 9324 16436 9380 19852
rect 9548 19684 9604 19694
rect 9548 19234 9604 19628
rect 9548 19182 9550 19234
rect 9602 19182 9604 19234
rect 9548 19170 9604 19182
rect 9660 18228 9716 18238
rect 9548 18226 9716 18228
rect 9548 18174 9662 18226
rect 9714 18174 9716 18226
rect 9548 18172 9716 18174
rect 9548 16436 9604 18172
rect 9660 18162 9716 18172
rect 9660 17554 9716 17566
rect 9660 17502 9662 17554
rect 9714 17502 9716 17554
rect 9660 16884 9716 17502
rect 9660 16818 9716 16828
rect 9324 16380 9492 16436
rect 9324 16100 9380 16110
rect 9324 16006 9380 16044
rect 9436 15148 9492 16380
rect 9548 16370 9604 16380
rect 9548 16210 9604 16222
rect 9548 16158 9550 16210
rect 9602 16158 9604 16210
rect 9548 15428 9604 16158
rect 9548 15334 9604 15372
rect 9660 15874 9716 15886
rect 9660 15822 9662 15874
rect 9714 15822 9716 15874
rect 9660 15316 9716 15822
rect 9660 15250 9716 15260
rect 8764 13570 8820 13580
rect 8876 14252 9268 14308
rect 9324 15092 9492 15148
rect 8764 12068 8820 12078
rect 8764 10610 8820 12012
rect 8876 11844 8932 14252
rect 9324 14084 9380 15092
rect 9436 14756 9492 14766
rect 9436 14642 9492 14700
rect 9436 14590 9438 14642
rect 9490 14590 9492 14642
rect 9436 14532 9492 14590
rect 9548 14644 9604 14654
rect 9548 14550 9604 14588
rect 9436 14466 9492 14476
rect 9772 14420 9828 20524
rect 9884 17556 9940 20636
rect 9996 19460 10052 20750
rect 9996 19394 10052 19404
rect 10108 20356 10164 20366
rect 9996 17892 10052 17902
rect 9996 17778 10052 17836
rect 9996 17726 9998 17778
rect 10050 17726 10052 17778
rect 9996 17714 10052 17726
rect 9884 17500 10052 17556
rect 9884 16770 9940 16782
rect 9884 16718 9886 16770
rect 9938 16718 9940 16770
rect 9884 16098 9940 16718
rect 9996 16548 10052 17500
rect 10108 16770 10164 20300
rect 10220 19348 10276 26852
rect 10332 25620 10388 25630
rect 10332 25172 10388 25564
rect 10444 25396 10500 25406
rect 10444 25394 10612 25396
rect 10444 25342 10446 25394
rect 10498 25342 10612 25394
rect 10444 25340 10612 25342
rect 10444 25330 10500 25340
rect 10556 25172 10612 25340
rect 10332 25116 10500 25172
rect 10332 22484 10388 22494
rect 10332 22390 10388 22428
rect 10444 21474 10500 25116
rect 10556 23604 10612 25116
rect 10668 25060 10724 35644
rect 10892 35634 10948 35644
rect 11004 35138 11060 35868
rect 11004 35086 11006 35138
rect 11058 35086 11060 35138
rect 11004 35074 11060 35086
rect 11228 36036 11284 36046
rect 11116 33124 11172 33134
rect 10892 33122 11172 33124
rect 10892 33070 11118 33122
rect 11170 33070 11172 33122
rect 10892 33068 11172 33070
rect 10780 31106 10836 31118
rect 10780 31054 10782 31106
rect 10834 31054 10836 31106
rect 10780 30436 10836 31054
rect 10892 30996 10948 33068
rect 11116 33058 11172 33068
rect 11228 32452 11284 35980
rect 11340 35812 11396 43596
rect 12236 42980 12292 42990
rect 12012 41748 12068 41758
rect 11788 40962 11844 40974
rect 11788 40910 11790 40962
rect 11842 40910 11844 40962
rect 11788 39844 11844 40910
rect 11788 39778 11844 39788
rect 11788 39620 11844 39630
rect 11788 39526 11844 39564
rect 11452 39506 11508 39518
rect 11452 39454 11454 39506
rect 11506 39454 11508 39506
rect 11452 38668 11508 39454
rect 11452 38612 11620 38668
rect 11564 37938 11620 38612
rect 11564 37886 11566 37938
rect 11618 37886 11620 37938
rect 11452 35812 11508 35822
rect 11340 35810 11508 35812
rect 11340 35758 11454 35810
rect 11506 35758 11508 35810
rect 11340 35756 11508 35758
rect 11452 35746 11508 35756
rect 11228 32396 11508 32452
rect 11004 32340 11060 32350
rect 11004 32338 11396 32340
rect 11004 32286 11006 32338
rect 11058 32286 11396 32338
rect 11004 32284 11396 32286
rect 11004 32274 11060 32284
rect 10892 30940 11060 30996
rect 10780 30370 10836 30380
rect 11004 30210 11060 30940
rect 11004 30158 11006 30210
rect 11058 30158 11060 30210
rect 11004 30146 11060 30158
rect 11340 30994 11396 32284
rect 11340 30942 11342 30994
rect 11394 30942 11396 30994
rect 11340 29652 11396 30942
rect 11340 29586 11396 29596
rect 11452 30210 11508 32396
rect 11452 30158 11454 30210
rect 11506 30158 11508 30210
rect 11340 29428 11396 29438
rect 11116 28868 11172 28878
rect 10892 28532 10948 28542
rect 10892 27076 10948 28476
rect 11004 27860 11060 27870
rect 11004 27766 11060 27804
rect 10892 27010 10948 27020
rect 10780 26962 10836 26974
rect 10780 26910 10782 26962
rect 10834 26910 10836 26962
rect 10780 25620 10836 26910
rect 10780 25554 10836 25564
rect 10892 25620 10948 25630
rect 11116 25620 11172 28812
rect 11340 28868 11396 29372
rect 11340 28774 11396 28812
rect 11452 27860 11508 30158
rect 11452 27794 11508 27804
rect 11564 27524 11620 37886
rect 11788 38164 11844 38174
rect 11788 37380 11844 38108
rect 11900 38052 11956 38062
rect 11900 37958 11956 37996
rect 11788 37314 11844 37324
rect 11788 36370 11844 36382
rect 11788 36318 11790 36370
rect 11842 36318 11844 36370
rect 11788 35700 11844 36318
rect 11900 35700 11956 35710
rect 11788 35698 11956 35700
rect 11788 35646 11902 35698
rect 11954 35646 11956 35698
rect 11788 35644 11956 35646
rect 11788 33348 11844 33358
rect 11900 33348 11956 35644
rect 12012 35140 12068 41692
rect 12124 38610 12180 38622
rect 12124 38558 12126 38610
rect 12178 38558 12180 38610
rect 12124 38052 12180 38558
rect 12124 37986 12180 37996
rect 12236 36820 12292 42924
rect 13020 42756 13076 42766
rect 12908 40180 12964 40190
rect 12460 40178 12964 40180
rect 12460 40126 12910 40178
rect 12962 40126 12964 40178
rect 12460 40124 12964 40126
rect 12460 39842 12516 40124
rect 12908 40114 12964 40124
rect 12460 39790 12462 39842
rect 12514 39790 12516 39842
rect 12460 39778 12516 39790
rect 12908 39844 12964 39854
rect 12908 39730 12964 39788
rect 12908 39678 12910 39730
rect 12962 39678 12964 39730
rect 12908 39666 12964 39678
rect 12348 39620 12404 39630
rect 12348 39618 12516 39620
rect 12348 39566 12350 39618
rect 12402 39566 12516 39618
rect 12348 39564 12516 39566
rect 12348 39554 12404 39564
rect 12460 38050 12516 39564
rect 12572 39004 12964 39060
rect 12572 38274 12628 39004
rect 12572 38222 12574 38274
rect 12626 38222 12628 38274
rect 12572 38210 12628 38222
rect 12684 38836 12740 38846
rect 12460 37998 12462 38050
rect 12514 37998 12516 38050
rect 12012 35074 12068 35084
rect 12124 36764 12292 36820
rect 12348 37828 12404 37838
rect 12124 34916 12180 36764
rect 12236 36596 12292 36606
rect 12348 36596 12404 37772
rect 12460 37268 12516 37998
rect 12460 37202 12516 37212
rect 12236 36594 12404 36596
rect 12236 36542 12238 36594
rect 12290 36542 12404 36594
rect 12236 36540 12404 36542
rect 12236 36530 12292 36540
rect 11788 33346 11956 33348
rect 11788 33294 11790 33346
rect 11842 33294 11956 33346
rect 11788 33292 11956 33294
rect 12012 34860 12180 34916
rect 11788 32564 11844 33292
rect 11788 32498 11844 32508
rect 12012 32116 12068 34860
rect 12572 34802 12628 34814
rect 12572 34750 12574 34802
rect 12626 34750 12628 34802
rect 12124 34692 12180 34702
rect 12124 34598 12180 34636
rect 12572 34244 12628 34750
rect 12572 34178 12628 34188
rect 12460 34020 12516 34030
rect 12236 33458 12292 33470
rect 12236 33406 12238 33458
rect 12290 33406 12292 33458
rect 12124 32340 12180 32350
rect 12124 32246 12180 32284
rect 12012 32060 12180 32116
rect 12012 31666 12068 31678
rect 12012 31614 12014 31666
rect 12066 31614 12068 31666
rect 11900 31444 11956 31454
rect 11900 31106 11956 31388
rect 11900 31054 11902 31106
rect 11954 31054 11956 31106
rect 11900 31042 11956 31054
rect 12012 31108 12068 31614
rect 12012 31042 12068 31052
rect 11900 30548 11956 30558
rect 11564 27458 11620 27468
rect 11676 29652 11732 29662
rect 10892 25618 11172 25620
rect 10892 25566 10894 25618
rect 10946 25566 11172 25618
rect 10892 25564 11172 25566
rect 11228 27188 11284 27198
rect 10668 24994 10724 25004
rect 10556 23538 10612 23548
rect 10668 24722 10724 24734
rect 10668 24670 10670 24722
rect 10722 24670 10724 24722
rect 10556 23044 10612 23054
rect 10556 22950 10612 22988
rect 10444 21422 10446 21474
rect 10498 21422 10500 21474
rect 10444 21410 10500 21422
rect 10444 20916 10500 20926
rect 10444 20802 10500 20860
rect 10444 20750 10446 20802
rect 10498 20750 10500 20802
rect 10444 20738 10500 20750
rect 10556 20244 10612 20254
rect 10556 20130 10612 20188
rect 10556 20078 10558 20130
rect 10610 20078 10612 20130
rect 10556 20066 10612 20078
rect 10220 19282 10276 19292
rect 10332 19236 10388 19246
rect 10332 19142 10388 19180
rect 10668 18788 10724 24670
rect 10892 24052 10948 25564
rect 10892 23986 10948 23996
rect 11228 24162 11284 27132
rect 11676 27188 11732 29596
rect 11788 29428 11844 29438
rect 11788 29334 11844 29372
rect 11676 27094 11732 27132
rect 11340 26964 11396 27002
rect 11340 26898 11396 26908
rect 11228 24110 11230 24162
rect 11282 24110 11284 24162
rect 10780 23826 10836 23838
rect 10780 23774 10782 23826
rect 10834 23774 10836 23826
rect 10780 23604 10836 23774
rect 11228 23548 11284 24110
rect 10780 23538 10836 23548
rect 11116 23492 11284 23548
rect 11452 26516 11508 26526
rect 10892 22372 10948 22382
rect 10892 22278 10948 22316
rect 11116 22148 11172 23492
rect 11452 23380 11508 26460
rect 11788 26068 11844 26078
rect 11676 23380 11732 23390
rect 10892 22092 11172 22148
rect 11228 23324 11508 23380
rect 11564 23378 11732 23380
rect 11564 23326 11678 23378
rect 11730 23326 11732 23378
rect 11564 23324 11732 23326
rect 10780 20692 10836 20702
rect 10780 20578 10836 20636
rect 10780 20526 10782 20578
rect 10834 20526 10836 20578
rect 10780 20514 10836 20526
rect 10668 18732 10836 18788
rect 10332 18564 10388 18574
rect 10332 17108 10388 18508
rect 10780 18452 10836 18732
rect 10780 18386 10836 18396
rect 10668 18340 10724 18350
rect 10668 18246 10724 18284
rect 10892 17556 10948 22092
rect 11004 20802 11060 20814
rect 11004 20750 11006 20802
rect 11058 20750 11060 20802
rect 11004 18564 11060 20750
rect 11116 20132 11172 20142
rect 11116 19346 11172 20076
rect 11116 19294 11118 19346
rect 11170 19294 11172 19346
rect 11116 19282 11172 19294
rect 11228 19236 11284 23324
rect 11452 23154 11508 23166
rect 11452 23102 11454 23154
rect 11506 23102 11508 23154
rect 11340 21812 11396 21822
rect 11340 20020 11396 21756
rect 11452 21364 11508 23102
rect 11452 21298 11508 21308
rect 11564 21140 11620 23324
rect 11676 23314 11732 23324
rect 11788 23156 11844 26012
rect 11676 23100 11844 23156
rect 11676 22932 11732 23100
rect 11676 22866 11732 22876
rect 11788 22930 11844 22942
rect 11788 22878 11790 22930
rect 11842 22878 11844 22930
rect 11676 21812 11732 21822
rect 11676 21718 11732 21756
rect 11564 21084 11732 21140
rect 11564 20804 11620 20814
rect 11564 20710 11620 20748
rect 11676 20468 11732 21084
rect 11788 20690 11844 22878
rect 11900 22708 11956 30492
rect 12124 29538 12180 32060
rect 12124 29486 12126 29538
rect 12178 29486 12180 29538
rect 12124 29474 12180 29486
rect 12236 29428 12292 33406
rect 12348 32340 12404 32350
rect 12348 31778 12404 32284
rect 12348 31726 12350 31778
rect 12402 31726 12404 31778
rect 12348 31714 12404 31726
rect 12460 30548 12516 33964
rect 12684 31332 12740 38780
rect 12908 38834 12964 39004
rect 12908 38782 12910 38834
rect 12962 38782 12964 38834
rect 12908 38770 12964 38782
rect 12796 38388 12852 38398
rect 12796 32004 12852 38332
rect 12908 35812 12964 35822
rect 13020 35812 13076 42700
rect 13132 38388 13188 44492
rect 13132 38322 13188 38332
rect 13244 38164 13300 50372
rect 13356 40514 13412 40526
rect 13356 40462 13358 40514
rect 13410 40462 13412 40514
rect 13356 39172 13412 40462
rect 13580 39618 13636 39630
rect 13580 39566 13582 39618
rect 13634 39566 13636 39618
rect 13356 39116 13524 39172
rect 13356 38946 13412 38958
rect 13356 38894 13358 38946
rect 13410 38894 13412 38946
rect 13356 38724 13412 38894
rect 13356 38658 13412 38668
rect 13468 38500 13524 39116
rect 13244 38098 13300 38108
rect 13356 38444 13524 38500
rect 13132 38052 13188 38062
rect 13132 37958 13188 37996
rect 13356 37828 13412 38444
rect 12908 35810 13076 35812
rect 12908 35758 12910 35810
rect 12962 35758 13076 35810
rect 12908 35756 13076 35758
rect 13132 37772 13412 37828
rect 13468 38052 13524 38062
rect 12908 35746 12964 35756
rect 12908 34914 12964 34926
rect 12908 34862 12910 34914
rect 12962 34862 12964 34914
rect 12908 34692 12964 34862
rect 12908 34626 12964 34636
rect 12796 31938 12852 31948
rect 12908 33012 12964 33022
rect 12908 31780 12964 32956
rect 13132 32900 13188 37772
rect 13468 37716 13524 37996
rect 13356 37660 13524 37716
rect 13580 38050 13636 39566
rect 13692 38668 13748 50372
rect 13692 38612 14196 38668
rect 13580 37998 13582 38050
rect 13634 37998 13636 38050
rect 13244 37604 13300 37614
rect 13244 35364 13300 37548
rect 13356 37268 13412 37660
rect 13356 37202 13412 37212
rect 13580 37156 13636 37998
rect 13580 37090 13636 37100
rect 13804 37940 13860 37950
rect 13356 36260 13412 36270
rect 13356 36166 13412 36204
rect 13356 35588 13412 35598
rect 13356 35586 13636 35588
rect 13356 35534 13358 35586
rect 13410 35534 13636 35586
rect 13356 35532 13636 35534
rect 13356 35522 13412 35532
rect 13244 35308 13412 35364
rect 13132 32834 13188 32844
rect 13244 35140 13300 35150
rect 13244 32676 13300 35084
rect 13356 34914 13412 35308
rect 13580 35138 13636 35532
rect 13580 35086 13582 35138
rect 13634 35086 13636 35138
rect 13580 35074 13636 35086
rect 13356 34862 13358 34914
rect 13410 34862 13412 34914
rect 13356 33012 13412 34862
rect 13356 32946 13412 32956
rect 13468 33122 13524 33134
rect 13468 33070 13470 33122
rect 13522 33070 13524 33122
rect 13356 32676 13412 32686
rect 13244 32674 13412 32676
rect 13244 32622 13358 32674
rect 13410 32622 13412 32674
rect 13244 32620 13412 32622
rect 13356 32610 13412 32620
rect 13020 32562 13076 32574
rect 13020 32510 13022 32562
rect 13074 32510 13076 32562
rect 13020 32002 13076 32510
rect 13020 31950 13022 32002
rect 13074 31950 13076 32002
rect 13020 31938 13076 31950
rect 13356 32004 13412 32014
rect 12460 30482 12516 30492
rect 12572 31276 12740 31332
rect 12796 31778 12964 31780
rect 12796 31726 12910 31778
rect 12962 31726 12964 31778
rect 12796 31724 12964 31726
rect 12460 30212 12516 30222
rect 12236 29362 12292 29372
rect 12348 30210 12516 30212
rect 12348 30158 12462 30210
rect 12514 30158 12516 30210
rect 12348 30156 12516 30158
rect 12124 27858 12180 27870
rect 12124 27806 12126 27858
rect 12178 27806 12180 27858
rect 12012 25284 12068 25294
rect 12012 25190 12068 25228
rect 12124 24948 12180 27806
rect 12124 24882 12180 24892
rect 12236 24610 12292 24622
rect 12236 24558 12238 24610
rect 12290 24558 12292 24610
rect 12012 24498 12068 24510
rect 12012 24446 12014 24498
rect 12066 24446 12068 24498
rect 12012 23268 12068 24446
rect 12012 23202 12068 23212
rect 12124 24498 12180 24510
rect 12124 24446 12126 24498
rect 12178 24446 12180 24498
rect 12012 23044 12068 23054
rect 12012 22950 12068 22988
rect 11900 22642 11956 22652
rect 11900 22372 11956 22382
rect 11900 22278 11956 22316
rect 12124 22260 12180 24446
rect 12236 23268 12292 24558
rect 12348 24052 12404 30156
rect 12460 30146 12516 30156
rect 12460 28644 12516 28654
rect 12460 28550 12516 28588
rect 12572 26068 12628 31276
rect 12572 26002 12628 26012
rect 12684 30660 12740 30670
rect 12572 25506 12628 25518
rect 12572 25454 12574 25506
rect 12626 25454 12628 25506
rect 12572 25172 12628 25454
rect 12572 25106 12628 25116
rect 12684 24724 12740 30604
rect 12796 26740 12852 31724
rect 12908 31714 12964 31724
rect 12908 28868 12964 28878
rect 12908 28754 12964 28812
rect 12908 28702 12910 28754
rect 12962 28702 12964 28754
rect 12908 28690 12964 28702
rect 13244 28644 13300 28654
rect 13020 28642 13300 28644
rect 13020 28590 13246 28642
rect 13298 28590 13300 28642
rect 13020 28588 13300 28590
rect 12908 27300 12964 27310
rect 13020 27300 13076 28588
rect 13244 28578 13300 28588
rect 13356 27748 13412 31948
rect 13468 31890 13524 33070
rect 13804 32564 13860 37884
rect 13804 32498 13860 32508
rect 13916 36370 13972 36382
rect 13916 36318 13918 36370
rect 13970 36318 13972 36370
rect 13804 32340 13860 32350
rect 13468 31838 13470 31890
rect 13522 31838 13524 31890
rect 13468 31826 13524 31838
rect 13692 32338 13860 32340
rect 13692 32286 13806 32338
rect 13858 32286 13860 32338
rect 13692 32284 13860 32286
rect 13692 31892 13748 32284
rect 13804 32274 13860 32284
rect 13916 32228 13972 36318
rect 14028 36260 14084 36270
rect 14028 35026 14084 36204
rect 14028 34974 14030 35026
rect 14082 34974 14084 35026
rect 14028 34962 14084 34974
rect 13916 32162 13972 32172
rect 14028 34244 14084 34254
rect 14028 32004 14084 34188
rect 13692 31826 13748 31836
rect 13804 31948 14084 32004
rect 13804 30436 13860 31948
rect 13692 30380 13860 30436
rect 14028 31778 14084 31790
rect 14028 31726 14030 31778
rect 14082 31726 14084 31778
rect 13580 29428 13636 29438
rect 13356 27682 13412 27692
rect 13468 29426 13636 29428
rect 13468 29374 13582 29426
rect 13634 29374 13636 29426
rect 13468 29372 13636 29374
rect 12908 27298 13076 27300
rect 12908 27246 12910 27298
rect 12962 27246 13076 27298
rect 12908 27244 13076 27246
rect 12908 27234 12964 27244
rect 13468 27074 13524 29372
rect 13580 29362 13636 29372
rect 13468 27022 13470 27074
rect 13522 27022 13524 27074
rect 12852 26684 12964 26740
rect 12796 26674 12852 26684
rect 12796 26066 12852 26078
rect 12796 26014 12798 26066
rect 12850 26014 12852 26066
rect 12796 25732 12852 26014
rect 12908 25844 12964 26684
rect 13356 26516 13412 26526
rect 13356 26402 13412 26460
rect 13356 26350 13358 26402
rect 13410 26350 13412 26402
rect 13356 26338 13412 26350
rect 13468 26292 13524 27022
rect 13468 26226 13524 26236
rect 13580 28868 13636 28878
rect 13580 27970 13636 28812
rect 13692 28642 13748 30380
rect 14028 30324 14084 31726
rect 14140 30436 14196 38612
rect 14252 35588 14308 50428
rect 14476 42532 14532 42542
rect 14364 36484 14420 36494
rect 14364 36390 14420 36428
rect 14252 35532 14420 35588
rect 14364 32674 14420 35532
rect 14364 32622 14366 32674
rect 14418 32622 14420 32674
rect 14364 32610 14420 32622
rect 14252 32564 14308 32574
rect 14252 31220 14308 32508
rect 14252 31164 14420 31220
rect 14252 30996 14308 31006
rect 14252 30902 14308 30940
rect 14140 30380 14308 30436
rect 13804 30268 14084 30324
rect 13804 28868 13860 30268
rect 14140 30212 14196 30222
rect 13804 28802 13860 28812
rect 13916 30210 14196 30212
rect 13916 30158 14142 30210
rect 14194 30158 14196 30210
rect 13916 30156 14196 30158
rect 13916 28866 13972 30156
rect 14140 30146 14196 30156
rect 14252 29428 14308 30380
rect 13916 28814 13918 28866
rect 13970 28814 13972 28866
rect 13916 28802 13972 28814
rect 14028 29372 14308 29428
rect 13692 28590 13694 28642
rect 13746 28590 13748 28642
rect 13692 28196 13748 28590
rect 14028 28308 14084 29372
rect 14140 29204 14196 29214
rect 14364 29204 14420 31164
rect 14140 29202 14364 29204
rect 14140 29150 14142 29202
rect 14194 29150 14364 29202
rect 14140 29148 14364 29150
rect 14140 29138 14196 29148
rect 14364 29110 14420 29148
rect 14476 28980 14532 42476
rect 14588 39618 14644 39630
rect 14588 39566 14590 39618
rect 14642 39566 14644 39618
rect 14588 38668 14644 39566
rect 14588 38612 14756 38668
rect 14700 38050 14756 38612
rect 15148 38274 15204 52892
rect 16716 52724 16772 52734
rect 16044 52164 16100 52174
rect 15820 48132 15876 48142
rect 15484 40514 15540 40526
rect 15484 40462 15486 40514
rect 15538 40462 15540 40514
rect 15372 40404 15428 40414
rect 15260 38836 15316 38846
rect 15260 38742 15316 38780
rect 15148 38222 15150 38274
rect 15202 38222 15204 38274
rect 15148 38210 15204 38222
rect 14700 37998 14702 38050
rect 14754 37998 14756 38050
rect 14700 36708 14756 37998
rect 14700 36652 14980 36708
rect 14812 36484 14868 36494
rect 14812 36390 14868 36428
rect 14700 34914 14756 34926
rect 14700 34862 14702 34914
rect 14754 34862 14756 34914
rect 14588 33460 14644 33470
rect 14588 33366 14644 33404
rect 14588 31892 14644 31902
rect 14588 30882 14644 31836
rect 14588 30830 14590 30882
rect 14642 30830 14644 30882
rect 14588 30818 14644 30830
rect 14700 30548 14756 34862
rect 14028 28242 14084 28252
rect 14140 28924 14532 28980
rect 14588 30492 14756 30548
rect 14812 32228 14868 32238
rect 13692 28130 13748 28140
rect 13580 27918 13582 27970
rect 13634 27918 13636 27970
rect 12908 25778 12964 25788
rect 12796 25666 12852 25676
rect 13132 25732 13188 25742
rect 13132 25638 13188 25676
rect 12684 24658 12740 24668
rect 13132 25284 13188 25294
rect 12908 24612 12964 24622
rect 12796 24610 12964 24612
rect 12796 24558 12910 24610
rect 12962 24558 12964 24610
rect 12796 24556 12964 24558
rect 12348 23996 12628 24052
rect 12348 23828 12404 23838
rect 12348 23734 12404 23772
rect 12236 23202 12292 23212
rect 12236 23044 12292 23054
rect 12236 23042 12516 23044
rect 12236 22990 12238 23042
rect 12290 22990 12516 23042
rect 12236 22988 12516 22990
rect 12236 22978 12292 22988
rect 12012 22204 12180 22260
rect 12236 22708 12292 22718
rect 11788 20638 11790 20690
rect 11842 20638 11844 20690
rect 11788 20626 11844 20638
rect 11900 20802 11956 20814
rect 11900 20750 11902 20802
rect 11954 20750 11956 20802
rect 11676 20412 11844 20468
rect 11452 20020 11508 20030
rect 11340 20018 11508 20020
rect 11340 19966 11454 20018
rect 11506 19966 11508 20018
rect 11340 19964 11508 19966
rect 11452 19954 11508 19964
rect 11676 19906 11732 19918
rect 11676 19854 11678 19906
rect 11730 19854 11732 19906
rect 11676 19572 11732 19854
rect 11788 19794 11844 20412
rect 11900 20244 11956 20750
rect 12012 20804 12068 22204
rect 12124 21924 12180 21934
rect 12124 21588 12180 21868
rect 12236 21700 12292 22652
rect 12236 21644 12404 21700
rect 12124 21532 12292 21588
rect 12236 21474 12292 21532
rect 12236 21422 12238 21474
rect 12290 21422 12292 21474
rect 12124 21364 12180 21374
rect 12124 21270 12180 21308
rect 12012 20738 12068 20748
rect 12236 20580 12292 21422
rect 12348 21028 12404 21644
rect 12460 21252 12516 22988
rect 12460 21186 12516 21196
rect 12348 20972 12516 21028
rect 12124 20524 12292 20580
rect 12348 20804 12404 20814
rect 11900 20178 11956 20188
rect 12012 20242 12068 20254
rect 12012 20190 12014 20242
rect 12066 20190 12068 20242
rect 12012 20132 12068 20190
rect 12012 20066 12068 20076
rect 12124 19908 12180 20524
rect 12236 20020 12292 20030
rect 12348 20020 12404 20748
rect 12236 20018 12404 20020
rect 12236 19966 12238 20018
rect 12290 19966 12404 20018
rect 12236 19964 12404 19966
rect 12236 19954 12292 19964
rect 12124 19842 12180 19852
rect 11788 19742 11790 19794
rect 11842 19742 11844 19794
rect 11788 19730 11844 19742
rect 11676 19506 11732 19516
rect 12348 19684 12404 19694
rect 11564 19460 11620 19470
rect 11564 19366 11620 19404
rect 11676 19348 11732 19358
rect 11228 19180 11620 19236
rect 11004 18498 11060 18508
rect 11564 18004 11620 19180
rect 10892 17490 10948 17500
rect 11228 17556 11284 17566
rect 11228 17462 11284 17500
rect 10332 17042 10388 17052
rect 10220 16994 10276 17006
rect 10220 16942 10222 16994
rect 10274 16942 10276 16994
rect 10220 16884 10276 16942
rect 10556 16884 10612 16894
rect 10220 16882 10612 16884
rect 10220 16830 10558 16882
rect 10610 16830 10612 16882
rect 10220 16828 10612 16830
rect 10556 16818 10612 16828
rect 10892 16882 10948 16894
rect 10892 16830 10894 16882
rect 10946 16830 10948 16882
rect 10108 16718 10110 16770
rect 10162 16718 10164 16770
rect 10108 16706 10164 16718
rect 9996 16482 10052 16492
rect 10780 16660 10836 16670
rect 10108 16212 10164 16222
rect 10108 16118 10164 16156
rect 10332 16210 10388 16222
rect 10332 16158 10334 16210
rect 10386 16158 10388 16210
rect 9884 16046 9886 16098
rect 9938 16046 9940 16098
rect 9884 15988 9940 16046
rect 9996 16100 10052 16110
rect 9996 16006 10052 16044
rect 9884 15876 9940 15932
rect 9884 15820 10164 15876
rect 10108 15204 10164 15820
rect 10108 15138 10164 15148
rect 10220 15764 10276 15774
rect 10332 15764 10388 16158
rect 10780 16210 10836 16604
rect 10780 16158 10782 16210
rect 10834 16158 10836 16210
rect 10780 16146 10836 16158
rect 10276 15708 10388 15764
rect 10892 15764 10948 16830
rect 11004 16882 11060 16894
rect 11004 16830 11006 16882
rect 11058 16830 11060 16882
rect 11004 15988 11060 16830
rect 11340 16770 11396 16782
rect 11340 16718 11342 16770
rect 11394 16718 11396 16770
rect 11228 16658 11284 16670
rect 11228 16606 11230 16658
rect 11282 16606 11284 16658
rect 11116 16324 11172 16334
rect 11116 16098 11172 16268
rect 11116 16046 11118 16098
rect 11170 16046 11172 16098
rect 11116 16034 11172 16046
rect 11004 15922 11060 15932
rect 9996 15090 10052 15102
rect 9996 15038 9998 15090
rect 10050 15038 10052 15090
rect 9996 14756 10052 15038
rect 9996 14700 10164 14756
rect 10108 14644 10164 14700
rect 10108 14550 10164 14588
rect 10220 14642 10276 15708
rect 10892 15698 10948 15708
rect 11116 15764 11172 15774
rect 11004 15428 11060 15438
rect 11004 15334 11060 15372
rect 10556 15316 10612 15326
rect 11116 15316 11172 15708
rect 11228 15538 11284 16606
rect 11228 15486 11230 15538
rect 11282 15486 11284 15538
rect 11228 15474 11284 15486
rect 11340 15316 11396 16718
rect 11116 15260 11284 15316
rect 10556 15222 10612 15260
rect 10668 15092 10724 15102
rect 10220 14590 10222 14642
rect 10274 14590 10276 14642
rect 10220 14578 10276 14590
rect 10556 15090 10724 15092
rect 10556 15038 10670 15090
rect 10722 15038 10724 15090
rect 10556 15036 10724 15038
rect 9996 14532 10052 14542
rect 9996 14438 10052 14476
rect 9548 14364 9828 14420
rect 9436 14308 9492 14318
rect 9436 14214 9492 14252
rect 9324 14028 9492 14084
rect 9324 13746 9380 13758
rect 9324 13694 9326 13746
rect 9378 13694 9380 13746
rect 9100 12852 9156 12862
rect 9324 12852 9380 13694
rect 9156 12796 9380 12852
rect 9436 13074 9492 14028
rect 9436 13022 9438 13074
rect 9490 13022 9492 13074
rect 9100 12758 9156 12796
rect 9324 12180 9380 12190
rect 9324 12086 9380 12124
rect 8988 12068 9044 12078
rect 8988 11974 9044 12012
rect 8876 11788 9044 11844
rect 8764 10558 8766 10610
rect 8818 10558 8820 10610
rect 8764 10546 8820 10558
rect 8876 9268 8932 9278
rect 8876 9174 8932 9212
rect 8652 8372 8820 8428
rect 3804 7868 4068 7878
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 3804 7802 4068 7812
rect 4464 7084 4728 7094
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4464 7018 4728 7028
rect 3804 6300 4068 6310
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 3804 6234 4068 6244
rect 2268 5906 2884 5908
rect 2268 5854 2270 5906
rect 2322 5854 2884 5906
rect 2268 5852 2884 5854
rect 2268 5842 2324 5852
rect 4464 5516 4728 5526
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4464 5450 4728 5460
rect 1260 5170 1316 5180
rect 3804 4732 4068 4742
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 3804 4666 4068 4676
rect 1484 4452 1540 4462
rect 1484 4358 1540 4396
rect 4464 3948 4728 3958
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4464 3882 4728 3892
rect 3804 3164 4068 3174
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 3804 3098 4068 3108
rect 1148 2706 1204 2716
rect 3388 2772 3444 2782
rect 2044 1428 2100 1438
rect 2044 112 2100 1372
rect 3388 112 3444 2716
rect 4464 2380 4728 2390
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4464 2314 4728 2324
rect 3804 1596 4068 1606
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 3804 1530 4068 1540
rect 5516 1314 5572 8372
rect 8316 8148 8372 8158
rect 8316 8054 8372 8092
rect 5516 1262 5518 1314
rect 5570 1262 5572 1314
rect 5516 1250 5572 1262
rect 7420 1652 7476 1662
rect 6860 1092 6916 1102
rect 6860 998 6916 1036
rect 4956 978 5012 990
rect 6300 980 6356 990
rect 4956 926 4958 978
rect 5010 926 5012 978
rect 4464 812 4728 822
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4464 746 4728 756
rect 4732 196 4788 206
rect 4732 112 4788 140
rect 4956 196 5012 926
rect 4956 130 5012 140
rect 6076 978 6356 980
rect 6076 926 6302 978
rect 6354 926 6356 978
rect 6076 924 6356 926
rect 6076 112 6132 924
rect 6300 914 6356 924
rect 7420 112 7476 1596
rect 8764 112 8820 8372
rect 8988 1652 9044 11788
rect 9436 11284 9492 13022
rect 9436 11218 9492 11228
rect 9548 11060 9604 14364
rect 9772 13860 9828 13870
rect 9772 13636 9828 13804
rect 9548 10994 9604 11004
rect 9660 13634 9828 13636
rect 9660 13582 9774 13634
rect 9826 13582 9828 13634
rect 9660 13580 9828 13582
rect 9660 10612 9716 13580
rect 9772 13570 9828 13580
rect 10108 12964 10164 12974
rect 9772 12178 9828 12190
rect 9772 12126 9774 12178
rect 9826 12126 9828 12178
rect 9772 11844 9828 12126
rect 9996 12068 10052 12078
rect 10108 12068 10164 12908
rect 9996 12066 10164 12068
rect 9996 12014 9998 12066
rect 10050 12014 10164 12066
rect 9996 12012 10164 12014
rect 9996 12002 10052 12012
rect 9772 11778 9828 11788
rect 9884 11956 9940 11966
rect 9884 11506 9940 11900
rect 9884 11454 9886 11506
rect 9938 11454 9940 11506
rect 9884 11442 9940 11454
rect 10108 11844 10164 11854
rect 9660 10546 9716 10556
rect 9884 10610 9940 10622
rect 9884 10558 9886 10610
rect 9938 10558 9940 10610
rect 9548 10388 9604 10398
rect 9548 9154 9604 10332
rect 9884 9828 9940 10558
rect 10108 9938 10164 11788
rect 10556 11620 10612 15036
rect 10668 15026 10724 15036
rect 10780 15092 10836 15102
rect 10780 15090 11172 15092
rect 10780 15038 10782 15090
rect 10834 15038 11172 15090
rect 10780 15036 11172 15038
rect 10780 15026 10836 15036
rect 11116 14754 11172 15036
rect 11116 14702 11118 14754
rect 11170 14702 11172 14754
rect 11116 14690 11172 14702
rect 11228 14754 11284 15260
rect 11340 15250 11396 15260
rect 11452 15314 11508 15326
rect 11452 15262 11454 15314
rect 11506 15262 11508 15314
rect 11452 15148 11508 15262
rect 11228 14702 11230 14754
rect 11282 14702 11284 14754
rect 11228 14690 11284 14702
rect 11340 15092 11508 15148
rect 10668 14532 10724 14542
rect 10668 14530 11172 14532
rect 10668 14478 10670 14530
rect 10722 14478 11172 14530
rect 10668 14476 11172 14478
rect 10668 14466 10724 14476
rect 11116 14420 11172 14476
rect 11340 14420 11396 15092
rect 11116 14364 11396 14420
rect 11004 14308 11060 14318
rect 11004 14214 11060 14252
rect 11004 13524 11060 13534
rect 11004 13522 11508 13524
rect 11004 13470 11006 13522
rect 11058 13470 11508 13522
rect 11004 13468 11508 13470
rect 11004 13458 11060 13468
rect 11340 12964 11396 12974
rect 10892 12962 11396 12964
rect 10892 12910 11342 12962
rect 11394 12910 11396 12962
rect 10892 12908 11396 12910
rect 10668 12738 10724 12750
rect 10668 12686 10670 12738
rect 10722 12686 10724 12738
rect 10668 12178 10724 12686
rect 10668 12126 10670 12178
rect 10722 12126 10724 12178
rect 10668 12114 10724 12126
rect 10556 11554 10612 11564
rect 10780 11844 10836 11854
rect 10220 11396 10276 11406
rect 10220 11302 10276 11340
rect 10780 11394 10836 11788
rect 10892 11618 10948 12908
rect 11340 12898 11396 12908
rect 10892 11566 10894 11618
rect 10946 11566 10948 11618
rect 10892 11554 10948 11566
rect 11228 12178 11284 12190
rect 11228 12126 11230 12178
rect 11282 12126 11284 12178
rect 10780 11342 10782 11394
rect 10834 11342 10836 11394
rect 10780 11330 10836 11342
rect 11228 11396 11284 12126
rect 11228 11330 11284 11340
rect 11452 11394 11508 13468
rect 11564 11844 11620 17948
rect 11676 16212 11732 19292
rect 11788 19234 11844 19246
rect 11788 19182 11790 19234
rect 11842 19182 11844 19234
rect 11788 17220 11844 19182
rect 12236 19236 12292 19246
rect 12236 19142 12292 19180
rect 11900 18340 11956 18350
rect 11900 18246 11956 18284
rect 12348 17668 12404 19628
rect 11788 17154 11844 17164
rect 12124 17666 12404 17668
rect 12124 17614 12350 17666
rect 12402 17614 12404 17666
rect 12124 17612 12404 17614
rect 11788 16882 11844 16894
rect 11788 16830 11790 16882
rect 11842 16830 11844 16882
rect 11788 16322 11844 16830
rect 12124 16660 12180 17612
rect 12348 17602 12404 17612
rect 12236 16996 12292 17006
rect 12460 16996 12516 20972
rect 12572 19684 12628 23996
rect 12796 23826 12852 24556
rect 12908 24546 12964 24556
rect 13132 23938 13188 25228
rect 13132 23886 13134 23938
rect 13186 23886 13188 23938
rect 13132 23874 13188 23886
rect 13244 24948 13300 24958
rect 12796 23774 12798 23826
rect 12850 23774 12852 23826
rect 12796 23044 12852 23774
rect 13132 23154 13188 23166
rect 13132 23102 13134 23154
rect 13186 23102 13188 23154
rect 12796 23042 12964 23044
rect 12796 22990 12798 23042
rect 12850 22990 12964 23042
rect 12796 22988 12964 22990
rect 12796 22978 12852 22988
rect 12796 21812 12852 21822
rect 12684 21810 12852 21812
rect 12684 21758 12798 21810
rect 12850 21758 12852 21810
rect 12684 21756 12852 21758
rect 12684 20804 12740 21756
rect 12796 21746 12852 21756
rect 12908 21588 12964 22988
rect 13020 22370 13076 22382
rect 13020 22318 13022 22370
rect 13074 22318 13076 22370
rect 13020 22148 13076 22318
rect 13020 22082 13076 22092
rect 12684 20738 12740 20748
rect 12796 21532 12964 21588
rect 13132 21812 13188 23102
rect 12796 20580 12852 21532
rect 12908 21364 12964 21374
rect 12908 21270 12964 21308
rect 13020 21252 13076 21262
rect 12908 20690 12964 20702
rect 12908 20638 12910 20690
rect 12962 20638 12964 20690
rect 12908 20580 12964 20638
rect 12572 19618 12628 19628
rect 12684 20524 12964 20580
rect 12572 19348 12628 19358
rect 12572 19254 12628 19292
rect 12236 16994 12516 16996
rect 12236 16942 12238 16994
rect 12290 16942 12516 16994
rect 12236 16940 12516 16942
rect 12236 16930 12292 16940
rect 11788 16270 11790 16322
rect 11842 16270 11844 16322
rect 11788 16258 11844 16270
rect 12012 16604 12124 16660
rect 11676 16098 11732 16156
rect 11676 16046 11678 16098
rect 11730 16046 11732 16098
rect 11676 16034 11732 16046
rect 11900 15540 11956 15550
rect 11900 15446 11956 15484
rect 11788 15204 11844 15242
rect 11788 15138 11844 15148
rect 11900 15204 11956 15214
rect 12012 15204 12068 16604
rect 12124 16594 12180 16604
rect 12236 16436 12292 16446
rect 12236 16210 12292 16380
rect 12236 16158 12238 16210
rect 12290 16158 12292 16210
rect 12236 16146 12292 16158
rect 11900 15202 12012 15204
rect 11900 15150 11902 15202
rect 11954 15150 12012 15202
rect 11900 15148 12012 15150
rect 11900 15138 11956 15148
rect 12012 15138 12068 15148
rect 12684 15148 12740 20524
rect 12908 20132 12964 20142
rect 13020 20132 13076 21196
rect 13132 20244 13188 21756
rect 13244 21364 13300 24892
rect 13356 24724 13412 24734
rect 13356 24630 13412 24668
rect 13580 24164 13636 27918
rect 14028 27860 14084 27870
rect 14028 27766 14084 27804
rect 14028 27300 14084 27310
rect 14140 27300 14196 28924
rect 14364 28644 14420 28654
rect 14364 28550 14420 28588
rect 14588 28532 14644 30492
rect 14588 28466 14644 28476
rect 14700 30098 14756 30110
rect 14700 30046 14702 30098
rect 14754 30046 14756 30098
rect 14028 27298 14196 27300
rect 14028 27246 14030 27298
rect 14082 27246 14196 27298
rect 14028 27244 14196 27246
rect 14028 27234 14084 27244
rect 14028 26066 14084 26078
rect 14028 26014 14030 26066
rect 14082 26014 14084 26066
rect 13468 24108 13636 24164
rect 13692 25060 13748 25070
rect 13692 24722 13748 25004
rect 13692 24670 13694 24722
rect 13746 24670 13748 24722
rect 13468 21364 13524 24108
rect 13692 23940 13748 24670
rect 13916 24612 13972 24622
rect 13916 24518 13972 24556
rect 13804 24164 13860 24174
rect 14028 24164 14084 26014
rect 13804 24162 14084 24164
rect 13804 24110 13806 24162
rect 13858 24110 14084 24162
rect 13804 24108 14084 24110
rect 14140 25732 14196 27244
rect 13804 24098 13860 24108
rect 13692 23938 14084 23940
rect 13692 23886 13694 23938
rect 13746 23886 14084 23938
rect 13692 23884 14084 23886
rect 13692 23874 13748 23884
rect 13804 23268 13860 23278
rect 13692 23154 13748 23166
rect 13692 23102 13694 23154
rect 13746 23102 13748 23154
rect 13692 22372 13748 23102
rect 13804 23042 13860 23212
rect 13804 22990 13806 23042
rect 13858 22990 13860 23042
rect 13804 22978 13860 22990
rect 13580 22148 13636 22158
rect 13580 21924 13636 22092
rect 13580 21586 13636 21868
rect 13692 21700 13748 22316
rect 13916 22370 13972 22382
rect 13916 22318 13918 22370
rect 13970 22318 13972 22370
rect 13916 22260 13972 22318
rect 13916 22194 13972 22204
rect 13804 21700 13860 21710
rect 13692 21644 13804 21700
rect 13580 21534 13582 21586
rect 13634 21534 13636 21586
rect 13580 21522 13636 21534
rect 13468 21308 13636 21364
rect 13244 20916 13300 21308
rect 13244 20850 13300 20860
rect 13356 20804 13412 20814
rect 13356 20710 13412 20748
rect 13132 20188 13412 20244
rect 12908 20130 13076 20132
rect 12908 20078 12910 20130
rect 12962 20078 13076 20130
rect 12908 20076 13076 20078
rect 12908 20066 12964 20076
rect 13244 20018 13300 20030
rect 13244 19966 13246 20018
rect 13298 19966 13300 20018
rect 13020 19908 13076 19918
rect 12908 19124 12964 19134
rect 12796 19122 12964 19124
rect 12796 19070 12910 19122
rect 12962 19070 12964 19122
rect 12796 19068 12964 19070
rect 12796 16098 12852 19068
rect 12908 19058 12964 19068
rect 12908 18564 12964 18574
rect 12908 16994 12964 18508
rect 12908 16942 12910 16994
rect 12962 16942 12964 16994
rect 12908 16930 12964 16942
rect 12908 16772 12964 16782
rect 13020 16772 13076 19852
rect 13244 19684 13300 19966
rect 13244 19618 13300 19628
rect 13356 19908 13412 20188
rect 13468 19908 13524 19918
rect 13356 19906 13524 19908
rect 13356 19854 13470 19906
rect 13522 19854 13524 19906
rect 13356 19852 13524 19854
rect 13132 19348 13188 19358
rect 13132 17106 13188 19292
rect 13356 19236 13412 19852
rect 13468 19842 13524 19852
rect 13356 19142 13412 19180
rect 13132 17054 13134 17106
rect 13186 17054 13188 17106
rect 13132 17042 13188 17054
rect 13244 19124 13300 19134
rect 13244 17666 13300 19068
rect 13244 17614 13246 17666
rect 13298 17614 13300 17666
rect 12908 16770 13076 16772
rect 12908 16718 12910 16770
rect 12962 16718 13076 16770
rect 12908 16716 13076 16718
rect 13132 16884 13188 16894
rect 12908 16706 12964 16716
rect 12796 16046 12798 16098
rect 12850 16046 12852 16098
rect 12796 16034 12852 16046
rect 13020 16098 13076 16110
rect 13020 16046 13022 16098
rect 13074 16046 13076 16098
rect 12684 15092 12964 15148
rect 12012 14644 12068 14654
rect 11900 12852 11956 12862
rect 11900 12758 11956 12796
rect 12012 12178 12068 14588
rect 12684 14532 12740 14542
rect 12236 12964 12292 12974
rect 12236 12870 12292 12908
rect 12012 12126 12014 12178
rect 12066 12126 12068 12178
rect 12012 12114 12068 12126
rect 11564 11778 11620 11788
rect 12124 12068 12180 12078
rect 12684 12068 12740 14476
rect 12796 13076 12852 13086
rect 12796 12982 12852 13020
rect 12796 12068 12852 12078
rect 12684 12066 12852 12068
rect 12684 12014 12798 12066
rect 12850 12014 12852 12066
rect 12684 12012 12852 12014
rect 11452 11342 11454 11394
rect 11506 11342 11508 11394
rect 11452 11330 11508 11342
rect 11676 11620 11732 11630
rect 10108 9886 10110 9938
rect 10162 9886 10164 9938
rect 10108 9874 10164 9886
rect 10220 10612 10276 10622
rect 9884 9762 9940 9772
rect 9548 9102 9550 9154
rect 9602 9102 9604 9154
rect 9548 9090 9604 9102
rect 9884 9380 9940 9390
rect 9660 9044 9716 9054
rect 9660 8258 9716 8988
rect 9884 8930 9940 9324
rect 9884 8878 9886 8930
rect 9938 8878 9940 8930
rect 9884 8866 9940 8878
rect 10220 8428 10276 10556
rect 10444 10610 10500 10622
rect 10444 10558 10446 10610
rect 10498 10558 10500 10610
rect 10444 10388 10500 10558
rect 10892 10612 10948 10622
rect 10892 10498 10948 10556
rect 10892 10446 10894 10498
rect 10946 10446 10948 10498
rect 10892 10434 10948 10446
rect 11228 10612 11284 10622
rect 10444 10322 10500 10332
rect 11116 9940 11172 9950
rect 11004 9938 11172 9940
rect 11004 9886 11118 9938
rect 11170 9886 11172 9938
rect 11004 9884 11172 9886
rect 10444 9826 10500 9838
rect 10444 9774 10446 9826
rect 10498 9774 10500 9826
rect 10444 9268 10500 9774
rect 10892 9826 10948 9838
rect 10892 9774 10894 9826
rect 10946 9774 10948 9826
rect 10892 9604 10948 9774
rect 10892 9538 10948 9548
rect 10444 9202 10500 9212
rect 9660 8206 9662 8258
rect 9714 8206 9716 8258
rect 9660 8194 9716 8206
rect 10108 8372 10276 8428
rect 10108 8370 10164 8372
rect 10108 8318 10110 8370
rect 10162 8318 10164 8370
rect 10108 7474 10164 8318
rect 10668 7700 10724 7710
rect 10668 7586 10724 7644
rect 10668 7534 10670 7586
rect 10722 7534 10724 7586
rect 10668 7522 10724 7534
rect 10108 7422 10110 7474
rect 10162 7422 10164 7474
rect 10108 7410 10164 7422
rect 11004 7474 11060 9884
rect 11116 9874 11172 9884
rect 11116 9268 11172 9278
rect 11228 9268 11284 10556
rect 11116 9266 11284 9268
rect 11116 9214 11118 9266
rect 11170 9214 11284 9266
rect 11116 9212 11284 9214
rect 11564 9826 11620 9838
rect 11564 9774 11566 9826
rect 11618 9774 11620 9826
rect 11116 9202 11172 9212
rect 11564 9156 11620 9774
rect 11340 9100 11620 9156
rect 11340 8482 11396 9100
rect 11340 8430 11342 8482
rect 11394 8430 11396 8482
rect 11340 8418 11396 8430
rect 11676 8428 11732 11564
rect 12012 11396 12068 11406
rect 12012 9940 12068 11340
rect 12124 10834 12180 12012
rect 12124 10782 12126 10834
rect 12178 10782 12180 10834
rect 12124 10770 12180 10782
rect 12012 9874 12068 9884
rect 12348 9940 12404 9950
rect 12348 9826 12404 9884
rect 12348 9774 12350 9826
rect 12402 9774 12404 9826
rect 12348 9762 12404 9774
rect 11004 7422 11006 7474
rect 11058 7422 11060 7474
rect 11004 7410 11060 7422
rect 11452 8372 11732 8428
rect 8988 1586 9044 1596
rect 10108 5236 10164 5246
rect 10108 112 10164 5180
rect 11452 112 11508 8372
rect 11564 7588 11620 7598
rect 11564 7494 11620 7532
rect 12796 7476 12852 12012
rect 12908 11394 12964 15092
rect 13020 14644 13076 16046
rect 13020 14578 13076 14588
rect 13132 13746 13188 16828
rect 13244 14532 13300 17614
rect 13356 18900 13412 18910
rect 13356 16884 13412 18844
rect 13580 18340 13636 21308
rect 13804 20802 13860 21644
rect 13804 20750 13806 20802
rect 13858 20750 13860 20802
rect 13804 20738 13860 20750
rect 13916 20914 13972 20926
rect 13916 20862 13918 20914
rect 13970 20862 13972 20914
rect 13804 20356 13860 20366
rect 13804 19906 13860 20300
rect 13804 19854 13806 19906
rect 13858 19854 13860 19906
rect 13804 19842 13860 19854
rect 13804 19684 13860 19694
rect 13692 19234 13748 19246
rect 13692 19182 13694 19234
rect 13746 19182 13748 19234
rect 13692 18676 13748 19182
rect 13692 18610 13748 18620
rect 13804 18674 13860 19628
rect 13916 19572 13972 20862
rect 14028 19908 14084 23884
rect 14028 19842 14084 19852
rect 13916 19506 13972 19516
rect 14028 19684 14084 19694
rect 13916 19348 13972 19358
rect 13916 19254 13972 19292
rect 13804 18622 13806 18674
rect 13858 18622 13860 18674
rect 13804 18564 13860 18622
rect 13804 18498 13860 18508
rect 14028 18340 14084 19628
rect 13580 18284 13972 18340
rect 13468 18228 13524 18238
rect 13468 18226 13748 18228
rect 13468 18174 13470 18226
rect 13522 18174 13748 18226
rect 13468 18172 13748 18174
rect 13468 18162 13524 18172
rect 13356 16818 13412 16828
rect 13580 16996 13636 17006
rect 13356 15652 13412 15662
rect 13356 15202 13412 15596
rect 13580 15314 13636 16940
rect 13692 16884 13748 18172
rect 13804 16884 13860 16894
rect 13692 16882 13860 16884
rect 13692 16830 13806 16882
rect 13858 16830 13860 16882
rect 13692 16828 13860 16830
rect 13804 16818 13860 16828
rect 13692 16660 13748 16670
rect 13692 15540 13748 16604
rect 13916 16660 13972 18284
rect 14028 17778 14084 18284
rect 14028 17726 14030 17778
rect 14082 17726 14084 17778
rect 14028 17108 14084 17726
rect 14028 16882 14084 17052
rect 14028 16830 14030 16882
rect 14082 16830 14084 16882
rect 14028 16818 14084 16830
rect 13916 16594 13972 16604
rect 13916 16100 13972 16110
rect 13916 16006 13972 16044
rect 13916 15540 13972 15550
rect 13692 15484 13916 15540
rect 13580 15262 13582 15314
rect 13634 15262 13636 15314
rect 13580 15250 13636 15262
rect 13356 15150 13358 15202
rect 13410 15150 13412 15202
rect 13356 15138 13412 15150
rect 13244 14466 13300 14476
rect 13580 15092 13636 15102
rect 13132 13694 13134 13746
rect 13186 13694 13188 13746
rect 13132 13682 13188 13694
rect 13580 13524 13636 15036
rect 13916 14418 13972 15484
rect 14140 14644 14196 25676
rect 14364 28196 14420 28206
rect 14364 27858 14420 28140
rect 14364 27806 14366 27858
rect 14418 27806 14420 27858
rect 14252 25282 14308 25294
rect 14252 25230 14254 25282
rect 14306 25230 14308 25282
rect 14252 24724 14308 25230
rect 14364 24948 14420 27806
rect 14476 27972 14532 27982
rect 14476 26402 14532 27916
rect 14588 27636 14644 27646
rect 14588 27542 14644 27580
rect 14700 27188 14756 30046
rect 14700 27122 14756 27132
rect 14476 26350 14478 26402
rect 14530 26350 14532 26402
rect 14476 26338 14532 26350
rect 14700 25506 14756 25518
rect 14700 25454 14702 25506
rect 14754 25454 14756 25506
rect 14364 24892 14644 24948
rect 14364 24724 14420 24734
rect 14252 24722 14420 24724
rect 14252 24670 14366 24722
rect 14418 24670 14420 24722
rect 14252 24668 14420 24670
rect 14364 24658 14420 24668
rect 14252 23938 14308 23950
rect 14252 23886 14254 23938
rect 14306 23886 14308 23938
rect 14252 23828 14308 23886
rect 14252 23762 14308 23772
rect 14364 23154 14420 23166
rect 14364 23102 14366 23154
rect 14418 23102 14420 23154
rect 14364 23044 14420 23102
rect 14364 20132 14420 22988
rect 14476 22260 14532 22270
rect 14476 21586 14532 22204
rect 14588 21812 14644 24892
rect 14700 24612 14756 25454
rect 14700 24546 14756 24556
rect 14812 24500 14868 32172
rect 14924 31780 14980 36652
rect 15148 36260 15204 36270
rect 15372 36260 15428 40348
rect 15484 38668 15540 40462
rect 15484 38612 15652 38668
rect 15148 36258 15428 36260
rect 15148 36206 15150 36258
rect 15202 36206 15428 36258
rect 15148 36204 15428 36206
rect 15484 38050 15540 38062
rect 15484 37998 15486 38050
rect 15538 37998 15540 38050
rect 15148 34468 15204 36204
rect 15484 35810 15540 37998
rect 15596 37492 15652 38612
rect 15596 37426 15652 37436
rect 15708 36596 15764 36606
rect 15484 35758 15486 35810
rect 15538 35758 15540 35810
rect 15484 35746 15540 35758
rect 15596 36594 15764 36596
rect 15596 36542 15710 36594
rect 15762 36542 15764 36594
rect 15596 36540 15764 36542
rect 15596 34916 15652 36540
rect 15708 36530 15764 36540
rect 15148 34402 15204 34412
rect 15484 34914 15652 34916
rect 15484 34862 15598 34914
rect 15650 34862 15652 34914
rect 15484 34860 15652 34862
rect 15148 33460 15204 33470
rect 15148 33366 15204 33404
rect 15148 32562 15204 32574
rect 15148 32510 15150 32562
rect 15202 32510 15204 32562
rect 14924 31714 14980 31724
rect 15036 31892 15092 31902
rect 15036 31778 15092 31836
rect 15036 31726 15038 31778
rect 15090 31726 15092 31778
rect 15036 31714 15092 31726
rect 15036 31556 15092 31566
rect 15036 30996 15092 31500
rect 15036 30930 15092 30940
rect 15148 31556 15204 32510
rect 15148 29428 15204 31500
rect 15148 29362 15204 29372
rect 15372 31892 15428 31902
rect 15484 31892 15540 34860
rect 15596 34850 15652 34860
rect 15708 34244 15764 34254
rect 15596 33348 15652 33358
rect 15596 32450 15652 33292
rect 15596 32398 15598 32450
rect 15650 32398 15652 32450
rect 15596 32386 15652 32398
rect 15428 31836 15540 31892
rect 15260 29202 15316 29214
rect 15260 29150 15262 29202
rect 15314 29150 15316 29202
rect 14924 28642 14980 28654
rect 14924 28590 14926 28642
rect 14978 28590 14980 28642
rect 14924 28532 14980 28590
rect 14924 27748 14980 28476
rect 14924 27682 14980 27692
rect 15148 27860 15204 27870
rect 15148 27298 15204 27804
rect 15260 27858 15316 29150
rect 15260 27806 15262 27858
rect 15314 27806 15316 27858
rect 15260 27794 15316 27806
rect 15148 27246 15150 27298
rect 15202 27246 15204 27298
rect 15148 27234 15204 27246
rect 15372 26908 15428 31836
rect 15708 30436 15764 34188
rect 15820 31556 15876 48076
rect 15932 36482 15988 36494
rect 15932 36430 15934 36482
rect 15986 36430 15988 36482
rect 15932 35140 15988 36430
rect 15932 35074 15988 35084
rect 16044 33460 16100 52108
rect 16044 33394 16100 33404
rect 16156 46788 16212 46798
rect 15820 31500 16100 31556
rect 15820 31220 15876 31230
rect 15820 31126 15876 31164
rect 15596 30380 15764 30436
rect 15596 29540 15652 30380
rect 15708 30210 15764 30222
rect 15708 30158 15710 30210
rect 15762 30158 15764 30210
rect 15708 29652 15764 30158
rect 16044 30098 16100 31500
rect 16156 31444 16212 46732
rect 16716 43708 16772 52668
rect 16492 43652 16772 43708
rect 17276 48020 17332 48030
rect 16268 41970 16324 41982
rect 16268 41918 16270 41970
rect 16322 41918 16324 41970
rect 16268 37378 16324 41918
rect 16268 37326 16270 37378
rect 16322 37326 16324 37378
rect 16268 37314 16324 37326
rect 16156 31378 16212 31388
rect 16044 30046 16046 30098
rect 16098 30046 16100 30098
rect 16044 30034 16100 30046
rect 15708 29596 16100 29652
rect 15596 29484 15764 29540
rect 15596 27636 15652 27646
rect 15596 27298 15652 27580
rect 15596 27246 15598 27298
rect 15650 27246 15652 27298
rect 15596 27234 15652 27246
rect 15148 26852 15428 26908
rect 15148 25396 15204 26852
rect 15260 25620 15316 25630
rect 15708 25620 15764 29484
rect 15820 29428 15876 29438
rect 15820 29334 15876 29372
rect 16044 29316 16100 29596
rect 16268 29316 16324 29326
rect 16044 29314 16324 29316
rect 16044 29262 16270 29314
rect 16322 29262 16324 29314
rect 16044 29260 16324 29262
rect 16156 28756 16212 28766
rect 16044 28642 16100 28654
rect 16044 28590 16046 28642
rect 16098 28590 16100 28642
rect 15820 27858 15876 27870
rect 15820 27806 15822 27858
rect 15874 27806 15876 27858
rect 15820 27748 15876 27806
rect 15820 27682 15876 27692
rect 15260 25618 15764 25620
rect 15260 25566 15262 25618
rect 15314 25566 15764 25618
rect 15260 25564 15764 25566
rect 15260 25554 15316 25564
rect 15148 25340 15316 25396
rect 14924 24948 14980 24958
rect 14924 24724 14980 24892
rect 14924 24722 15092 24724
rect 14924 24670 14926 24722
rect 14978 24670 15092 24722
rect 14924 24668 15092 24670
rect 14924 24658 14980 24668
rect 14812 24444 14980 24500
rect 14700 23716 14756 23726
rect 14700 22482 14756 23660
rect 14700 22430 14702 22482
rect 14754 22430 14756 22482
rect 14700 22418 14756 22430
rect 14812 23156 14868 23166
rect 14812 21924 14868 23100
rect 14924 22484 14980 24444
rect 15036 23938 15092 24668
rect 15036 23886 15038 23938
rect 15090 23886 15092 23938
rect 15036 23874 15092 23886
rect 15148 22932 15204 22942
rect 15148 22594 15204 22876
rect 15148 22542 15150 22594
rect 15202 22542 15204 22594
rect 15148 22530 15204 22542
rect 14924 22418 14980 22428
rect 15260 22372 15316 25340
rect 15932 24722 15988 24734
rect 15932 24670 15934 24722
rect 15986 24670 15988 24722
rect 15932 23938 15988 24670
rect 15932 23886 15934 23938
rect 15986 23886 15988 23938
rect 15932 23380 15988 23886
rect 15932 23154 15988 23324
rect 15932 23102 15934 23154
rect 15986 23102 15988 23154
rect 15148 22316 15316 22372
rect 15372 22370 15428 22382
rect 15372 22318 15374 22370
rect 15426 22318 15428 22370
rect 14924 21924 14980 21934
rect 14812 21868 14924 21924
rect 14588 21756 14868 21812
rect 14476 21534 14478 21586
rect 14530 21534 14532 21586
rect 14476 21522 14532 21534
rect 14700 21364 14756 21374
rect 14252 19796 14308 19806
rect 14252 17106 14308 19740
rect 14364 19346 14420 20076
rect 14588 20802 14644 20814
rect 14588 20750 14590 20802
rect 14642 20750 14644 20802
rect 14364 19294 14366 19346
rect 14418 19294 14420 19346
rect 14364 19282 14420 19294
rect 14476 19908 14532 19918
rect 14476 18338 14532 19852
rect 14588 19684 14644 20750
rect 14700 20018 14756 21308
rect 14700 19966 14702 20018
rect 14754 19966 14756 20018
rect 14700 19954 14756 19966
rect 14812 21140 14868 21756
rect 14588 19618 14644 19628
rect 14812 19348 14868 21084
rect 14812 19282 14868 19292
rect 14924 20802 14980 21868
rect 14924 20750 14926 20802
rect 14978 20750 14980 20802
rect 14924 19124 14980 20750
rect 15036 20130 15092 20142
rect 15036 20078 15038 20130
rect 15090 20078 15092 20130
rect 15036 19908 15092 20078
rect 15036 19842 15092 19852
rect 15036 19236 15092 19246
rect 15036 19142 15092 19180
rect 14700 19068 14980 19124
rect 14588 18452 14644 18462
rect 14588 18358 14644 18396
rect 14476 18286 14478 18338
rect 14530 18286 14532 18338
rect 14252 17054 14254 17106
rect 14306 17054 14308 17106
rect 14252 17042 14308 17054
rect 14364 18116 14420 18126
rect 14476 18116 14532 18286
rect 14588 18116 14644 18126
rect 14476 18060 14588 18116
rect 14364 16882 14420 18060
rect 14588 18050 14644 18060
rect 14588 17892 14644 17902
rect 14476 17780 14532 17790
rect 14588 17780 14644 17836
rect 14476 17778 14644 17780
rect 14476 17726 14478 17778
rect 14530 17726 14644 17778
rect 14476 17724 14644 17726
rect 14476 17714 14532 17724
rect 14588 17654 14644 17666
rect 14588 17602 14590 17654
rect 14642 17602 14644 17654
rect 14588 17556 14644 17602
rect 14476 17500 14644 17556
rect 14476 17220 14532 17500
rect 14476 17154 14532 17164
rect 14364 16830 14366 16882
rect 14418 16830 14420 16882
rect 14364 16818 14420 16830
rect 14588 16772 14644 16782
rect 14588 16658 14644 16716
rect 14588 16606 14590 16658
rect 14642 16606 14644 16658
rect 14588 16594 14644 16606
rect 14364 16436 14420 16446
rect 14252 14644 14308 14654
rect 13916 14366 13918 14418
rect 13970 14366 13972 14418
rect 13916 14354 13972 14366
rect 14028 14642 14308 14644
rect 14028 14590 14254 14642
rect 14306 14590 14308 14642
rect 14028 14588 14308 14590
rect 14028 14196 14084 14588
rect 14252 14578 14308 14588
rect 13692 14140 14084 14196
rect 13692 13634 13748 14140
rect 13692 13582 13694 13634
rect 13746 13582 13748 13634
rect 13692 13570 13748 13582
rect 13580 13458 13636 13468
rect 14140 13524 14196 13534
rect 13580 12740 13636 12750
rect 12908 11342 12910 11394
rect 12962 11342 12964 11394
rect 12908 8428 12964 11342
rect 13132 12178 13188 12190
rect 13132 12126 13134 12178
rect 13186 12126 13188 12178
rect 13132 10612 13188 12126
rect 13580 12178 13636 12684
rect 13580 12126 13582 12178
rect 13634 12126 13636 12178
rect 13580 11788 13636 12126
rect 13804 11954 13860 11966
rect 13804 11902 13806 11954
rect 13858 11902 13860 11954
rect 13580 11732 13748 11788
rect 13132 10546 13188 10556
rect 13468 11620 13524 11630
rect 13468 10500 13524 11564
rect 13580 10612 13636 10622
rect 13580 10518 13636 10556
rect 13468 10434 13524 10444
rect 13244 9828 13300 9838
rect 13244 9734 13300 9772
rect 13692 8428 13748 11732
rect 13804 10612 13860 11902
rect 14140 11396 14196 13468
rect 14252 12068 14308 12078
rect 14252 11974 14308 12012
rect 14364 11396 14420 16380
rect 14700 15148 14756 19068
rect 14924 18452 14980 18462
rect 15148 18452 15204 22316
rect 15372 21588 15428 22318
rect 15820 22372 15876 22382
rect 15820 22278 15876 22316
rect 15820 21588 15876 21598
rect 15372 21586 15876 21588
rect 15372 21534 15822 21586
rect 15874 21534 15876 21586
rect 15372 21532 15876 21534
rect 15260 21476 15316 21486
rect 15260 21382 15316 21420
rect 15596 20188 15652 21532
rect 15820 21522 15876 21532
rect 15708 21364 15764 21374
rect 15708 21270 15764 21308
rect 15372 20132 15652 20188
rect 15820 20804 15876 20814
rect 15372 18564 15428 20132
rect 15820 20018 15876 20748
rect 15932 20802 15988 23102
rect 16044 23156 16100 28590
rect 16156 27186 16212 28700
rect 16156 27134 16158 27186
rect 16210 27134 16212 27186
rect 16156 27122 16212 27134
rect 16268 26628 16324 29260
rect 16268 26562 16324 26572
rect 16380 27972 16436 27982
rect 16380 27076 16436 27916
rect 16380 26290 16436 27020
rect 16492 26964 16548 43652
rect 16716 39618 16772 39630
rect 16716 39566 16718 39618
rect 16770 39566 16772 39618
rect 16716 38836 16772 39566
rect 16716 38770 16772 38780
rect 17276 38668 17332 47964
rect 17276 38612 17444 38668
rect 16716 38050 16772 38062
rect 16716 37998 16718 38050
rect 16770 37998 16772 38050
rect 16604 37154 16660 37166
rect 16604 37102 16606 37154
rect 16658 37102 16660 37154
rect 16604 34132 16660 37102
rect 16716 34242 16772 37998
rect 17276 37492 17332 37502
rect 17164 36484 17220 36494
rect 17052 36372 17108 36382
rect 17052 35812 17108 36316
rect 17052 35746 17108 35756
rect 16940 35588 16996 35598
rect 16828 35140 16884 35150
rect 16828 35046 16884 35084
rect 16940 34916 16996 35532
rect 16716 34190 16718 34242
rect 16770 34190 16772 34242
rect 16716 34178 16772 34190
rect 16828 34860 16996 34916
rect 16604 34066 16660 34076
rect 16828 33458 16884 34860
rect 16828 33406 16830 33458
rect 16882 33406 16884 33458
rect 16828 33394 16884 33406
rect 16940 33684 16996 33694
rect 16828 32338 16884 32350
rect 16828 32286 16830 32338
rect 16882 32286 16884 32338
rect 16828 31892 16884 32286
rect 16828 31826 16884 31836
rect 16716 31780 16772 31790
rect 16716 31686 16772 31724
rect 16828 31668 16884 31678
rect 16716 30882 16772 30894
rect 16716 30830 16718 30882
rect 16770 30830 16772 30882
rect 16716 29988 16772 30830
rect 16828 30660 16884 31612
rect 16940 30772 16996 33628
rect 17052 31778 17108 31790
rect 17052 31726 17054 31778
rect 17106 31726 17108 31778
rect 17052 31220 17108 31726
rect 17164 31668 17220 36428
rect 17276 32564 17332 37436
rect 17388 33796 17444 38612
rect 17500 38052 17556 38062
rect 17500 37958 17556 37996
rect 17388 33730 17444 33740
rect 17612 33684 17668 54124
rect 18284 53172 18340 55246
rect 19404 55298 19460 55310
rect 19404 55246 19406 55298
rect 19458 55246 19460 55298
rect 18956 54292 19012 54302
rect 18956 54198 19012 54236
rect 18284 53106 18340 53116
rect 17836 51268 17892 51278
rect 17724 40404 17780 40414
rect 17724 40310 17780 40348
rect 17836 38612 17892 51212
rect 19404 43708 19460 55246
rect 19516 54628 19572 54638
rect 19516 54534 19572 54572
rect 19628 53284 19684 55412
rect 20188 55412 20244 56030
rect 20188 55346 20244 55356
rect 21084 55972 21140 55982
rect 20076 55298 20132 55310
rect 20076 55246 20078 55298
rect 20130 55246 20132 55298
rect 19628 53218 19684 53228
rect 19964 53618 20020 53630
rect 19964 53566 19966 53618
rect 20018 53566 20020 53618
rect 19068 43652 19460 43708
rect 19628 53060 19684 53070
rect 17836 38546 17892 38556
rect 17948 42868 18004 42878
rect 17612 33618 17668 33628
rect 17836 36482 17892 36494
rect 17836 36430 17838 36482
rect 17890 36430 17892 36482
rect 17388 33348 17444 33358
rect 17388 33346 17780 33348
rect 17388 33294 17390 33346
rect 17442 33294 17780 33346
rect 17388 33292 17780 33294
rect 17388 33282 17444 33292
rect 17388 33012 17444 33022
rect 17388 32674 17444 32956
rect 17388 32622 17390 32674
rect 17442 32622 17444 32674
rect 17388 32610 17444 32622
rect 17276 31780 17332 32508
rect 17612 32116 17668 32126
rect 17500 31780 17556 31790
rect 17276 31778 17556 31780
rect 17276 31726 17502 31778
rect 17554 31726 17556 31778
rect 17276 31724 17556 31726
rect 17164 31602 17220 31612
rect 17052 31154 17108 31164
rect 17164 30996 17220 31006
rect 17164 30994 17444 30996
rect 17164 30942 17166 30994
rect 17218 30942 17444 30994
rect 17164 30940 17444 30942
rect 17164 30930 17220 30940
rect 17276 30772 17332 30782
rect 16940 30716 17220 30772
rect 16828 30604 16996 30660
rect 16716 29922 16772 29932
rect 16828 30210 16884 30222
rect 16828 30158 16830 30210
rect 16882 30158 16884 30210
rect 16828 29428 16884 30158
rect 16828 29362 16884 29372
rect 16828 29092 16884 29102
rect 16492 26898 16548 26908
rect 16604 27858 16660 27870
rect 16604 27806 16606 27858
rect 16658 27806 16660 27858
rect 16380 26238 16382 26290
rect 16434 26238 16436 26290
rect 16380 26226 16436 26238
rect 16604 24948 16660 27806
rect 16044 23090 16100 23100
rect 16492 24892 16660 24948
rect 16380 22932 16436 22942
rect 16380 22838 16436 22876
rect 16156 22258 16212 22270
rect 16156 22206 16158 22258
rect 16210 22206 16212 22258
rect 16156 21700 16212 22206
rect 16156 21634 16212 21644
rect 16380 21588 16436 21598
rect 16380 21494 16436 21532
rect 15932 20750 15934 20802
rect 15986 20750 15988 20802
rect 15932 20738 15988 20750
rect 16044 20244 16100 20282
rect 16044 20178 16100 20188
rect 15820 19966 15822 20018
rect 15874 19966 15876 20018
rect 15820 19954 15876 19966
rect 16044 20018 16100 20030
rect 16044 19966 16046 20018
rect 16098 19966 16100 20018
rect 15484 19906 15540 19918
rect 15484 19854 15486 19906
rect 15538 19854 15540 19906
rect 15484 19460 15540 19854
rect 15708 19906 15764 19918
rect 15708 19854 15710 19906
rect 15762 19854 15764 19906
rect 15596 19796 15652 19806
rect 15596 19702 15652 19740
rect 15484 19394 15540 19404
rect 15372 18498 15428 18508
rect 14812 18340 14868 18350
rect 14812 17220 14868 18284
rect 14924 17668 14980 18396
rect 15036 18396 15204 18452
rect 15596 18450 15652 18462
rect 15596 18398 15598 18450
rect 15650 18398 15652 18450
rect 15036 18004 15092 18396
rect 15260 18338 15316 18350
rect 15260 18286 15262 18338
rect 15314 18286 15316 18338
rect 15148 18228 15204 18238
rect 15148 18134 15204 18172
rect 15036 17948 15204 18004
rect 15036 17668 15092 17678
rect 14924 17666 15092 17668
rect 14924 17614 15038 17666
rect 15090 17614 15092 17666
rect 14924 17612 15092 17614
rect 14812 17154 14868 17164
rect 15036 16884 15092 17612
rect 15036 16818 15092 16828
rect 14924 16772 14980 16782
rect 14588 15092 14756 15148
rect 14812 16770 14980 16772
rect 14812 16718 14926 16770
rect 14978 16718 14980 16770
rect 14812 16716 14980 16718
rect 14476 13074 14532 13086
rect 14476 13022 14478 13074
rect 14530 13022 14532 13074
rect 14476 11620 14532 13022
rect 14588 12628 14644 15092
rect 14812 14644 14868 16716
rect 14924 16706 14980 16716
rect 15148 15428 15204 17948
rect 15260 17556 15316 18286
rect 15260 17490 15316 17500
rect 15372 18340 15428 18350
rect 15260 16884 15316 16894
rect 15260 16790 15316 16828
rect 15260 16212 15316 16222
rect 15372 16212 15428 18284
rect 15260 16210 15428 16212
rect 15260 16158 15262 16210
rect 15314 16158 15428 16210
rect 15260 16156 15428 16158
rect 15484 17554 15540 17566
rect 15484 17502 15486 17554
rect 15538 17502 15540 17554
rect 15260 16100 15316 16156
rect 15260 16034 15316 16044
rect 15484 16100 15540 17502
rect 15596 17108 15652 18398
rect 15708 18452 15764 19854
rect 16044 19684 16100 19966
rect 16044 19618 16100 19628
rect 15932 19234 15988 19246
rect 15932 19182 15934 19234
rect 15986 19182 15988 19234
rect 15820 18676 15876 18686
rect 15820 18582 15876 18620
rect 15932 18452 15988 19182
rect 16492 19236 16548 24892
rect 16604 24724 16660 24734
rect 16604 24630 16660 24668
rect 16828 23940 16884 29036
rect 16940 26852 16996 30604
rect 16940 26786 16996 26796
rect 16940 26628 16996 26638
rect 16940 26178 16996 26572
rect 17164 26516 17220 30716
rect 17164 26450 17220 26460
rect 16940 26126 16942 26178
rect 16994 26126 16996 26178
rect 16940 25284 16996 26126
rect 16940 25218 16996 25228
rect 16828 23884 16996 23940
rect 16828 23716 16884 23726
rect 16828 23622 16884 23660
rect 16940 23266 16996 23884
rect 16940 23214 16942 23266
rect 16994 23214 16996 23266
rect 16940 23202 16996 23214
rect 16828 22370 16884 22382
rect 16828 22318 16830 22370
rect 16882 22318 16884 22370
rect 16716 22148 16772 22158
rect 16604 22146 16772 22148
rect 16604 22094 16718 22146
rect 16770 22094 16772 22146
rect 16604 22092 16772 22094
rect 16604 19460 16660 22092
rect 16716 22082 16772 22092
rect 16828 22148 16884 22318
rect 16828 22082 16884 22092
rect 16716 21700 16772 21710
rect 16716 21606 16772 21644
rect 17164 21476 17220 21486
rect 17164 21382 17220 21420
rect 16940 21364 16996 21374
rect 16716 20804 16772 20842
rect 16716 20738 16772 20748
rect 16716 20578 16772 20590
rect 16716 20526 16718 20578
rect 16770 20526 16772 20578
rect 16716 20244 16772 20526
rect 16940 20468 16996 21308
rect 17052 20916 17108 20926
rect 17052 20692 17108 20860
rect 17052 20626 17108 20636
rect 16940 20402 16996 20412
rect 16716 20178 16772 20188
rect 16604 19394 16660 19404
rect 16716 19572 16772 19582
rect 16716 19346 16772 19516
rect 16716 19294 16718 19346
rect 16770 19294 16772 19346
rect 16716 19282 16772 19294
rect 16940 19346 16996 19358
rect 16940 19294 16942 19346
rect 16994 19294 16996 19346
rect 16604 19236 16660 19246
rect 16492 19180 16604 19236
rect 15708 18386 15764 18396
rect 15820 18396 15932 18452
rect 15820 18340 15876 18396
rect 15932 18386 15988 18396
rect 16044 18562 16100 18574
rect 16044 18510 16046 18562
rect 16098 18510 16100 18562
rect 15820 18274 15876 18284
rect 16044 18340 16100 18510
rect 16492 18564 16548 18574
rect 16492 18450 16548 18508
rect 16492 18398 16494 18450
rect 16546 18398 16548 18450
rect 16492 18386 16548 18398
rect 16044 18004 16100 18284
rect 16268 18228 16324 18238
rect 15708 17948 16100 18004
rect 16156 18226 16324 18228
rect 16156 18174 16270 18226
rect 16322 18174 16324 18226
rect 16156 18172 16324 18174
rect 15708 17332 15764 17948
rect 16044 17778 16100 17790
rect 16044 17726 16046 17778
rect 16098 17726 16100 17778
rect 16044 17556 16100 17726
rect 16044 17490 16100 17500
rect 16156 17554 16212 18172
rect 16268 18162 16324 18172
rect 16380 18226 16436 18238
rect 16380 18174 16382 18226
rect 16434 18174 16436 18226
rect 16156 17502 16158 17554
rect 16210 17502 16212 17554
rect 16156 17490 16212 17502
rect 15820 17444 15876 17454
rect 15820 17442 15988 17444
rect 15820 17390 15822 17442
rect 15874 17390 15988 17442
rect 15820 17388 15988 17390
rect 15820 17378 15876 17388
rect 15708 17266 15764 17276
rect 15820 17220 15876 17230
rect 15596 17052 15764 17108
rect 15484 16034 15540 16044
rect 15596 16884 15652 16894
rect 15372 15988 15428 15998
rect 15372 15894 15428 15932
rect 15036 15372 15204 15428
rect 15260 15652 15316 15662
rect 15260 15426 15316 15596
rect 15260 15374 15262 15426
rect 15314 15374 15316 15426
rect 14924 15204 14980 15242
rect 14924 15138 14980 15148
rect 15036 14868 15092 15372
rect 15260 15362 15316 15374
rect 15372 15428 15428 15438
rect 15372 15314 15428 15372
rect 15372 15262 15374 15314
rect 15426 15262 15428 15314
rect 15372 15250 15428 15262
rect 15148 15202 15204 15214
rect 15148 15150 15150 15202
rect 15202 15150 15204 15202
rect 15148 15092 15204 15150
rect 15596 15092 15652 16828
rect 15708 16772 15764 17052
rect 15708 16706 15764 16716
rect 15820 16882 15876 17164
rect 15820 16830 15822 16882
rect 15874 16830 15876 16882
rect 15148 15026 15204 15036
rect 15260 15036 15652 15092
rect 15708 16210 15764 16222
rect 15708 16158 15710 16210
rect 15762 16158 15764 16210
rect 15036 14812 15204 14868
rect 14812 14578 14868 14588
rect 14924 14756 14980 14766
rect 14924 14420 14980 14700
rect 14924 14364 15092 14420
rect 14924 13972 14980 13982
rect 14812 13524 14868 13534
rect 14588 12562 14644 12572
rect 14700 13522 14868 13524
rect 14700 13470 14814 13522
rect 14866 13470 14868 13522
rect 14700 13468 14868 13470
rect 14476 11554 14532 11564
rect 14700 11506 14756 13468
rect 14812 13458 14868 13468
rect 14812 13076 14868 13086
rect 14924 13076 14980 13916
rect 14812 13074 14980 13076
rect 14812 13022 14814 13074
rect 14866 13022 14980 13074
rect 14812 13020 14980 13022
rect 14812 13010 14868 13020
rect 14924 12740 14980 12750
rect 14700 11454 14702 11506
rect 14754 11454 14756 11506
rect 14700 11442 14756 11454
rect 14812 12628 14868 12638
rect 14140 11340 14308 11396
rect 14364 11340 14644 11396
rect 14252 11284 14308 11340
rect 14252 11228 14532 11284
rect 14140 11172 14196 11182
rect 14140 11170 14420 11172
rect 14140 11118 14142 11170
rect 14194 11118 14420 11170
rect 14140 11116 14420 11118
rect 14140 11106 14196 11116
rect 14028 10836 14084 10846
rect 14028 10722 14084 10780
rect 14028 10670 14030 10722
rect 14082 10670 14084 10722
rect 14028 10658 14084 10670
rect 13804 10546 13860 10556
rect 14364 10610 14420 11116
rect 14476 11170 14532 11228
rect 14476 11118 14478 11170
rect 14530 11118 14532 11170
rect 14476 11106 14532 11118
rect 14364 10558 14366 10610
rect 14418 10558 14420 10610
rect 14364 10546 14420 10558
rect 12908 8372 13412 8428
rect 12796 7410 12852 7420
rect 12796 5124 12852 5134
rect 12796 112 12852 5068
rect 13356 3444 13412 8372
rect 13580 8372 13748 8428
rect 13580 8036 13636 8372
rect 13580 7970 13636 7980
rect 14588 6020 14644 11340
rect 14812 8428 14868 12572
rect 14924 10722 14980 12684
rect 15036 12180 15092 14364
rect 15148 12852 15204 14812
rect 15260 13636 15316 15036
rect 15708 14980 15764 16158
rect 15484 14924 15764 14980
rect 15484 14754 15540 14924
rect 15484 14702 15486 14754
rect 15538 14702 15540 14754
rect 15484 14690 15540 14702
rect 15708 14532 15764 14924
rect 15820 15202 15876 16830
rect 15932 16770 15988 17388
rect 16380 16996 16436 18174
rect 16380 16930 16436 16940
rect 16492 17108 16548 17118
rect 16492 16882 16548 17052
rect 16492 16830 16494 16882
rect 16546 16830 16548 16882
rect 16492 16818 16548 16830
rect 16604 16884 16660 19180
rect 16828 19122 16884 19134
rect 16828 19070 16830 19122
rect 16882 19070 16884 19122
rect 16828 18676 16884 19070
rect 16828 18610 16884 18620
rect 16940 18452 16996 19294
rect 17052 18564 17108 18574
rect 17052 18470 17108 18508
rect 16828 18396 16996 18452
rect 16828 17556 16884 18396
rect 16940 18226 16996 18238
rect 16940 18174 16942 18226
rect 16994 18174 16996 18226
rect 16940 17892 16996 18174
rect 17164 18228 17220 18238
rect 17164 18134 17220 18172
rect 16940 17826 16996 17836
rect 16828 17490 16884 17500
rect 16604 16818 16660 16828
rect 16940 16884 16996 16894
rect 16940 16790 16996 16828
rect 15932 16718 15934 16770
rect 15986 16718 15988 16770
rect 15932 16706 15988 16718
rect 15932 16098 15988 16110
rect 15932 16046 15934 16098
rect 15986 16046 15988 16098
rect 15932 15652 15988 16046
rect 16268 16098 16324 16110
rect 16268 16046 16270 16098
rect 16322 16046 16324 16098
rect 16044 15876 16100 15886
rect 16044 15782 16100 15820
rect 15932 15586 15988 15596
rect 15820 15150 15822 15202
rect 15874 15150 15876 15202
rect 15820 14756 15876 15150
rect 15932 15202 15988 15214
rect 15932 15150 15934 15202
rect 15986 15150 15988 15202
rect 15932 14868 15988 15150
rect 16044 15204 16100 15214
rect 16044 15110 16100 15148
rect 15932 14812 16212 14868
rect 15820 14690 15876 14700
rect 16044 14644 16100 14654
rect 16044 14550 16100 14588
rect 15708 14466 15764 14476
rect 15932 14530 15988 14542
rect 15932 14478 15934 14530
rect 15986 14478 15988 14530
rect 15932 14420 15988 14478
rect 15932 14354 15988 14364
rect 16156 14084 16212 14812
rect 16268 14754 16324 16046
rect 16828 15876 16884 15886
rect 16380 15874 16884 15876
rect 16380 15822 16830 15874
rect 16882 15822 16884 15874
rect 16380 15820 16884 15822
rect 16380 15428 16436 15820
rect 16828 15810 16884 15820
rect 16380 14868 16436 15372
rect 16940 15204 16996 15214
rect 16828 15148 16940 15204
rect 16492 15092 16548 15102
rect 16492 15090 16772 15092
rect 16492 15038 16494 15090
rect 16546 15038 16772 15090
rect 16492 15036 16772 15038
rect 16492 15026 16548 15036
rect 16380 14812 16548 14868
rect 16268 14702 16270 14754
rect 16322 14702 16324 14754
rect 16268 14690 16324 14702
rect 16492 14420 16548 14812
rect 16716 14530 16772 15036
rect 16716 14478 16718 14530
rect 16770 14478 16772 14530
rect 16716 14466 16772 14478
rect 16380 14308 16436 14318
rect 16156 14028 16324 14084
rect 15372 13972 15428 13982
rect 15372 13970 16212 13972
rect 15372 13918 15374 13970
rect 15426 13918 16212 13970
rect 15372 13916 16212 13918
rect 15372 13906 15428 13916
rect 15708 13748 15764 13758
rect 15260 13570 15316 13580
rect 15372 13746 15764 13748
rect 15372 13694 15710 13746
rect 15762 13694 15764 13746
rect 15372 13692 15764 13694
rect 15260 13412 15316 13422
rect 15260 13074 15316 13356
rect 15372 13186 15428 13692
rect 15708 13682 15764 13692
rect 16044 13748 16100 13758
rect 16044 13654 16100 13692
rect 16156 13746 16212 13916
rect 16156 13694 16158 13746
rect 16210 13694 16212 13746
rect 16156 13682 16212 13694
rect 15372 13134 15374 13186
rect 15426 13134 15428 13186
rect 15372 13122 15428 13134
rect 15820 13636 15876 13646
rect 15260 13022 15262 13074
rect 15314 13022 15316 13074
rect 15260 12964 15316 13022
rect 15484 12964 15540 12974
rect 15260 12908 15428 12964
rect 15148 12796 15316 12852
rect 15036 12086 15092 12124
rect 14924 10670 14926 10722
rect 14978 10670 14980 10722
rect 14924 10658 14980 10670
rect 15148 11506 15204 11518
rect 15148 11454 15150 11506
rect 15202 11454 15204 11506
rect 15148 9828 15204 11454
rect 15148 9268 15204 9772
rect 15148 9202 15204 9212
rect 14588 5954 14644 5964
rect 14700 8372 14868 8428
rect 15148 9044 15204 9054
rect 14700 4452 14756 8372
rect 15148 5796 15204 8988
rect 15260 8428 15316 12796
rect 15372 9044 15428 12908
rect 15484 12870 15540 12908
rect 15372 8978 15428 8988
rect 15820 12178 15876 13580
rect 16044 13188 16100 13198
rect 16268 13188 16324 14028
rect 16380 13858 16436 14252
rect 16380 13806 16382 13858
rect 16434 13806 16436 13858
rect 16380 13794 16436 13806
rect 16492 13748 16548 14364
rect 16828 13748 16884 15148
rect 16940 15110 16996 15148
rect 17164 14532 17220 14542
rect 17164 14438 17220 14476
rect 17052 14420 17108 14430
rect 16940 14308 16996 14318
rect 16940 14214 16996 14252
rect 17052 13972 17108 14364
rect 17276 14196 17332 30716
rect 17388 30548 17444 30940
rect 17500 30994 17556 31724
rect 17500 30942 17502 30994
rect 17554 30942 17556 30994
rect 17500 30930 17556 30942
rect 17388 30492 17556 30548
rect 17388 30322 17444 30334
rect 17388 30270 17390 30322
rect 17442 30270 17444 30322
rect 17388 27076 17444 30270
rect 17500 29650 17556 30492
rect 17500 29598 17502 29650
rect 17554 29598 17556 29650
rect 17500 29586 17556 29598
rect 17612 29652 17668 32060
rect 17724 32002 17780 33292
rect 17836 33236 17892 36430
rect 17948 35140 18004 42812
rect 18396 41858 18452 41870
rect 18396 41806 18398 41858
rect 18450 41806 18452 41858
rect 18396 40402 18452 41806
rect 18396 40350 18398 40402
rect 18450 40350 18452 40402
rect 18396 40338 18452 40350
rect 18844 39844 18900 39854
rect 18732 39508 18788 39518
rect 18396 39506 18788 39508
rect 18396 39454 18734 39506
rect 18786 39454 18788 39506
rect 18396 39452 18788 39454
rect 17948 35046 18004 35084
rect 18172 38276 18228 38286
rect 18060 35026 18116 35038
rect 18060 34974 18062 35026
rect 18114 34974 18116 35026
rect 17948 33236 18004 33246
rect 17836 33234 18004 33236
rect 17836 33182 17950 33234
rect 18002 33182 18004 33234
rect 17836 33180 18004 33182
rect 17724 31950 17726 32002
rect 17778 31950 17780 32002
rect 17724 31938 17780 31950
rect 17836 32338 17892 32350
rect 17836 32286 17838 32338
rect 17890 32286 17892 32338
rect 17724 30884 17780 30894
rect 17836 30884 17892 32286
rect 17724 30882 17892 30884
rect 17724 30830 17726 30882
rect 17778 30830 17892 30882
rect 17724 30828 17892 30830
rect 17724 30818 17780 30828
rect 17948 30772 18004 33180
rect 17948 30706 18004 30716
rect 18060 29652 18116 34974
rect 18172 33460 18228 38220
rect 18284 36482 18340 36494
rect 18284 36430 18286 36482
rect 18338 36430 18340 36482
rect 18284 36372 18340 36430
rect 18284 34804 18340 36316
rect 18396 35698 18452 39452
rect 18732 39442 18788 39452
rect 18620 38722 18676 38734
rect 18620 38670 18622 38722
rect 18674 38670 18676 38722
rect 18620 37266 18676 38670
rect 18620 37214 18622 37266
rect 18674 37214 18676 37266
rect 18620 37202 18676 37214
rect 18844 36594 18900 39788
rect 18844 36542 18846 36594
rect 18898 36542 18900 36594
rect 18844 36530 18900 36542
rect 18396 35646 18398 35698
rect 18450 35646 18452 35698
rect 18396 35634 18452 35646
rect 18956 34914 19012 34926
rect 18956 34862 18958 34914
rect 19010 34862 19012 34914
rect 18396 34804 18452 34814
rect 18284 34802 18452 34804
rect 18284 34750 18398 34802
rect 18450 34750 18452 34802
rect 18284 34748 18452 34750
rect 18284 33460 18340 33470
rect 18172 33458 18340 33460
rect 18172 33406 18286 33458
rect 18338 33406 18340 33458
rect 18172 33404 18340 33406
rect 18172 32116 18228 33404
rect 18284 33394 18340 33404
rect 18284 32788 18340 32798
rect 18284 32694 18340 32732
rect 18396 32564 18452 34748
rect 18508 34132 18564 34142
rect 18508 34038 18564 34076
rect 18956 32788 19012 34862
rect 18956 32722 19012 32732
rect 18172 32050 18228 32060
rect 18284 32508 18452 32564
rect 18620 32564 18676 32574
rect 19068 32564 19124 43652
rect 18172 31892 18228 31902
rect 18172 31798 18228 31836
rect 18060 29596 18228 29652
rect 17612 29586 17668 29596
rect 18060 29428 18116 29438
rect 17500 29426 18116 29428
rect 17500 29374 18062 29426
rect 18114 29374 18116 29426
rect 17500 29372 18116 29374
rect 17500 27972 17556 29372
rect 18060 29362 18116 29372
rect 17500 27878 17556 27916
rect 17724 29204 17780 29214
rect 18172 29204 18228 29596
rect 17388 27010 17444 27020
rect 17500 27636 17556 27646
rect 17388 26852 17444 26862
rect 17388 23604 17444 26796
rect 17388 23538 17444 23548
rect 17500 25394 17556 27580
rect 17500 25342 17502 25394
rect 17554 25342 17556 25394
rect 17388 22930 17444 22942
rect 17388 22878 17390 22930
rect 17442 22878 17444 22930
rect 17388 22372 17444 22878
rect 17388 22306 17444 22316
rect 17388 22146 17444 22158
rect 17388 22094 17390 22146
rect 17442 22094 17444 22146
rect 17388 20804 17444 22094
rect 17388 20738 17444 20748
rect 17388 18340 17444 18350
rect 17388 18246 17444 18284
rect 17500 17668 17556 25342
rect 17612 26964 17668 26974
rect 17612 24276 17668 26908
rect 17724 26908 17780 29148
rect 17948 29148 18228 29204
rect 17836 27972 17892 27982
rect 17836 27074 17892 27916
rect 17948 27746 18004 29148
rect 17948 27694 17950 27746
rect 18002 27694 18004 27746
rect 17948 27412 18004 27694
rect 18284 27412 18340 32508
rect 18620 32470 18676 32508
rect 18844 32508 19124 32564
rect 19292 40516 19348 40526
rect 18396 30996 18452 31006
rect 18732 30996 18788 31006
rect 18396 30994 18564 30996
rect 18396 30942 18398 30994
rect 18450 30942 18564 30994
rect 18396 30940 18564 30942
rect 18396 30930 18452 30940
rect 18508 30210 18564 30940
rect 18508 30158 18510 30210
rect 18562 30158 18564 30210
rect 18508 30146 18564 30158
rect 18620 30994 18788 30996
rect 18620 30942 18734 30994
rect 18786 30942 18788 30994
rect 18620 30940 18788 30942
rect 18620 29988 18676 30940
rect 18732 30930 18788 30940
rect 18844 30772 18900 32508
rect 19180 32452 19236 32462
rect 19180 32358 19236 32396
rect 18396 29932 18676 29988
rect 18732 30716 18900 30772
rect 18956 31778 19012 31790
rect 18956 31726 18958 31778
rect 19010 31726 19012 31778
rect 18396 28754 18452 29932
rect 18396 28702 18398 28754
rect 18450 28702 18452 28754
rect 18396 27636 18452 28702
rect 18396 27570 18452 27580
rect 18508 29652 18564 29662
rect 18508 29314 18564 29596
rect 18508 29262 18510 29314
rect 18562 29262 18564 29314
rect 17948 27356 18228 27412
rect 18284 27356 18452 27412
rect 17836 27022 17838 27074
rect 17890 27022 17892 27074
rect 17836 27010 17892 27022
rect 18060 27076 18116 27086
rect 17724 26796 17892 26908
rect 17724 24612 17780 26796
rect 18060 26292 18116 27020
rect 17724 24518 17780 24556
rect 17836 26236 18116 26292
rect 17612 24220 17780 24276
rect 17612 21588 17668 21598
rect 17612 21026 17668 21532
rect 17724 21252 17780 24220
rect 17724 21186 17780 21196
rect 17612 20974 17614 21026
rect 17666 20974 17668 21026
rect 17612 20962 17668 20974
rect 17724 20916 17780 20926
rect 17724 18228 17780 20860
rect 17836 20132 17892 26236
rect 18060 26066 18116 26078
rect 18060 26014 18062 26066
rect 18114 26014 18116 26066
rect 17948 25508 18004 25518
rect 18060 25508 18116 26014
rect 17948 25506 18116 25508
rect 17948 25454 17950 25506
rect 18002 25454 18116 25506
rect 17948 25452 18116 25454
rect 17948 25442 18004 25452
rect 17948 25284 18004 25294
rect 18172 25284 18228 27356
rect 18284 27186 18340 27198
rect 18284 27134 18286 27186
rect 18338 27134 18340 27186
rect 18284 26852 18340 27134
rect 18396 27076 18452 27356
rect 18396 27010 18452 27020
rect 18284 26786 18340 26796
rect 18284 26516 18340 26526
rect 18284 25506 18340 26460
rect 18508 26292 18564 29262
rect 18508 25844 18564 26236
rect 18620 28980 18676 28990
rect 18620 25956 18676 28924
rect 18732 26068 18788 30716
rect 18956 28868 19012 31726
rect 18956 28802 19012 28812
rect 19180 31780 19236 31790
rect 18844 28644 18900 28654
rect 18844 28642 19124 28644
rect 18844 28590 18846 28642
rect 18898 28590 19124 28642
rect 18844 28588 19124 28590
rect 18844 28578 18900 28588
rect 19068 28082 19124 28588
rect 19068 28030 19070 28082
rect 19122 28030 19124 28082
rect 19068 28018 19124 28030
rect 19180 28642 19236 31724
rect 19180 28590 19182 28642
rect 19234 28590 19236 28642
rect 19180 26516 19236 28590
rect 19180 26450 19236 26460
rect 19180 26292 19236 26302
rect 19180 26198 19236 26236
rect 18732 26012 19124 26068
rect 18620 25900 18900 25956
rect 18284 25454 18286 25506
rect 18338 25454 18340 25506
rect 18284 25442 18340 25454
rect 18396 25788 18564 25844
rect 18396 25396 18452 25788
rect 18508 25620 18564 25630
rect 18508 25618 18788 25620
rect 18508 25566 18510 25618
rect 18562 25566 18788 25618
rect 18508 25564 18788 25566
rect 18508 25554 18564 25564
rect 18396 25340 18676 25396
rect 18172 25228 18340 25284
rect 17948 24162 18004 25228
rect 18060 25172 18116 25182
rect 18060 24836 18116 25116
rect 18172 24836 18228 24846
rect 18060 24834 18228 24836
rect 18060 24782 18174 24834
rect 18226 24782 18228 24834
rect 18060 24780 18228 24782
rect 17948 24110 17950 24162
rect 18002 24110 18004 24162
rect 17948 24098 18004 24110
rect 18060 24612 18116 24622
rect 18060 23940 18116 24556
rect 17948 23884 18116 23940
rect 18172 23940 18228 24780
rect 17948 20916 18004 23884
rect 18172 23874 18228 23884
rect 18284 21476 18340 25228
rect 18508 24388 18564 24398
rect 18396 23940 18452 23950
rect 18396 23846 18452 23884
rect 18508 23828 18564 24332
rect 18508 23762 18564 23772
rect 18508 23604 18564 23614
rect 18508 22932 18564 23548
rect 17948 20850 18004 20860
rect 18060 21474 18340 21476
rect 18060 21422 18286 21474
rect 18338 21422 18340 21474
rect 18060 21420 18340 21422
rect 17836 18900 17892 20076
rect 17836 18834 17892 18844
rect 17948 18340 18004 18350
rect 17836 18228 17892 18238
rect 17724 18172 17836 18228
rect 17500 17602 17556 17612
rect 17836 16324 17892 18172
rect 17948 16882 18004 18284
rect 17948 16830 17950 16882
rect 18002 16830 18004 16882
rect 17948 16818 18004 16830
rect 17948 16324 18004 16334
rect 17836 16322 18004 16324
rect 17836 16270 17950 16322
rect 18002 16270 18004 16322
rect 17836 16268 18004 16270
rect 17948 16258 18004 16268
rect 17724 15988 17780 15998
rect 17612 15876 17668 15886
rect 17612 14754 17668 15820
rect 17612 14702 17614 14754
rect 17666 14702 17668 14754
rect 17612 14690 17668 14702
rect 17052 13906 17108 13916
rect 17164 14140 17332 14196
rect 17388 14530 17444 14542
rect 17388 14478 17390 14530
rect 17442 14478 17444 14530
rect 16492 13746 16772 13748
rect 16492 13694 16494 13746
rect 16546 13694 16772 13746
rect 16492 13692 16772 13694
rect 16492 13188 16548 13692
rect 16716 13524 16772 13692
rect 16828 13654 16884 13692
rect 17052 13746 17108 13758
rect 17052 13694 17054 13746
rect 17106 13694 17108 13746
rect 17052 13524 17108 13694
rect 16716 13468 17108 13524
rect 16044 13186 16324 13188
rect 16044 13134 16046 13186
rect 16098 13134 16324 13186
rect 16044 13132 16324 13134
rect 16380 13132 16548 13188
rect 16044 13122 16100 13132
rect 16380 13076 16436 13132
rect 16156 13020 16436 13076
rect 16156 12964 16212 13020
rect 16156 12870 16212 12908
rect 15820 12126 15822 12178
rect 15874 12126 15876 12178
rect 15260 8372 15540 8428
rect 15148 5730 15204 5740
rect 14700 4386 14756 4396
rect 13356 3378 13412 3388
rect 15484 1204 15540 8372
rect 15820 6580 15876 12126
rect 15820 6514 15876 6524
rect 15484 1138 15540 1148
rect 16828 4228 16884 4238
rect 14140 980 14196 990
rect 14140 112 14196 924
rect 15484 644 15540 654
rect 15484 112 15540 588
rect 16828 112 16884 4172
rect 17164 1092 17220 14140
rect 17388 13970 17444 14478
rect 17500 14420 17556 14430
rect 17500 14326 17556 14364
rect 17724 14084 17780 15932
rect 18060 15202 18116 21420
rect 18284 21410 18340 21420
rect 18396 22930 18564 22932
rect 18396 22878 18510 22930
rect 18562 22878 18564 22930
rect 18396 22876 18564 22878
rect 18396 21364 18452 22876
rect 18508 22866 18564 22876
rect 18396 21298 18452 21308
rect 18620 22482 18676 25340
rect 18732 24724 18788 25564
rect 18732 24658 18788 24668
rect 18620 22430 18622 22482
rect 18674 22430 18676 22482
rect 18284 21252 18340 21262
rect 18172 20132 18228 20142
rect 18172 20038 18228 20076
rect 18060 15150 18062 15202
rect 18114 15150 18116 15202
rect 18060 15138 18116 15150
rect 17388 13918 17390 13970
rect 17442 13918 17444 13970
rect 17388 13906 17444 13918
rect 17500 14028 17780 14084
rect 17276 13748 17332 13758
rect 17500 13748 17556 14028
rect 17276 13746 17556 13748
rect 17276 13694 17278 13746
rect 17330 13694 17556 13746
rect 17276 13692 17556 13694
rect 17276 13682 17332 13692
rect 18284 8428 18340 21196
rect 18620 21028 18676 22430
rect 18732 23940 18788 23950
rect 18732 21698 18788 23884
rect 18732 21646 18734 21698
rect 18786 21646 18788 21698
rect 18732 21634 18788 21646
rect 18732 21028 18788 21038
rect 18620 21026 18788 21028
rect 18620 20974 18734 21026
rect 18786 20974 18788 21026
rect 18620 20972 18788 20974
rect 18732 20962 18788 20972
rect 18396 20692 18452 20702
rect 18396 16212 18452 20636
rect 18620 19794 18676 19806
rect 18620 19742 18622 19794
rect 18674 19742 18676 19794
rect 18620 18228 18676 19742
rect 18620 18162 18676 18172
rect 18396 16156 18564 16212
rect 18396 15988 18452 15998
rect 18396 15894 18452 15932
rect 18508 15764 18564 16156
rect 18396 15708 18564 15764
rect 18620 15988 18676 15998
rect 18396 13972 18452 15708
rect 18620 15540 18676 15932
rect 18620 15314 18676 15484
rect 18620 15262 18622 15314
rect 18674 15262 18676 15314
rect 18620 15250 18676 15262
rect 18396 13906 18452 13916
rect 18844 8428 18900 25900
rect 19068 25284 19124 26012
rect 19180 25508 19236 25518
rect 19180 25414 19236 25452
rect 19068 25228 19236 25284
rect 18956 24724 19012 24734
rect 18956 24630 19012 24668
rect 18956 23940 19012 23950
rect 18956 23266 19012 23884
rect 18956 23214 18958 23266
rect 19010 23214 19012 23266
rect 18956 20692 19012 23214
rect 18956 20626 19012 20636
rect 19068 22370 19124 22382
rect 19068 22318 19070 22370
rect 19122 22318 19124 22370
rect 18956 18228 19012 18238
rect 18956 18134 19012 18172
rect 19068 15988 19124 22318
rect 19180 20916 19236 25228
rect 19292 23716 19348 40460
rect 19628 38668 19684 53004
rect 19964 52612 20020 53566
rect 19964 52546 20020 52556
rect 20076 49476 20132 55246
rect 20524 55300 20580 55310
rect 20524 55206 20580 55244
rect 20748 55300 20804 55310
rect 20636 54290 20692 54302
rect 20636 54238 20638 54290
rect 20690 54238 20692 54290
rect 20636 54068 20692 54238
rect 20636 54002 20692 54012
rect 20524 53732 20580 53742
rect 20524 53638 20580 53676
rect 19964 49420 20132 49476
rect 19852 46900 19908 46910
rect 19852 45444 19908 46844
rect 19852 45378 19908 45388
rect 19404 38612 19684 38668
rect 19404 32788 19460 38612
rect 19740 37940 19796 37950
rect 19740 37846 19796 37884
rect 19852 35140 19908 35150
rect 19852 35046 19908 35084
rect 19516 34802 19572 34814
rect 19516 34750 19518 34802
rect 19570 34750 19572 34802
rect 19516 33460 19572 34750
rect 19516 33404 19796 33460
rect 19516 33124 19572 33134
rect 19516 33030 19572 33068
rect 19404 32732 19684 32788
rect 19404 32564 19460 32574
rect 19404 32470 19460 32508
rect 19404 28754 19460 28766
rect 19404 28702 19406 28754
rect 19458 28702 19460 28754
rect 19404 27860 19460 28702
rect 19516 27860 19572 27870
rect 19404 27858 19572 27860
rect 19404 27806 19518 27858
rect 19570 27806 19572 27858
rect 19404 27804 19572 27806
rect 19516 27794 19572 27804
rect 19404 26850 19460 26862
rect 19404 26798 19406 26850
rect 19458 26798 19460 26850
rect 19404 25508 19460 26798
rect 19404 25442 19460 25452
rect 19516 26068 19572 26078
rect 19516 24834 19572 26012
rect 19516 24782 19518 24834
rect 19570 24782 19572 24834
rect 19516 24770 19572 24782
rect 19516 23938 19572 23950
rect 19516 23886 19518 23938
rect 19570 23886 19572 23938
rect 19292 23660 19460 23716
rect 19292 21476 19348 21486
rect 19292 21382 19348 21420
rect 19404 21252 19460 23660
rect 19516 23604 19572 23886
rect 19516 23538 19572 23548
rect 19180 20850 19236 20860
rect 19292 21196 19460 21252
rect 19180 20692 19236 20702
rect 19180 20598 19236 20636
rect 19068 15922 19124 15932
rect 17164 1026 17220 1036
rect 18172 8372 18340 8428
rect 18620 8372 18900 8428
rect 18172 112 18228 8372
rect 18620 1092 18676 8372
rect 19292 7588 19348 21196
rect 19404 20916 19460 20926
rect 19404 8428 19460 20860
rect 19516 18452 19572 18462
rect 19516 18358 19572 18396
rect 19404 8372 19572 8428
rect 19292 7522 19348 7532
rect 18620 1026 18676 1036
rect 19516 112 19572 8372
rect 19628 5124 19684 32732
rect 19740 30100 19796 33404
rect 19740 30034 19796 30044
rect 19852 32452 19908 32462
rect 19852 31778 19908 32396
rect 19852 31726 19854 31778
rect 19906 31726 19908 31778
rect 19852 30994 19908 31726
rect 19852 30942 19854 30994
rect 19906 30942 19908 30994
rect 19740 29202 19796 29214
rect 19740 29150 19742 29202
rect 19794 29150 19796 29202
rect 19740 28756 19796 29150
rect 19852 28980 19908 30942
rect 19852 28914 19908 28924
rect 19852 28756 19908 28766
rect 19740 28754 19908 28756
rect 19740 28702 19854 28754
rect 19906 28702 19908 28754
rect 19740 28700 19908 28702
rect 19852 28690 19908 28700
rect 19964 28532 20020 49420
rect 20300 48692 20356 48702
rect 19740 28476 20020 28532
rect 20076 45444 20132 45454
rect 19740 26404 19796 28476
rect 20076 28308 20132 45388
rect 19964 28252 20132 28308
rect 19964 26908 20020 28252
rect 20076 28084 20132 28094
rect 20076 27970 20132 28028
rect 20076 27918 20078 27970
rect 20130 27918 20132 27970
rect 20076 27906 20132 27918
rect 19964 26852 20132 26908
rect 19740 26348 19908 26404
rect 19740 26180 19796 26190
rect 19740 26086 19796 26124
rect 19740 25732 19796 25742
rect 19740 25506 19796 25676
rect 19740 25454 19742 25506
rect 19794 25454 19796 25506
rect 19740 25442 19796 25454
rect 19852 23828 19908 26348
rect 19964 24052 20020 24062
rect 20076 24052 20132 26852
rect 19964 24050 20132 24052
rect 19964 23998 19966 24050
rect 20018 23998 20132 24050
rect 19964 23996 20132 23998
rect 20188 25844 20244 25854
rect 19964 23986 20020 23996
rect 20076 23828 20132 23838
rect 19852 23772 20020 23828
rect 19852 21362 19908 21374
rect 19852 21310 19854 21362
rect 19906 21310 19908 21362
rect 19852 21026 19908 21310
rect 19852 20974 19854 21026
rect 19906 20974 19908 21026
rect 19852 20962 19908 20974
rect 19740 20916 19796 20926
rect 19740 20130 19796 20860
rect 19740 20078 19742 20130
rect 19794 20078 19796 20130
rect 19740 20066 19796 20078
rect 19964 5236 20020 23772
rect 20076 15988 20132 23772
rect 20188 20802 20244 25788
rect 20188 20750 20190 20802
rect 20242 20750 20244 20802
rect 20188 20738 20244 20750
rect 20076 15922 20132 15932
rect 19964 5170 20020 5180
rect 19628 5058 19684 5068
rect 20300 644 20356 48636
rect 20748 43708 20804 55244
rect 20972 55298 21028 55310
rect 20972 55246 20974 55298
rect 21026 55246 21028 55298
rect 20860 53730 20916 53742
rect 20860 53678 20862 53730
rect 20914 53678 20916 53730
rect 20860 48692 20916 53678
rect 20860 48626 20916 48636
rect 20412 43652 20804 43708
rect 20412 35026 20468 43652
rect 20972 35476 21028 55246
rect 21084 54626 21140 55916
rect 21980 55972 22036 55982
rect 21644 55860 21700 55870
rect 21644 55410 21700 55804
rect 21644 55358 21646 55410
rect 21698 55358 21700 55410
rect 21644 55346 21700 55358
rect 21084 54574 21086 54626
rect 21138 54574 21140 54626
rect 21084 54562 21140 54574
rect 21532 54402 21588 54414
rect 21532 54350 21534 54402
rect 21586 54350 21588 54402
rect 21532 53956 21588 54350
rect 21532 53890 21588 53900
rect 21532 53732 21588 53742
rect 21308 53620 21364 53630
rect 21308 53526 21364 53564
rect 20972 35410 21028 35420
rect 21084 53508 21140 53518
rect 20412 34974 20414 35026
rect 20466 34974 20468 35026
rect 20412 34962 20468 34974
rect 20412 28868 20468 28878
rect 20412 28642 20468 28812
rect 20412 28590 20414 28642
rect 20466 28590 20468 28642
rect 20412 25732 20468 28590
rect 20412 25666 20468 25676
rect 20972 25732 21028 25742
rect 20636 25506 20692 25518
rect 20636 25454 20638 25506
rect 20690 25454 20692 25506
rect 20636 23380 20692 25454
rect 20636 23314 20692 23324
rect 20748 22036 20804 22046
rect 20412 20916 20468 20926
rect 20412 20822 20468 20860
rect 20748 20914 20804 21980
rect 20748 20862 20750 20914
rect 20802 20862 20804 20914
rect 20748 4900 20804 20862
rect 20972 10052 21028 25676
rect 21084 18452 21140 53452
rect 21308 52836 21364 52846
rect 21308 52742 21364 52780
rect 21420 28642 21476 28654
rect 21420 28590 21422 28642
rect 21474 28590 21476 28642
rect 21084 18386 21140 18396
rect 21196 23380 21252 23390
rect 20972 9986 21028 9996
rect 20748 4834 20804 4844
rect 20300 578 20356 588
rect 20860 3332 20916 3342
rect 20860 112 20916 3276
rect 21196 2884 21252 23324
rect 21420 20188 21476 28590
rect 21308 20132 21476 20188
rect 21308 18340 21364 20132
rect 21308 17108 21364 18284
rect 21308 17042 21364 17052
rect 21532 5124 21588 53676
rect 21868 53730 21924 53742
rect 21868 53678 21870 53730
rect 21922 53678 21924 53730
rect 21756 53172 21812 53182
rect 21756 53058 21812 53116
rect 21756 53006 21758 53058
rect 21810 53006 21812 53058
rect 21756 52994 21812 53006
rect 21868 53060 21924 53678
rect 21868 52994 21924 53004
rect 21868 52276 21924 52286
rect 21980 52276 22036 55916
rect 22540 54738 22596 56140
rect 22652 55186 22708 57148
rect 23548 56308 23604 57344
rect 24220 57204 24276 57214
rect 23804 56476 24068 56486
rect 23860 56420 23908 56476
rect 23964 56420 24012 56476
rect 23804 56410 24068 56420
rect 23548 56242 23604 56252
rect 23548 56084 23604 56094
rect 22876 55970 22932 55982
rect 22876 55918 22878 55970
rect 22930 55918 22932 55970
rect 22876 55468 22932 55918
rect 23212 55524 23268 55534
rect 22876 55412 23044 55468
rect 22652 55134 22654 55186
rect 22706 55134 22708 55186
rect 22652 55122 22708 55134
rect 22540 54686 22542 54738
rect 22594 54686 22596 54738
rect 22540 54674 22596 54686
rect 22204 53844 22260 53854
rect 22204 53618 22260 53788
rect 22204 53566 22206 53618
rect 22258 53566 22260 53618
rect 22204 53554 22260 53566
rect 22876 53730 22932 53742
rect 22876 53678 22878 53730
rect 22930 53678 22932 53730
rect 22652 53284 22708 53294
rect 22652 53058 22708 53228
rect 22652 53006 22654 53058
rect 22706 53006 22708 53058
rect 22652 52994 22708 53006
rect 22204 52724 22260 52734
rect 22204 52630 22260 52668
rect 21868 52274 22036 52276
rect 21868 52222 21870 52274
rect 21922 52222 22036 52274
rect 21868 52220 22036 52222
rect 22764 52612 22820 52622
rect 22764 52274 22820 52556
rect 22764 52222 22766 52274
rect 22818 52222 22820 52274
rect 21868 52210 21924 52220
rect 22764 52210 22820 52222
rect 22428 52162 22484 52174
rect 22428 52110 22430 52162
rect 22482 52110 22484 52162
rect 21868 38052 21924 38062
rect 21868 29876 21924 37996
rect 21868 29810 21924 29820
rect 22204 33796 22260 33806
rect 21532 5058 21588 5068
rect 21196 2818 21252 2828
rect 22204 112 22260 33740
rect 22428 1652 22484 52110
rect 22876 51380 22932 53678
rect 22876 51314 22932 51324
rect 22428 1586 22484 1596
rect 22764 51154 22820 51166
rect 22764 51102 22766 51154
rect 22818 51102 22820 51154
rect 22764 980 22820 51102
rect 22988 49924 23044 55412
rect 23100 54404 23156 54414
rect 23100 54310 23156 54348
rect 22988 49858 23044 49868
rect 23100 52834 23156 52846
rect 23100 52782 23102 52834
rect 23154 52782 23156 52834
rect 23100 12404 23156 52782
rect 23212 51490 23268 55468
rect 23548 52274 23604 56028
rect 23884 55972 23940 55982
rect 23884 55878 23940 55916
rect 23548 52222 23550 52274
rect 23602 52222 23604 52274
rect 23548 52210 23604 52222
rect 23660 55298 23716 55310
rect 23660 55246 23662 55298
rect 23714 55246 23716 55298
rect 23212 51438 23214 51490
rect 23266 51438 23268 51490
rect 23212 51426 23268 51438
rect 23548 52052 23604 52062
rect 23436 50708 23492 50718
rect 23548 50708 23604 51996
rect 23660 51604 23716 55246
rect 23804 54908 24068 54918
rect 23860 54852 23908 54908
rect 23964 54852 24012 54908
rect 23804 54842 24068 54852
rect 24108 54740 24164 54750
rect 24108 54646 24164 54684
rect 23772 54516 23828 54526
rect 23772 53618 23828 54460
rect 23772 53566 23774 53618
rect 23826 53566 23828 53618
rect 23772 53554 23828 53566
rect 23804 53340 24068 53350
rect 23860 53284 23908 53340
rect 23964 53284 24012 53340
rect 23804 53274 24068 53284
rect 24108 53172 24164 53182
rect 24220 53172 24276 57148
rect 24444 56308 24500 56318
rect 24444 56214 24500 56252
rect 24892 56308 24948 57344
rect 25452 57316 25508 57326
rect 24892 56242 24948 56252
rect 25340 56756 25396 56766
rect 24464 55692 24728 55702
rect 24520 55636 24568 55692
rect 24624 55636 24672 55692
rect 24464 55626 24728 55636
rect 25004 55412 25060 55422
rect 24892 55298 24948 55310
rect 24892 55246 24894 55298
rect 24946 55246 24948 55298
rect 24668 54404 24724 54414
rect 24108 53170 24276 53172
rect 24108 53118 24110 53170
rect 24162 53118 24276 53170
rect 24108 53116 24276 53118
rect 24332 54402 24724 54404
rect 24332 54350 24670 54402
rect 24722 54350 24724 54402
rect 24332 54348 24724 54350
rect 24108 53106 24164 53116
rect 24220 52948 24276 52958
rect 24220 51828 24276 52892
rect 24332 52052 24388 54348
rect 24668 54338 24724 54348
rect 24464 54124 24728 54134
rect 24520 54068 24568 54124
rect 24624 54068 24672 54124
rect 24464 54058 24728 54068
rect 24668 53730 24724 53742
rect 24668 53678 24670 53730
rect 24722 53678 24724 53730
rect 24668 53508 24724 53678
rect 24668 53442 24724 53452
rect 24668 52836 24724 52846
rect 24668 52742 24724 52780
rect 24464 52556 24728 52566
rect 24520 52500 24568 52556
rect 24624 52500 24672 52556
rect 24464 52490 24728 52500
rect 24668 52276 24724 52286
rect 24668 52182 24724 52220
rect 24332 51986 24388 51996
rect 23804 51772 24068 51782
rect 24220 51772 24388 51828
rect 23860 51716 23908 51772
rect 23964 51716 24012 51772
rect 23804 51706 24068 51716
rect 23660 51548 24276 51604
rect 23772 51156 23828 51166
rect 23772 51062 23828 51100
rect 23436 50706 23604 50708
rect 23436 50654 23438 50706
rect 23490 50654 23604 50706
rect 23436 50652 23604 50654
rect 23436 50642 23492 50652
rect 23884 50596 23940 50606
rect 23548 50594 23940 50596
rect 23548 50542 23886 50594
rect 23938 50542 23940 50594
rect 23548 50540 23940 50542
rect 23548 50260 23604 50540
rect 23884 50530 23940 50540
rect 23100 12338 23156 12348
rect 23436 50204 23604 50260
rect 23804 50204 24068 50214
rect 23436 6804 23492 50204
rect 23860 50148 23908 50204
rect 23964 50148 24012 50204
rect 23804 50138 24068 50148
rect 24220 50148 24276 51548
rect 24332 51490 24388 51772
rect 24892 51604 24948 55246
rect 25004 54516 25060 55356
rect 25004 54450 25060 54460
rect 24332 51438 24334 51490
rect 24386 51438 24388 51490
rect 24332 51426 24388 51438
rect 24780 51548 24948 51604
rect 24780 51156 24836 51548
rect 25340 51490 25396 56700
rect 25452 54626 25508 57260
rect 26236 57316 26292 57344
rect 26236 57250 26292 57260
rect 26012 56308 26068 56318
rect 26012 56214 26068 56252
rect 25676 56082 25732 56094
rect 25676 56030 25678 56082
rect 25730 56030 25732 56082
rect 25452 54574 25454 54626
rect 25506 54574 25508 54626
rect 25452 54562 25508 54574
rect 25564 55186 25620 55198
rect 25564 55134 25566 55186
rect 25618 55134 25620 55186
rect 25564 54516 25620 55134
rect 25564 54450 25620 54460
rect 25564 53620 25620 53630
rect 25564 53526 25620 53564
rect 25452 52834 25508 52846
rect 25452 52782 25454 52834
rect 25506 52782 25508 52834
rect 25452 52724 25508 52782
rect 25452 52658 25508 52668
rect 25564 52050 25620 52062
rect 25564 51998 25566 52050
rect 25618 51998 25620 52050
rect 25564 51828 25620 51998
rect 25564 51762 25620 51772
rect 25340 51438 25342 51490
rect 25394 51438 25396 51490
rect 25340 51426 25396 51438
rect 24892 51380 24948 51390
rect 24892 51378 25172 51380
rect 24892 51326 24894 51378
rect 24946 51326 25172 51378
rect 24892 51324 25172 51326
rect 24892 51314 24948 51324
rect 24780 51100 25060 51156
rect 24464 50988 24728 50998
rect 24520 50932 24568 50988
rect 24624 50932 24672 50988
rect 24464 50922 24728 50932
rect 24668 50594 24724 50606
rect 24668 50542 24670 50594
rect 24722 50542 24724 50594
rect 24668 50484 24724 50542
rect 24668 50418 24724 50428
rect 24220 50092 24388 50148
rect 24220 49924 24276 49934
rect 24220 49830 24276 49868
rect 23772 49586 23828 49598
rect 23772 49534 23774 49586
rect 23826 49534 23828 49586
rect 23772 49252 23828 49534
rect 23772 49186 23828 49196
rect 23804 48636 24068 48646
rect 23860 48580 23908 48636
rect 23964 48580 24012 48636
rect 23804 48570 24068 48580
rect 24332 48468 24388 50092
rect 24892 49810 24948 49822
rect 24892 49758 24894 49810
rect 24946 49758 24948 49810
rect 24464 49420 24728 49430
rect 24520 49364 24568 49420
rect 24624 49364 24672 49420
rect 24464 49354 24728 49364
rect 24668 49026 24724 49038
rect 24668 48974 24670 49026
rect 24722 48974 24724 49026
rect 24668 48916 24724 48974
rect 24668 48850 24724 48860
rect 24892 48580 24948 49758
rect 24892 48514 24948 48524
rect 24332 48412 24724 48468
rect 24444 48020 24500 48058
rect 24444 47954 24500 47964
rect 24668 48020 24724 48412
rect 25004 48356 25060 51100
rect 24780 48300 25060 48356
rect 24780 48020 24836 48300
rect 25004 48130 25060 48142
rect 25004 48078 25006 48130
rect 25058 48078 25060 48130
rect 25004 48020 25060 48078
rect 24780 47964 24948 48020
rect 24668 47954 24724 47964
rect 24464 47852 24728 47862
rect 24520 47796 24568 47852
rect 24624 47796 24672 47852
rect 24464 47786 24728 47796
rect 24668 47458 24724 47470
rect 24668 47406 24670 47458
rect 24722 47406 24724 47458
rect 23804 47068 24068 47078
rect 23860 47012 23908 47068
rect 23964 47012 24012 47068
rect 23804 47002 24068 47012
rect 24668 46900 24724 47406
rect 24668 46834 24724 46844
rect 24668 46564 24724 46574
rect 24220 46562 24724 46564
rect 24220 46510 24670 46562
rect 24722 46510 24724 46562
rect 24220 46508 24724 46510
rect 23804 45500 24068 45510
rect 23860 45444 23908 45500
rect 23964 45444 24012 45500
rect 23804 45434 24068 45444
rect 23804 43932 24068 43942
rect 23860 43876 23908 43932
rect 23964 43876 24012 43932
rect 23804 43866 24068 43876
rect 24220 42980 24276 46508
rect 24668 46498 24724 46508
rect 24464 46284 24728 46294
rect 24520 46228 24568 46284
rect 24624 46228 24672 46284
rect 24464 46218 24728 46228
rect 24780 45892 24836 45902
rect 24780 45798 24836 45836
rect 24464 44716 24728 44726
rect 24520 44660 24568 44716
rect 24624 44660 24672 44716
rect 24464 44650 24728 44660
rect 24668 44324 24724 44334
rect 24668 44230 24724 44268
rect 24892 43708 24948 47964
rect 25004 47954 25060 47964
rect 24892 43652 25060 43708
rect 24892 43538 24948 43550
rect 24892 43486 24894 43538
rect 24946 43486 24948 43538
rect 24464 43148 24728 43158
rect 24520 43092 24568 43148
rect 24624 43092 24672 43148
rect 24464 43082 24728 43092
rect 24220 42914 24276 42924
rect 24668 42756 24724 42766
rect 24668 42662 24724 42700
rect 23804 42364 24068 42374
rect 23860 42308 23908 42364
rect 23964 42308 24012 42364
rect 23804 42298 24068 42308
rect 24892 41972 24948 43486
rect 24892 41906 24948 41916
rect 24464 41580 24728 41590
rect 24520 41524 24568 41580
rect 24624 41524 24672 41580
rect 24464 41514 24728 41524
rect 24668 41188 24724 41198
rect 23660 41186 24724 41188
rect 23660 41134 24670 41186
rect 24722 41134 24724 41186
rect 23660 41132 24724 41134
rect 23660 33012 23716 41132
rect 24668 41122 24724 41132
rect 23804 40796 24068 40806
rect 23860 40740 23908 40796
rect 23964 40740 24012 40796
rect 23804 40730 24068 40740
rect 24892 40628 24948 40638
rect 24668 40516 24724 40526
rect 24668 40402 24724 40460
rect 24668 40350 24670 40402
rect 24722 40350 24724 40402
rect 24668 40338 24724 40350
rect 24464 40012 24728 40022
rect 24520 39956 24568 40012
rect 24624 39956 24672 40012
rect 24464 39946 24728 39956
rect 24892 39618 24948 40572
rect 24892 39566 24894 39618
rect 24946 39566 24948 39618
rect 24892 39554 24948 39566
rect 23804 39228 24068 39238
rect 23860 39172 23908 39228
rect 23964 39172 24012 39228
rect 23804 39162 24068 39172
rect 24464 38444 24728 38454
rect 24520 38388 24568 38444
rect 24624 38388 24672 38444
rect 24464 38378 24728 38388
rect 24668 38052 24724 38062
rect 24220 38050 24724 38052
rect 24220 37998 24670 38050
rect 24722 37998 24724 38050
rect 24220 37996 24724 37998
rect 23804 37660 24068 37670
rect 23860 37604 23908 37660
rect 23964 37604 24012 37660
rect 23804 37594 24068 37604
rect 23804 36092 24068 36102
rect 23860 36036 23908 36092
rect 23964 36036 24012 36092
rect 23804 36026 24068 36036
rect 23804 34524 24068 34534
rect 23860 34468 23908 34524
rect 23964 34468 24012 34524
rect 23804 34458 24068 34468
rect 23660 32946 23716 32956
rect 23804 32956 24068 32966
rect 23860 32900 23908 32956
rect 23964 32900 24012 32956
rect 23804 32890 24068 32900
rect 23804 31388 24068 31398
rect 23860 31332 23908 31388
rect 23964 31332 24012 31388
rect 23804 31322 24068 31332
rect 23804 29820 24068 29830
rect 23860 29764 23908 29820
rect 23964 29764 24012 29820
rect 23804 29754 24068 29764
rect 24220 28644 24276 37996
rect 24668 37986 24724 37996
rect 24892 37266 24948 37278
rect 24892 37214 24894 37266
rect 24946 37214 24948 37266
rect 24464 36876 24728 36886
rect 24520 36820 24568 36876
rect 24624 36820 24672 36876
rect 24464 36810 24728 36820
rect 24668 36484 24724 36494
rect 24668 36390 24724 36428
rect 24464 35308 24728 35318
rect 24520 35252 24568 35308
rect 24624 35252 24672 35308
rect 24464 35242 24728 35252
rect 24780 34914 24836 34926
rect 24780 34862 24782 34914
rect 24834 34862 24836 34914
rect 24668 34020 24724 34030
rect 24332 34018 24724 34020
rect 24332 33966 24670 34018
rect 24722 33966 24724 34018
rect 24332 33964 24724 33966
rect 24332 29092 24388 33964
rect 24668 33954 24724 33964
rect 24780 33908 24836 34862
rect 24892 34244 24948 37214
rect 24892 34178 24948 34188
rect 24780 33842 24836 33852
rect 24464 33740 24728 33750
rect 24520 33684 24568 33740
rect 24624 33684 24672 33740
rect 24464 33674 24728 33684
rect 24892 33348 24948 33358
rect 24892 33254 24948 33292
rect 24892 32788 24948 32798
rect 24464 32172 24728 32182
rect 24520 32116 24568 32172
rect 24624 32116 24672 32172
rect 24464 32106 24728 32116
rect 24780 31778 24836 31790
rect 24780 31726 24782 31778
rect 24834 31726 24836 31778
rect 24780 30772 24836 31726
rect 24892 30994 24948 32732
rect 24892 30942 24894 30994
rect 24946 30942 24948 30994
rect 24892 30930 24948 30942
rect 24780 30706 24836 30716
rect 24464 30604 24728 30614
rect 24520 30548 24568 30604
rect 24624 30548 24672 30604
rect 24464 30538 24728 30548
rect 24892 30100 24948 30110
rect 24332 29026 24388 29036
rect 24464 29036 24728 29046
rect 24520 28980 24568 29036
rect 24624 28980 24672 29036
rect 24464 28970 24728 28980
rect 24220 28578 24276 28588
rect 24668 28420 24724 28430
rect 23804 28252 24068 28262
rect 23860 28196 23908 28252
rect 23964 28196 24012 28252
rect 23804 28186 24068 28196
rect 24668 27858 24724 28364
rect 24668 27806 24670 27858
rect 24722 27806 24724 27858
rect 24668 27794 24724 27806
rect 24464 27468 24728 27478
rect 24520 27412 24568 27468
rect 24624 27412 24672 27468
rect 24464 27402 24728 27412
rect 24668 27188 24724 27198
rect 24668 27094 24724 27132
rect 23804 26684 24068 26694
rect 23860 26628 23908 26684
rect 23964 26628 24012 26684
rect 23804 26618 24068 26628
rect 24464 25900 24728 25910
rect 24520 25844 24568 25900
rect 24624 25844 24672 25900
rect 24464 25834 24728 25844
rect 24668 25620 24724 25630
rect 24668 25526 24724 25564
rect 23804 25116 24068 25126
rect 23860 25060 23908 25116
rect 23964 25060 24012 25116
rect 23804 25050 24068 25060
rect 24668 24610 24724 24622
rect 24668 24558 24670 24610
rect 24722 24558 24724 24610
rect 24668 24500 24724 24558
rect 24668 24434 24724 24444
rect 24464 24332 24728 24342
rect 24520 24276 24568 24332
rect 24624 24276 24672 24332
rect 24464 24266 24728 24276
rect 24892 23938 24948 30044
rect 25004 26180 25060 43652
rect 25004 26114 25060 26124
rect 24892 23886 24894 23938
rect 24946 23886 24948 23938
rect 24892 23874 24948 23886
rect 23804 23548 24068 23558
rect 23860 23492 23908 23548
rect 23964 23492 24012 23548
rect 23804 23482 24068 23492
rect 24464 22764 24728 22774
rect 24520 22708 24568 22764
rect 24624 22708 24672 22764
rect 24464 22698 24728 22708
rect 24892 22370 24948 22382
rect 24892 22318 24894 22370
rect 24946 22318 24948 22370
rect 23804 21980 24068 21990
rect 23860 21924 23908 21980
rect 23964 21924 24012 21980
rect 23804 21914 24068 21924
rect 24464 21196 24728 21206
rect 24520 21140 24568 21196
rect 24624 21140 24672 21196
rect 24464 21130 24728 21140
rect 23804 20412 24068 20422
rect 23860 20356 23908 20412
rect 23964 20356 24012 20412
rect 23804 20346 24068 20356
rect 24464 19628 24728 19638
rect 24520 19572 24568 19628
rect 24624 19572 24672 19628
rect 24464 19562 24728 19572
rect 23804 18844 24068 18854
rect 23860 18788 23908 18844
rect 23964 18788 24012 18844
rect 23804 18778 24068 18788
rect 24464 18060 24728 18070
rect 24520 18004 24568 18060
rect 24624 18004 24672 18060
rect 24464 17994 24728 18004
rect 23804 17276 24068 17286
rect 23860 17220 23908 17276
rect 23964 17220 24012 17276
rect 23804 17210 24068 17220
rect 24464 16492 24728 16502
rect 24520 16436 24568 16492
rect 24624 16436 24672 16492
rect 24464 16426 24728 16436
rect 23804 15708 24068 15718
rect 23860 15652 23908 15708
rect 23964 15652 24012 15708
rect 23804 15642 24068 15652
rect 24464 14924 24728 14934
rect 24520 14868 24568 14924
rect 24624 14868 24672 14924
rect 24464 14858 24728 14868
rect 23804 14140 24068 14150
rect 23860 14084 23908 14140
rect 23964 14084 24012 14140
rect 23804 14074 24068 14084
rect 23884 13636 23940 13646
rect 23884 13412 23940 13580
rect 23884 13346 23940 13356
rect 24464 13356 24728 13366
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24464 13290 24728 13300
rect 24892 12740 24948 22318
rect 25116 14756 25172 51324
rect 25564 50484 25620 50494
rect 25564 50390 25620 50428
rect 25452 49698 25508 49710
rect 25452 49646 25454 49698
rect 25506 49646 25508 49698
rect 25452 49588 25508 49646
rect 25452 49522 25508 49532
rect 25564 48914 25620 48926
rect 25564 48862 25566 48914
rect 25618 48862 25620 48914
rect 25564 48692 25620 48862
rect 25564 48626 25620 48636
rect 25676 48356 25732 56030
rect 27580 56084 27636 57344
rect 27580 56018 27636 56028
rect 26236 55300 26292 55310
rect 26236 55206 26292 55244
rect 27244 55074 27300 55086
rect 27244 55022 27246 55074
rect 27298 55022 27300 55074
rect 26236 54402 26292 54414
rect 26236 54350 26238 54402
rect 26290 54350 26292 54402
rect 26236 54292 26292 54350
rect 26236 54226 26292 54236
rect 27020 54402 27076 54414
rect 27020 54350 27022 54402
rect 27074 54350 27076 54402
rect 26236 53732 26292 53742
rect 26236 53638 26292 53676
rect 27020 53172 27076 54350
rect 27244 54068 27300 55022
rect 27244 54002 27300 54012
rect 27020 53106 27076 53116
rect 27244 53506 27300 53518
rect 27244 53454 27246 53506
rect 27298 53454 27300 53506
rect 27132 53058 27188 53070
rect 27132 53006 27134 53058
rect 27186 53006 27188 53058
rect 26236 52834 26292 52846
rect 26236 52782 26238 52834
rect 26290 52782 26292 52834
rect 26236 52388 26292 52782
rect 26236 52322 26292 52332
rect 26236 52164 26292 52174
rect 26236 52070 26292 52108
rect 27132 51380 27188 53006
rect 27244 52276 27300 53454
rect 27244 52210 27300 52220
rect 27356 52948 27412 52958
rect 27132 51314 27188 51324
rect 27244 51938 27300 51950
rect 27244 51886 27246 51938
rect 27298 51886 27300 51938
rect 26236 51268 26292 51278
rect 26236 51174 26292 51212
rect 27020 51266 27076 51278
rect 27020 51214 27022 51266
rect 27074 51214 27076 51266
rect 26236 50708 26292 50718
rect 26236 50614 26292 50652
rect 27020 50036 27076 51214
rect 27244 50932 27300 51886
rect 27244 50866 27300 50876
rect 27020 49970 27076 49980
rect 27244 50370 27300 50382
rect 27244 50318 27246 50370
rect 27298 50318 27300 50370
rect 27132 49922 27188 49934
rect 27132 49870 27134 49922
rect 27186 49870 27188 49922
rect 26348 49810 26404 49822
rect 26348 49758 26350 49810
rect 26402 49758 26404 49810
rect 26236 49028 26292 49038
rect 26236 48934 26292 48972
rect 26348 48804 26404 49758
rect 26348 48738 26404 48748
rect 25788 48356 25844 48366
rect 25676 48354 25844 48356
rect 25676 48302 25790 48354
rect 25842 48302 25844 48354
rect 25676 48300 25844 48302
rect 25788 48290 25844 48300
rect 27132 48244 27188 49870
rect 27244 49140 27300 50318
rect 27244 49074 27300 49084
rect 27132 48178 27188 48188
rect 27244 48802 27300 48814
rect 27244 48750 27246 48802
rect 27298 48750 27300 48802
rect 26236 48132 26292 48142
rect 26236 48038 26292 48076
rect 27020 48130 27076 48142
rect 27020 48078 27022 48130
rect 27074 48078 27076 48130
rect 25340 48020 25396 48030
rect 25340 47926 25396 47964
rect 26236 47458 26292 47470
rect 26236 47406 26238 47458
rect 26290 47406 26292 47458
rect 25676 47348 25732 47358
rect 25676 47254 25732 47292
rect 25676 46786 25732 46798
rect 25676 46734 25678 46786
rect 25730 46734 25732 46786
rect 25676 46452 25732 46734
rect 26236 46788 26292 47406
rect 27020 46900 27076 48078
rect 27244 47796 27300 48750
rect 27244 47730 27300 47740
rect 27020 46834 27076 46844
rect 27244 47234 27300 47246
rect 27244 47182 27246 47234
rect 27298 47182 27300 47234
rect 26236 46722 26292 46732
rect 27132 46786 27188 46798
rect 27132 46734 27134 46786
rect 27186 46734 27188 46786
rect 26236 46564 26292 46574
rect 26236 46470 26292 46508
rect 25676 46386 25732 46396
rect 26460 45890 26516 45902
rect 26460 45838 26462 45890
rect 26514 45838 26516 45890
rect 25676 45666 25732 45678
rect 25676 45614 25678 45666
rect 25730 45614 25732 45666
rect 25676 45556 25732 45614
rect 25676 45490 25732 45500
rect 26348 45106 26404 45118
rect 26348 45054 26350 45106
rect 26402 45054 26404 45106
rect 26236 44324 26292 44334
rect 25788 44322 26292 44324
rect 25788 44270 26238 44322
rect 26290 44270 26292 44322
rect 25788 44268 26292 44270
rect 25676 44212 25732 44222
rect 25676 44118 25732 44156
rect 25788 43988 25844 44268
rect 26236 44258 26292 44268
rect 25564 43932 25844 43988
rect 25564 43708 25620 43932
rect 25340 43652 25620 43708
rect 25340 35588 25396 43652
rect 25676 43650 25732 43662
rect 25676 43598 25678 43650
rect 25730 43598 25732 43650
rect 25676 43316 25732 43598
rect 25676 43250 25732 43260
rect 26236 43426 26292 43438
rect 26236 43374 26238 43426
rect 26290 43374 26292 43426
rect 26236 43092 26292 43374
rect 25452 43036 26292 43092
rect 25452 38612 25508 43036
rect 26236 42756 26292 42766
rect 25900 42754 26292 42756
rect 25900 42702 26238 42754
rect 26290 42702 26292 42754
rect 25900 42700 26292 42702
rect 25676 42530 25732 42542
rect 25676 42478 25678 42530
rect 25730 42478 25732 42530
rect 25676 42420 25732 42478
rect 25676 42354 25732 42364
rect 25676 41076 25732 41086
rect 25676 40982 25732 41020
rect 25676 40514 25732 40526
rect 25676 40462 25678 40514
rect 25730 40462 25732 40514
rect 25676 40180 25732 40462
rect 25676 40114 25732 40124
rect 25676 39394 25732 39406
rect 25676 39342 25678 39394
rect 25730 39342 25732 39394
rect 25676 39284 25732 39342
rect 25676 39218 25732 39228
rect 25452 38546 25508 38556
rect 25676 37940 25732 37950
rect 25676 37846 25732 37884
rect 25452 37154 25508 37166
rect 25452 37102 25454 37154
rect 25506 37102 25508 37154
rect 25452 37044 25508 37102
rect 25452 36978 25508 36988
rect 25788 37156 25844 37166
rect 25676 36258 25732 36270
rect 25676 36206 25678 36258
rect 25730 36206 25732 36258
rect 25676 36148 25732 36206
rect 25676 36082 25732 36092
rect 25340 35522 25396 35532
rect 25228 34916 25284 34926
rect 25228 27860 25284 34860
rect 25676 34804 25732 34814
rect 25676 34710 25732 34748
rect 25676 34242 25732 34254
rect 25676 34190 25678 34242
rect 25730 34190 25732 34242
rect 25676 33908 25732 34190
rect 25676 33842 25732 33852
rect 25788 33572 25844 37100
rect 25788 33506 25844 33516
rect 25676 33122 25732 33134
rect 25676 33070 25678 33122
rect 25730 33070 25732 33122
rect 25676 33012 25732 33070
rect 25676 32946 25732 32956
rect 25228 27794 25284 27804
rect 25340 32900 25396 32910
rect 25228 26404 25284 26414
rect 25228 24724 25284 26348
rect 25228 24658 25284 24668
rect 25340 23828 25396 32844
rect 25564 32788 25620 32798
rect 25452 30882 25508 30894
rect 25452 30830 25454 30882
rect 25506 30830 25508 30882
rect 25452 30772 25508 30830
rect 25452 30706 25508 30716
rect 25452 29988 25508 29998
rect 25452 24836 25508 29932
rect 25564 26404 25620 32732
rect 25676 31668 25732 31678
rect 25676 31574 25732 31612
rect 25676 27970 25732 27982
rect 25676 27918 25678 27970
rect 25730 27918 25732 27970
rect 25676 27188 25732 27918
rect 25676 27122 25732 27132
rect 25564 26338 25620 26348
rect 25676 26850 25732 26862
rect 25676 26798 25678 26850
rect 25730 26798 25732 26850
rect 25676 26292 25732 26798
rect 25676 26226 25732 26236
rect 25452 24770 25508 24780
rect 25564 25956 25620 25966
rect 25452 24610 25508 24622
rect 25452 24558 25454 24610
rect 25506 24558 25508 24610
rect 25452 24052 25508 24558
rect 25452 23986 25508 23996
rect 25340 23772 25508 23828
rect 25340 21474 25396 21486
rect 25340 21422 25342 21474
rect 25394 21422 25396 21474
rect 25340 20244 25396 21422
rect 25340 20178 25396 20188
rect 25116 14690 25172 14700
rect 24892 12674 24948 12684
rect 23804 12572 24068 12582
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 23804 12506 24068 12516
rect 25452 12404 25508 23772
rect 25564 19908 25620 25900
rect 25676 25282 25732 25294
rect 25676 25230 25678 25282
rect 25730 25230 25732 25282
rect 25676 24948 25732 25230
rect 25676 24882 25732 24892
rect 25788 25172 25844 25182
rect 25676 23714 25732 23726
rect 25676 23662 25678 23714
rect 25730 23662 25732 23714
rect 25676 23156 25732 23662
rect 25676 23090 25732 23100
rect 25676 22146 25732 22158
rect 25676 22094 25678 22146
rect 25730 22094 25732 22146
rect 25676 21812 25732 22094
rect 25676 21746 25732 21756
rect 25788 20188 25844 25116
rect 25900 22596 25956 42700
rect 26236 42690 26292 42700
rect 26236 41860 26292 41870
rect 26236 41766 26292 41804
rect 26348 41412 26404 45054
rect 26460 43708 26516 45838
rect 26796 45892 26852 45902
rect 26460 43652 26628 43708
rect 26348 41346 26404 41356
rect 26236 41188 26292 41198
rect 26236 41094 26292 41132
rect 26460 40402 26516 40414
rect 26460 40350 26462 40402
rect 26514 40350 26516 40402
rect 26236 39620 26292 39630
rect 26236 39526 26292 39564
rect 26236 38724 26292 38734
rect 26012 38722 26292 38724
rect 26012 38670 26238 38722
rect 26290 38670 26292 38722
rect 26012 38668 26292 38670
rect 26012 26180 26068 38668
rect 26236 38658 26292 38668
rect 26348 38724 26404 38734
rect 26236 38052 26292 38062
rect 26236 37958 26292 37996
rect 26236 37156 26292 37166
rect 26236 37062 26292 37100
rect 26348 36482 26404 38668
rect 26348 36430 26350 36482
rect 26402 36430 26404 36482
rect 26348 36418 26404 36430
rect 26348 35698 26404 35710
rect 26348 35646 26350 35698
rect 26402 35646 26404 35698
rect 26124 35028 26180 35038
rect 26124 32452 26180 34972
rect 26236 34916 26292 34926
rect 26236 34822 26292 34860
rect 26348 34356 26404 35646
rect 26348 34290 26404 34300
rect 26236 34020 26292 34030
rect 26236 33926 26292 33964
rect 26236 33346 26292 33358
rect 26236 33294 26238 33346
rect 26290 33294 26292 33346
rect 26236 32676 26292 33294
rect 26460 32900 26516 40350
rect 26460 32834 26516 32844
rect 26572 32788 26628 43652
rect 26572 32722 26628 32732
rect 26684 33348 26740 33358
rect 26236 32610 26292 32620
rect 26236 32452 26292 32462
rect 26124 32450 26292 32452
rect 26124 32398 26238 32450
rect 26290 32398 26292 32450
rect 26124 32396 26292 32398
rect 26236 32386 26292 32396
rect 26348 31778 26404 31790
rect 26348 31726 26350 31778
rect 26402 31726 26404 31778
rect 26124 30436 26180 30446
rect 26124 28756 26180 30380
rect 26236 29316 26292 29326
rect 26236 29222 26292 29260
rect 26236 28756 26292 28766
rect 26124 28754 26292 28756
rect 26124 28702 26238 28754
rect 26290 28702 26292 28754
rect 26124 28700 26292 28702
rect 26236 28690 26292 28700
rect 26348 28084 26404 31726
rect 26460 30996 26516 31006
rect 26460 30994 26628 30996
rect 26460 30942 26462 30994
rect 26514 30942 26628 30994
rect 26460 30940 26628 30942
rect 26460 30930 26516 30940
rect 26348 28018 26404 28028
rect 26460 30210 26516 30222
rect 26460 30158 26462 30210
rect 26514 30158 26516 30210
rect 26348 27858 26404 27870
rect 26348 27806 26350 27858
rect 26402 27806 26404 27858
rect 26236 27636 26292 27646
rect 26236 27186 26292 27580
rect 26236 27134 26238 27186
rect 26290 27134 26292 27186
rect 26236 27122 26292 27134
rect 26012 26124 26180 26180
rect 26124 25956 26180 26124
rect 26236 26178 26292 26190
rect 26236 26126 26238 26178
rect 26290 26126 26292 26178
rect 26236 26068 26292 26126
rect 26236 26002 26292 26012
rect 26124 25890 26180 25900
rect 26236 25508 26292 25518
rect 26236 25414 26292 25452
rect 26348 25060 26404 27806
rect 26460 25172 26516 30158
rect 26572 28756 26628 30940
rect 26572 28690 26628 28700
rect 26460 25106 26516 25116
rect 26348 24994 26404 25004
rect 25900 22530 25956 22540
rect 26012 24836 26068 24846
rect 25900 21362 25956 21374
rect 25900 21310 25902 21362
rect 25954 21310 25956 21362
rect 25900 20916 25956 21310
rect 25900 20850 25956 20860
rect 26012 20914 26068 24780
rect 26236 24610 26292 24622
rect 26236 24558 26238 24610
rect 26290 24558 26292 24610
rect 26236 24164 26292 24558
rect 26236 24098 26292 24108
rect 26236 23938 26292 23950
rect 26236 23886 26238 23938
rect 26290 23886 26292 23938
rect 26236 23268 26292 23886
rect 26236 23202 26292 23212
rect 26348 23154 26404 23166
rect 26348 23102 26350 23154
rect 26402 23102 26404 23154
rect 26236 22484 26292 22494
rect 26236 22390 26292 22428
rect 26012 20862 26014 20914
rect 26066 20862 26068 20914
rect 26012 20850 26068 20862
rect 26124 21700 26180 21710
rect 25564 19842 25620 19852
rect 25676 20132 25844 20188
rect 26012 20132 26068 20142
rect 25676 13076 25732 20132
rect 25900 19348 25956 19358
rect 25900 17780 25956 19292
rect 26012 19346 26068 20076
rect 26012 19294 26014 19346
rect 26066 19294 26068 19346
rect 26012 19282 26068 19294
rect 26124 18562 26180 21644
rect 26236 21474 26292 21486
rect 26236 21422 26238 21474
rect 26290 21422 26292 21474
rect 26236 21364 26292 21422
rect 26236 21298 26292 21308
rect 26348 21028 26404 23102
rect 26348 20962 26404 20972
rect 26460 22148 26516 22158
rect 26124 18510 26126 18562
rect 26178 18510 26180 18562
rect 26124 18498 26180 18510
rect 26348 18452 26404 18462
rect 26124 17892 26180 17902
rect 26012 17780 26068 17790
rect 25900 17778 26068 17780
rect 25900 17726 26014 17778
rect 26066 17726 26068 17778
rect 25900 17724 26068 17726
rect 26012 17714 26068 17724
rect 25900 16212 25956 16222
rect 25676 13010 25732 13020
rect 25788 16100 25844 16110
rect 25452 12338 25508 12348
rect 24464 11788 24728 11798
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24464 11722 24728 11732
rect 23804 11004 24068 11014
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 23804 10938 24068 10948
rect 24464 10220 24728 10230
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24464 10154 24728 10164
rect 25788 9716 25844 16044
rect 25900 11508 25956 16156
rect 26012 15988 26068 15998
rect 26012 15894 26068 15932
rect 26124 15426 26180 17836
rect 26124 15374 26126 15426
rect 26178 15374 26180 15426
rect 26124 15362 26180 15374
rect 26236 15316 26292 15326
rect 26124 14418 26180 14430
rect 26124 14366 26126 14418
rect 26178 14366 26180 14418
rect 26012 13188 26068 13198
rect 26012 13074 26068 13132
rect 26012 13022 26014 13074
rect 26066 13022 26068 13074
rect 26012 13010 26068 13022
rect 26012 12292 26068 12302
rect 26012 12198 26068 12236
rect 26124 11956 26180 14366
rect 26124 11890 26180 11900
rect 26012 11508 26068 11518
rect 25900 11506 26068 11508
rect 25900 11454 26014 11506
rect 26066 11454 26068 11506
rect 25900 11452 26068 11454
rect 26012 11442 26068 11452
rect 26012 10052 26068 10062
rect 26012 9938 26068 9996
rect 26012 9886 26014 9938
rect 26066 9886 26068 9938
rect 26012 9874 26068 9886
rect 25788 9660 26068 9716
rect 23804 9436 24068 9446
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 23804 9370 24068 9380
rect 25788 9268 25844 9278
rect 24464 8652 24728 8662
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24464 8586 24728 8596
rect 23804 7868 24068 7878
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 23804 7802 24068 7812
rect 24464 7084 24728 7094
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 24464 7018 24728 7028
rect 23436 6738 23492 6748
rect 23804 6300 24068 6310
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 23804 6234 24068 6244
rect 24464 5516 24728 5526
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24464 5450 24728 5460
rect 23804 4732 24068 4742
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 23804 4666 24068 4676
rect 24464 3948 24728 3958
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24464 3882 24728 3892
rect 23804 3164 24068 3174
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 23804 3098 24068 3108
rect 24464 2380 24728 2390
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24464 2314 24728 2324
rect 25788 2100 25844 9212
rect 26012 9154 26068 9660
rect 26012 9102 26014 9154
rect 26066 9102 26068 9154
rect 26012 9090 26068 9102
rect 26236 8932 26292 15260
rect 26348 10836 26404 18396
rect 26348 10770 26404 10780
rect 26012 8876 26292 8932
rect 26012 8370 26068 8876
rect 26460 8428 26516 22092
rect 26572 20802 26628 20814
rect 26572 20750 26574 20802
rect 26626 20750 26628 20802
rect 26572 20020 26628 20750
rect 26572 19954 26628 19964
rect 26572 19234 26628 19246
rect 26572 19182 26574 19234
rect 26626 19182 26628 19234
rect 26572 18676 26628 19182
rect 26572 18610 26628 18620
rect 26684 18452 26740 33292
rect 26684 18386 26740 18396
rect 26572 18228 26628 18238
rect 26572 18226 26740 18228
rect 26572 18174 26574 18226
rect 26626 18174 26740 18226
rect 26572 18172 26740 18174
rect 26572 18162 26628 18172
rect 26684 17780 26740 18172
rect 26684 17714 26740 17724
rect 26572 17666 26628 17678
rect 26572 17614 26574 17666
rect 26626 17614 26628 17666
rect 26572 16884 26628 17614
rect 26572 16818 26628 16828
rect 26572 16098 26628 16110
rect 26572 16046 26574 16098
rect 26626 16046 26628 16098
rect 26572 15540 26628 16046
rect 26572 15474 26628 15484
rect 26572 15092 26628 15102
rect 26572 15090 26740 15092
rect 26572 15038 26574 15090
rect 26626 15038 26740 15090
rect 26572 15036 26740 15038
rect 26572 15026 26628 15036
rect 26684 14644 26740 15036
rect 26684 14578 26740 14588
rect 26572 14530 26628 14542
rect 26572 14478 26574 14530
rect 26626 14478 26628 14530
rect 26572 13748 26628 14478
rect 26572 13682 26628 13692
rect 26572 12962 26628 12974
rect 26572 12910 26574 12962
rect 26626 12910 26628 12962
rect 26572 12404 26628 12910
rect 26572 12338 26628 12348
rect 26572 11956 26628 11966
rect 26572 11954 26740 11956
rect 26572 11902 26574 11954
rect 26626 11902 26740 11954
rect 26572 11900 26740 11902
rect 26572 11890 26628 11900
rect 26684 11508 26740 11900
rect 26684 11442 26740 11452
rect 26572 11394 26628 11406
rect 26572 11342 26574 11394
rect 26626 11342 26628 11394
rect 26572 10612 26628 11342
rect 26572 10546 26628 10556
rect 26572 9826 26628 9838
rect 26572 9774 26574 9826
rect 26626 9774 26628 9826
rect 26572 9268 26628 9774
rect 26572 9202 26628 9212
rect 26012 8318 26014 8370
rect 26066 8318 26068 8370
rect 26012 8306 26068 8318
rect 26124 8372 26516 8428
rect 26572 8818 26628 8830
rect 26572 8766 26574 8818
rect 26626 8766 26628 8818
rect 26572 8428 26628 8766
rect 26572 8372 26740 8428
rect 26012 6580 26068 6590
rect 26012 6486 26068 6524
rect 26012 5796 26068 5806
rect 26012 5702 26068 5740
rect 26012 5236 26068 5246
rect 26124 5236 26180 8372
rect 26684 8306 26740 8316
rect 26572 8258 26628 8270
rect 26572 8206 26574 8258
rect 26626 8206 26628 8258
rect 26572 7588 26628 8206
rect 26796 7700 26852 45836
rect 27132 45108 27188 46734
rect 27244 46004 27300 47182
rect 27244 45938 27300 45948
rect 27132 45042 27188 45052
rect 27244 45666 27300 45678
rect 27244 45614 27246 45666
rect 27298 45614 27300 45666
rect 27020 44994 27076 45006
rect 27020 44942 27022 44994
rect 27074 44942 27076 44994
rect 27020 43764 27076 44942
rect 27244 44660 27300 45614
rect 27244 44594 27300 44604
rect 27020 43698 27076 43708
rect 27244 44098 27300 44110
rect 27244 44046 27246 44098
rect 27298 44046 27300 44098
rect 27132 43650 27188 43662
rect 27132 43598 27134 43650
rect 27186 43598 27188 43650
rect 27132 41972 27188 43598
rect 27244 42868 27300 44046
rect 27244 42802 27300 42812
rect 27132 41906 27188 41916
rect 27244 42530 27300 42542
rect 27244 42478 27246 42530
rect 27298 42478 27300 42530
rect 27020 41858 27076 41870
rect 27020 41806 27022 41858
rect 27074 41806 27076 41858
rect 27020 40628 27076 41806
rect 27244 41524 27300 42478
rect 27244 41458 27300 41468
rect 27020 40562 27076 40572
rect 27244 40962 27300 40974
rect 27244 40910 27246 40962
rect 27298 40910 27300 40962
rect 27132 40514 27188 40526
rect 27132 40462 27134 40514
rect 27186 40462 27188 40514
rect 27132 38836 27188 40462
rect 27244 39732 27300 40910
rect 27244 39666 27300 39676
rect 27132 38770 27188 38780
rect 27244 39394 27300 39406
rect 27244 39342 27246 39394
rect 27298 39342 27300 39394
rect 27020 38722 27076 38734
rect 27020 38670 27022 38722
rect 27074 38670 27076 38722
rect 27020 37492 27076 38670
rect 27244 38388 27300 39342
rect 27244 38322 27300 38332
rect 27020 37426 27076 37436
rect 27244 37826 27300 37838
rect 27244 37774 27246 37826
rect 27298 37774 27300 37826
rect 27132 37378 27188 37390
rect 27132 37326 27134 37378
rect 27186 37326 27188 37378
rect 27132 35700 27188 37326
rect 27244 36596 27300 37774
rect 27244 36530 27300 36540
rect 27132 35634 27188 35644
rect 27244 36258 27300 36270
rect 27244 36206 27246 36258
rect 27298 36206 27300 36258
rect 27020 35586 27076 35598
rect 27020 35534 27022 35586
rect 27074 35534 27076 35586
rect 27020 34356 27076 35534
rect 27244 35252 27300 36206
rect 27244 35186 27300 35196
rect 27020 34290 27076 34300
rect 27244 34690 27300 34702
rect 27244 34638 27246 34690
rect 27298 34638 27300 34690
rect 27132 34242 27188 34254
rect 27132 34190 27134 34242
rect 27186 34190 27188 34242
rect 27132 32564 27188 34190
rect 27244 33460 27300 34638
rect 27244 33394 27300 33404
rect 27132 32498 27188 32508
rect 27244 33122 27300 33134
rect 27244 33070 27246 33122
rect 27298 33070 27300 33122
rect 27020 32450 27076 32462
rect 27020 32398 27022 32450
rect 27074 32398 27076 32450
rect 27020 31220 27076 32398
rect 27244 32116 27300 33070
rect 27244 32050 27300 32060
rect 27020 31154 27076 31164
rect 27244 31554 27300 31566
rect 27244 31502 27246 31554
rect 27298 31502 27300 31554
rect 27020 30882 27076 30894
rect 27020 30830 27022 30882
rect 27074 30830 27076 30882
rect 27020 29876 27076 30830
rect 27244 30324 27300 31502
rect 27244 30258 27300 30268
rect 27020 29810 27076 29820
rect 27132 30098 27188 30110
rect 27132 30046 27134 30098
rect 27186 30046 27188 30098
rect 27132 29428 27188 30046
rect 27132 29362 27188 29372
rect 27244 29538 27300 29550
rect 27244 29486 27246 29538
rect 27298 29486 27300 29538
rect 27244 28980 27300 29486
rect 27244 28914 27300 28924
rect 27244 28532 27300 28542
rect 27244 28438 27300 28476
rect 27244 28084 27300 28094
rect 27244 27990 27300 28028
rect 27244 27636 27300 27646
rect 26908 27300 26964 27310
rect 26908 20914 26964 27244
rect 27244 26962 27300 27580
rect 27244 26910 27246 26962
rect 27298 26910 27300 26962
rect 27244 26898 27300 26910
rect 27244 26740 27300 26750
rect 27244 26514 27300 26684
rect 27244 26462 27246 26514
rect 27298 26462 27300 26514
rect 27244 26450 27300 26462
rect 26908 20862 26910 20914
rect 26962 20862 26964 20914
rect 26908 20850 26964 20862
rect 27020 26180 27076 26190
rect 27020 20692 27076 26124
rect 27244 25844 27300 25854
rect 27132 25396 27188 25406
rect 27132 24834 27188 25340
rect 27244 25394 27300 25788
rect 27244 25342 27246 25394
rect 27298 25342 27300 25394
rect 27244 25330 27300 25342
rect 27132 24782 27134 24834
rect 27186 24782 27188 24834
rect 27132 24770 27188 24782
rect 27244 24500 27300 24510
rect 27244 23826 27300 24444
rect 27244 23774 27246 23826
rect 27298 23774 27300 23826
rect 27244 23762 27300 23774
rect 27132 23604 27188 23614
rect 27132 23266 27188 23548
rect 27132 23214 27134 23266
rect 27186 23214 27188 23266
rect 27132 23202 27188 23214
rect 27244 22708 27300 22718
rect 27132 22260 27188 22270
rect 27132 21698 27188 22204
rect 27244 22258 27300 22652
rect 27244 22206 27246 22258
rect 27298 22206 27300 22258
rect 27244 22194 27300 22206
rect 27132 21646 27134 21698
rect 27186 21646 27188 21698
rect 27132 21634 27188 21646
rect 26908 20636 27076 20692
rect 26908 18900 26964 20636
rect 27020 20132 27076 20142
rect 27020 20038 27076 20076
rect 27020 19124 27076 19134
rect 27020 19122 27300 19124
rect 27020 19070 27022 19122
rect 27074 19070 27300 19122
rect 27020 19068 27300 19070
rect 27020 19058 27076 19068
rect 26908 18844 27188 18900
rect 26908 18452 26964 18462
rect 26908 18358 26964 18396
rect 26908 17892 26964 17902
rect 26908 17778 26964 17836
rect 26908 17726 26910 17778
rect 26962 17726 26964 17778
rect 26908 17714 26964 17726
rect 27020 17556 27076 17566
rect 27020 16994 27076 17500
rect 27020 16942 27022 16994
rect 27074 16942 27076 16994
rect 27020 16930 27076 16942
rect 27132 16772 27188 18844
rect 27020 16716 27188 16772
rect 27020 15986 27076 16716
rect 27020 15934 27022 15986
rect 27074 15934 27076 15986
rect 27020 15922 27076 15934
rect 27132 16324 27188 16334
rect 27020 15426 27076 15438
rect 27020 15374 27022 15426
rect 27074 15374 27076 15426
rect 26908 14418 26964 14430
rect 26908 14366 26910 14418
rect 26962 14366 26964 14418
rect 26908 13860 26964 14366
rect 27020 14308 27076 15374
rect 27020 14242 27076 14252
rect 26908 13794 26964 13804
rect 26908 13636 26964 13646
rect 26908 13542 26964 13580
rect 27020 12852 27076 12862
rect 27132 12852 27188 16268
rect 27244 15092 27300 19068
rect 27244 15026 27300 15036
rect 27020 12850 27188 12852
rect 27020 12798 27022 12850
rect 27074 12798 27188 12850
rect 27020 12796 27188 12798
rect 27244 13524 27300 13534
rect 27020 12786 27076 12796
rect 27244 12740 27300 13468
rect 27132 12684 27300 12740
rect 26908 12292 26964 12302
rect 26908 12198 26964 12236
rect 27020 12068 27076 12078
rect 26908 11284 26964 11294
rect 26908 11190 26964 11228
rect 26908 10724 26964 10734
rect 26908 10630 26964 10668
rect 26908 9940 26964 9950
rect 26908 9846 26964 9884
rect 27020 9154 27076 12012
rect 27020 9102 27022 9154
rect 27074 9102 27076 9154
rect 27020 9090 27076 9102
rect 27020 8932 27076 8942
rect 26908 8146 26964 8158
rect 26908 8094 26910 8146
rect 26962 8094 26964 8146
rect 26908 8036 26964 8094
rect 26908 7970 26964 7980
rect 26796 7634 26852 7644
rect 26572 7522 26628 7532
rect 26908 7476 26964 7486
rect 26908 7382 26964 7420
rect 27020 6916 27076 8876
rect 26796 6860 27076 6916
rect 26012 5234 26180 5236
rect 26012 5182 26014 5234
rect 26066 5182 26180 5234
rect 26012 5180 26180 5182
rect 26236 6804 26292 6814
rect 26012 5170 26068 5180
rect 26012 3444 26068 3454
rect 26012 3350 26068 3388
rect 26012 2884 26068 2894
rect 26012 2790 26068 2828
rect 26012 2100 26068 2110
rect 25788 2098 26068 2100
rect 25788 2046 26014 2098
rect 26066 2046 26068 2098
rect 25788 2044 26068 2046
rect 26012 2034 26068 2044
rect 22764 914 22820 924
rect 23548 1652 23604 1662
rect 23548 112 23604 1596
rect 23804 1596 24068 1606
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 23804 1530 24068 1540
rect 24892 1540 24948 1550
rect 24780 1204 24836 1214
rect 24780 1110 24836 1148
rect 24464 812 24728 822
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24464 746 24728 756
rect 24892 112 24948 1484
rect 26124 1202 26180 1214
rect 26124 1150 26126 1202
rect 26178 1150 26180 1202
rect 25676 1092 25732 1102
rect 25676 998 25732 1036
rect 25340 978 25396 990
rect 25340 926 25342 978
rect 25394 926 25396 978
rect 25340 756 25396 926
rect 25340 690 25396 700
rect 26124 308 26180 1150
rect 26124 242 26180 252
rect 26236 112 26292 6748
rect 26572 6690 26628 6702
rect 26572 6638 26574 6690
rect 26626 6638 26628 6690
rect 26572 6132 26628 6638
rect 26572 6066 26628 6076
rect 26796 5796 26852 6860
rect 26908 6692 26964 6702
rect 26908 6598 26964 6636
rect 27132 6356 27188 12684
rect 27244 12180 27300 12190
rect 27244 6692 27300 12124
rect 27244 6626 27300 6636
rect 26908 6300 27188 6356
rect 26908 6018 26964 6300
rect 26908 5966 26910 6018
rect 26962 5966 26964 6018
rect 26908 5954 26964 5966
rect 27132 5796 27188 5806
rect 26796 5740 26964 5796
rect 26572 5684 26628 5694
rect 26572 5682 26740 5684
rect 26572 5630 26574 5682
rect 26626 5630 26740 5682
rect 26572 5628 26740 5630
rect 26572 5618 26628 5628
rect 26684 5236 26740 5628
rect 26684 5170 26740 5180
rect 26908 5234 26964 5740
rect 26908 5182 26910 5234
rect 26962 5182 26964 5234
rect 26908 5170 26964 5182
rect 26572 5122 26628 5134
rect 26572 5070 26574 5122
rect 26626 5070 26628 5122
rect 26460 4900 26516 4910
rect 26460 1316 26516 4844
rect 26572 4340 26628 5070
rect 26572 4274 26628 4284
rect 26796 5124 26852 5134
rect 26572 3554 26628 3566
rect 26572 3502 26574 3554
rect 26626 3502 26628 3554
rect 26572 2996 26628 3502
rect 26572 2930 26628 2940
rect 26572 2548 26628 2558
rect 26572 2546 26740 2548
rect 26572 2494 26574 2546
rect 26626 2494 26740 2546
rect 26572 2492 26740 2494
rect 26572 2482 26628 2492
rect 26684 2100 26740 2492
rect 26684 2034 26740 2044
rect 26572 1986 26628 1998
rect 26572 1934 26574 1986
rect 26626 1934 26628 1986
rect 26572 1652 26628 1934
rect 26572 1586 26628 1596
rect 26572 1316 26628 1326
rect 26460 1314 26628 1316
rect 26460 1262 26574 1314
rect 26626 1262 26628 1314
rect 26460 1260 26628 1262
rect 26572 1250 26628 1260
rect 26796 196 26852 5068
rect 26908 4452 26964 4462
rect 26908 3668 26964 4396
rect 27020 4452 27076 4462
rect 27132 4452 27188 5740
rect 27020 4450 27188 4452
rect 27020 4398 27022 4450
rect 27074 4398 27188 4450
rect 27020 4396 27188 4398
rect 27020 4386 27076 4396
rect 27356 4228 27412 52892
rect 27580 49252 27636 49262
rect 27468 21364 27524 21374
rect 27468 21026 27524 21308
rect 27468 20974 27470 21026
rect 27522 20974 27524 21026
rect 27468 20962 27524 20974
rect 27468 20468 27524 20478
rect 27468 20018 27524 20412
rect 27468 19966 27470 20018
rect 27522 19966 27524 20018
rect 27468 19954 27524 19966
rect 27468 19572 27524 19582
rect 27468 19458 27524 19516
rect 27468 19406 27470 19458
rect 27522 19406 27524 19458
rect 27468 19394 27524 19406
rect 27468 19124 27524 19134
rect 27468 18450 27524 19068
rect 27468 18398 27470 18450
rect 27522 18398 27524 18450
rect 27468 18386 27524 18398
rect 27468 18004 27524 18014
rect 27468 17890 27524 17948
rect 27468 17838 27470 17890
rect 27522 17838 27524 17890
rect 27468 17826 27524 17838
rect 27468 17332 27524 17342
rect 27468 16882 27524 17276
rect 27468 16830 27470 16882
rect 27522 16830 27524 16882
rect 27468 16818 27524 16830
rect 27468 16436 27524 16446
rect 27468 16322 27524 16380
rect 27468 16270 27470 16322
rect 27522 16270 27524 16322
rect 27468 16258 27524 16270
rect 27468 15988 27524 15998
rect 27468 15314 27524 15932
rect 27468 15262 27470 15314
rect 27522 15262 27524 15314
rect 27468 15250 27524 15262
rect 27468 14868 27524 14878
rect 27468 14754 27524 14812
rect 27468 14702 27470 14754
rect 27522 14702 27524 14754
rect 27468 14690 27524 14702
rect 27580 14420 27636 49196
rect 28140 48020 28196 48030
rect 27916 31108 27972 31118
rect 27804 29540 27860 29550
rect 27580 14354 27636 14364
rect 27692 27860 27748 27870
rect 27468 14196 27524 14206
rect 27692 14196 27748 27804
rect 27804 18452 27860 29484
rect 27916 20132 27972 31052
rect 27916 20066 27972 20076
rect 28028 30212 28084 30222
rect 27804 18386 27860 18396
rect 28028 17892 28084 30156
rect 28028 17826 28084 17836
rect 27916 17668 27972 17678
rect 27468 13746 27524 14140
rect 27468 13694 27470 13746
rect 27522 13694 27524 13746
rect 27468 13682 27524 13694
rect 27580 14140 27748 14196
rect 27804 14420 27860 14430
rect 27468 13300 27524 13310
rect 27468 13186 27524 13244
rect 27468 13134 27470 13186
rect 27522 13134 27524 13186
rect 27468 13122 27524 13134
rect 27468 12852 27524 12862
rect 27468 12178 27524 12796
rect 27468 12126 27470 12178
rect 27522 12126 27524 12178
rect 27468 12114 27524 12126
rect 27580 12180 27636 14140
rect 27580 12114 27636 12124
rect 27692 13860 27748 13870
rect 27580 11956 27636 11966
rect 27468 11620 27524 11630
rect 27580 11620 27636 11900
rect 27468 11618 27636 11620
rect 27468 11566 27470 11618
rect 27522 11566 27636 11618
rect 27468 11564 27636 11566
rect 27468 11554 27524 11564
rect 27468 11060 27524 11070
rect 27468 10610 27524 11004
rect 27468 10558 27470 10610
rect 27522 10558 27524 10610
rect 27468 10546 27524 10558
rect 27468 10164 27524 10174
rect 27468 10050 27524 10108
rect 27468 9998 27470 10050
rect 27522 9998 27524 10050
rect 27468 9986 27524 9998
rect 27468 9716 27524 9726
rect 27468 9042 27524 9660
rect 27468 8990 27470 9042
rect 27522 8990 27524 9042
rect 27468 8978 27524 8990
rect 27580 8820 27636 8830
rect 27468 8484 27524 8494
rect 27580 8484 27636 8764
rect 27468 8482 27636 8484
rect 27468 8430 27470 8482
rect 27522 8430 27636 8482
rect 27468 8428 27636 8430
rect 27468 8418 27524 8428
rect 27468 7924 27524 7934
rect 27468 7474 27524 7868
rect 27468 7422 27470 7474
rect 27522 7422 27524 7474
rect 27468 7410 27524 7422
rect 27468 7028 27524 7038
rect 27468 6914 27524 6972
rect 27468 6862 27470 6914
rect 27522 6862 27524 6914
rect 27468 6850 27524 6862
rect 27468 6580 27524 6590
rect 27468 5906 27524 6524
rect 27468 5854 27470 5906
rect 27522 5854 27524 5906
rect 27468 5842 27524 5854
rect 27580 5684 27636 5694
rect 27468 5348 27524 5358
rect 27580 5348 27636 5628
rect 27468 5346 27636 5348
rect 27468 5294 27470 5346
rect 27522 5294 27636 5346
rect 27468 5292 27636 5294
rect 27468 5282 27524 5292
rect 27468 4788 27524 4798
rect 27468 4338 27524 4732
rect 27468 4286 27470 4338
rect 27522 4286 27524 4338
rect 27468 4274 27524 4286
rect 27356 4162 27412 4172
rect 27468 3892 27524 3902
rect 27468 3778 27524 3836
rect 27468 3726 27470 3778
rect 27522 3726 27524 3778
rect 27468 3714 27524 3726
rect 26908 3612 27076 3668
rect 26908 3444 26964 3454
rect 26908 3350 26964 3388
rect 26908 2884 26964 2894
rect 26908 2790 26964 2828
rect 27020 1874 27076 3612
rect 27468 3444 27524 3454
rect 27468 2770 27524 3388
rect 27692 3332 27748 13804
rect 27692 3266 27748 3276
rect 27804 2884 27860 14364
rect 27916 12292 27972 17612
rect 27916 12226 27972 12236
rect 28028 13972 28084 13982
rect 28028 8428 28084 13916
rect 27916 8372 28084 8428
rect 27916 3556 27972 8372
rect 27916 3490 27972 3500
rect 27804 2818 27860 2828
rect 27468 2718 27470 2770
rect 27522 2718 27524 2770
rect 27468 2706 27524 2718
rect 27580 2548 27636 2558
rect 27468 2212 27524 2222
rect 27580 2212 27636 2492
rect 27468 2210 27636 2212
rect 27468 2158 27470 2210
rect 27522 2158 27636 2210
rect 27468 2156 27636 2158
rect 27468 2146 27524 2156
rect 27020 1822 27022 1874
rect 27074 1822 27076 1874
rect 27020 1810 27076 1822
rect 28140 1540 28196 47964
rect 28252 21476 28308 21486
rect 28308 21420 28420 21476
rect 28252 21410 28308 21420
rect 28252 17108 28308 17118
rect 28252 8932 28308 17052
rect 28364 14420 28420 21420
rect 28364 14354 28420 14364
rect 28252 8866 28308 8876
rect 28140 1474 28196 1484
rect 27132 1204 27188 1214
rect 27132 1110 27188 1148
rect 26796 130 26852 140
rect 27580 196 27636 206
rect 27580 112 27636 140
rect 672 0 784 112
rect 2016 0 2128 112
rect 3360 0 3472 112
rect 4704 0 4816 112
rect 6048 0 6160 112
rect 7392 0 7504 112
rect 8736 0 8848 112
rect 10080 0 10192 112
rect 11424 0 11536 112
rect 12768 0 12880 112
rect 14112 0 14224 112
rect 15456 0 15568 112
rect 16800 0 16912 112
rect 18144 0 18256 112
rect 19488 0 19600 112
rect 20832 0 20944 112
rect 22176 0 22288 112
rect 23520 0 23632 112
rect 24864 0 24976 112
rect 26208 0 26320 112
rect 27552 0 27664 112
<< via2 >>
rect 1036 53564 1092 53620
rect 4732 57260 4788 57316
rect 5516 57260 5572 57316
rect 3804 56474 3860 56476
rect 3804 56422 3806 56474
rect 3806 56422 3858 56474
rect 3858 56422 3860 56474
rect 3804 56420 3860 56422
rect 3908 56474 3964 56476
rect 3908 56422 3910 56474
rect 3910 56422 3962 56474
rect 3962 56422 3964 56474
rect 3908 56420 3964 56422
rect 4012 56474 4068 56476
rect 4012 56422 4014 56474
rect 4014 56422 4066 56474
rect 4066 56422 4068 56474
rect 4012 56420 4068 56422
rect 3052 55970 3108 55972
rect 3052 55918 3054 55970
rect 3054 55918 3106 55970
rect 3106 55918 3108 55970
rect 3052 55916 3108 55918
rect 4464 55690 4520 55692
rect 4464 55638 4466 55690
rect 4466 55638 4518 55690
rect 4518 55638 4520 55690
rect 4464 55636 4520 55638
rect 4568 55690 4624 55692
rect 4568 55638 4570 55690
rect 4570 55638 4622 55690
rect 4622 55638 4624 55690
rect 4568 55636 4624 55638
rect 4672 55690 4728 55692
rect 4672 55638 4674 55690
rect 4674 55638 4726 55690
rect 4726 55638 4728 55690
rect 4672 55636 4728 55638
rect 8092 55970 8148 55972
rect 8092 55918 8094 55970
rect 8094 55918 8146 55970
rect 8146 55918 8148 55970
rect 8092 55916 8148 55918
rect 1372 52892 1428 52948
rect 252 52780 308 52836
rect 140 28700 196 28756
rect 1036 52220 1092 52276
rect 1596 52834 1652 52836
rect 1596 52782 1598 52834
rect 1598 52782 1650 52834
rect 1650 52782 1652 52834
rect 1596 52780 1652 52782
rect 476 49868 532 49924
rect 588 41804 644 41860
rect 364 27580 420 27636
rect 476 30940 532 30996
rect 252 26572 308 26628
rect 364 27020 420 27076
rect 140 19740 196 19796
rect 252 26348 308 26404
rect 364 20636 420 20692
rect 252 17724 308 17780
rect 364 17052 420 17108
rect 700 41020 756 41076
rect 1036 50876 1092 50932
rect 1596 49868 1652 49924
rect 1596 49698 1652 49700
rect 1596 49646 1598 49698
rect 1598 49646 1650 49698
rect 1650 49646 1652 49698
rect 1596 49644 1652 49646
rect 1036 49586 1092 49588
rect 1036 49534 1038 49586
rect 1038 49534 1090 49586
rect 1090 49534 1092 49586
rect 1036 49532 1092 49534
rect 1596 48914 1652 48916
rect 1596 48862 1598 48914
rect 1598 48862 1650 48914
rect 1650 48862 1652 48914
rect 1596 48860 1652 48862
rect 1036 48188 1092 48244
rect 1036 46844 1092 46900
rect 1484 45778 1540 45780
rect 1484 45726 1486 45778
rect 1486 45726 1538 45778
rect 1538 45726 1540 45778
rect 1484 45724 1540 45726
rect 1036 45500 1092 45556
rect 1036 44156 1092 44212
rect 1596 43708 1652 43764
rect 1484 43596 1540 43652
rect 3804 54906 3860 54908
rect 3804 54854 3806 54906
rect 3806 54854 3858 54906
rect 3858 54854 3860 54906
rect 3804 54852 3860 54854
rect 3908 54906 3964 54908
rect 3908 54854 3910 54906
rect 3910 54854 3962 54906
rect 3962 54854 3964 54906
rect 3908 54852 3964 54854
rect 4012 54906 4068 54908
rect 4012 54854 4014 54906
rect 4014 54854 4066 54906
rect 4066 54854 4068 54906
rect 4012 54852 4068 54854
rect 4464 54122 4520 54124
rect 4464 54070 4466 54122
rect 4466 54070 4518 54122
rect 4518 54070 4520 54122
rect 4464 54068 4520 54070
rect 4568 54122 4624 54124
rect 4568 54070 4570 54122
rect 4570 54070 4622 54122
rect 4622 54070 4624 54122
rect 4568 54068 4624 54070
rect 4672 54122 4728 54124
rect 4672 54070 4674 54122
rect 4674 54070 4726 54122
rect 4726 54070 4728 54122
rect 4672 54068 4728 54070
rect 3804 53338 3860 53340
rect 3804 53286 3806 53338
rect 3806 53286 3858 53338
rect 3858 53286 3860 53338
rect 3804 53284 3860 53286
rect 3908 53338 3964 53340
rect 3908 53286 3910 53338
rect 3910 53286 3962 53338
rect 3962 53286 3964 53338
rect 3908 53284 3964 53286
rect 4012 53338 4068 53340
rect 4012 53286 4014 53338
rect 4014 53286 4066 53338
rect 4066 53286 4068 53338
rect 4012 53284 4068 53286
rect 4464 52554 4520 52556
rect 4464 52502 4466 52554
rect 4466 52502 4518 52554
rect 4518 52502 4520 52554
rect 4464 52500 4520 52502
rect 4568 52554 4624 52556
rect 4568 52502 4570 52554
rect 4570 52502 4622 52554
rect 4622 52502 4624 52554
rect 4568 52500 4624 52502
rect 4672 52554 4728 52556
rect 4672 52502 4674 52554
rect 4674 52502 4726 52554
rect 4726 52502 4728 52554
rect 4672 52500 4728 52502
rect 3804 51770 3860 51772
rect 3804 51718 3806 51770
rect 3806 51718 3858 51770
rect 3858 51718 3860 51770
rect 3804 51716 3860 51718
rect 3908 51770 3964 51772
rect 3908 51718 3910 51770
rect 3910 51718 3962 51770
rect 3962 51718 3964 51770
rect 3908 51716 3964 51718
rect 4012 51770 4068 51772
rect 4012 51718 4014 51770
rect 4014 51718 4066 51770
rect 4066 51718 4068 51770
rect 4012 51716 4068 51718
rect 4464 50986 4520 50988
rect 4464 50934 4466 50986
rect 4466 50934 4518 50986
rect 4518 50934 4520 50986
rect 4464 50932 4520 50934
rect 4568 50986 4624 50988
rect 4568 50934 4570 50986
rect 4570 50934 4622 50986
rect 4622 50934 4624 50986
rect 4568 50932 4624 50934
rect 4672 50986 4728 50988
rect 4672 50934 4674 50986
rect 4674 50934 4726 50986
rect 4726 50934 4728 50986
rect 4672 50932 4728 50934
rect 3804 50202 3860 50204
rect 3804 50150 3806 50202
rect 3806 50150 3858 50202
rect 3858 50150 3860 50202
rect 3804 50148 3860 50150
rect 3908 50202 3964 50204
rect 3908 50150 3910 50202
rect 3910 50150 3962 50202
rect 3962 50150 3964 50202
rect 3908 50148 3964 50150
rect 4012 50202 4068 50204
rect 4012 50150 4014 50202
rect 4014 50150 4066 50202
rect 4066 50150 4068 50202
rect 4012 50148 4068 50150
rect 4464 49418 4520 49420
rect 4464 49366 4466 49418
rect 4466 49366 4518 49418
rect 4518 49366 4520 49418
rect 4464 49364 4520 49366
rect 4568 49418 4624 49420
rect 4568 49366 4570 49418
rect 4570 49366 4622 49418
rect 4622 49366 4624 49418
rect 4568 49364 4624 49366
rect 4672 49418 4728 49420
rect 4672 49366 4674 49418
rect 4674 49366 4726 49418
rect 4726 49366 4728 49418
rect 4672 49364 4728 49366
rect 3804 48634 3860 48636
rect 3804 48582 3806 48634
rect 3806 48582 3858 48634
rect 3858 48582 3860 48634
rect 3804 48580 3860 48582
rect 3908 48634 3964 48636
rect 3908 48582 3910 48634
rect 3910 48582 3962 48634
rect 3962 48582 3964 48634
rect 3908 48580 3964 48582
rect 4012 48634 4068 48636
rect 4012 48582 4014 48634
rect 4014 48582 4066 48634
rect 4066 48582 4068 48634
rect 4012 48580 4068 48582
rect 4464 47850 4520 47852
rect 4464 47798 4466 47850
rect 4466 47798 4518 47850
rect 4518 47798 4520 47850
rect 4464 47796 4520 47798
rect 4568 47850 4624 47852
rect 4568 47798 4570 47850
rect 4570 47798 4622 47850
rect 4622 47798 4624 47850
rect 4568 47796 4624 47798
rect 4672 47850 4728 47852
rect 4672 47798 4674 47850
rect 4674 47798 4726 47850
rect 4726 47798 4728 47850
rect 4672 47796 4728 47798
rect 3804 47066 3860 47068
rect 3804 47014 3806 47066
rect 3806 47014 3858 47066
rect 3858 47014 3860 47066
rect 3804 47012 3860 47014
rect 3908 47066 3964 47068
rect 3908 47014 3910 47066
rect 3910 47014 3962 47066
rect 3962 47014 3964 47066
rect 3908 47012 3964 47014
rect 4012 47066 4068 47068
rect 4012 47014 4014 47066
rect 4014 47014 4066 47066
rect 4066 47014 4068 47066
rect 4012 47012 4068 47014
rect 4464 46282 4520 46284
rect 4464 46230 4466 46282
rect 4466 46230 4518 46282
rect 4518 46230 4520 46282
rect 4464 46228 4520 46230
rect 4568 46282 4624 46284
rect 4568 46230 4570 46282
rect 4570 46230 4622 46282
rect 4622 46230 4624 46282
rect 4568 46228 4624 46230
rect 4672 46282 4728 46284
rect 4672 46230 4674 46282
rect 4674 46230 4726 46282
rect 4726 46230 4728 46282
rect 4672 46228 4728 46230
rect 3804 45498 3860 45500
rect 3804 45446 3806 45498
rect 3806 45446 3858 45498
rect 3858 45446 3860 45498
rect 3804 45444 3860 45446
rect 3908 45498 3964 45500
rect 3908 45446 3910 45498
rect 3910 45446 3962 45498
rect 3962 45446 3964 45498
rect 3908 45444 3964 45446
rect 4012 45498 4068 45500
rect 4012 45446 4014 45498
rect 4014 45446 4066 45498
rect 4066 45446 4068 45498
rect 4012 45444 4068 45446
rect 4464 44714 4520 44716
rect 4464 44662 4466 44714
rect 4466 44662 4518 44714
rect 4518 44662 4520 44714
rect 4464 44660 4520 44662
rect 4568 44714 4624 44716
rect 4568 44662 4570 44714
rect 4570 44662 4622 44714
rect 4622 44662 4624 44714
rect 4568 44660 4624 44662
rect 4672 44714 4728 44716
rect 4672 44662 4674 44714
rect 4674 44662 4726 44714
rect 4726 44662 4728 44714
rect 4672 44660 4728 44662
rect 3804 43930 3860 43932
rect 3804 43878 3806 43930
rect 3806 43878 3858 43930
rect 3858 43878 3860 43930
rect 3804 43876 3860 43878
rect 3908 43930 3964 43932
rect 3908 43878 3910 43930
rect 3910 43878 3962 43930
rect 3962 43878 3964 43930
rect 3908 43876 3964 43878
rect 4012 43930 4068 43932
rect 4012 43878 4014 43930
rect 4014 43878 4066 43930
rect 4066 43878 4068 43930
rect 4012 43876 4068 43878
rect 3500 43596 3556 43652
rect 3612 43708 3668 43764
rect 1596 43426 1652 43428
rect 1596 43374 1598 43426
rect 1598 43374 1650 43426
rect 1650 43374 1652 43426
rect 1596 43372 1652 43374
rect 924 42812 980 42868
rect 1820 42476 1876 42532
rect 2156 42028 2212 42084
rect 1596 41858 1652 41860
rect 1596 41806 1598 41858
rect 1598 41806 1650 41858
rect 1650 41806 1652 41858
rect 1596 41804 1652 41806
rect 1148 41468 1204 41524
rect 2044 41298 2100 41300
rect 2044 41246 2046 41298
rect 2046 41246 2098 41298
rect 2098 41246 2100 41298
rect 2044 41244 2100 41246
rect 924 40124 980 40180
rect 812 40012 868 40068
rect 1484 41074 1540 41076
rect 1484 41022 1486 41074
rect 1486 41022 1538 41074
rect 1538 41022 1540 41074
rect 1484 41020 1540 41022
rect 4464 43146 4520 43148
rect 4464 43094 4466 43146
rect 4466 43094 4518 43146
rect 4518 43094 4520 43146
rect 4464 43092 4520 43094
rect 4568 43146 4624 43148
rect 4568 43094 4570 43146
rect 4570 43094 4622 43146
rect 4622 43094 4624 43146
rect 4568 43092 4624 43094
rect 4672 43146 4728 43148
rect 4672 43094 4674 43146
rect 4674 43094 4726 43146
rect 4726 43094 4728 43146
rect 4672 43092 4728 43094
rect 3804 42362 3860 42364
rect 3804 42310 3806 42362
rect 3806 42310 3858 42362
rect 3858 42310 3860 42362
rect 3804 42308 3860 42310
rect 3908 42362 3964 42364
rect 3908 42310 3910 42362
rect 3910 42310 3962 42362
rect 3962 42310 3964 42362
rect 3908 42308 3964 42310
rect 4012 42362 4068 42364
rect 4012 42310 4014 42362
rect 4014 42310 4066 42362
rect 4066 42310 4068 42362
rect 4012 42308 4068 42310
rect 2604 41804 2660 41860
rect 2492 41356 2548 41412
rect 2380 41244 2436 41300
rect 1708 40236 1764 40292
rect 2268 40236 2324 40292
rect 1932 40012 1988 40068
rect 1036 38780 1092 38836
rect 700 32956 756 33012
rect 812 36764 868 36820
rect 1036 37436 1092 37492
rect 924 36092 980 36148
rect 1036 37212 1092 37268
rect 1484 37324 1540 37380
rect 1596 37154 1652 37156
rect 1596 37102 1598 37154
rect 1598 37102 1650 37154
rect 1650 37102 1652 37154
rect 1596 37100 1652 37102
rect 1260 36764 1316 36820
rect 924 33404 980 33460
rect 1372 34748 1428 34804
rect 2044 39618 2100 39620
rect 2044 39566 2046 39618
rect 2046 39566 2098 39618
rect 2098 39566 2100 39618
rect 2044 39564 2100 39566
rect 1708 36706 1764 36708
rect 1708 36654 1710 36706
rect 1710 36654 1762 36706
rect 1762 36654 1764 36706
rect 1708 36652 1764 36654
rect 1708 36204 1764 36260
rect 1596 35586 1652 35588
rect 1596 35534 1598 35586
rect 1598 35534 1650 35586
rect 1650 35534 1652 35586
rect 1596 35532 1652 35534
rect 1932 36316 1988 36372
rect 1036 32060 1092 32116
rect 1260 32620 1316 32676
rect 812 30044 868 30100
rect 588 29260 644 29316
rect 1036 29372 1092 29428
rect 588 29036 644 29092
rect 1260 31612 1316 31668
rect 1260 30994 1316 30996
rect 1260 30942 1262 30994
rect 1262 30942 1314 30994
rect 1314 30942 1316 30994
rect 1260 30940 1316 30942
rect 1036 27580 1092 27636
rect 1260 30098 1316 30100
rect 1260 30046 1262 30098
rect 1262 30046 1314 30098
rect 1314 30046 1316 30098
rect 1260 30044 1316 30046
rect 1260 28476 1316 28532
rect 1148 27132 1204 27188
rect 1036 26684 1092 26740
rect 700 26572 756 26628
rect 1036 25340 1092 25396
rect 700 23100 756 23156
rect 924 23996 980 24052
rect 588 20412 644 20468
rect 700 22876 756 22932
rect 812 22652 868 22708
rect 1372 25564 1428 25620
rect 1596 33458 1652 33460
rect 1596 33406 1598 33458
rect 1598 33406 1650 33458
rect 1650 33406 1652 33458
rect 1596 33404 1652 33406
rect 1596 32956 1652 33012
rect 1708 32844 1764 32900
rect 1708 32674 1764 32676
rect 1708 32622 1710 32674
rect 1710 32622 1762 32674
rect 1762 32622 1764 32674
rect 1708 32620 1764 32622
rect 2156 33516 2212 33572
rect 1708 31612 1764 31668
rect 1820 30828 1876 30884
rect 1708 29314 1764 29316
rect 1708 29262 1710 29314
rect 1710 29262 1762 29314
rect 1762 29262 1764 29314
rect 1708 29260 1764 29262
rect 1596 28754 1652 28756
rect 1596 28702 1598 28754
rect 1598 28702 1650 28754
rect 1650 28702 1652 28754
rect 1596 28700 1652 28702
rect 4172 41858 4228 41860
rect 4172 41806 4174 41858
rect 4174 41806 4226 41858
rect 4226 41806 4228 41858
rect 4172 41804 4228 41806
rect 4464 41578 4520 41580
rect 4464 41526 4466 41578
rect 4466 41526 4518 41578
rect 4518 41526 4520 41578
rect 4464 41524 4520 41526
rect 4568 41578 4624 41580
rect 4568 41526 4570 41578
rect 4570 41526 4622 41578
rect 4622 41526 4624 41578
rect 4568 41524 4624 41526
rect 4672 41578 4728 41580
rect 4672 41526 4674 41578
rect 4674 41526 4726 41578
rect 4726 41526 4728 41578
rect 4672 41524 4728 41526
rect 4284 41298 4340 41300
rect 4284 41246 4286 41298
rect 4286 41246 4338 41298
rect 4338 41246 4340 41298
rect 4284 41244 4340 41246
rect 3500 41020 3556 41076
rect 2492 37378 2548 37380
rect 2492 37326 2494 37378
rect 2494 37326 2546 37378
rect 2546 37326 2548 37378
rect 2492 37324 2548 37326
rect 3052 40290 3108 40292
rect 3052 40238 3054 40290
rect 3054 40238 3106 40290
rect 3106 40238 3108 40290
rect 3052 40236 3108 40238
rect 2940 39564 2996 39620
rect 2940 38892 2996 38948
rect 2716 38834 2772 38836
rect 2716 38782 2718 38834
rect 2718 38782 2770 38834
rect 2770 38782 2772 38834
rect 2716 38780 2772 38782
rect 3276 37772 3332 37828
rect 2716 36764 2772 36820
rect 2828 36876 2884 36932
rect 2828 36652 2884 36708
rect 2940 36764 2996 36820
rect 2604 35196 2660 35252
rect 2044 32844 2100 32900
rect 1820 27580 1876 27636
rect 1708 27132 1764 27188
rect 1708 26908 1764 26964
rect 1484 26124 1540 26180
rect 1596 25394 1652 25396
rect 1596 25342 1598 25394
rect 1598 25342 1650 25394
rect 1650 25342 1652 25394
rect 1596 25340 1652 25342
rect 2268 32060 2324 32116
rect 2380 31052 2436 31108
rect 2716 36540 2772 36596
rect 2716 33404 2772 33460
rect 2156 28700 2212 28756
rect 2268 27020 2324 27076
rect 2156 26066 2212 26068
rect 2156 26014 2158 26066
rect 2158 26014 2210 26066
rect 2210 26014 2212 26066
rect 2156 26012 2212 26014
rect 1372 24892 1428 24948
rect 1372 24108 1428 24164
rect 1148 22482 1204 22484
rect 1148 22430 1150 22482
rect 1150 22430 1202 22482
rect 1202 22430 1204 22482
rect 1148 22428 1204 22430
rect 1148 21308 1204 21364
rect 1036 20636 1092 20692
rect 700 17836 756 17892
rect 924 18620 980 18676
rect 700 17388 756 17444
rect 476 14364 532 14420
rect 588 15932 644 15988
rect 364 10780 420 10836
rect 476 13692 532 13748
rect 588 10668 644 10724
rect 476 4396 532 4452
rect 1596 23826 1652 23828
rect 1596 23774 1598 23826
rect 1598 23774 1650 23826
rect 1650 23774 1652 23826
rect 1596 23772 1652 23774
rect 1596 23324 1652 23380
rect 1708 22594 1764 22596
rect 1708 22542 1710 22594
rect 1710 22542 1762 22594
rect 1762 22542 1764 22594
rect 1708 22540 1764 22542
rect 1372 20914 1428 20916
rect 1372 20862 1374 20914
rect 1374 20862 1426 20914
rect 1426 20862 1428 20914
rect 1372 20860 1428 20862
rect 1260 20188 1316 20244
rect 1372 20412 1428 20468
rect 1148 16604 1204 16660
rect 1260 14476 1316 14532
rect 1148 13634 1204 13636
rect 1148 13582 1150 13634
rect 1150 13582 1202 13634
rect 1202 13582 1204 13634
rect 1148 13580 1204 13582
rect 1036 13468 1092 13524
rect 1260 13468 1316 13524
rect 1148 13244 1204 13300
rect 924 11900 980 11956
rect 1036 10668 1092 10724
rect 1036 9324 1092 9380
rect 1260 10556 1316 10612
rect 1260 9212 1316 9268
rect 1596 20524 1652 20580
rect 1596 20076 1652 20132
rect 1596 19628 1652 19684
rect 1596 19458 1652 19460
rect 1596 19406 1598 19458
rect 1598 19406 1650 19458
rect 1650 19406 1652 19458
rect 1596 19404 1652 19406
rect 1708 18396 1764 18452
rect 2044 25618 2100 25620
rect 2044 25566 2046 25618
rect 2046 25566 2098 25618
rect 2098 25566 2100 25618
rect 2044 25564 2100 25566
rect 2828 32060 2884 32116
rect 2828 31890 2884 31892
rect 2828 31838 2830 31890
rect 2830 31838 2882 31890
rect 2882 31838 2884 31890
rect 2828 31836 2884 31838
rect 3052 36540 3108 36596
rect 3388 36988 3444 37044
rect 3276 36316 3332 36372
rect 3164 35308 3220 35364
rect 3804 40794 3860 40796
rect 3804 40742 3806 40794
rect 3806 40742 3858 40794
rect 3858 40742 3860 40794
rect 3804 40740 3860 40742
rect 3908 40794 3964 40796
rect 3908 40742 3910 40794
rect 3910 40742 3962 40794
rect 3962 40742 3964 40794
rect 3908 40740 3964 40742
rect 4012 40794 4068 40796
rect 4012 40742 4014 40794
rect 4014 40742 4066 40794
rect 4066 40742 4068 40794
rect 4012 40740 4068 40742
rect 4284 40402 4340 40404
rect 4284 40350 4286 40402
rect 4286 40350 4338 40402
rect 4338 40350 4340 40402
rect 4284 40348 4340 40350
rect 4464 40010 4520 40012
rect 4464 39958 4466 40010
rect 4466 39958 4518 40010
rect 4518 39958 4520 40010
rect 4464 39956 4520 39958
rect 4568 40010 4624 40012
rect 4568 39958 4570 40010
rect 4570 39958 4622 40010
rect 4622 39958 4624 40010
rect 4568 39956 4624 39958
rect 4672 40010 4728 40012
rect 4672 39958 4674 40010
rect 4674 39958 4726 40010
rect 4726 39958 4728 40010
rect 4672 39956 4728 39958
rect 5068 39730 5124 39732
rect 5068 39678 5070 39730
rect 5070 39678 5122 39730
rect 5122 39678 5124 39730
rect 5068 39676 5124 39678
rect 3804 39226 3860 39228
rect 3804 39174 3806 39226
rect 3806 39174 3858 39226
rect 3858 39174 3860 39226
rect 3804 39172 3860 39174
rect 3908 39226 3964 39228
rect 3908 39174 3910 39226
rect 3910 39174 3962 39226
rect 3962 39174 3964 39226
rect 3908 39172 3964 39174
rect 4012 39226 4068 39228
rect 4012 39174 4014 39226
rect 4014 39174 4066 39226
rect 4066 39174 4068 39226
rect 4012 39172 4068 39174
rect 3612 38780 3668 38836
rect 4284 38722 4340 38724
rect 4284 38670 4286 38722
rect 4286 38670 4338 38722
rect 4338 38670 4340 38722
rect 4284 38668 4340 38670
rect 3836 38556 3892 38612
rect 4464 38442 4520 38444
rect 4464 38390 4466 38442
rect 4466 38390 4518 38442
rect 4518 38390 4520 38442
rect 4464 38388 4520 38390
rect 4568 38442 4624 38444
rect 4568 38390 4570 38442
rect 4570 38390 4622 38442
rect 4622 38390 4624 38442
rect 4568 38388 4624 38390
rect 4672 38442 4728 38444
rect 4672 38390 4674 38442
rect 4674 38390 4726 38442
rect 4726 38390 4728 38442
rect 4672 38388 4728 38390
rect 3804 37658 3860 37660
rect 3804 37606 3806 37658
rect 3806 37606 3858 37658
rect 3858 37606 3860 37658
rect 3804 37604 3860 37606
rect 3908 37658 3964 37660
rect 3908 37606 3910 37658
rect 3910 37606 3962 37658
rect 3962 37606 3964 37658
rect 3908 37604 3964 37606
rect 4012 37658 4068 37660
rect 4012 37606 4014 37658
rect 4014 37606 4066 37658
rect 4066 37606 4068 37658
rect 4012 37604 4068 37606
rect 3948 36988 4004 37044
rect 3500 36764 3556 36820
rect 3612 36876 3668 36932
rect 3612 36652 3668 36708
rect 3388 36204 3444 36260
rect 2716 30940 2772 30996
rect 2828 30268 2884 30324
rect 2716 29932 2772 29988
rect 2828 30044 2884 30100
rect 2604 29260 2660 29316
rect 2604 29036 2660 29092
rect 2716 28476 2772 28532
rect 3388 35868 3444 35924
rect 3388 35308 3444 35364
rect 3276 33570 3332 33572
rect 3276 33518 3278 33570
rect 3278 33518 3330 33570
rect 3330 33518 3332 33570
rect 3276 33516 3332 33518
rect 3500 35196 3556 35252
rect 3500 34076 3556 34132
rect 3804 36090 3860 36092
rect 3804 36038 3806 36090
rect 3806 36038 3858 36090
rect 3858 36038 3860 36090
rect 3804 36036 3860 36038
rect 3908 36090 3964 36092
rect 3908 36038 3910 36090
rect 3910 36038 3962 36090
rect 3962 36038 3964 36090
rect 3908 36036 3964 36038
rect 4012 36090 4068 36092
rect 4012 36038 4014 36090
rect 4014 36038 4066 36090
rect 4066 36038 4068 36090
rect 4012 36036 4068 36038
rect 3804 34522 3860 34524
rect 3804 34470 3806 34522
rect 3806 34470 3858 34522
rect 3858 34470 3860 34522
rect 3804 34468 3860 34470
rect 3908 34522 3964 34524
rect 3908 34470 3910 34522
rect 3910 34470 3962 34522
rect 3962 34470 3964 34522
rect 3908 34468 3964 34470
rect 4012 34522 4068 34524
rect 4012 34470 4014 34522
rect 4014 34470 4066 34522
rect 4066 34470 4068 34522
rect 4012 34468 4068 34470
rect 4844 37436 4900 37492
rect 4464 36874 4520 36876
rect 4464 36822 4466 36874
rect 4466 36822 4518 36874
rect 4518 36822 4520 36874
rect 4464 36820 4520 36822
rect 4568 36874 4624 36876
rect 4568 36822 4570 36874
rect 4570 36822 4622 36874
rect 4622 36822 4624 36874
rect 4568 36820 4624 36822
rect 4672 36874 4728 36876
rect 4672 36822 4674 36874
rect 4674 36822 4726 36874
rect 4726 36822 4728 36874
rect 4672 36820 4728 36822
rect 4464 35306 4520 35308
rect 4464 35254 4466 35306
rect 4466 35254 4518 35306
rect 4518 35254 4520 35306
rect 4464 35252 4520 35254
rect 4568 35306 4624 35308
rect 4568 35254 4570 35306
rect 4570 35254 4622 35306
rect 4622 35254 4624 35306
rect 4568 35252 4624 35254
rect 4672 35306 4728 35308
rect 4672 35254 4674 35306
rect 4674 35254 4726 35306
rect 4726 35254 4728 35306
rect 4672 35252 4728 35254
rect 4284 35084 4340 35140
rect 4284 34914 4340 34916
rect 4284 34862 4286 34914
rect 4286 34862 4338 34914
rect 4338 34862 4340 34914
rect 4284 34860 4340 34862
rect 4060 34188 4116 34244
rect 3836 33852 3892 33908
rect 3804 32954 3860 32956
rect 3804 32902 3806 32954
rect 3806 32902 3858 32954
rect 3858 32902 3860 32954
rect 3804 32900 3860 32902
rect 3908 32954 3964 32956
rect 3908 32902 3910 32954
rect 3910 32902 3962 32954
rect 3962 32902 3964 32954
rect 3908 32900 3964 32902
rect 4012 32954 4068 32956
rect 4012 32902 4014 32954
rect 4014 32902 4066 32954
rect 4066 32902 4068 32954
rect 4012 32900 4068 32902
rect 4464 33738 4520 33740
rect 4464 33686 4466 33738
rect 4466 33686 4518 33738
rect 4518 33686 4520 33738
rect 4464 33684 4520 33686
rect 4568 33738 4624 33740
rect 4568 33686 4570 33738
rect 4570 33686 4622 33738
rect 4622 33686 4624 33738
rect 4568 33684 4624 33686
rect 4672 33738 4728 33740
rect 4672 33686 4674 33738
rect 4674 33686 4726 33738
rect 4726 33686 4728 33738
rect 4672 33684 4728 33686
rect 4396 32620 4452 32676
rect 3724 31836 3780 31892
rect 4060 31778 4116 31780
rect 4060 31726 4062 31778
rect 4062 31726 4114 31778
rect 4114 31726 4116 31778
rect 4060 31724 4116 31726
rect 3612 31500 3668 31556
rect 3804 31386 3860 31388
rect 3804 31334 3806 31386
rect 3806 31334 3858 31386
rect 3858 31334 3860 31386
rect 3804 31332 3860 31334
rect 3908 31386 3964 31388
rect 3908 31334 3910 31386
rect 3910 31334 3962 31386
rect 3962 31334 3964 31386
rect 3908 31332 3964 31334
rect 4012 31386 4068 31388
rect 4012 31334 4014 31386
rect 4014 31334 4066 31386
rect 4066 31334 4068 31386
rect 4012 31332 4068 31334
rect 3500 30994 3556 30996
rect 3500 30942 3502 30994
rect 3502 30942 3554 30994
rect 3554 30942 3556 30994
rect 3500 30940 3556 30942
rect 3164 30434 3220 30436
rect 3164 30382 3166 30434
rect 3166 30382 3218 30434
rect 3218 30382 3220 30434
rect 3164 30380 3220 30382
rect 3164 30156 3220 30212
rect 3164 27580 3220 27636
rect 3388 30380 3444 30436
rect 3500 30716 3556 30772
rect 3948 30044 4004 30100
rect 3804 29818 3860 29820
rect 3804 29766 3806 29818
rect 3806 29766 3858 29818
rect 3858 29766 3860 29818
rect 3804 29764 3860 29766
rect 3908 29818 3964 29820
rect 3908 29766 3910 29818
rect 3910 29766 3962 29818
rect 3962 29766 3964 29818
rect 3908 29764 3964 29766
rect 4012 29818 4068 29820
rect 4012 29766 4014 29818
rect 4014 29766 4066 29818
rect 4066 29766 4068 29818
rect 4012 29764 4068 29766
rect 3724 29538 3780 29540
rect 3724 29486 3726 29538
rect 3726 29486 3778 29538
rect 3778 29486 3780 29538
rect 3724 29484 3780 29486
rect 3500 28530 3556 28532
rect 3500 28478 3502 28530
rect 3502 28478 3554 28530
rect 3554 28478 3556 28530
rect 3500 28476 3556 28478
rect 3388 28028 3444 28084
rect 3052 27132 3108 27188
rect 2940 26460 2996 26516
rect 2828 26236 2884 26292
rect 2828 26012 2884 26068
rect 2268 24668 2324 24724
rect 2380 23996 2436 24052
rect 2380 23772 2436 23828
rect 2268 23436 2324 23492
rect 2156 21756 2212 21812
rect 2716 23100 2772 23156
rect 2044 21644 2100 21700
rect 1708 18060 1764 18116
rect 1596 17778 1652 17780
rect 1596 17726 1598 17778
rect 1598 17726 1650 17778
rect 1650 17726 1652 17778
rect 1596 17724 1652 17726
rect 2044 20972 2100 21028
rect 2156 21532 2212 21588
rect 1932 20914 1988 20916
rect 1932 20862 1934 20914
rect 1934 20862 1986 20914
rect 1986 20862 1988 20914
rect 1932 20860 1988 20862
rect 2044 20130 2100 20132
rect 2044 20078 2046 20130
rect 2046 20078 2098 20130
rect 2098 20078 2100 20130
rect 2044 20076 2100 20078
rect 1932 19964 1988 20020
rect 2044 18172 2100 18228
rect 1708 16604 1764 16660
rect 2268 20972 2324 21028
rect 2156 17724 2212 17780
rect 2268 19068 2324 19124
rect 3052 25730 3108 25732
rect 3052 25678 3054 25730
rect 3054 25678 3106 25730
rect 3106 25678 3108 25730
rect 3052 25676 3108 25678
rect 3052 25228 3108 25284
rect 2492 21868 2548 21924
rect 2940 25004 2996 25060
rect 2604 21586 2660 21588
rect 2604 21534 2606 21586
rect 2606 21534 2658 21586
rect 2658 21534 2660 21586
rect 2604 21532 2660 21534
rect 2492 20748 2548 20804
rect 2828 21756 2884 21812
rect 2940 20748 2996 20804
rect 3388 27074 3444 27076
rect 3388 27022 3390 27074
rect 3390 27022 3442 27074
rect 3442 27022 3444 27074
rect 3388 27020 3444 27022
rect 3276 25452 3332 25508
rect 3804 28250 3860 28252
rect 3804 28198 3806 28250
rect 3806 28198 3858 28250
rect 3858 28198 3860 28250
rect 3804 28196 3860 28198
rect 3908 28250 3964 28252
rect 3908 28198 3910 28250
rect 3910 28198 3962 28250
rect 3962 28198 3964 28250
rect 3908 28196 3964 28198
rect 4012 28250 4068 28252
rect 4012 28198 4014 28250
rect 4014 28198 4066 28250
rect 4066 28198 4068 28250
rect 4012 28196 4068 28198
rect 4464 32170 4520 32172
rect 4464 32118 4466 32170
rect 4466 32118 4518 32170
rect 4518 32118 4520 32170
rect 4464 32116 4520 32118
rect 4568 32170 4624 32172
rect 4568 32118 4570 32170
rect 4570 32118 4622 32170
rect 4622 32118 4624 32170
rect 4568 32116 4624 32118
rect 4672 32170 4728 32172
rect 4672 32118 4674 32170
rect 4674 32118 4726 32170
rect 4726 32118 4728 32170
rect 4672 32116 4728 32118
rect 5068 36652 5124 36708
rect 5180 37548 5236 37604
rect 5068 36258 5124 36260
rect 5068 36206 5070 36258
rect 5070 36206 5122 36258
rect 5122 36206 5124 36258
rect 5068 36204 5124 36206
rect 4956 35084 5012 35140
rect 4396 31106 4452 31108
rect 4396 31054 4398 31106
rect 4398 31054 4450 31106
rect 4450 31054 4452 31106
rect 4396 31052 4452 31054
rect 4732 31724 4788 31780
rect 4844 31612 4900 31668
rect 4620 30940 4676 30996
rect 4844 31164 4900 31220
rect 4396 30828 4452 30884
rect 4464 30602 4520 30604
rect 4464 30550 4466 30602
rect 4466 30550 4518 30602
rect 4518 30550 4520 30602
rect 4464 30548 4520 30550
rect 4568 30602 4624 30604
rect 4568 30550 4570 30602
rect 4570 30550 4622 30602
rect 4622 30550 4624 30602
rect 4568 30548 4624 30550
rect 4672 30602 4728 30604
rect 4672 30550 4674 30602
rect 4674 30550 4726 30602
rect 4726 30550 4728 30602
rect 4672 30548 4728 30550
rect 4464 29034 4520 29036
rect 4464 28982 4466 29034
rect 4466 28982 4518 29034
rect 4518 28982 4520 29034
rect 4464 28980 4520 28982
rect 4568 29034 4624 29036
rect 4568 28982 4570 29034
rect 4570 28982 4622 29034
rect 4622 28982 4624 29034
rect 4568 28980 4624 28982
rect 4672 29034 4728 29036
rect 4672 28982 4674 29034
rect 4674 28982 4726 29034
rect 4726 28982 4728 29034
rect 4672 28980 4728 28982
rect 4732 28476 4788 28532
rect 4284 27858 4340 27860
rect 4284 27806 4286 27858
rect 4286 27806 4338 27858
rect 4338 27806 4340 27858
rect 4284 27804 4340 27806
rect 5068 34802 5124 34804
rect 5068 34750 5070 34802
rect 5070 34750 5122 34802
rect 5122 34750 5124 34802
rect 5068 34748 5124 34750
rect 5180 34130 5236 34132
rect 5180 34078 5182 34130
rect 5182 34078 5234 34130
rect 5234 34078 5236 34130
rect 5180 34076 5236 34078
rect 5180 33628 5236 33684
rect 5068 31500 5124 31556
rect 5180 32956 5236 33012
rect 5068 29484 5124 29540
rect 5068 29036 5124 29092
rect 4172 27132 4228 27188
rect 3724 26962 3780 26964
rect 3724 26910 3726 26962
rect 3726 26910 3778 26962
rect 3778 26910 3780 26962
rect 3724 26908 3780 26910
rect 3804 26682 3860 26684
rect 3804 26630 3806 26682
rect 3806 26630 3858 26682
rect 3858 26630 3860 26682
rect 3804 26628 3860 26630
rect 3908 26682 3964 26684
rect 3908 26630 3910 26682
rect 3910 26630 3962 26682
rect 3962 26630 3964 26682
rect 3908 26628 3964 26630
rect 4012 26682 4068 26684
rect 4012 26630 4014 26682
rect 4014 26630 4066 26682
rect 4066 26630 4068 26682
rect 4012 26628 4068 26630
rect 4464 27466 4520 27468
rect 4464 27414 4466 27466
rect 4466 27414 4518 27466
rect 4518 27414 4520 27466
rect 4464 27412 4520 27414
rect 4568 27466 4624 27468
rect 4568 27414 4570 27466
rect 4570 27414 4622 27466
rect 4622 27414 4624 27466
rect 4568 27412 4624 27414
rect 4672 27466 4728 27468
rect 4672 27414 4674 27466
rect 4674 27414 4726 27466
rect 4726 27414 4728 27466
rect 4672 27412 4728 27414
rect 4956 27356 5012 27412
rect 4956 26908 5012 26964
rect 4284 26572 4340 26628
rect 4396 26796 4452 26852
rect 3724 25676 3780 25732
rect 3612 25340 3668 25396
rect 3276 25004 3332 25060
rect 3500 25228 3556 25284
rect 4464 25898 4520 25900
rect 4464 25846 4466 25898
rect 4466 25846 4518 25898
rect 4518 25846 4520 25898
rect 4464 25844 4520 25846
rect 4568 25898 4624 25900
rect 4568 25846 4570 25898
rect 4570 25846 4622 25898
rect 4622 25846 4624 25898
rect 4568 25844 4624 25846
rect 4672 25898 4728 25900
rect 4672 25846 4674 25898
rect 4674 25846 4726 25898
rect 4726 25846 4728 25898
rect 4672 25844 4728 25846
rect 3804 25114 3860 25116
rect 3804 25062 3806 25114
rect 3806 25062 3858 25114
rect 3858 25062 3860 25114
rect 3804 25060 3860 25062
rect 3908 25114 3964 25116
rect 3908 25062 3910 25114
rect 3910 25062 3962 25114
rect 3962 25062 3964 25114
rect 3908 25060 3964 25062
rect 4012 25114 4068 25116
rect 4012 25062 4014 25114
rect 4014 25062 4066 25114
rect 4066 25062 4068 25114
rect 4012 25060 4068 25062
rect 3276 22540 3332 22596
rect 3164 21868 3220 21924
rect 3276 20914 3332 20916
rect 3276 20862 3278 20914
rect 3278 20862 3330 20914
rect 3330 20862 3332 20914
rect 3276 20860 3332 20862
rect 2604 19404 2660 19460
rect 2716 19628 2772 19684
rect 2716 19292 2772 19348
rect 2492 18060 2548 18116
rect 2604 18396 2660 18452
rect 3388 19292 3444 19348
rect 3164 19122 3220 19124
rect 3164 19070 3166 19122
rect 3166 19070 3218 19122
rect 3218 19070 3220 19122
rect 3164 19068 3220 19070
rect 3164 18450 3220 18452
rect 3164 18398 3166 18450
rect 3166 18398 3218 18450
rect 3218 18398 3220 18450
rect 3164 18396 3220 18398
rect 4060 24444 4116 24500
rect 3612 23436 3668 23492
rect 3804 23546 3860 23548
rect 3804 23494 3806 23546
rect 3806 23494 3858 23546
rect 3858 23494 3860 23546
rect 3804 23492 3860 23494
rect 3908 23546 3964 23548
rect 3908 23494 3910 23546
rect 3910 23494 3962 23546
rect 3962 23494 3964 23546
rect 3908 23492 3964 23494
rect 4012 23546 4068 23548
rect 4012 23494 4014 23546
rect 4014 23494 4066 23546
rect 4066 23494 4068 23546
rect 4012 23492 4068 23494
rect 5180 28476 5236 28532
rect 6524 52220 6580 52276
rect 5740 49644 5796 49700
rect 5516 38834 5572 38836
rect 5516 38782 5518 38834
rect 5518 38782 5570 38834
rect 5570 38782 5572 38834
rect 5516 38780 5572 38782
rect 5516 37548 5572 37604
rect 5516 36652 5572 36708
rect 5516 36204 5572 36260
rect 5404 34914 5460 34916
rect 5404 34862 5406 34914
rect 5406 34862 5458 34914
rect 5458 34862 5460 34914
rect 5404 34860 5460 34862
rect 5404 29036 5460 29092
rect 6076 48860 6132 48916
rect 5852 39900 5908 39956
rect 6188 39900 6244 39956
rect 5964 38892 6020 38948
rect 6300 39452 6356 39508
rect 5852 35810 5908 35812
rect 5852 35758 5854 35810
rect 5854 35758 5906 35810
rect 5906 35758 5908 35810
rect 5852 35756 5908 35758
rect 5740 35308 5796 35364
rect 6636 51324 6692 51380
rect 7420 48860 7476 48916
rect 7084 48188 7140 48244
rect 6636 40572 6692 40628
rect 6972 40514 7028 40516
rect 6972 40462 6974 40514
rect 6974 40462 7026 40514
rect 7026 40462 7028 40514
rect 6972 40460 7028 40462
rect 6636 39452 6692 39508
rect 6748 39004 6804 39060
rect 5852 34412 5908 34468
rect 5628 32956 5684 33012
rect 5852 30210 5908 30212
rect 5852 30158 5854 30210
rect 5854 30158 5906 30210
rect 5906 30158 5908 30210
rect 5852 30156 5908 30158
rect 5292 27858 5348 27860
rect 5292 27806 5294 27858
rect 5294 27806 5346 27858
rect 5346 27806 5348 27858
rect 5292 27804 5348 27806
rect 4956 24444 5012 24500
rect 4464 24330 4520 24332
rect 4464 24278 4466 24330
rect 4466 24278 4518 24330
rect 4518 24278 4520 24330
rect 4464 24276 4520 24278
rect 4568 24330 4624 24332
rect 4568 24278 4570 24330
rect 4570 24278 4622 24330
rect 4622 24278 4624 24330
rect 4568 24276 4624 24278
rect 4672 24330 4728 24332
rect 4672 24278 4674 24330
rect 4674 24278 4726 24330
rect 4726 24278 4728 24330
rect 4672 24276 4728 24278
rect 4284 23884 4340 23940
rect 4620 23996 4676 24052
rect 4284 23548 4340 23604
rect 3804 21978 3860 21980
rect 3804 21926 3806 21978
rect 3806 21926 3858 21978
rect 3858 21926 3860 21978
rect 3804 21924 3860 21926
rect 3908 21978 3964 21980
rect 3908 21926 3910 21978
rect 3910 21926 3962 21978
rect 3962 21926 3964 21978
rect 3908 21924 3964 21926
rect 4012 21978 4068 21980
rect 4012 21926 4014 21978
rect 4014 21926 4066 21978
rect 4066 21926 4068 21978
rect 4012 21924 4068 21926
rect 3804 20410 3860 20412
rect 3804 20358 3806 20410
rect 3806 20358 3858 20410
rect 3858 20358 3860 20410
rect 3804 20356 3860 20358
rect 3908 20410 3964 20412
rect 3908 20358 3910 20410
rect 3910 20358 3962 20410
rect 3962 20358 3964 20410
rect 3908 20356 3964 20358
rect 4012 20410 4068 20412
rect 4012 20358 4014 20410
rect 4014 20358 4066 20410
rect 4066 20358 4068 20410
rect 4012 20356 4068 20358
rect 3836 20076 3892 20132
rect 3612 19068 3668 19124
rect 4464 22762 4520 22764
rect 4464 22710 4466 22762
rect 4466 22710 4518 22762
rect 4518 22710 4520 22762
rect 4464 22708 4520 22710
rect 4568 22762 4624 22764
rect 4568 22710 4570 22762
rect 4570 22710 4622 22762
rect 4622 22710 4624 22762
rect 4568 22708 4624 22710
rect 4672 22762 4728 22764
rect 4672 22710 4674 22762
rect 4674 22710 4726 22762
rect 4726 22710 4728 22762
rect 4672 22708 4728 22710
rect 4284 21810 4340 21812
rect 4284 21758 4286 21810
rect 4286 21758 4338 21810
rect 4338 21758 4340 21810
rect 4284 21756 4340 21758
rect 4464 21194 4520 21196
rect 4464 21142 4466 21194
rect 4466 21142 4518 21194
rect 4518 21142 4520 21194
rect 4464 21140 4520 21142
rect 4568 21194 4624 21196
rect 4568 21142 4570 21194
rect 4570 21142 4622 21194
rect 4622 21142 4624 21194
rect 4568 21140 4624 21142
rect 4672 21194 4728 21196
rect 4672 21142 4674 21194
rect 4674 21142 4726 21194
rect 4726 21142 4728 21194
rect 4672 21140 4728 21142
rect 4172 20076 4228 20132
rect 4508 19964 4564 20020
rect 4464 19626 4520 19628
rect 4464 19574 4466 19626
rect 4466 19574 4518 19626
rect 4518 19574 4520 19626
rect 4464 19572 4520 19574
rect 4568 19626 4624 19628
rect 4568 19574 4570 19626
rect 4570 19574 4622 19626
rect 4622 19574 4624 19626
rect 4568 19572 4624 19574
rect 4672 19626 4728 19628
rect 4672 19574 4674 19626
rect 4674 19574 4726 19626
rect 4726 19574 4728 19626
rect 4672 19572 4728 19574
rect 4508 19346 4564 19348
rect 4508 19294 4510 19346
rect 4510 19294 4562 19346
rect 4562 19294 4564 19346
rect 4508 19292 4564 19294
rect 3836 18956 3892 19012
rect 3500 18620 3556 18676
rect 3612 18844 3668 18900
rect 3804 18842 3860 18844
rect 3804 18790 3806 18842
rect 3806 18790 3858 18842
rect 3858 18790 3860 18842
rect 3804 18788 3860 18790
rect 3908 18842 3964 18844
rect 3908 18790 3910 18842
rect 3910 18790 3962 18842
rect 3962 18790 3964 18842
rect 3908 18788 3964 18790
rect 4012 18842 4068 18844
rect 4012 18790 4014 18842
rect 4014 18790 4066 18842
rect 4066 18790 4068 18842
rect 4012 18788 4068 18790
rect 4284 18844 4340 18900
rect 4172 18620 4228 18676
rect 2492 17612 2548 17668
rect 2268 16604 2324 16660
rect 1932 15874 1988 15876
rect 1932 15822 1934 15874
rect 1934 15822 1986 15874
rect 1986 15822 1988 15874
rect 1932 15820 1988 15822
rect 1708 15708 1764 15764
rect 2156 15708 2212 15764
rect 1484 15036 1540 15092
rect 1932 15090 1988 15092
rect 1932 15038 1934 15090
rect 1934 15038 1986 15090
rect 1986 15038 1988 15090
rect 1932 15036 1988 15038
rect 2044 14924 2100 14980
rect 1820 14812 1876 14868
rect 1708 14588 1764 14644
rect 1596 13804 1652 13860
rect 1932 14530 1988 14532
rect 1932 14478 1934 14530
rect 1934 14478 1986 14530
rect 1986 14478 1988 14530
rect 1932 14476 1988 14478
rect 1932 13746 1988 13748
rect 1932 13694 1934 13746
rect 1934 13694 1986 13746
rect 1986 13694 1988 13746
rect 1932 13692 1988 13694
rect 1932 12178 1988 12180
rect 1932 12126 1934 12178
rect 1934 12126 1986 12178
rect 1986 12126 1988 12178
rect 1932 12124 1988 12126
rect 1596 11340 1652 11396
rect 1596 10780 1652 10836
rect 2156 13692 2212 13748
rect 2156 13244 2212 13300
rect 2268 12124 2324 12180
rect 2268 11564 2324 11620
rect 2604 15820 2660 15876
rect 2492 14642 2548 14644
rect 2492 14590 2494 14642
rect 2494 14590 2546 14642
rect 2546 14590 2548 14642
rect 2492 14588 2548 14590
rect 2492 13916 2548 13972
rect 2828 16604 2884 16660
rect 2940 16828 2996 16884
rect 2828 15148 2884 15204
rect 2492 12066 2548 12068
rect 2492 12014 2494 12066
rect 2494 12014 2546 12066
rect 2546 12014 2548 12066
rect 2492 12012 2548 12014
rect 2156 10444 2212 10500
rect 1484 9324 1540 9380
rect 1596 9548 1652 9604
rect 812 8204 868 8260
rect 1036 7868 1092 7924
rect 1036 3836 1092 3892
rect 2044 9100 2100 9156
rect 1596 8258 1652 8260
rect 1596 8206 1598 8258
rect 1598 8206 1650 8258
rect 1650 8206 1652 8258
rect 1596 8204 1652 8206
rect 3052 16268 3108 16324
rect 3276 16994 3332 16996
rect 3276 16942 3278 16994
rect 3278 16942 3330 16994
rect 3330 16942 3332 16994
rect 3276 16940 3332 16942
rect 3052 16044 3108 16100
rect 3052 15202 3108 15204
rect 3052 15150 3054 15202
rect 3054 15150 3106 15202
rect 3106 15150 3108 15202
rect 3052 15148 3108 15150
rect 3836 18226 3892 18228
rect 3836 18174 3838 18226
rect 3838 18174 3890 18226
rect 3890 18174 3892 18226
rect 3836 18172 3892 18174
rect 3724 17890 3780 17892
rect 3724 17838 3726 17890
rect 3726 17838 3778 17890
rect 3778 17838 3780 17890
rect 3724 17836 3780 17838
rect 3500 16098 3556 16100
rect 3500 16046 3502 16098
rect 3502 16046 3554 16098
rect 3554 16046 3556 16098
rect 3500 16044 3556 16046
rect 3612 17612 3668 17668
rect 3804 17274 3860 17276
rect 3804 17222 3806 17274
rect 3806 17222 3858 17274
rect 3858 17222 3860 17274
rect 3804 17220 3860 17222
rect 3908 17274 3964 17276
rect 3908 17222 3910 17274
rect 3910 17222 3962 17274
rect 3962 17222 3964 17274
rect 3908 17220 3964 17222
rect 4012 17274 4068 17276
rect 4012 17222 4014 17274
rect 4014 17222 4066 17274
rect 4066 17222 4068 17274
rect 4012 17220 4068 17222
rect 3836 16882 3892 16884
rect 3836 16830 3838 16882
rect 3838 16830 3890 16882
rect 3890 16830 3892 16882
rect 3836 16828 3892 16830
rect 3804 15706 3860 15708
rect 3804 15654 3806 15706
rect 3806 15654 3858 15706
rect 3858 15654 3860 15706
rect 3804 15652 3860 15654
rect 3908 15706 3964 15708
rect 3908 15654 3910 15706
rect 3910 15654 3962 15706
rect 3962 15654 3964 15706
rect 3908 15652 3964 15654
rect 4012 15706 4068 15708
rect 4012 15654 4014 15706
rect 4014 15654 4066 15706
rect 4066 15654 4068 15706
rect 4012 15652 4068 15654
rect 3276 15148 3332 15204
rect 2492 8930 2548 8932
rect 2492 8878 2494 8930
rect 2494 8878 2546 8930
rect 2546 8878 2548 8930
rect 2492 8876 2548 8878
rect 1260 6578 1316 6580
rect 1260 6526 1262 6578
rect 1262 6526 1314 6578
rect 1314 6526 1316 6578
rect 1260 6524 1316 6526
rect 3276 14700 3332 14756
rect 3388 13580 3444 13636
rect 3276 12348 3332 12404
rect 3276 11452 3332 11508
rect 2940 11228 2996 11284
rect 3164 11116 3220 11172
rect 4396 18450 4452 18452
rect 4396 18398 4398 18450
rect 4398 18398 4450 18450
rect 4450 18398 4452 18450
rect 4396 18396 4452 18398
rect 4464 18058 4520 18060
rect 4464 18006 4466 18058
rect 4466 18006 4518 18058
rect 4518 18006 4520 18058
rect 4464 18004 4520 18006
rect 4568 18058 4624 18060
rect 4568 18006 4570 18058
rect 4570 18006 4622 18058
rect 4622 18006 4624 18058
rect 4568 18004 4624 18006
rect 4672 18058 4728 18060
rect 4672 18006 4674 18058
rect 4674 18006 4726 18058
rect 4726 18006 4728 18058
rect 4672 18004 4728 18006
rect 4284 17724 4340 17780
rect 4620 17836 4676 17892
rect 4844 17890 4900 17892
rect 4844 17838 4846 17890
rect 4846 17838 4898 17890
rect 4898 17838 4900 17890
rect 4844 17836 4900 17838
rect 5516 28642 5572 28644
rect 5516 28590 5518 28642
rect 5518 28590 5570 28642
rect 5570 28590 5572 28642
rect 5516 28588 5572 28590
rect 5404 27298 5460 27300
rect 5404 27246 5406 27298
rect 5406 27246 5458 27298
rect 5458 27246 5460 27298
rect 5404 27244 5460 27246
rect 5516 27132 5572 27188
rect 5740 27858 5796 27860
rect 5740 27806 5742 27858
rect 5742 27806 5794 27858
rect 5794 27806 5796 27858
rect 5740 27804 5796 27806
rect 5404 24892 5460 24948
rect 5516 24668 5572 24724
rect 5740 26684 5796 26740
rect 5068 21084 5124 21140
rect 5404 23938 5460 23940
rect 5404 23886 5406 23938
rect 5406 23886 5458 23938
rect 5458 23886 5460 23938
rect 5404 23884 5460 23886
rect 5404 22316 5460 22372
rect 5292 21756 5348 21812
rect 6300 35308 6356 35364
rect 6300 34748 6356 34804
rect 6076 33570 6132 33572
rect 6076 33518 6078 33570
rect 6078 33518 6130 33570
rect 6130 33518 6132 33570
rect 6076 33516 6132 33518
rect 6300 30828 6356 30884
rect 7196 39058 7252 39060
rect 7196 39006 7198 39058
rect 7198 39006 7250 39058
rect 7250 39006 7252 39058
rect 7196 39004 7252 39006
rect 15484 56252 15540 56308
rect 16492 56306 16548 56308
rect 16492 56254 16494 56306
rect 16494 56254 16546 56306
rect 16546 56254 16548 56306
rect 16492 56252 16548 56254
rect 11564 55356 11620 55412
rect 9996 54572 10052 54628
rect 10892 54348 10948 54404
rect 9212 54012 9268 54068
rect 7644 40572 7700 40628
rect 7532 39900 7588 39956
rect 8988 41132 9044 41188
rect 8652 40572 8708 40628
rect 8092 39676 8148 39732
rect 7756 38444 7812 38500
rect 7420 37772 7476 37828
rect 6524 37100 6580 37156
rect 6748 35868 6804 35924
rect 6972 37100 7028 37156
rect 7532 37154 7588 37156
rect 7532 37102 7534 37154
rect 7534 37102 7586 37154
rect 7586 37102 7588 37154
rect 7532 37100 7588 37102
rect 6636 34972 6692 35028
rect 6524 33516 6580 33572
rect 6636 34300 6692 34356
rect 6524 31500 6580 31556
rect 5964 27244 6020 27300
rect 5964 26684 6020 26740
rect 6076 27132 6132 27188
rect 5964 26236 6020 26292
rect 5964 25564 6020 25620
rect 6748 32562 6804 32564
rect 6748 32510 6750 32562
rect 6750 32510 6802 32562
rect 6802 32510 6804 32562
rect 6748 32508 6804 32510
rect 6636 30828 6692 30884
rect 6636 30044 6692 30100
rect 6636 28530 6692 28532
rect 6636 28478 6638 28530
rect 6638 28478 6690 28530
rect 6690 28478 6692 28530
rect 6636 28476 6692 28478
rect 6300 26908 6356 26964
rect 6412 28364 6468 28420
rect 6300 26572 6356 26628
rect 6300 26236 6356 26292
rect 6300 25506 6356 25508
rect 6300 25454 6302 25506
rect 6302 25454 6354 25506
rect 6354 25454 6356 25506
rect 6300 25452 6356 25454
rect 6188 24834 6244 24836
rect 6188 24782 6190 24834
rect 6190 24782 6242 24834
rect 6242 24782 6244 24834
rect 6188 24780 6244 24782
rect 6300 23324 6356 23380
rect 5292 21084 5348 21140
rect 5740 22370 5796 22372
rect 5740 22318 5742 22370
rect 5742 22318 5794 22370
rect 5794 22318 5796 22370
rect 5740 22316 5796 22318
rect 5180 18508 5236 18564
rect 5628 20860 5684 20916
rect 5964 21362 6020 21364
rect 5964 21310 5966 21362
rect 5966 21310 6018 21362
rect 6018 21310 6020 21362
rect 5964 21308 6020 21310
rect 6188 23154 6244 23156
rect 6188 23102 6190 23154
rect 6190 23102 6242 23154
rect 6242 23102 6244 23154
rect 6188 23100 6244 23102
rect 6300 21698 6356 21700
rect 6300 21646 6302 21698
rect 6302 21646 6354 21698
rect 6354 21646 6356 21698
rect 6300 21644 6356 21646
rect 6300 20972 6356 21028
rect 5740 19964 5796 20020
rect 5852 20748 5908 20804
rect 5404 17836 5460 17892
rect 5740 19458 5796 19460
rect 5740 19406 5742 19458
rect 5742 19406 5794 19458
rect 5794 19406 5796 19458
rect 5740 19404 5796 19406
rect 6188 20802 6244 20804
rect 6188 20750 6190 20802
rect 6190 20750 6242 20802
rect 6242 20750 6244 20802
rect 6188 20748 6244 20750
rect 6188 20130 6244 20132
rect 6188 20078 6190 20130
rect 6190 20078 6242 20130
rect 6242 20078 6244 20130
rect 6188 20076 6244 20078
rect 5964 19292 6020 19348
rect 5516 18396 5572 18452
rect 5516 17388 5572 17444
rect 4956 16882 5012 16884
rect 4956 16830 4958 16882
rect 4958 16830 5010 16882
rect 5010 16830 5012 16882
rect 4956 16828 5012 16830
rect 4464 16490 4520 16492
rect 4464 16438 4466 16490
rect 4466 16438 4518 16490
rect 4518 16438 4520 16490
rect 4464 16436 4520 16438
rect 4568 16490 4624 16492
rect 4568 16438 4570 16490
rect 4570 16438 4622 16490
rect 4622 16438 4624 16490
rect 4568 16436 4624 16438
rect 4672 16490 4728 16492
rect 4672 16438 4674 16490
rect 4674 16438 4726 16490
rect 4726 16438 4728 16490
rect 4672 16436 4728 16438
rect 4284 16268 4340 16324
rect 4732 16210 4788 16212
rect 4732 16158 4734 16210
rect 4734 16158 4786 16210
rect 4786 16158 4788 16210
rect 4732 16156 4788 16158
rect 4284 16098 4340 16100
rect 4284 16046 4286 16098
rect 4286 16046 4338 16098
rect 4338 16046 4340 16098
rect 4284 16044 4340 16046
rect 3804 14138 3860 14140
rect 3804 14086 3806 14138
rect 3806 14086 3858 14138
rect 3858 14086 3860 14138
rect 3804 14084 3860 14086
rect 3908 14138 3964 14140
rect 3908 14086 3910 14138
rect 3910 14086 3962 14138
rect 3962 14086 3964 14138
rect 3908 14084 3964 14086
rect 4012 14138 4068 14140
rect 4012 14086 4014 14138
rect 4014 14086 4066 14138
rect 4066 14086 4068 14138
rect 4012 14084 4068 14086
rect 4172 14140 4228 14196
rect 4464 14922 4520 14924
rect 4464 14870 4466 14922
rect 4466 14870 4518 14922
rect 4518 14870 4520 14922
rect 4464 14868 4520 14870
rect 4568 14922 4624 14924
rect 4568 14870 4570 14922
rect 4570 14870 4622 14922
rect 4622 14870 4624 14922
rect 4568 14868 4624 14870
rect 4672 14922 4728 14924
rect 4672 14870 4674 14922
rect 4674 14870 4726 14922
rect 4726 14870 4728 14922
rect 4672 14868 4728 14870
rect 5180 16716 5236 16772
rect 4508 14140 4564 14196
rect 4844 14252 4900 14308
rect 4284 13916 4340 13972
rect 4284 13746 4340 13748
rect 4284 13694 4286 13746
rect 4286 13694 4338 13746
rect 4338 13694 4340 13746
rect 4284 13692 4340 13694
rect 4172 13580 4228 13636
rect 3724 12962 3780 12964
rect 3724 12910 3726 12962
rect 3726 12910 3778 12962
rect 3778 12910 3780 12962
rect 3724 12908 3780 12910
rect 4464 13354 4520 13356
rect 4464 13302 4466 13354
rect 4466 13302 4518 13354
rect 4518 13302 4520 13354
rect 4464 13300 4520 13302
rect 4568 13354 4624 13356
rect 4568 13302 4570 13354
rect 4570 13302 4622 13354
rect 4622 13302 4624 13354
rect 4568 13300 4624 13302
rect 4672 13354 4728 13356
rect 4672 13302 4674 13354
rect 4674 13302 4726 13354
rect 4726 13302 4728 13354
rect 4672 13300 4728 13302
rect 4508 12962 4564 12964
rect 4508 12910 4510 12962
rect 4510 12910 4562 12962
rect 4562 12910 4564 12962
rect 4508 12908 4564 12910
rect 4956 14028 5012 14084
rect 5404 16604 5460 16660
rect 3804 12570 3860 12572
rect 3804 12518 3806 12570
rect 3806 12518 3858 12570
rect 3858 12518 3860 12570
rect 3804 12516 3860 12518
rect 3908 12570 3964 12572
rect 3908 12518 3910 12570
rect 3910 12518 3962 12570
rect 3962 12518 3964 12570
rect 3908 12516 3964 12518
rect 4012 12570 4068 12572
rect 4012 12518 4014 12570
rect 4014 12518 4066 12570
rect 4066 12518 4068 12570
rect 4012 12516 4068 12518
rect 4284 12460 4340 12516
rect 3724 12178 3780 12180
rect 3724 12126 3726 12178
rect 3726 12126 3778 12178
rect 3778 12126 3780 12178
rect 3724 12124 3780 12126
rect 4464 11786 4520 11788
rect 4464 11734 4466 11786
rect 4466 11734 4518 11786
rect 4518 11734 4520 11786
rect 4464 11732 4520 11734
rect 4568 11786 4624 11788
rect 4568 11734 4570 11786
rect 4570 11734 4622 11786
rect 4622 11734 4624 11786
rect 4568 11732 4624 11734
rect 4672 11786 4728 11788
rect 4672 11734 4674 11786
rect 4674 11734 4726 11786
rect 4726 11734 4728 11786
rect 4672 11732 4728 11734
rect 5292 14924 5348 14980
rect 5292 14364 5348 14420
rect 5180 13244 5236 13300
rect 3612 11340 3668 11396
rect 4396 11340 4452 11396
rect 3804 11002 3860 11004
rect 3804 10950 3806 11002
rect 3806 10950 3858 11002
rect 3858 10950 3860 11002
rect 3804 10948 3860 10950
rect 3908 11002 3964 11004
rect 3908 10950 3910 11002
rect 3910 10950 3962 11002
rect 3962 10950 3964 11002
rect 3908 10948 3964 10950
rect 4012 11002 4068 11004
rect 4012 10950 4014 11002
rect 4014 10950 4066 11002
rect 4066 10950 4068 11002
rect 4012 10948 4068 10950
rect 5068 10556 5124 10612
rect 4396 10332 4452 10388
rect 4464 10218 4520 10220
rect 4464 10166 4466 10218
rect 4466 10166 4518 10218
rect 4518 10166 4520 10218
rect 4464 10164 4520 10166
rect 4568 10218 4624 10220
rect 4568 10166 4570 10218
rect 4570 10166 4622 10218
rect 4622 10166 4624 10218
rect 4568 10164 4624 10166
rect 4672 10218 4728 10220
rect 4672 10166 4674 10218
rect 4674 10166 4726 10218
rect 4726 10166 4728 10218
rect 4672 10164 4728 10166
rect 3164 9996 3220 10052
rect 4732 9938 4788 9940
rect 4732 9886 4734 9938
rect 4734 9886 4786 9938
rect 4786 9886 4788 9938
rect 4732 9884 4788 9886
rect 5292 10610 5348 10612
rect 5292 10558 5294 10610
rect 5294 10558 5346 10610
rect 5346 10558 5348 10610
rect 5292 10556 5348 10558
rect 3804 9434 3860 9436
rect 3804 9382 3806 9434
rect 3806 9382 3858 9434
rect 3858 9382 3860 9434
rect 3804 9380 3860 9382
rect 3908 9434 3964 9436
rect 3908 9382 3910 9434
rect 3910 9382 3962 9434
rect 3962 9382 3964 9434
rect 3908 9380 3964 9382
rect 4012 9434 4068 9436
rect 4012 9382 4014 9434
rect 4014 9382 4066 9434
rect 4066 9382 4068 9434
rect 4012 9380 4068 9382
rect 4464 8650 4520 8652
rect 4464 8598 4466 8650
rect 4466 8598 4518 8650
rect 4518 8598 4520 8650
rect 4464 8596 4520 8598
rect 4568 8650 4624 8652
rect 4568 8598 4570 8650
rect 4570 8598 4622 8650
rect 4622 8598 4624 8650
rect 4568 8596 4624 8598
rect 4672 8650 4728 8652
rect 4672 8598 4674 8650
rect 4674 8598 4726 8650
rect 4726 8598 4728 8650
rect 4672 8596 4728 8598
rect 6076 18226 6132 18228
rect 6076 18174 6078 18226
rect 6078 18174 6130 18226
rect 6130 18174 6132 18226
rect 6076 18172 6132 18174
rect 5628 16268 5684 16324
rect 5740 16828 5796 16884
rect 5628 13916 5684 13972
rect 6188 16716 6244 16772
rect 5852 13468 5908 13524
rect 6188 15202 6244 15204
rect 6188 15150 6190 15202
rect 6190 15150 6242 15202
rect 6242 15150 6244 15202
rect 6188 15148 6244 15150
rect 7420 35308 7476 35364
rect 7084 34412 7140 34468
rect 7196 33292 7252 33348
rect 7196 32508 7252 32564
rect 7420 33068 7476 33124
rect 7420 32508 7476 32564
rect 7084 32284 7140 32340
rect 7308 31778 7364 31780
rect 7308 31726 7310 31778
rect 7310 31726 7362 31778
rect 7362 31726 7364 31778
rect 7308 31724 7364 31726
rect 7084 30044 7140 30100
rect 6972 28754 7028 28756
rect 6972 28702 6974 28754
rect 6974 28702 7026 28754
rect 7026 28702 7028 28754
rect 6972 28700 7028 28702
rect 6972 27804 7028 27860
rect 6636 25618 6692 25620
rect 6636 25566 6638 25618
rect 6638 25566 6690 25618
rect 6690 25566 6692 25618
rect 6636 25564 6692 25566
rect 6748 25116 6804 25172
rect 6860 25004 6916 25060
rect 6860 23660 6916 23716
rect 7084 25004 7140 25060
rect 7308 30716 7364 30772
rect 7196 23212 7252 23268
rect 7756 32284 7812 32340
rect 7644 31554 7700 31556
rect 7644 31502 7646 31554
rect 7646 31502 7698 31554
rect 7698 31502 7700 31554
rect 7644 31500 7700 31502
rect 7644 30940 7700 30996
rect 7644 30770 7700 30772
rect 7644 30718 7646 30770
rect 7646 30718 7698 30770
rect 7698 30718 7700 30770
rect 7644 30716 7700 30718
rect 7308 30156 7364 30212
rect 7420 28476 7476 28532
rect 7644 26290 7700 26292
rect 7644 26238 7646 26290
rect 7646 26238 7698 26290
rect 7698 26238 7700 26290
rect 7644 26236 7700 26238
rect 7420 25116 7476 25172
rect 7532 25004 7588 25060
rect 6972 22370 7028 22372
rect 6972 22318 6974 22370
rect 6974 22318 7026 22370
rect 7026 22318 7028 22370
rect 6972 22316 7028 22318
rect 7084 21586 7140 21588
rect 7084 21534 7086 21586
rect 7086 21534 7138 21586
rect 7138 21534 7140 21586
rect 7084 21532 7140 21534
rect 6636 20914 6692 20916
rect 6636 20862 6638 20914
rect 6638 20862 6690 20914
rect 6690 20862 6692 20914
rect 6636 20860 6692 20862
rect 6748 20130 6804 20132
rect 6748 20078 6750 20130
rect 6750 20078 6802 20130
rect 6802 20078 6804 20130
rect 6748 20076 6804 20078
rect 6524 19404 6580 19460
rect 6636 19292 6692 19348
rect 6636 19122 6692 19124
rect 6636 19070 6638 19122
rect 6638 19070 6690 19122
rect 6690 19070 6692 19122
rect 6636 19068 6692 19070
rect 7308 21362 7364 21364
rect 7308 21310 7310 21362
rect 7310 21310 7362 21362
rect 7362 21310 7364 21362
rect 7308 21308 7364 21310
rect 7196 20860 7252 20916
rect 7644 23938 7700 23940
rect 7644 23886 7646 23938
rect 7646 23886 7698 23938
rect 7698 23886 7700 23938
rect 7644 23884 7700 23886
rect 7532 22988 7588 23044
rect 7644 23660 7700 23716
rect 7420 20412 7476 20468
rect 7196 19906 7252 19908
rect 7196 19854 7198 19906
rect 7198 19854 7250 19906
rect 7250 19854 7252 19906
rect 7196 19852 7252 19854
rect 6860 19068 6916 19124
rect 6972 19292 7028 19348
rect 6636 18508 6692 18564
rect 6636 17666 6692 17668
rect 6636 17614 6638 17666
rect 6638 17614 6690 17666
rect 6690 17614 6692 17666
rect 6636 17612 6692 17614
rect 6636 16882 6692 16884
rect 6636 16830 6638 16882
rect 6638 16830 6690 16882
rect 6690 16830 6692 16882
rect 6636 16828 6692 16830
rect 6972 18172 7028 18228
rect 7084 16770 7140 16772
rect 7084 16718 7086 16770
rect 7086 16718 7138 16770
rect 7138 16718 7140 16770
rect 7084 16716 7140 16718
rect 7420 19292 7476 19348
rect 7532 22316 7588 22372
rect 6860 15260 6916 15316
rect 7420 19068 7476 19124
rect 5740 10668 5796 10724
rect 5852 11676 5908 11732
rect 5964 10556 6020 10612
rect 6412 13692 6468 13748
rect 6748 13522 6804 13524
rect 6748 13470 6750 13522
rect 6750 13470 6802 13522
rect 6802 13470 6804 13522
rect 6748 13468 6804 13470
rect 6412 13132 6468 13188
rect 6636 12124 6692 12180
rect 6972 12178 7028 12180
rect 6972 12126 6974 12178
rect 6974 12126 7026 12178
rect 7026 12126 7028 12178
rect 6972 12124 7028 12126
rect 7084 12012 7140 12068
rect 7308 15708 7364 15764
rect 7308 12962 7364 12964
rect 7308 12910 7310 12962
rect 7310 12910 7362 12962
rect 7362 12910 7364 12962
rect 7308 12908 7364 12910
rect 7644 14700 7700 14756
rect 8204 39618 8260 39620
rect 8204 39566 8206 39618
rect 8206 39566 8258 39618
rect 8258 39566 8260 39618
rect 8204 39564 8260 39566
rect 8316 37436 8372 37492
rect 8204 37100 8260 37156
rect 8092 35644 8148 35700
rect 8316 35532 8372 35588
rect 8764 40402 8820 40404
rect 8764 40350 8766 40402
rect 8766 40350 8818 40402
rect 8818 40350 8820 40402
rect 8764 40348 8820 40350
rect 8204 35308 8260 35364
rect 8204 33740 8260 33796
rect 8092 33628 8148 33684
rect 8204 33516 8260 33572
rect 8428 32562 8484 32564
rect 8428 32510 8430 32562
rect 8430 32510 8482 32562
rect 8482 32510 8484 32562
rect 8428 32508 8484 32510
rect 8652 35698 8708 35700
rect 8652 35646 8654 35698
rect 8654 35646 8706 35698
rect 8706 35646 8708 35698
rect 8652 35644 8708 35646
rect 8652 35420 8708 35476
rect 8988 38668 9044 38724
rect 9996 48972 10052 49028
rect 9324 40572 9380 40628
rect 9436 40348 9492 40404
rect 9884 39842 9940 39844
rect 9884 39790 9886 39842
rect 9886 39790 9938 39842
rect 9938 39790 9940 39842
rect 9884 39788 9940 39790
rect 9436 38050 9492 38052
rect 9436 37998 9438 38050
rect 9438 37998 9490 38050
rect 9490 37998 9492 38050
rect 9436 37996 9492 37998
rect 9212 36092 9268 36148
rect 8988 35644 9044 35700
rect 9324 35698 9380 35700
rect 9324 35646 9326 35698
rect 9326 35646 9378 35698
rect 9378 35646 9380 35698
rect 9324 35644 9380 35646
rect 8876 35586 8932 35588
rect 8876 35534 8878 35586
rect 8878 35534 8930 35586
rect 8930 35534 8932 35586
rect 8876 35532 8932 35534
rect 9212 35532 9268 35588
rect 9100 35420 9156 35476
rect 9100 32956 9156 33012
rect 9772 39564 9828 39620
rect 13580 54236 13636 54292
rect 12908 53340 12964 53396
rect 13020 53900 13076 53956
rect 12796 52332 12852 52388
rect 11004 50652 11060 50708
rect 15596 55468 15652 55524
rect 19516 56252 19572 56308
rect 20636 56306 20692 56308
rect 20636 56254 20638 56306
rect 20638 56254 20690 56306
rect 20690 56254 20692 56306
rect 20636 56252 20692 56254
rect 20860 56252 20916 56308
rect 21868 56306 21924 56308
rect 21868 56254 21870 56306
rect 21870 56254 21922 56306
rect 21922 56254 21924 56306
rect 21868 56252 21924 56254
rect 22540 56140 22596 56196
rect 14028 53788 14084 53844
rect 18844 55410 18900 55412
rect 18844 55358 18846 55410
rect 18846 55358 18898 55410
rect 18898 55358 18900 55410
rect 18844 55356 18900 55358
rect 17500 53564 17556 53620
rect 17612 54124 17668 54180
rect 15148 52892 15204 52948
rect 14252 50428 14308 50484
rect 11004 42028 11060 42084
rect 11340 43596 11396 43652
rect 10892 41804 10948 41860
rect 10556 41020 10612 41076
rect 10108 40348 10164 40404
rect 9548 33628 9604 33684
rect 9996 37772 10052 37828
rect 9996 36988 10052 37044
rect 10108 36316 10164 36372
rect 9660 35644 9716 35700
rect 8764 32732 8820 32788
rect 9548 32732 9604 32788
rect 8652 31836 8708 31892
rect 8876 31778 8932 31780
rect 8876 31726 8878 31778
rect 8878 31726 8930 31778
rect 8930 31726 8932 31778
rect 8876 31724 8932 31726
rect 8316 30156 8372 30212
rect 7980 26178 8036 26180
rect 7980 26126 7982 26178
rect 7982 26126 8034 26178
rect 8034 26126 8036 26178
rect 7980 26124 8036 26126
rect 7980 24444 8036 24500
rect 7868 23884 7924 23940
rect 8204 27804 8260 27860
rect 8428 29148 8484 29204
rect 8204 24332 8260 24388
rect 8092 23436 8148 23492
rect 7868 21756 7924 21812
rect 8316 22428 8372 22484
rect 8092 22204 8148 22260
rect 8204 22316 8260 22372
rect 7980 21644 8036 21700
rect 8092 21756 8148 21812
rect 8316 21868 8372 21924
rect 8316 20018 8372 20020
rect 8316 19966 8318 20018
rect 8318 19966 8370 20018
rect 8370 19966 8372 20018
rect 8316 19964 8372 19966
rect 8540 28476 8596 28532
rect 8876 29314 8932 29316
rect 8876 29262 8878 29314
rect 8878 29262 8930 29314
rect 8930 29262 8932 29314
rect 8876 29260 8932 29262
rect 9212 32396 9268 32452
rect 9212 29484 9268 29540
rect 9436 32508 9492 32564
rect 9100 28252 9156 28308
rect 8988 28028 9044 28084
rect 8652 27356 8708 27412
rect 8428 19852 8484 19908
rect 8540 24220 8596 24276
rect 9324 28028 9380 28084
rect 9436 29260 9492 29316
rect 9324 27858 9380 27860
rect 9324 27806 9326 27858
rect 9326 27806 9378 27858
rect 9378 27806 9380 27858
rect 9324 27804 9380 27806
rect 8092 19180 8148 19236
rect 8092 18562 8148 18564
rect 8092 18510 8094 18562
rect 8094 18510 8146 18562
rect 8146 18510 8148 18562
rect 8092 18508 8148 18510
rect 7868 16828 7924 16884
rect 7980 16268 8036 16324
rect 7532 12236 7588 12292
rect 7084 10610 7140 10612
rect 7084 10558 7086 10610
rect 7086 10558 7138 10610
rect 7138 10558 7140 10610
rect 7084 10556 7140 10558
rect 6300 9884 6356 9940
rect 7084 9714 7140 9716
rect 7084 9662 7086 9714
rect 7086 9662 7138 9714
rect 7138 9662 7140 9714
rect 7084 9660 7140 9662
rect 7420 12012 7476 12068
rect 7196 9100 7252 9156
rect 7756 13244 7812 13300
rect 8316 17276 8372 17332
rect 8204 16268 8260 16324
rect 8316 16156 8372 16212
rect 8092 15986 8148 15988
rect 8092 15934 8094 15986
rect 8094 15934 8146 15986
rect 8146 15934 8148 15986
rect 8092 15932 8148 15934
rect 8204 12850 8260 12852
rect 8204 12798 8206 12850
rect 8206 12798 8258 12850
rect 8258 12798 8260 12850
rect 8204 12796 8260 12798
rect 8204 12124 8260 12180
rect 7980 9548 8036 9604
rect 7420 9324 7476 9380
rect 7308 9042 7364 9044
rect 7308 8990 7310 9042
rect 7310 8990 7362 9042
rect 7362 8990 7364 9042
rect 7308 8988 7364 8990
rect 8204 11394 8260 11396
rect 8204 11342 8206 11394
rect 8206 11342 8258 11394
rect 8258 11342 8260 11394
rect 8204 11340 8260 11342
rect 8204 10668 8260 10724
rect 8540 18396 8596 18452
rect 8540 12178 8596 12180
rect 8540 12126 8542 12178
rect 8542 12126 8594 12178
rect 8594 12126 8596 12178
rect 8540 12124 8596 12126
rect 8428 9996 8484 10052
rect 8092 8988 8148 9044
rect 8764 22988 8820 23044
rect 8988 21532 9044 21588
rect 9324 26124 9380 26180
rect 9324 24108 9380 24164
rect 9324 23436 9380 23492
rect 9212 22370 9268 22372
rect 9212 22318 9214 22370
rect 9214 22318 9266 22370
rect 9266 22318 9268 22370
rect 9212 22316 9268 22318
rect 9548 24892 9604 24948
rect 9884 35698 9940 35700
rect 9884 35646 9886 35698
rect 9886 35646 9938 35698
rect 9938 35646 9940 35698
rect 9884 35644 9940 35646
rect 9884 33458 9940 33460
rect 9884 33406 9886 33458
rect 9886 33406 9938 33458
rect 9938 33406 9940 33458
rect 9884 33404 9940 33406
rect 9772 29372 9828 29428
rect 11004 39618 11060 39620
rect 11004 39566 11006 39618
rect 11006 39566 11058 39618
rect 11058 39566 11060 39618
rect 11004 39564 11060 39566
rect 10556 37996 10612 38052
rect 10668 35980 10724 36036
rect 10556 35756 10612 35812
rect 11116 38050 11172 38052
rect 11116 37998 11118 38050
rect 11118 37998 11170 38050
rect 11170 37998 11172 38050
rect 11116 37996 11172 37998
rect 11004 35868 11060 35924
rect 10556 32562 10612 32564
rect 10556 32510 10558 32562
rect 10558 32510 10610 32562
rect 10610 32510 10612 32562
rect 10556 32508 10612 32510
rect 10220 30210 10276 30212
rect 10220 30158 10222 30210
rect 10222 30158 10274 30210
rect 10274 30158 10276 30210
rect 10220 30156 10276 30158
rect 10220 29372 10276 29428
rect 9884 24220 9940 24276
rect 9436 22316 9492 22372
rect 9436 21980 9492 22036
rect 8988 20076 9044 20132
rect 8988 18508 9044 18564
rect 9100 15484 9156 15540
rect 9660 22316 9716 22372
rect 9660 21868 9716 21924
rect 9772 21644 9828 21700
rect 10108 21586 10164 21588
rect 10108 21534 10110 21586
rect 10110 21534 10162 21586
rect 10162 21534 10164 21586
rect 10108 21532 10164 21534
rect 9772 21308 9828 21364
rect 9884 20914 9940 20916
rect 9884 20862 9886 20914
rect 9886 20862 9938 20914
rect 9938 20862 9940 20914
rect 9884 20860 9940 20862
rect 9436 20188 9492 20244
rect 9324 19906 9380 19908
rect 9324 19854 9326 19906
rect 9326 19854 9378 19906
rect 9378 19854 9380 19906
rect 9324 19852 9380 19854
rect 9548 19628 9604 19684
rect 9660 16828 9716 16884
rect 9324 16098 9380 16100
rect 9324 16046 9326 16098
rect 9326 16046 9378 16098
rect 9378 16046 9380 16098
rect 9324 16044 9380 16046
rect 9548 16380 9604 16436
rect 9548 15426 9604 15428
rect 9548 15374 9550 15426
rect 9550 15374 9602 15426
rect 9602 15374 9604 15426
rect 9548 15372 9604 15374
rect 9660 15260 9716 15316
rect 8764 13580 8820 13636
rect 8764 12012 8820 12068
rect 9436 14700 9492 14756
rect 9548 14642 9604 14644
rect 9548 14590 9550 14642
rect 9550 14590 9602 14642
rect 9602 14590 9604 14642
rect 9548 14588 9604 14590
rect 9436 14476 9492 14532
rect 9996 19404 10052 19460
rect 10108 20300 10164 20356
rect 9996 17836 10052 17892
rect 10332 25564 10388 25620
rect 10332 22482 10388 22484
rect 10332 22430 10334 22482
rect 10334 22430 10386 22482
rect 10386 22430 10388 22482
rect 10332 22428 10388 22430
rect 10556 25116 10612 25172
rect 11228 35980 11284 36036
rect 12236 42924 12292 42980
rect 12012 41692 12068 41748
rect 11788 39788 11844 39844
rect 11788 39618 11844 39620
rect 11788 39566 11790 39618
rect 11790 39566 11842 39618
rect 11842 39566 11844 39618
rect 11788 39564 11844 39566
rect 10780 30380 10836 30436
rect 11340 29596 11396 29652
rect 11340 29372 11396 29428
rect 11116 28812 11172 28868
rect 10892 28530 10948 28532
rect 10892 28478 10894 28530
rect 10894 28478 10946 28530
rect 10946 28478 10948 28530
rect 10892 28476 10948 28478
rect 11004 27858 11060 27860
rect 11004 27806 11006 27858
rect 11006 27806 11058 27858
rect 11058 27806 11060 27858
rect 11004 27804 11060 27806
rect 10892 27020 10948 27076
rect 10780 25564 10836 25620
rect 11340 28866 11396 28868
rect 11340 28814 11342 28866
rect 11342 28814 11394 28866
rect 11394 28814 11396 28866
rect 11340 28812 11396 28814
rect 11452 27804 11508 27860
rect 11788 38108 11844 38164
rect 11900 38050 11956 38052
rect 11900 37998 11902 38050
rect 11902 37998 11954 38050
rect 11954 37998 11956 38050
rect 11900 37996 11956 37998
rect 11788 37324 11844 37380
rect 12124 37996 12180 38052
rect 13020 42700 13076 42756
rect 12908 39788 12964 39844
rect 12684 38780 12740 38836
rect 12012 35084 12068 35140
rect 12348 37772 12404 37828
rect 12460 37212 12516 37268
rect 11788 32508 11844 32564
rect 12124 34690 12180 34692
rect 12124 34638 12126 34690
rect 12126 34638 12178 34690
rect 12178 34638 12180 34690
rect 12124 34636 12180 34638
rect 12572 34188 12628 34244
rect 12460 33964 12516 34020
rect 12124 32338 12180 32340
rect 12124 32286 12126 32338
rect 12126 32286 12178 32338
rect 12178 32286 12180 32338
rect 12124 32284 12180 32286
rect 11900 31388 11956 31444
rect 12012 31052 12068 31108
rect 11900 30492 11956 30548
rect 11564 27468 11620 27524
rect 11676 29596 11732 29652
rect 11228 27132 11284 27188
rect 10668 25004 10724 25060
rect 10556 23548 10612 23604
rect 10556 23042 10612 23044
rect 10556 22990 10558 23042
rect 10558 22990 10610 23042
rect 10610 22990 10612 23042
rect 10556 22988 10612 22990
rect 10444 20860 10500 20916
rect 10556 20188 10612 20244
rect 10220 19292 10276 19348
rect 10332 19234 10388 19236
rect 10332 19182 10334 19234
rect 10334 19182 10386 19234
rect 10386 19182 10388 19234
rect 10332 19180 10388 19182
rect 10892 23996 10948 24052
rect 11788 29426 11844 29428
rect 11788 29374 11790 29426
rect 11790 29374 11842 29426
rect 11842 29374 11844 29426
rect 11788 29372 11844 29374
rect 11676 27186 11732 27188
rect 11676 27134 11678 27186
rect 11678 27134 11730 27186
rect 11730 27134 11732 27186
rect 11676 27132 11732 27134
rect 11340 26962 11396 26964
rect 11340 26910 11342 26962
rect 11342 26910 11394 26962
rect 11394 26910 11396 26962
rect 11340 26908 11396 26910
rect 10780 23548 10836 23604
rect 11452 26460 11508 26516
rect 10892 22370 10948 22372
rect 10892 22318 10894 22370
rect 10894 22318 10946 22370
rect 10946 22318 10948 22370
rect 10892 22316 10948 22318
rect 11788 26012 11844 26068
rect 10780 20636 10836 20692
rect 10332 18562 10388 18564
rect 10332 18510 10334 18562
rect 10334 18510 10386 18562
rect 10386 18510 10388 18562
rect 10332 18508 10388 18510
rect 10780 18396 10836 18452
rect 10668 18338 10724 18340
rect 10668 18286 10670 18338
rect 10670 18286 10722 18338
rect 10722 18286 10724 18338
rect 10668 18284 10724 18286
rect 11116 20076 11172 20132
rect 11340 21756 11396 21812
rect 11452 21308 11508 21364
rect 11676 22876 11732 22932
rect 11676 21810 11732 21812
rect 11676 21758 11678 21810
rect 11678 21758 11730 21810
rect 11730 21758 11732 21810
rect 11676 21756 11732 21758
rect 11564 20802 11620 20804
rect 11564 20750 11566 20802
rect 11566 20750 11618 20802
rect 11618 20750 11620 20802
rect 11564 20748 11620 20750
rect 12348 32284 12404 32340
rect 12796 38332 12852 38388
rect 13132 38332 13188 38388
rect 13356 38668 13412 38724
rect 13244 38108 13300 38164
rect 13132 38050 13188 38052
rect 13132 37998 13134 38050
rect 13134 37998 13186 38050
rect 13186 37998 13188 38050
rect 13132 37996 13188 37998
rect 13468 37996 13524 38052
rect 12908 34636 12964 34692
rect 12796 31948 12852 32004
rect 12908 32956 12964 33012
rect 13244 37548 13300 37604
rect 13356 37212 13412 37268
rect 13580 37100 13636 37156
rect 13804 37884 13860 37940
rect 13356 36258 13412 36260
rect 13356 36206 13358 36258
rect 13358 36206 13410 36258
rect 13410 36206 13412 36258
rect 13356 36204 13412 36206
rect 13132 32844 13188 32900
rect 13244 35084 13300 35140
rect 13356 32956 13412 33012
rect 13356 31948 13412 32004
rect 12460 30492 12516 30548
rect 12236 29372 12292 29428
rect 12012 25282 12068 25284
rect 12012 25230 12014 25282
rect 12014 25230 12066 25282
rect 12066 25230 12068 25282
rect 12012 25228 12068 25230
rect 12124 24892 12180 24948
rect 12012 23212 12068 23268
rect 12012 23042 12068 23044
rect 12012 22990 12014 23042
rect 12014 22990 12066 23042
rect 12066 22990 12068 23042
rect 12012 22988 12068 22990
rect 11900 22652 11956 22708
rect 11900 22370 11956 22372
rect 11900 22318 11902 22370
rect 11902 22318 11954 22370
rect 11954 22318 11956 22370
rect 11900 22316 11956 22318
rect 12460 28642 12516 28644
rect 12460 28590 12462 28642
rect 12462 28590 12514 28642
rect 12514 28590 12516 28642
rect 12460 28588 12516 28590
rect 12572 26012 12628 26068
rect 12684 30604 12740 30660
rect 12572 25116 12628 25172
rect 12908 28812 12964 28868
rect 13804 32508 13860 32564
rect 14028 36204 14084 36260
rect 13916 32172 13972 32228
rect 14028 34188 14084 34244
rect 13692 31836 13748 31892
rect 13356 27692 13412 27748
rect 12796 26684 12852 26740
rect 13356 26460 13412 26516
rect 13468 26236 13524 26292
rect 13580 28812 13636 28868
rect 14476 42476 14532 42532
rect 14364 36482 14420 36484
rect 14364 36430 14366 36482
rect 14366 36430 14418 36482
rect 14418 36430 14420 36482
rect 14364 36428 14420 36430
rect 14252 32508 14308 32564
rect 14252 30994 14308 30996
rect 14252 30942 14254 30994
rect 14254 30942 14306 30994
rect 14306 30942 14308 30994
rect 14252 30940 14308 30942
rect 13804 28812 13860 28868
rect 14364 29148 14420 29204
rect 16716 52668 16772 52724
rect 16044 52108 16100 52164
rect 15820 48076 15876 48132
rect 15372 40348 15428 40404
rect 15260 38834 15316 38836
rect 15260 38782 15262 38834
rect 15262 38782 15314 38834
rect 15314 38782 15316 38834
rect 15260 38780 15316 38782
rect 14812 36482 14868 36484
rect 14812 36430 14814 36482
rect 14814 36430 14866 36482
rect 14866 36430 14868 36482
rect 14812 36428 14868 36430
rect 14588 33458 14644 33460
rect 14588 33406 14590 33458
rect 14590 33406 14642 33458
rect 14642 33406 14644 33458
rect 14588 33404 14644 33406
rect 14588 31836 14644 31892
rect 14028 28252 14084 28308
rect 14812 32172 14868 32228
rect 13692 28140 13748 28196
rect 12908 25788 12964 25844
rect 12796 25676 12852 25732
rect 13132 25730 13188 25732
rect 13132 25678 13134 25730
rect 13134 25678 13186 25730
rect 13186 25678 13188 25730
rect 13132 25676 13188 25678
rect 12684 24668 12740 24724
rect 13132 25228 13188 25284
rect 12348 23826 12404 23828
rect 12348 23774 12350 23826
rect 12350 23774 12402 23826
rect 12402 23774 12404 23826
rect 12348 23772 12404 23774
rect 12236 23212 12292 23268
rect 12236 22652 12292 22708
rect 12124 21868 12180 21924
rect 12124 21362 12180 21364
rect 12124 21310 12126 21362
rect 12126 21310 12178 21362
rect 12178 21310 12180 21362
rect 12124 21308 12180 21310
rect 12012 20748 12068 20804
rect 12460 21196 12516 21252
rect 12348 20748 12404 20804
rect 11900 20188 11956 20244
rect 12012 20076 12068 20132
rect 12124 19852 12180 19908
rect 11676 19516 11732 19572
rect 12348 19628 12404 19684
rect 11564 19458 11620 19460
rect 11564 19406 11566 19458
rect 11566 19406 11618 19458
rect 11618 19406 11620 19458
rect 11564 19404 11620 19406
rect 11676 19292 11732 19348
rect 11004 18508 11060 18564
rect 11564 17948 11620 18004
rect 10892 17500 10948 17556
rect 11228 17554 11284 17556
rect 11228 17502 11230 17554
rect 11230 17502 11282 17554
rect 11282 17502 11284 17554
rect 11228 17500 11284 17502
rect 10332 17052 10388 17108
rect 9996 16492 10052 16548
rect 10780 16604 10836 16660
rect 10108 16210 10164 16212
rect 10108 16158 10110 16210
rect 10110 16158 10162 16210
rect 10162 16158 10164 16210
rect 10108 16156 10164 16158
rect 9996 16098 10052 16100
rect 9996 16046 9998 16098
rect 9998 16046 10050 16098
rect 10050 16046 10052 16098
rect 9996 16044 10052 16046
rect 9884 15932 9940 15988
rect 10108 15202 10164 15204
rect 10108 15150 10110 15202
rect 10110 15150 10162 15202
rect 10162 15150 10164 15202
rect 10108 15148 10164 15150
rect 10220 15708 10276 15764
rect 11116 16268 11172 16324
rect 11004 15932 11060 15988
rect 10892 15708 10948 15764
rect 10108 14642 10164 14644
rect 10108 14590 10110 14642
rect 10110 14590 10162 14642
rect 10162 14590 10164 14642
rect 10108 14588 10164 14590
rect 11116 15708 11172 15764
rect 11004 15426 11060 15428
rect 11004 15374 11006 15426
rect 11006 15374 11058 15426
rect 11058 15374 11060 15426
rect 11004 15372 11060 15374
rect 10556 15314 10612 15316
rect 10556 15262 10558 15314
rect 10558 15262 10610 15314
rect 10610 15262 10612 15314
rect 10556 15260 10612 15262
rect 9996 14530 10052 14532
rect 9996 14478 9998 14530
rect 9998 14478 10050 14530
rect 10050 14478 10052 14530
rect 9996 14476 10052 14478
rect 9436 14306 9492 14308
rect 9436 14254 9438 14306
rect 9438 14254 9490 14306
rect 9490 14254 9492 14306
rect 9436 14252 9492 14254
rect 9100 12850 9156 12852
rect 9100 12798 9102 12850
rect 9102 12798 9154 12850
rect 9154 12798 9156 12850
rect 9100 12796 9156 12798
rect 9324 12178 9380 12180
rect 9324 12126 9326 12178
rect 9326 12126 9378 12178
rect 9378 12126 9380 12178
rect 9324 12124 9380 12126
rect 8988 12066 9044 12068
rect 8988 12014 8990 12066
rect 8990 12014 9042 12066
rect 9042 12014 9044 12066
rect 8988 12012 9044 12014
rect 8876 9266 8932 9268
rect 8876 9214 8878 9266
rect 8878 9214 8930 9266
rect 8930 9214 8932 9266
rect 8876 9212 8932 9214
rect 3804 7866 3860 7868
rect 3804 7814 3806 7866
rect 3806 7814 3858 7866
rect 3858 7814 3860 7866
rect 3804 7812 3860 7814
rect 3908 7866 3964 7868
rect 3908 7814 3910 7866
rect 3910 7814 3962 7866
rect 3962 7814 3964 7866
rect 3908 7812 3964 7814
rect 4012 7866 4068 7868
rect 4012 7814 4014 7866
rect 4014 7814 4066 7866
rect 4066 7814 4068 7866
rect 4012 7812 4068 7814
rect 4464 7082 4520 7084
rect 4464 7030 4466 7082
rect 4466 7030 4518 7082
rect 4518 7030 4520 7082
rect 4464 7028 4520 7030
rect 4568 7082 4624 7084
rect 4568 7030 4570 7082
rect 4570 7030 4622 7082
rect 4622 7030 4624 7082
rect 4568 7028 4624 7030
rect 4672 7082 4728 7084
rect 4672 7030 4674 7082
rect 4674 7030 4726 7082
rect 4726 7030 4728 7082
rect 4672 7028 4728 7030
rect 3804 6298 3860 6300
rect 3804 6246 3806 6298
rect 3806 6246 3858 6298
rect 3858 6246 3860 6298
rect 3804 6244 3860 6246
rect 3908 6298 3964 6300
rect 3908 6246 3910 6298
rect 3910 6246 3962 6298
rect 3962 6246 3964 6298
rect 3908 6244 3964 6246
rect 4012 6298 4068 6300
rect 4012 6246 4014 6298
rect 4014 6246 4066 6298
rect 4066 6246 4068 6298
rect 4012 6244 4068 6246
rect 4464 5514 4520 5516
rect 4464 5462 4466 5514
rect 4466 5462 4518 5514
rect 4518 5462 4520 5514
rect 4464 5460 4520 5462
rect 4568 5514 4624 5516
rect 4568 5462 4570 5514
rect 4570 5462 4622 5514
rect 4622 5462 4624 5514
rect 4568 5460 4624 5462
rect 4672 5514 4728 5516
rect 4672 5462 4674 5514
rect 4674 5462 4726 5514
rect 4726 5462 4728 5514
rect 4672 5460 4728 5462
rect 1260 5180 1316 5236
rect 3804 4730 3860 4732
rect 3804 4678 3806 4730
rect 3806 4678 3858 4730
rect 3858 4678 3860 4730
rect 3804 4676 3860 4678
rect 3908 4730 3964 4732
rect 3908 4678 3910 4730
rect 3910 4678 3962 4730
rect 3962 4678 3964 4730
rect 3908 4676 3964 4678
rect 4012 4730 4068 4732
rect 4012 4678 4014 4730
rect 4014 4678 4066 4730
rect 4066 4678 4068 4730
rect 4012 4676 4068 4678
rect 1484 4450 1540 4452
rect 1484 4398 1486 4450
rect 1486 4398 1538 4450
rect 1538 4398 1540 4450
rect 1484 4396 1540 4398
rect 4464 3946 4520 3948
rect 4464 3894 4466 3946
rect 4466 3894 4518 3946
rect 4518 3894 4520 3946
rect 4464 3892 4520 3894
rect 4568 3946 4624 3948
rect 4568 3894 4570 3946
rect 4570 3894 4622 3946
rect 4622 3894 4624 3946
rect 4568 3892 4624 3894
rect 4672 3946 4728 3948
rect 4672 3894 4674 3946
rect 4674 3894 4726 3946
rect 4726 3894 4728 3946
rect 4672 3892 4728 3894
rect 3804 3162 3860 3164
rect 3804 3110 3806 3162
rect 3806 3110 3858 3162
rect 3858 3110 3860 3162
rect 3804 3108 3860 3110
rect 3908 3162 3964 3164
rect 3908 3110 3910 3162
rect 3910 3110 3962 3162
rect 3962 3110 3964 3162
rect 3908 3108 3964 3110
rect 4012 3162 4068 3164
rect 4012 3110 4014 3162
rect 4014 3110 4066 3162
rect 4066 3110 4068 3162
rect 4012 3108 4068 3110
rect 1148 2716 1204 2772
rect 3388 2716 3444 2772
rect 2044 1372 2100 1428
rect 4464 2378 4520 2380
rect 4464 2326 4466 2378
rect 4466 2326 4518 2378
rect 4518 2326 4520 2378
rect 4464 2324 4520 2326
rect 4568 2378 4624 2380
rect 4568 2326 4570 2378
rect 4570 2326 4622 2378
rect 4622 2326 4624 2378
rect 4568 2324 4624 2326
rect 4672 2378 4728 2380
rect 4672 2326 4674 2378
rect 4674 2326 4726 2378
rect 4726 2326 4728 2378
rect 4672 2324 4728 2326
rect 3804 1594 3860 1596
rect 3804 1542 3806 1594
rect 3806 1542 3858 1594
rect 3858 1542 3860 1594
rect 3804 1540 3860 1542
rect 3908 1594 3964 1596
rect 3908 1542 3910 1594
rect 3910 1542 3962 1594
rect 3962 1542 3964 1594
rect 3908 1540 3964 1542
rect 4012 1594 4068 1596
rect 4012 1542 4014 1594
rect 4014 1542 4066 1594
rect 4066 1542 4068 1594
rect 4012 1540 4068 1542
rect 8316 8146 8372 8148
rect 8316 8094 8318 8146
rect 8318 8094 8370 8146
rect 8370 8094 8372 8146
rect 8316 8092 8372 8094
rect 7420 1596 7476 1652
rect 6860 1090 6916 1092
rect 6860 1038 6862 1090
rect 6862 1038 6914 1090
rect 6914 1038 6916 1090
rect 6860 1036 6916 1038
rect 4464 810 4520 812
rect 4464 758 4466 810
rect 4466 758 4518 810
rect 4518 758 4520 810
rect 4464 756 4520 758
rect 4568 810 4624 812
rect 4568 758 4570 810
rect 4570 758 4622 810
rect 4622 758 4624 810
rect 4568 756 4624 758
rect 4672 810 4728 812
rect 4672 758 4674 810
rect 4674 758 4726 810
rect 4726 758 4728 810
rect 4672 756 4728 758
rect 4732 140 4788 196
rect 4956 140 5012 196
rect 9436 11228 9492 11284
rect 9772 13804 9828 13860
rect 9548 11004 9604 11060
rect 10108 12908 10164 12964
rect 9772 11788 9828 11844
rect 9884 11900 9940 11956
rect 10108 11788 10164 11844
rect 9660 10556 9716 10612
rect 9548 10332 9604 10388
rect 11340 15260 11396 15316
rect 11004 14306 11060 14308
rect 11004 14254 11006 14306
rect 11006 14254 11058 14306
rect 11058 14254 11060 14306
rect 11004 14252 11060 14254
rect 10556 11564 10612 11620
rect 10780 11788 10836 11844
rect 10220 11394 10276 11396
rect 10220 11342 10222 11394
rect 10222 11342 10274 11394
rect 10274 11342 10276 11394
rect 10220 11340 10276 11342
rect 11228 11340 11284 11396
rect 12236 19234 12292 19236
rect 12236 19182 12238 19234
rect 12238 19182 12290 19234
rect 12290 19182 12292 19234
rect 12236 19180 12292 19182
rect 11900 18338 11956 18340
rect 11900 18286 11902 18338
rect 11902 18286 11954 18338
rect 11954 18286 11956 18338
rect 11900 18284 11956 18286
rect 11788 17164 11844 17220
rect 13244 24892 13300 24948
rect 13020 22092 13076 22148
rect 12684 20748 12740 20804
rect 13132 21810 13188 21812
rect 13132 21758 13134 21810
rect 13134 21758 13186 21810
rect 13186 21758 13188 21810
rect 13132 21756 13188 21758
rect 12908 21362 12964 21364
rect 12908 21310 12910 21362
rect 12910 21310 12962 21362
rect 12962 21310 12964 21362
rect 12908 21308 12964 21310
rect 13020 21196 13076 21252
rect 12572 19628 12628 19684
rect 12572 19346 12628 19348
rect 12572 19294 12574 19346
rect 12574 19294 12626 19346
rect 12626 19294 12628 19346
rect 12572 19292 12628 19294
rect 12124 16604 12180 16660
rect 11676 16156 11732 16212
rect 11900 15538 11956 15540
rect 11900 15486 11902 15538
rect 11902 15486 11954 15538
rect 11954 15486 11956 15538
rect 11900 15484 11956 15486
rect 11788 15202 11844 15204
rect 11788 15150 11790 15202
rect 11790 15150 11842 15202
rect 11842 15150 11844 15202
rect 11788 15148 11844 15150
rect 12236 16380 12292 16436
rect 12012 15148 12068 15204
rect 13356 24722 13412 24724
rect 13356 24670 13358 24722
rect 13358 24670 13410 24722
rect 13410 24670 13412 24722
rect 13356 24668 13412 24670
rect 14028 27858 14084 27860
rect 14028 27806 14030 27858
rect 14030 27806 14082 27858
rect 14082 27806 14084 27858
rect 14028 27804 14084 27806
rect 14364 28642 14420 28644
rect 14364 28590 14366 28642
rect 14366 28590 14418 28642
rect 14418 28590 14420 28642
rect 14364 28588 14420 28590
rect 14588 28476 14644 28532
rect 13244 21308 13300 21364
rect 13692 25004 13748 25060
rect 13916 24610 13972 24612
rect 13916 24558 13918 24610
rect 13918 24558 13970 24610
rect 13970 24558 13972 24610
rect 13916 24556 13972 24558
rect 14140 25676 14196 25732
rect 13804 23212 13860 23268
rect 13692 22316 13748 22372
rect 13580 22092 13636 22148
rect 13580 21868 13636 21924
rect 13916 22204 13972 22260
rect 13804 21644 13860 21700
rect 13244 20860 13300 20916
rect 13356 20802 13412 20804
rect 13356 20750 13358 20802
rect 13358 20750 13410 20802
rect 13410 20750 13412 20802
rect 13356 20748 13412 20750
rect 13020 19852 13076 19908
rect 12908 18508 12964 18564
rect 13244 19628 13300 19684
rect 13132 19292 13188 19348
rect 13356 19234 13412 19236
rect 13356 19182 13358 19234
rect 13358 19182 13410 19234
rect 13410 19182 13412 19234
rect 13356 19180 13412 19182
rect 13244 19068 13300 19124
rect 13132 16828 13188 16884
rect 12012 14588 12068 14644
rect 11900 12850 11956 12852
rect 11900 12798 11902 12850
rect 11902 12798 11954 12850
rect 11954 12798 11956 12850
rect 11900 12796 11956 12798
rect 12684 14476 12740 14532
rect 12236 12962 12292 12964
rect 12236 12910 12238 12962
rect 12238 12910 12290 12962
rect 12290 12910 12292 12962
rect 12236 12908 12292 12910
rect 11564 11788 11620 11844
rect 12124 12012 12180 12068
rect 12796 13074 12852 13076
rect 12796 13022 12798 13074
rect 12798 13022 12850 13074
rect 12850 13022 12852 13074
rect 12796 13020 12852 13022
rect 11676 11564 11732 11620
rect 10220 10556 10276 10612
rect 9884 9772 9940 9828
rect 9884 9324 9940 9380
rect 9660 8988 9716 9044
rect 10892 10556 10948 10612
rect 11228 10556 11284 10612
rect 10444 10332 10500 10388
rect 10892 9548 10948 9604
rect 10444 9212 10500 9268
rect 10668 7644 10724 7700
rect 12012 11394 12068 11396
rect 12012 11342 12014 11394
rect 12014 11342 12066 11394
rect 12066 11342 12068 11394
rect 12012 11340 12068 11342
rect 12012 9884 12068 9940
rect 12348 9884 12404 9940
rect 8988 1596 9044 1652
rect 10108 5180 10164 5236
rect 11564 7586 11620 7588
rect 11564 7534 11566 7586
rect 11566 7534 11618 7586
rect 11618 7534 11620 7586
rect 11564 7532 11620 7534
rect 13020 14588 13076 14644
rect 13356 18844 13412 18900
rect 13804 20300 13860 20356
rect 13804 19628 13860 19684
rect 13692 18620 13748 18676
rect 14028 19906 14084 19908
rect 14028 19854 14030 19906
rect 14030 19854 14082 19906
rect 14082 19854 14084 19906
rect 14028 19852 14084 19854
rect 13916 19516 13972 19572
rect 14028 19628 14084 19684
rect 13916 19346 13972 19348
rect 13916 19294 13918 19346
rect 13918 19294 13970 19346
rect 13970 19294 13972 19346
rect 13916 19292 13972 19294
rect 13804 18508 13860 18564
rect 13356 16828 13412 16884
rect 13580 16940 13636 16996
rect 13356 15596 13412 15652
rect 13692 16604 13748 16660
rect 14028 18284 14084 18340
rect 14028 17052 14084 17108
rect 13916 16604 13972 16660
rect 13916 16098 13972 16100
rect 13916 16046 13918 16098
rect 13918 16046 13970 16098
rect 13970 16046 13972 16098
rect 13916 16044 13972 16046
rect 13916 15484 13972 15540
rect 13244 14476 13300 14532
rect 13580 15036 13636 15092
rect 14364 28140 14420 28196
rect 14476 27916 14532 27972
rect 14588 27634 14644 27636
rect 14588 27582 14590 27634
rect 14590 27582 14642 27634
rect 14642 27582 14644 27634
rect 14588 27580 14644 27582
rect 14700 27132 14756 27188
rect 14252 23772 14308 23828
rect 14364 22988 14420 23044
rect 14476 22204 14532 22260
rect 14700 24556 14756 24612
rect 15596 37436 15652 37492
rect 15148 34412 15204 34468
rect 15148 33458 15204 33460
rect 15148 33406 15150 33458
rect 15150 33406 15202 33458
rect 15202 33406 15204 33458
rect 15148 33404 15204 33406
rect 14924 31724 14980 31780
rect 15036 31836 15092 31892
rect 15036 31500 15092 31556
rect 15036 30940 15092 30996
rect 15148 31500 15204 31556
rect 15148 29372 15204 29428
rect 15708 34188 15764 34244
rect 15596 33292 15652 33348
rect 15372 31836 15428 31892
rect 14924 28476 14980 28532
rect 14924 27692 14980 27748
rect 15148 27804 15204 27860
rect 15932 35084 15988 35140
rect 16044 33404 16100 33460
rect 16156 46732 16212 46788
rect 15820 31218 15876 31220
rect 15820 31166 15822 31218
rect 15822 31166 15874 31218
rect 15874 31166 15876 31218
rect 15820 31164 15876 31166
rect 17276 47964 17332 48020
rect 16156 31388 16212 31444
rect 15596 27580 15652 27636
rect 15820 29426 15876 29428
rect 15820 29374 15822 29426
rect 15822 29374 15874 29426
rect 15874 29374 15876 29426
rect 15820 29372 15876 29374
rect 16156 28700 16212 28756
rect 15820 27692 15876 27748
rect 14924 24892 14980 24948
rect 14700 23660 14756 23716
rect 14812 23154 14868 23156
rect 14812 23102 14814 23154
rect 14814 23102 14866 23154
rect 14866 23102 14868 23154
rect 14812 23100 14868 23102
rect 15148 22876 15204 22932
rect 14924 22428 14980 22484
rect 15932 23324 15988 23380
rect 14924 21868 14980 21924
rect 14700 21308 14756 21364
rect 14364 20076 14420 20132
rect 14252 19740 14308 19796
rect 14476 19852 14532 19908
rect 14812 21084 14868 21140
rect 14588 19628 14644 19684
rect 14812 19292 14868 19348
rect 15036 19852 15092 19908
rect 15036 19234 15092 19236
rect 15036 19182 15038 19234
rect 15038 19182 15090 19234
rect 15090 19182 15092 19234
rect 15036 19180 15092 19182
rect 14588 18450 14644 18452
rect 14588 18398 14590 18450
rect 14590 18398 14642 18450
rect 14642 18398 14644 18450
rect 14588 18396 14644 18398
rect 14364 18060 14420 18116
rect 14588 18060 14644 18116
rect 14588 17836 14644 17892
rect 14476 17164 14532 17220
rect 14588 16716 14644 16772
rect 14364 16380 14420 16436
rect 13580 13468 13636 13524
rect 14140 13468 14196 13524
rect 13580 12684 13636 12740
rect 13132 10556 13188 10612
rect 13468 11564 13524 11620
rect 13580 10610 13636 10612
rect 13580 10558 13582 10610
rect 13582 10558 13634 10610
rect 13634 10558 13636 10610
rect 13580 10556 13636 10558
rect 13468 10444 13524 10500
rect 13244 9826 13300 9828
rect 13244 9774 13246 9826
rect 13246 9774 13298 9826
rect 13298 9774 13300 9826
rect 13244 9772 13300 9774
rect 14252 12066 14308 12068
rect 14252 12014 14254 12066
rect 14254 12014 14306 12066
rect 14306 12014 14308 12066
rect 14252 12012 14308 12014
rect 15820 22370 15876 22372
rect 15820 22318 15822 22370
rect 15822 22318 15874 22370
rect 15874 22318 15876 22370
rect 15820 22316 15876 22318
rect 15260 21474 15316 21476
rect 15260 21422 15262 21474
rect 15262 21422 15314 21474
rect 15314 21422 15316 21474
rect 15260 21420 15316 21422
rect 15708 21362 15764 21364
rect 15708 21310 15710 21362
rect 15710 21310 15762 21362
rect 15762 21310 15764 21362
rect 15708 21308 15764 21310
rect 15820 20748 15876 20804
rect 16268 26572 16324 26628
rect 16380 27916 16436 27972
rect 16380 27020 16436 27076
rect 16716 38780 16772 38836
rect 17276 37436 17332 37492
rect 17164 36428 17220 36484
rect 17052 36370 17108 36372
rect 17052 36318 17054 36370
rect 17054 36318 17106 36370
rect 17106 36318 17108 36370
rect 17052 36316 17108 36318
rect 17052 35756 17108 35812
rect 16940 35532 16996 35588
rect 16828 35138 16884 35140
rect 16828 35086 16830 35138
rect 16830 35086 16882 35138
rect 16882 35086 16884 35138
rect 16828 35084 16884 35086
rect 16604 34076 16660 34132
rect 16940 33628 16996 33684
rect 16828 31836 16884 31892
rect 16716 31778 16772 31780
rect 16716 31726 16718 31778
rect 16718 31726 16770 31778
rect 16770 31726 16772 31778
rect 16716 31724 16772 31726
rect 16828 31612 16884 31668
rect 17500 38050 17556 38052
rect 17500 37998 17502 38050
rect 17502 37998 17554 38050
rect 17554 37998 17556 38050
rect 17500 37996 17556 37998
rect 17388 33740 17444 33796
rect 18956 54290 19012 54292
rect 18956 54238 18958 54290
rect 18958 54238 19010 54290
rect 19010 54238 19012 54290
rect 18956 54236 19012 54238
rect 18284 53116 18340 53172
rect 17836 51212 17892 51268
rect 17724 40402 17780 40404
rect 17724 40350 17726 40402
rect 17726 40350 17778 40402
rect 17778 40350 17780 40402
rect 17724 40348 17780 40350
rect 19516 54626 19572 54628
rect 19516 54574 19518 54626
rect 19518 54574 19570 54626
rect 19570 54574 19572 54626
rect 19516 54572 19572 54574
rect 20188 55356 20244 55412
rect 21084 55916 21140 55972
rect 19628 53228 19684 53284
rect 19628 53004 19684 53060
rect 17836 38556 17892 38612
rect 17948 42812 18004 42868
rect 17612 33628 17668 33684
rect 17388 32956 17444 33012
rect 17276 32508 17332 32564
rect 17612 32060 17668 32116
rect 17164 31612 17220 31668
rect 17052 31164 17108 31220
rect 16716 29932 16772 29988
rect 16828 29372 16884 29428
rect 16828 29036 16884 29092
rect 16492 26908 16548 26964
rect 16044 23100 16100 23156
rect 16380 22930 16436 22932
rect 16380 22878 16382 22930
rect 16382 22878 16434 22930
rect 16434 22878 16436 22930
rect 16380 22876 16436 22878
rect 16156 21644 16212 21700
rect 16380 21586 16436 21588
rect 16380 21534 16382 21586
rect 16382 21534 16434 21586
rect 16434 21534 16436 21586
rect 16380 21532 16436 21534
rect 16044 20242 16100 20244
rect 16044 20190 16046 20242
rect 16046 20190 16098 20242
rect 16098 20190 16100 20242
rect 16044 20188 16100 20190
rect 15596 19794 15652 19796
rect 15596 19742 15598 19794
rect 15598 19742 15650 19794
rect 15650 19742 15652 19794
rect 15596 19740 15652 19742
rect 15484 19404 15540 19460
rect 15372 18508 15428 18564
rect 14924 18396 14980 18452
rect 14812 18284 14868 18340
rect 15148 18226 15204 18228
rect 15148 18174 15150 18226
rect 15150 18174 15202 18226
rect 15202 18174 15204 18226
rect 15148 18172 15204 18174
rect 14812 17164 14868 17220
rect 15036 16828 15092 16884
rect 15260 17500 15316 17556
rect 15372 18284 15428 18340
rect 15260 16882 15316 16884
rect 15260 16830 15262 16882
rect 15262 16830 15314 16882
rect 15314 16830 15316 16882
rect 15260 16828 15316 16830
rect 15260 16044 15316 16100
rect 16044 19628 16100 19684
rect 15820 18674 15876 18676
rect 15820 18622 15822 18674
rect 15822 18622 15874 18674
rect 15874 18622 15876 18674
rect 15820 18620 15876 18622
rect 16604 24722 16660 24724
rect 16604 24670 16606 24722
rect 16606 24670 16658 24722
rect 16658 24670 16660 24722
rect 16604 24668 16660 24670
rect 16940 26796 16996 26852
rect 16940 26572 16996 26628
rect 17164 26460 17220 26516
rect 17276 30716 17332 30772
rect 16940 25228 16996 25284
rect 16828 23714 16884 23716
rect 16828 23662 16830 23714
rect 16830 23662 16882 23714
rect 16882 23662 16884 23714
rect 16828 23660 16884 23662
rect 16828 22092 16884 22148
rect 16716 21698 16772 21700
rect 16716 21646 16718 21698
rect 16718 21646 16770 21698
rect 16770 21646 16772 21698
rect 16716 21644 16772 21646
rect 17164 21474 17220 21476
rect 17164 21422 17166 21474
rect 17166 21422 17218 21474
rect 17218 21422 17220 21474
rect 17164 21420 17220 21422
rect 16940 21308 16996 21364
rect 16716 20802 16772 20804
rect 16716 20750 16718 20802
rect 16718 20750 16770 20802
rect 16770 20750 16772 20802
rect 16716 20748 16772 20750
rect 17052 20914 17108 20916
rect 17052 20862 17054 20914
rect 17054 20862 17106 20914
rect 17106 20862 17108 20914
rect 17052 20860 17108 20862
rect 17052 20636 17108 20692
rect 16940 20412 16996 20468
rect 16716 20188 16772 20244
rect 16604 19404 16660 19460
rect 16716 19516 16772 19572
rect 16604 19180 16660 19236
rect 15708 18396 15764 18452
rect 15932 18396 15988 18452
rect 15820 18284 15876 18340
rect 16492 18508 16548 18564
rect 16044 18284 16100 18340
rect 16044 17500 16100 17556
rect 15708 17276 15764 17332
rect 15820 17164 15876 17220
rect 15484 16044 15540 16100
rect 15596 16828 15652 16884
rect 15372 15986 15428 15988
rect 15372 15934 15374 15986
rect 15374 15934 15426 15986
rect 15426 15934 15428 15986
rect 15372 15932 15428 15934
rect 15260 15596 15316 15652
rect 14924 15202 14980 15204
rect 14924 15150 14926 15202
rect 14926 15150 14978 15202
rect 14978 15150 14980 15202
rect 14924 15148 14980 15150
rect 15372 15372 15428 15428
rect 15708 16716 15764 16772
rect 15148 15036 15204 15092
rect 14812 14588 14868 14644
rect 14924 14700 14980 14756
rect 14924 13916 14980 13972
rect 14588 12572 14644 12628
rect 14476 11564 14532 11620
rect 14924 12684 14980 12740
rect 14812 12572 14868 12628
rect 14028 10780 14084 10836
rect 13804 10556 13860 10612
rect 12796 7420 12852 7476
rect 12796 5068 12852 5124
rect 13580 7980 13636 8036
rect 16380 16940 16436 16996
rect 16492 17052 16548 17108
rect 16828 18620 16884 18676
rect 17052 18562 17108 18564
rect 17052 18510 17054 18562
rect 17054 18510 17106 18562
rect 17106 18510 17108 18562
rect 17052 18508 17108 18510
rect 17164 18226 17220 18228
rect 17164 18174 17166 18226
rect 17166 18174 17218 18226
rect 17218 18174 17220 18226
rect 17164 18172 17220 18174
rect 16940 17836 16996 17892
rect 16828 17500 16884 17556
rect 16604 16828 16660 16884
rect 16940 16882 16996 16884
rect 16940 16830 16942 16882
rect 16942 16830 16994 16882
rect 16994 16830 16996 16882
rect 16940 16828 16996 16830
rect 16044 15874 16100 15876
rect 16044 15822 16046 15874
rect 16046 15822 16098 15874
rect 16098 15822 16100 15874
rect 16044 15820 16100 15822
rect 15932 15596 15988 15652
rect 16044 15202 16100 15204
rect 16044 15150 16046 15202
rect 16046 15150 16098 15202
rect 16098 15150 16100 15202
rect 16044 15148 16100 15150
rect 15820 14700 15876 14756
rect 16044 14642 16100 14644
rect 16044 14590 16046 14642
rect 16046 14590 16098 14642
rect 16098 14590 16100 14642
rect 16044 14588 16100 14590
rect 15708 14476 15764 14532
rect 15932 14364 15988 14420
rect 16380 15372 16436 15428
rect 16940 15202 16996 15204
rect 16940 15150 16942 15202
rect 16942 15150 16994 15202
rect 16994 15150 16996 15202
rect 16940 15148 16996 15150
rect 16492 14364 16548 14420
rect 16380 14252 16436 14308
rect 15260 13634 15316 13636
rect 15260 13582 15262 13634
rect 15262 13582 15314 13634
rect 15314 13582 15316 13634
rect 15260 13580 15316 13582
rect 15260 13356 15316 13412
rect 16044 13746 16100 13748
rect 16044 13694 16046 13746
rect 16046 13694 16098 13746
rect 16098 13694 16100 13746
rect 16044 13692 16100 13694
rect 15820 13580 15876 13636
rect 15036 12178 15092 12180
rect 15036 12126 15038 12178
rect 15038 12126 15090 12178
rect 15090 12126 15092 12178
rect 15036 12124 15092 12126
rect 15148 9772 15204 9828
rect 15148 9212 15204 9268
rect 14588 5964 14644 6020
rect 15148 8988 15204 9044
rect 15484 12962 15540 12964
rect 15484 12910 15486 12962
rect 15486 12910 15538 12962
rect 15538 12910 15540 12962
rect 15484 12908 15540 12910
rect 15372 8988 15428 9044
rect 17164 14530 17220 14532
rect 17164 14478 17166 14530
rect 17166 14478 17218 14530
rect 17218 14478 17220 14530
rect 17164 14476 17220 14478
rect 17052 14364 17108 14420
rect 16940 14306 16996 14308
rect 16940 14254 16942 14306
rect 16942 14254 16994 14306
rect 16994 14254 16996 14306
rect 16940 14252 16996 14254
rect 18844 39788 18900 39844
rect 17948 35138 18004 35140
rect 17948 35086 17950 35138
rect 17950 35086 18002 35138
rect 18002 35086 18004 35138
rect 17948 35084 18004 35086
rect 18172 38220 18228 38276
rect 17948 30716 18004 30772
rect 17612 29596 17668 29652
rect 18284 36316 18340 36372
rect 18284 32786 18340 32788
rect 18284 32734 18286 32786
rect 18286 32734 18338 32786
rect 18338 32734 18340 32786
rect 18284 32732 18340 32734
rect 18508 34130 18564 34132
rect 18508 34078 18510 34130
rect 18510 34078 18562 34130
rect 18562 34078 18564 34130
rect 18508 34076 18564 34078
rect 18956 32732 19012 32788
rect 18172 32060 18228 32116
rect 18620 32562 18676 32564
rect 18620 32510 18622 32562
rect 18622 32510 18674 32562
rect 18674 32510 18676 32562
rect 18620 32508 18676 32510
rect 18172 31890 18228 31892
rect 18172 31838 18174 31890
rect 18174 31838 18226 31890
rect 18226 31838 18228 31890
rect 18172 31836 18228 31838
rect 17500 27970 17556 27972
rect 17500 27918 17502 27970
rect 17502 27918 17554 27970
rect 17554 27918 17556 27970
rect 17500 27916 17556 27918
rect 17724 29148 17780 29204
rect 17388 27020 17444 27076
rect 17500 27580 17556 27636
rect 17388 26796 17444 26852
rect 17388 23548 17444 23604
rect 17388 22316 17444 22372
rect 17388 20748 17444 20804
rect 17388 18338 17444 18340
rect 17388 18286 17390 18338
rect 17390 18286 17442 18338
rect 17442 18286 17444 18338
rect 17388 18284 17444 18286
rect 17612 26908 17668 26964
rect 17836 27916 17892 27972
rect 19292 40460 19348 40516
rect 19180 32450 19236 32452
rect 19180 32398 19182 32450
rect 19182 32398 19234 32450
rect 19234 32398 19236 32450
rect 19180 32396 19236 32398
rect 18396 27580 18452 27636
rect 18508 29596 18564 29652
rect 18060 27020 18116 27076
rect 17724 24610 17780 24612
rect 17724 24558 17726 24610
rect 17726 24558 17778 24610
rect 17778 24558 17780 24610
rect 17724 24556 17780 24558
rect 17612 21532 17668 21588
rect 17724 21196 17780 21252
rect 17724 20860 17780 20916
rect 17948 25228 18004 25284
rect 18396 27020 18452 27076
rect 18284 26796 18340 26852
rect 18284 26460 18340 26516
rect 18508 26236 18564 26292
rect 18620 28924 18676 28980
rect 18956 28812 19012 28868
rect 19180 31724 19236 31780
rect 19180 26460 19236 26516
rect 19180 26290 19236 26292
rect 19180 26238 19182 26290
rect 19182 26238 19234 26290
rect 19234 26238 19236 26290
rect 19180 26236 19236 26238
rect 18060 25116 18116 25172
rect 18060 24556 18116 24612
rect 18172 23884 18228 23940
rect 18508 24332 18564 24388
rect 18396 23938 18452 23940
rect 18396 23886 18398 23938
rect 18398 23886 18450 23938
rect 18450 23886 18452 23938
rect 18396 23884 18452 23886
rect 18508 23772 18564 23828
rect 18508 23548 18564 23604
rect 17948 20860 18004 20916
rect 17836 20076 17892 20132
rect 17836 18844 17892 18900
rect 17948 18284 18004 18340
rect 17836 18172 17892 18228
rect 17500 17612 17556 17668
rect 17724 15932 17780 15988
rect 17612 15820 17668 15876
rect 17052 13916 17108 13972
rect 16828 13746 16884 13748
rect 16828 13694 16830 13746
rect 16830 13694 16882 13746
rect 16882 13694 16884 13746
rect 16828 13692 16884 13694
rect 16156 12962 16212 12964
rect 16156 12910 16158 12962
rect 16158 12910 16210 12962
rect 16210 12910 16212 12962
rect 16156 12908 16212 12910
rect 15148 5740 15204 5796
rect 14700 4396 14756 4452
rect 13356 3388 13412 3444
rect 15820 6524 15876 6580
rect 15484 1148 15540 1204
rect 16828 4172 16884 4228
rect 14140 924 14196 980
rect 15484 588 15540 644
rect 17500 14418 17556 14420
rect 17500 14366 17502 14418
rect 17502 14366 17554 14418
rect 17554 14366 17556 14418
rect 17500 14364 17556 14366
rect 18396 21308 18452 21364
rect 18732 24668 18788 24724
rect 18284 21196 18340 21252
rect 18172 20130 18228 20132
rect 18172 20078 18174 20130
rect 18174 20078 18226 20130
rect 18226 20078 18228 20130
rect 18172 20076 18228 20078
rect 18732 23884 18788 23940
rect 18396 20636 18452 20692
rect 18620 18172 18676 18228
rect 18396 15986 18452 15988
rect 18396 15934 18398 15986
rect 18398 15934 18450 15986
rect 18450 15934 18452 15986
rect 18396 15932 18452 15934
rect 18620 15932 18676 15988
rect 18620 15484 18676 15540
rect 18396 13916 18452 13972
rect 19180 25506 19236 25508
rect 19180 25454 19182 25506
rect 19182 25454 19234 25506
rect 19234 25454 19236 25506
rect 19180 25452 19236 25454
rect 18956 24722 19012 24724
rect 18956 24670 18958 24722
rect 18958 24670 19010 24722
rect 19010 24670 19012 24722
rect 18956 24668 19012 24670
rect 18956 23884 19012 23940
rect 18956 20636 19012 20692
rect 18956 18226 19012 18228
rect 18956 18174 18958 18226
rect 18958 18174 19010 18226
rect 19010 18174 19012 18226
rect 18956 18172 19012 18174
rect 19964 52556 20020 52612
rect 20524 55298 20580 55300
rect 20524 55246 20526 55298
rect 20526 55246 20578 55298
rect 20578 55246 20580 55298
rect 20524 55244 20580 55246
rect 20748 55244 20804 55300
rect 20636 54012 20692 54068
rect 20524 53730 20580 53732
rect 20524 53678 20526 53730
rect 20526 53678 20578 53730
rect 20578 53678 20580 53730
rect 20524 53676 20580 53678
rect 19852 46844 19908 46900
rect 19852 45388 19908 45444
rect 19740 37938 19796 37940
rect 19740 37886 19742 37938
rect 19742 37886 19794 37938
rect 19794 37886 19796 37938
rect 19740 37884 19796 37886
rect 19852 35138 19908 35140
rect 19852 35086 19854 35138
rect 19854 35086 19906 35138
rect 19906 35086 19908 35138
rect 19852 35084 19908 35086
rect 19516 33122 19572 33124
rect 19516 33070 19518 33122
rect 19518 33070 19570 33122
rect 19570 33070 19572 33122
rect 19516 33068 19572 33070
rect 19404 32562 19460 32564
rect 19404 32510 19406 32562
rect 19406 32510 19458 32562
rect 19458 32510 19460 32562
rect 19404 32508 19460 32510
rect 19404 25452 19460 25508
rect 19516 26012 19572 26068
rect 19292 21474 19348 21476
rect 19292 21422 19294 21474
rect 19294 21422 19346 21474
rect 19346 21422 19348 21474
rect 19292 21420 19348 21422
rect 19516 23548 19572 23604
rect 19180 20860 19236 20916
rect 19180 20690 19236 20692
rect 19180 20638 19182 20690
rect 19182 20638 19234 20690
rect 19234 20638 19236 20690
rect 19180 20636 19236 20638
rect 19068 15932 19124 15988
rect 17164 1036 17220 1092
rect 19404 20860 19460 20916
rect 19516 18450 19572 18452
rect 19516 18398 19518 18450
rect 19518 18398 19570 18450
rect 19570 18398 19572 18450
rect 19516 18396 19572 18398
rect 19292 7532 19348 7588
rect 18620 1036 18676 1092
rect 19740 30044 19796 30100
rect 19852 32396 19908 32452
rect 19852 28924 19908 28980
rect 20300 48636 20356 48692
rect 20076 45388 20132 45444
rect 20076 28028 20132 28084
rect 19740 26178 19796 26180
rect 19740 26126 19742 26178
rect 19742 26126 19794 26178
rect 19794 26126 19796 26178
rect 19740 26124 19796 26126
rect 19740 25676 19796 25732
rect 20188 25788 20244 25844
rect 19740 20860 19796 20916
rect 20076 23772 20132 23828
rect 20076 15932 20132 15988
rect 19964 5180 20020 5236
rect 19628 5068 19684 5124
rect 20860 48636 20916 48692
rect 21980 55916 22036 55972
rect 21644 55804 21700 55860
rect 21532 53900 21588 53956
rect 21532 53676 21588 53732
rect 21308 53618 21364 53620
rect 21308 53566 21310 53618
rect 21310 53566 21362 53618
rect 21362 53566 21364 53618
rect 21308 53564 21364 53566
rect 20972 35420 21028 35476
rect 21084 53452 21140 53508
rect 20412 28812 20468 28868
rect 20412 25676 20468 25732
rect 20972 25676 21028 25732
rect 20636 23324 20692 23380
rect 20748 21980 20804 22036
rect 20412 20914 20468 20916
rect 20412 20862 20414 20914
rect 20414 20862 20466 20914
rect 20466 20862 20468 20914
rect 20412 20860 20468 20862
rect 21308 52834 21364 52836
rect 21308 52782 21310 52834
rect 21310 52782 21362 52834
rect 21362 52782 21364 52834
rect 21308 52780 21364 52782
rect 21084 18396 21140 18452
rect 21196 23324 21252 23380
rect 20972 9996 21028 10052
rect 20748 4844 20804 4900
rect 20300 588 20356 644
rect 20860 3276 20916 3332
rect 21308 18284 21364 18340
rect 21308 17052 21364 17108
rect 21756 53116 21812 53172
rect 21868 53004 21924 53060
rect 24220 57148 24276 57204
rect 23804 56474 23860 56476
rect 23804 56422 23806 56474
rect 23806 56422 23858 56474
rect 23858 56422 23860 56474
rect 23804 56420 23860 56422
rect 23908 56474 23964 56476
rect 23908 56422 23910 56474
rect 23910 56422 23962 56474
rect 23962 56422 23964 56474
rect 23908 56420 23964 56422
rect 24012 56474 24068 56476
rect 24012 56422 24014 56474
rect 24014 56422 24066 56474
rect 24066 56422 24068 56474
rect 24012 56420 24068 56422
rect 23548 56252 23604 56308
rect 23548 56028 23604 56084
rect 23212 55468 23268 55524
rect 22204 53788 22260 53844
rect 22652 53228 22708 53284
rect 22204 52722 22260 52724
rect 22204 52670 22206 52722
rect 22206 52670 22258 52722
rect 22258 52670 22260 52722
rect 22204 52668 22260 52670
rect 22764 52556 22820 52612
rect 21868 37996 21924 38052
rect 21868 29820 21924 29876
rect 22204 33740 22260 33796
rect 21532 5068 21588 5124
rect 21196 2828 21252 2884
rect 22876 51324 22932 51380
rect 22428 1596 22484 1652
rect 23100 54402 23156 54404
rect 23100 54350 23102 54402
rect 23102 54350 23154 54402
rect 23154 54350 23156 54402
rect 23100 54348 23156 54350
rect 22988 49868 23044 49924
rect 23884 55970 23940 55972
rect 23884 55918 23886 55970
rect 23886 55918 23938 55970
rect 23938 55918 23940 55970
rect 23884 55916 23940 55918
rect 23548 51996 23604 52052
rect 23804 54906 23860 54908
rect 23804 54854 23806 54906
rect 23806 54854 23858 54906
rect 23858 54854 23860 54906
rect 23804 54852 23860 54854
rect 23908 54906 23964 54908
rect 23908 54854 23910 54906
rect 23910 54854 23962 54906
rect 23962 54854 23964 54906
rect 23908 54852 23964 54854
rect 24012 54906 24068 54908
rect 24012 54854 24014 54906
rect 24014 54854 24066 54906
rect 24066 54854 24068 54906
rect 24012 54852 24068 54854
rect 24108 54738 24164 54740
rect 24108 54686 24110 54738
rect 24110 54686 24162 54738
rect 24162 54686 24164 54738
rect 24108 54684 24164 54686
rect 23772 54460 23828 54516
rect 23804 53338 23860 53340
rect 23804 53286 23806 53338
rect 23806 53286 23858 53338
rect 23858 53286 23860 53338
rect 23804 53284 23860 53286
rect 23908 53338 23964 53340
rect 23908 53286 23910 53338
rect 23910 53286 23962 53338
rect 23962 53286 23964 53338
rect 23908 53284 23964 53286
rect 24012 53338 24068 53340
rect 24012 53286 24014 53338
rect 24014 53286 24066 53338
rect 24066 53286 24068 53338
rect 24012 53284 24068 53286
rect 24444 56306 24500 56308
rect 24444 56254 24446 56306
rect 24446 56254 24498 56306
rect 24498 56254 24500 56306
rect 24444 56252 24500 56254
rect 25452 57260 25508 57316
rect 24892 56252 24948 56308
rect 25340 56700 25396 56756
rect 24464 55690 24520 55692
rect 24464 55638 24466 55690
rect 24466 55638 24518 55690
rect 24518 55638 24520 55690
rect 24464 55636 24520 55638
rect 24568 55690 24624 55692
rect 24568 55638 24570 55690
rect 24570 55638 24622 55690
rect 24622 55638 24624 55690
rect 24568 55636 24624 55638
rect 24672 55690 24728 55692
rect 24672 55638 24674 55690
rect 24674 55638 24726 55690
rect 24726 55638 24728 55690
rect 24672 55636 24728 55638
rect 25004 55356 25060 55412
rect 24220 52892 24276 52948
rect 24464 54122 24520 54124
rect 24464 54070 24466 54122
rect 24466 54070 24518 54122
rect 24518 54070 24520 54122
rect 24464 54068 24520 54070
rect 24568 54122 24624 54124
rect 24568 54070 24570 54122
rect 24570 54070 24622 54122
rect 24622 54070 24624 54122
rect 24568 54068 24624 54070
rect 24672 54122 24728 54124
rect 24672 54070 24674 54122
rect 24674 54070 24726 54122
rect 24726 54070 24728 54122
rect 24672 54068 24728 54070
rect 24668 53452 24724 53508
rect 24668 52834 24724 52836
rect 24668 52782 24670 52834
rect 24670 52782 24722 52834
rect 24722 52782 24724 52834
rect 24668 52780 24724 52782
rect 24464 52554 24520 52556
rect 24464 52502 24466 52554
rect 24466 52502 24518 52554
rect 24518 52502 24520 52554
rect 24464 52500 24520 52502
rect 24568 52554 24624 52556
rect 24568 52502 24570 52554
rect 24570 52502 24622 52554
rect 24622 52502 24624 52554
rect 24568 52500 24624 52502
rect 24672 52554 24728 52556
rect 24672 52502 24674 52554
rect 24674 52502 24726 52554
rect 24726 52502 24728 52554
rect 24672 52500 24728 52502
rect 24668 52274 24724 52276
rect 24668 52222 24670 52274
rect 24670 52222 24722 52274
rect 24722 52222 24724 52274
rect 24668 52220 24724 52222
rect 24332 51996 24388 52052
rect 23804 51770 23860 51772
rect 23804 51718 23806 51770
rect 23806 51718 23858 51770
rect 23858 51718 23860 51770
rect 23804 51716 23860 51718
rect 23908 51770 23964 51772
rect 23908 51718 23910 51770
rect 23910 51718 23962 51770
rect 23962 51718 23964 51770
rect 23908 51716 23964 51718
rect 24012 51770 24068 51772
rect 24012 51718 24014 51770
rect 24014 51718 24066 51770
rect 24066 51718 24068 51770
rect 24012 51716 24068 51718
rect 23772 51154 23828 51156
rect 23772 51102 23774 51154
rect 23774 51102 23826 51154
rect 23826 51102 23828 51154
rect 23772 51100 23828 51102
rect 23100 12348 23156 12404
rect 23804 50202 23860 50204
rect 23804 50150 23806 50202
rect 23806 50150 23858 50202
rect 23858 50150 23860 50202
rect 23804 50148 23860 50150
rect 23908 50202 23964 50204
rect 23908 50150 23910 50202
rect 23910 50150 23962 50202
rect 23962 50150 23964 50202
rect 23908 50148 23964 50150
rect 24012 50202 24068 50204
rect 24012 50150 24014 50202
rect 24014 50150 24066 50202
rect 24066 50150 24068 50202
rect 24012 50148 24068 50150
rect 25004 54460 25060 54516
rect 26236 57260 26292 57316
rect 26012 56306 26068 56308
rect 26012 56254 26014 56306
rect 26014 56254 26066 56306
rect 26066 56254 26068 56306
rect 26012 56252 26068 56254
rect 25564 54460 25620 54516
rect 25564 53618 25620 53620
rect 25564 53566 25566 53618
rect 25566 53566 25618 53618
rect 25618 53566 25620 53618
rect 25564 53564 25620 53566
rect 25452 52668 25508 52724
rect 25564 51772 25620 51828
rect 24464 50986 24520 50988
rect 24464 50934 24466 50986
rect 24466 50934 24518 50986
rect 24518 50934 24520 50986
rect 24464 50932 24520 50934
rect 24568 50986 24624 50988
rect 24568 50934 24570 50986
rect 24570 50934 24622 50986
rect 24622 50934 24624 50986
rect 24568 50932 24624 50934
rect 24672 50986 24728 50988
rect 24672 50934 24674 50986
rect 24674 50934 24726 50986
rect 24726 50934 24728 50986
rect 24672 50932 24728 50934
rect 24668 50428 24724 50484
rect 24220 49922 24276 49924
rect 24220 49870 24222 49922
rect 24222 49870 24274 49922
rect 24274 49870 24276 49922
rect 24220 49868 24276 49870
rect 23772 49196 23828 49252
rect 23804 48634 23860 48636
rect 23804 48582 23806 48634
rect 23806 48582 23858 48634
rect 23858 48582 23860 48634
rect 23804 48580 23860 48582
rect 23908 48634 23964 48636
rect 23908 48582 23910 48634
rect 23910 48582 23962 48634
rect 23962 48582 23964 48634
rect 23908 48580 23964 48582
rect 24012 48634 24068 48636
rect 24012 48582 24014 48634
rect 24014 48582 24066 48634
rect 24066 48582 24068 48634
rect 24012 48580 24068 48582
rect 24464 49418 24520 49420
rect 24464 49366 24466 49418
rect 24466 49366 24518 49418
rect 24518 49366 24520 49418
rect 24464 49364 24520 49366
rect 24568 49418 24624 49420
rect 24568 49366 24570 49418
rect 24570 49366 24622 49418
rect 24622 49366 24624 49418
rect 24568 49364 24624 49366
rect 24672 49418 24728 49420
rect 24672 49366 24674 49418
rect 24674 49366 24726 49418
rect 24726 49366 24728 49418
rect 24672 49364 24728 49366
rect 24668 48860 24724 48916
rect 24892 48524 24948 48580
rect 24444 48018 24500 48020
rect 24444 47966 24446 48018
rect 24446 47966 24498 48018
rect 24498 47966 24500 48018
rect 24444 47964 24500 47966
rect 24668 47964 24724 48020
rect 24464 47850 24520 47852
rect 24464 47798 24466 47850
rect 24466 47798 24518 47850
rect 24518 47798 24520 47850
rect 24464 47796 24520 47798
rect 24568 47850 24624 47852
rect 24568 47798 24570 47850
rect 24570 47798 24622 47850
rect 24622 47798 24624 47850
rect 24568 47796 24624 47798
rect 24672 47850 24728 47852
rect 24672 47798 24674 47850
rect 24674 47798 24726 47850
rect 24726 47798 24728 47850
rect 24672 47796 24728 47798
rect 23804 47066 23860 47068
rect 23804 47014 23806 47066
rect 23806 47014 23858 47066
rect 23858 47014 23860 47066
rect 23804 47012 23860 47014
rect 23908 47066 23964 47068
rect 23908 47014 23910 47066
rect 23910 47014 23962 47066
rect 23962 47014 23964 47066
rect 23908 47012 23964 47014
rect 24012 47066 24068 47068
rect 24012 47014 24014 47066
rect 24014 47014 24066 47066
rect 24066 47014 24068 47066
rect 24012 47012 24068 47014
rect 24668 46844 24724 46900
rect 23804 45498 23860 45500
rect 23804 45446 23806 45498
rect 23806 45446 23858 45498
rect 23858 45446 23860 45498
rect 23804 45444 23860 45446
rect 23908 45498 23964 45500
rect 23908 45446 23910 45498
rect 23910 45446 23962 45498
rect 23962 45446 23964 45498
rect 23908 45444 23964 45446
rect 24012 45498 24068 45500
rect 24012 45446 24014 45498
rect 24014 45446 24066 45498
rect 24066 45446 24068 45498
rect 24012 45444 24068 45446
rect 23804 43930 23860 43932
rect 23804 43878 23806 43930
rect 23806 43878 23858 43930
rect 23858 43878 23860 43930
rect 23804 43876 23860 43878
rect 23908 43930 23964 43932
rect 23908 43878 23910 43930
rect 23910 43878 23962 43930
rect 23962 43878 23964 43930
rect 23908 43876 23964 43878
rect 24012 43930 24068 43932
rect 24012 43878 24014 43930
rect 24014 43878 24066 43930
rect 24066 43878 24068 43930
rect 24012 43876 24068 43878
rect 24464 46282 24520 46284
rect 24464 46230 24466 46282
rect 24466 46230 24518 46282
rect 24518 46230 24520 46282
rect 24464 46228 24520 46230
rect 24568 46282 24624 46284
rect 24568 46230 24570 46282
rect 24570 46230 24622 46282
rect 24622 46230 24624 46282
rect 24568 46228 24624 46230
rect 24672 46282 24728 46284
rect 24672 46230 24674 46282
rect 24674 46230 24726 46282
rect 24726 46230 24728 46282
rect 24672 46228 24728 46230
rect 24780 45890 24836 45892
rect 24780 45838 24782 45890
rect 24782 45838 24834 45890
rect 24834 45838 24836 45890
rect 24780 45836 24836 45838
rect 24464 44714 24520 44716
rect 24464 44662 24466 44714
rect 24466 44662 24518 44714
rect 24518 44662 24520 44714
rect 24464 44660 24520 44662
rect 24568 44714 24624 44716
rect 24568 44662 24570 44714
rect 24570 44662 24622 44714
rect 24622 44662 24624 44714
rect 24568 44660 24624 44662
rect 24672 44714 24728 44716
rect 24672 44662 24674 44714
rect 24674 44662 24726 44714
rect 24726 44662 24728 44714
rect 24672 44660 24728 44662
rect 24668 44322 24724 44324
rect 24668 44270 24670 44322
rect 24670 44270 24722 44322
rect 24722 44270 24724 44322
rect 24668 44268 24724 44270
rect 25004 47964 25060 48020
rect 24464 43146 24520 43148
rect 24464 43094 24466 43146
rect 24466 43094 24518 43146
rect 24518 43094 24520 43146
rect 24464 43092 24520 43094
rect 24568 43146 24624 43148
rect 24568 43094 24570 43146
rect 24570 43094 24622 43146
rect 24622 43094 24624 43146
rect 24568 43092 24624 43094
rect 24672 43146 24728 43148
rect 24672 43094 24674 43146
rect 24674 43094 24726 43146
rect 24726 43094 24728 43146
rect 24672 43092 24728 43094
rect 24220 42924 24276 42980
rect 24668 42754 24724 42756
rect 24668 42702 24670 42754
rect 24670 42702 24722 42754
rect 24722 42702 24724 42754
rect 24668 42700 24724 42702
rect 23804 42362 23860 42364
rect 23804 42310 23806 42362
rect 23806 42310 23858 42362
rect 23858 42310 23860 42362
rect 23804 42308 23860 42310
rect 23908 42362 23964 42364
rect 23908 42310 23910 42362
rect 23910 42310 23962 42362
rect 23962 42310 23964 42362
rect 23908 42308 23964 42310
rect 24012 42362 24068 42364
rect 24012 42310 24014 42362
rect 24014 42310 24066 42362
rect 24066 42310 24068 42362
rect 24012 42308 24068 42310
rect 24892 41916 24948 41972
rect 24464 41578 24520 41580
rect 24464 41526 24466 41578
rect 24466 41526 24518 41578
rect 24518 41526 24520 41578
rect 24464 41524 24520 41526
rect 24568 41578 24624 41580
rect 24568 41526 24570 41578
rect 24570 41526 24622 41578
rect 24622 41526 24624 41578
rect 24568 41524 24624 41526
rect 24672 41578 24728 41580
rect 24672 41526 24674 41578
rect 24674 41526 24726 41578
rect 24726 41526 24728 41578
rect 24672 41524 24728 41526
rect 23804 40794 23860 40796
rect 23804 40742 23806 40794
rect 23806 40742 23858 40794
rect 23858 40742 23860 40794
rect 23804 40740 23860 40742
rect 23908 40794 23964 40796
rect 23908 40742 23910 40794
rect 23910 40742 23962 40794
rect 23962 40742 23964 40794
rect 23908 40740 23964 40742
rect 24012 40794 24068 40796
rect 24012 40742 24014 40794
rect 24014 40742 24066 40794
rect 24066 40742 24068 40794
rect 24012 40740 24068 40742
rect 24892 40572 24948 40628
rect 24668 40460 24724 40516
rect 24464 40010 24520 40012
rect 24464 39958 24466 40010
rect 24466 39958 24518 40010
rect 24518 39958 24520 40010
rect 24464 39956 24520 39958
rect 24568 40010 24624 40012
rect 24568 39958 24570 40010
rect 24570 39958 24622 40010
rect 24622 39958 24624 40010
rect 24568 39956 24624 39958
rect 24672 40010 24728 40012
rect 24672 39958 24674 40010
rect 24674 39958 24726 40010
rect 24726 39958 24728 40010
rect 24672 39956 24728 39958
rect 23804 39226 23860 39228
rect 23804 39174 23806 39226
rect 23806 39174 23858 39226
rect 23858 39174 23860 39226
rect 23804 39172 23860 39174
rect 23908 39226 23964 39228
rect 23908 39174 23910 39226
rect 23910 39174 23962 39226
rect 23962 39174 23964 39226
rect 23908 39172 23964 39174
rect 24012 39226 24068 39228
rect 24012 39174 24014 39226
rect 24014 39174 24066 39226
rect 24066 39174 24068 39226
rect 24012 39172 24068 39174
rect 24464 38442 24520 38444
rect 24464 38390 24466 38442
rect 24466 38390 24518 38442
rect 24518 38390 24520 38442
rect 24464 38388 24520 38390
rect 24568 38442 24624 38444
rect 24568 38390 24570 38442
rect 24570 38390 24622 38442
rect 24622 38390 24624 38442
rect 24568 38388 24624 38390
rect 24672 38442 24728 38444
rect 24672 38390 24674 38442
rect 24674 38390 24726 38442
rect 24726 38390 24728 38442
rect 24672 38388 24728 38390
rect 23804 37658 23860 37660
rect 23804 37606 23806 37658
rect 23806 37606 23858 37658
rect 23858 37606 23860 37658
rect 23804 37604 23860 37606
rect 23908 37658 23964 37660
rect 23908 37606 23910 37658
rect 23910 37606 23962 37658
rect 23962 37606 23964 37658
rect 23908 37604 23964 37606
rect 24012 37658 24068 37660
rect 24012 37606 24014 37658
rect 24014 37606 24066 37658
rect 24066 37606 24068 37658
rect 24012 37604 24068 37606
rect 23804 36090 23860 36092
rect 23804 36038 23806 36090
rect 23806 36038 23858 36090
rect 23858 36038 23860 36090
rect 23804 36036 23860 36038
rect 23908 36090 23964 36092
rect 23908 36038 23910 36090
rect 23910 36038 23962 36090
rect 23962 36038 23964 36090
rect 23908 36036 23964 36038
rect 24012 36090 24068 36092
rect 24012 36038 24014 36090
rect 24014 36038 24066 36090
rect 24066 36038 24068 36090
rect 24012 36036 24068 36038
rect 23804 34522 23860 34524
rect 23804 34470 23806 34522
rect 23806 34470 23858 34522
rect 23858 34470 23860 34522
rect 23804 34468 23860 34470
rect 23908 34522 23964 34524
rect 23908 34470 23910 34522
rect 23910 34470 23962 34522
rect 23962 34470 23964 34522
rect 23908 34468 23964 34470
rect 24012 34522 24068 34524
rect 24012 34470 24014 34522
rect 24014 34470 24066 34522
rect 24066 34470 24068 34522
rect 24012 34468 24068 34470
rect 23660 32956 23716 33012
rect 23804 32954 23860 32956
rect 23804 32902 23806 32954
rect 23806 32902 23858 32954
rect 23858 32902 23860 32954
rect 23804 32900 23860 32902
rect 23908 32954 23964 32956
rect 23908 32902 23910 32954
rect 23910 32902 23962 32954
rect 23962 32902 23964 32954
rect 23908 32900 23964 32902
rect 24012 32954 24068 32956
rect 24012 32902 24014 32954
rect 24014 32902 24066 32954
rect 24066 32902 24068 32954
rect 24012 32900 24068 32902
rect 23804 31386 23860 31388
rect 23804 31334 23806 31386
rect 23806 31334 23858 31386
rect 23858 31334 23860 31386
rect 23804 31332 23860 31334
rect 23908 31386 23964 31388
rect 23908 31334 23910 31386
rect 23910 31334 23962 31386
rect 23962 31334 23964 31386
rect 23908 31332 23964 31334
rect 24012 31386 24068 31388
rect 24012 31334 24014 31386
rect 24014 31334 24066 31386
rect 24066 31334 24068 31386
rect 24012 31332 24068 31334
rect 23804 29818 23860 29820
rect 23804 29766 23806 29818
rect 23806 29766 23858 29818
rect 23858 29766 23860 29818
rect 23804 29764 23860 29766
rect 23908 29818 23964 29820
rect 23908 29766 23910 29818
rect 23910 29766 23962 29818
rect 23962 29766 23964 29818
rect 23908 29764 23964 29766
rect 24012 29818 24068 29820
rect 24012 29766 24014 29818
rect 24014 29766 24066 29818
rect 24066 29766 24068 29818
rect 24012 29764 24068 29766
rect 24464 36874 24520 36876
rect 24464 36822 24466 36874
rect 24466 36822 24518 36874
rect 24518 36822 24520 36874
rect 24464 36820 24520 36822
rect 24568 36874 24624 36876
rect 24568 36822 24570 36874
rect 24570 36822 24622 36874
rect 24622 36822 24624 36874
rect 24568 36820 24624 36822
rect 24672 36874 24728 36876
rect 24672 36822 24674 36874
rect 24674 36822 24726 36874
rect 24726 36822 24728 36874
rect 24672 36820 24728 36822
rect 24668 36482 24724 36484
rect 24668 36430 24670 36482
rect 24670 36430 24722 36482
rect 24722 36430 24724 36482
rect 24668 36428 24724 36430
rect 24464 35306 24520 35308
rect 24464 35254 24466 35306
rect 24466 35254 24518 35306
rect 24518 35254 24520 35306
rect 24464 35252 24520 35254
rect 24568 35306 24624 35308
rect 24568 35254 24570 35306
rect 24570 35254 24622 35306
rect 24622 35254 24624 35306
rect 24568 35252 24624 35254
rect 24672 35306 24728 35308
rect 24672 35254 24674 35306
rect 24674 35254 24726 35306
rect 24726 35254 24728 35306
rect 24672 35252 24728 35254
rect 24892 34188 24948 34244
rect 24780 33852 24836 33908
rect 24464 33738 24520 33740
rect 24464 33686 24466 33738
rect 24466 33686 24518 33738
rect 24518 33686 24520 33738
rect 24464 33684 24520 33686
rect 24568 33738 24624 33740
rect 24568 33686 24570 33738
rect 24570 33686 24622 33738
rect 24622 33686 24624 33738
rect 24568 33684 24624 33686
rect 24672 33738 24728 33740
rect 24672 33686 24674 33738
rect 24674 33686 24726 33738
rect 24726 33686 24728 33738
rect 24672 33684 24728 33686
rect 24892 33346 24948 33348
rect 24892 33294 24894 33346
rect 24894 33294 24946 33346
rect 24946 33294 24948 33346
rect 24892 33292 24948 33294
rect 24892 32732 24948 32788
rect 24464 32170 24520 32172
rect 24464 32118 24466 32170
rect 24466 32118 24518 32170
rect 24518 32118 24520 32170
rect 24464 32116 24520 32118
rect 24568 32170 24624 32172
rect 24568 32118 24570 32170
rect 24570 32118 24622 32170
rect 24622 32118 24624 32170
rect 24568 32116 24624 32118
rect 24672 32170 24728 32172
rect 24672 32118 24674 32170
rect 24674 32118 24726 32170
rect 24726 32118 24728 32170
rect 24672 32116 24728 32118
rect 24780 30716 24836 30772
rect 24464 30602 24520 30604
rect 24464 30550 24466 30602
rect 24466 30550 24518 30602
rect 24518 30550 24520 30602
rect 24464 30548 24520 30550
rect 24568 30602 24624 30604
rect 24568 30550 24570 30602
rect 24570 30550 24622 30602
rect 24622 30550 24624 30602
rect 24568 30548 24624 30550
rect 24672 30602 24728 30604
rect 24672 30550 24674 30602
rect 24674 30550 24726 30602
rect 24726 30550 24728 30602
rect 24672 30548 24728 30550
rect 24332 29036 24388 29092
rect 24892 30044 24948 30100
rect 24464 29034 24520 29036
rect 24464 28982 24466 29034
rect 24466 28982 24518 29034
rect 24518 28982 24520 29034
rect 24464 28980 24520 28982
rect 24568 29034 24624 29036
rect 24568 28982 24570 29034
rect 24570 28982 24622 29034
rect 24622 28982 24624 29034
rect 24568 28980 24624 28982
rect 24672 29034 24728 29036
rect 24672 28982 24674 29034
rect 24674 28982 24726 29034
rect 24726 28982 24728 29034
rect 24672 28980 24728 28982
rect 24220 28588 24276 28644
rect 24668 28364 24724 28420
rect 23804 28250 23860 28252
rect 23804 28198 23806 28250
rect 23806 28198 23858 28250
rect 23858 28198 23860 28250
rect 23804 28196 23860 28198
rect 23908 28250 23964 28252
rect 23908 28198 23910 28250
rect 23910 28198 23962 28250
rect 23962 28198 23964 28250
rect 23908 28196 23964 28198
rect 24012 28250 24068 28252
rect 24012 28198 24014 28250
rect 24014 28198 24066 28250
rect 24066 28198 24068 28250
rect 24012 28196 24068 28198
rect 24464 27466 24520 27468
rect 24464 27414 24466 27466
rect 24466 27414 24518 27466
rect 24518 27414 24520 27466
rect 24464 27412 24520 27414
rect 24568 27466 24624 27468
rect 24568 27414 24570 27466
rect 24570 27414 24622 27466
rect 24622 27414 24624 27466
rect 24568 27412 24624 27414
rect 24672 27466 24728 27468
rect 24672 27414 24674 27466
rect 24674 27414 24726 27466
rect 24726 27414 24728 27466
rect 24672 27412 24728 27414
rect 24668 27186 24724 27188
rect 24668 27134 24670 27186
rect 24670 27134 24722 27186
rect 24722 27134 24724 27186
rect 24668 27132 24724 27134
rect 23804 26682 23860 26684
rect 23804 26630 23806 26682
rect 23806 26630 23858 26682
rect 23858 26630 23860 26682
rect 23804 26628 23860 26630
rect 23908 26682 23964 26684
rect 23908 26630 23910 26682
rect 23910 26630 23962 26682
rect 23962 26630 23964 26682
rect 23908 26628 23964 26630
rect 24012 26682 24068 26684
rect 24012 26630 24014 26682
rect 24014 26630 24066 26682
rect 24066 26630 24068 26682
rect 24012 26628 24068 26630
rect 24464 25898 24520 25900
rect 24464 25846 24466 25898
rect 24466 25846 24518 25898
rect 24518 25846 24520 25898
rect 24464 25844 24520 25846
rect 24568 25898 24624 25900
rect 24568 25846 24570 25898
rect 24570 25846 24622 25898
rect 24622 25846 24624 25898
rect 24568 25844 24624 25846
rect 24672 25898 24728 25900
rect 24672 25846 24674 25898
rect 24674 25846 24726 25898
rect 24726 25846 24728 25898
rect 24672 25844 24728 25846
rect 24668 25618 24724 25620
rect 24668 25566 24670 25618
rect 24670 25566 24722 25618
rect 24722 25566 24724 25618
rect 24668 25564 24724 25566
rect 23804 25114 23860 25116
rect 23804 25062 23806 25114
rect 23806 25062 23858 25114
rect 23858 25062 23860 25114
rect 23804 25060 23860 25062
rect 23908 25114 23964 25116
rect 23908 25062 23910 25114
rect 23910 25062 23962 25114
rect 23962 25062 23964 25114
rect 23908 25060 23964 25062
rect 24012 25114 24068 25116
rect 24012 25062 24014 25114
rect 24014 25062 24066 25114
rect 24066 25062 24068 25114
rect 24012 25060 24068 25062
rect 24668 24444 24724 24500
rect 24464 24330 24520 24332
rect 24464 24278 24466 24330
rect 24466 24278 24518 24330
rect 24518 24278 24520 24330
rect 24464 24276 24520 24278
rect 24568 24330 24624 24332
rect 24568 24278 24570 24330
rect 24570 24278 24622 24330
rect 24622 24278 24624 24330
rect 24568 24276 24624 24278
rect 24672 24330 24728 24332
rect 24672 24278 24674 24330
rect 24674 24278 24726 24330
rect 24726 24278 24728 24330
rect 24672 24276 24728 24278
rect 25004 26124 25060 26180
rect 23804 23546 23860 23548
rect 23804 23494 23806 23546
rect 23806 23494 23858 23546
rect 23858 23494 23860 23546
rect 23804 23492 23860 23494
rect 23908 23546 23964 23548
rect 23908 23494 23910 23546
rect 23910 23494 23962 23546
rect 23962 23494 23964 23546
rect 23908 23492 23964 23494
rect 24012 23546 24068 23548
rect 24012 23494 24014 23546
rect 24014 23494 24066 23546
rect 24066 23494 24068 23546
rect 24012 23492 24068 23494
rect 24464 22762 24520 22764
rect 24464 22710 24466 22762
rect 24466 22710 24518 22762
rect 24518 22710 24520 22762
rect 24464 22708 24520 22710
rect 24568 22762 24624 22764
rect 24568 22710 24570 22762
rect 24570 22710 24622 22762
rect 24622 22710 24624 22762
rect 24568 22708 24624 22710
rect 24672 22762 24728 22764
rect 24672 22710 24674 22762
rect 24674 22710 24726 22762
rect 24726 22710 24728 22762
rect 24672 22708 24728 22710
rect 23804 21978 23860 21980
rect 23804 21926 23806 21978
rect 23806 21926 23858 21978
rect 23858 21926 23860 21978
rect 23804 21924 23860 21926
rect 23908 21978 23964 21980
rect 23908 21926 23910 21978
rect 23910 21926 23962 21978
rect 23962 21926 23964 21978
rect 23908 21924 23964 21926
rect 24012 21978 24068 21980
rect 24012 21926 24014 21978
rect 24014 21926 24066 21978
rect 24066 21926 24068 21978
rect 24012 21924 24068 21926
rect 24464 21194 24520 21196
rect 24464 21142 24466 21194
rect 24466 21142 24518 21194
rect 24518 21142 24520 21194
rect 24464 21140 24520 21142
rect 24568 21194 24624 21196
rect 24568 21142 24570 21194
rect 24570 21142 24622 21194
rect 24622 21142 24624 21194
rect 24568 21140 24624 21142
rect 24672 21194 24728 21196
rect 24672 21142 24674 21194
rect 24674 21142 24726 21194
rect 24726 21142 24728 21194
rect 24672 21140 24728 21142
rect 23804 20410 23860 20412
rect 23804 20358 23806 20410
rect 23806 20358 23858 20410
rect 23858 20358 23860 20410
rect 23804 20356 23860 20358
rect 23908 20410 23964 20412
rect 23908 20358 23910 20410
rect 23910 20358 23962 20410
rect 23962 20358 23964 20410
rect 23908 20356 23964 20358
rect 24012 20410 24068 20412
rect 24012 20358 24014 20410
rect 24014 20358 24066 20410
rect 24066 20358 24068 20410
rect 24012 20356 24068 20358
rect 24464 19626 24520 19628
rect 24464 19574 24466 19626
rect 24466 19574 24518 19626
rect 24518 19574 24520 19626
rect 24464 19572 24520 19574
rect 24568 19626 24624 19628
rect 24568 19574 24570 19626
rect 24570 19574 24622 19626
rect 24622 19574 24624 19626
rect 24568 19572 24624 19574
rect 24672 19626 24728 19628
rect 24672 19574 24674 19626
rect 24674 19574 24726 19626
rect 24726 19574 24728 19626
rect 24672 19572 24728 19574
rect 23804 18842 23860 18844
rect 23804 18790 23806 18842
rect 23806 18790 23858 18842
rect 23858 18790 23860 18842
rect 23804 18788 23860 18790
rect 23908 18842 23964 18844
rect 23908 18790 23910 18842
rect 23910 18790 23962 18842
rect 23962 18790 23964 18842
rect 23908 18788 23964 18790
rect 24012 18842 24068 18844
rect 24012 18790 24014 18842
rect 24014 18790 24066 18842
rect 24066 18790 24068 18842
rect 24012 18788 24068 18790
rect 24464 18058 24520 18060
rect 24464 18006 24466 18058
rect 24466 18006 24518 18058
rect 24518 18006 24520 18058
rect 24464 18004 24520 18006
rect 24568 18058 24624 18060
rect 24568 18006 24570 18058
rect 24570 18006 24622 18058
rect 24622 18006 24624 18058
rect 24568 18004 24624 18006
rect 24672 18058 24728 18060
rect 24672 18006 24674 18058
rect 24674 18006 24726 18058
rect 24726 18006 24728 18058
rect 24672 18004 24728 18006
rect 23804 17274 23860 17276
rect 23804 17222 23806 17274
rect 23806 17222 23858 17274
rect 23858 17222 23860 17274
rect 23804 17220 23860 17222
rect 23908 17274 23964 17276
rect 23908 17222 23910 17274
rect 23910 17222 23962 17274
rect 23962 17222 23964 17274
rect 23908 17220 23964 17222
rect 24012 17274 24068 17276
rect 24012 17222 24014 17274
rect 24014 17222 24066 17274
rect 24066 17222 24068 17274
rect 24012 17220 24068 17222
rect 24464 16490 24520 16492
rect 24464 16438 24466 16490
rect 24466 16438 24518 16490
rect 24518 16438 24520 16490
rect 24464 16436 24520 16438
rect 24568 16490 24624 16492
rect 24568 16438 24570 16490
rect 24570 16438 24622 16490
rect 24622 16438 24624 16490
rect 24568 16436 24624 16438
rect 24672 16490 24728 16492
rect 24672 16438 24674 16490
rect 24674 16438 24726 16490
rect 24726 16438 24728 16490
rect 24672 16436 24728 16438
rect 23804 15706 23860 15708
rect 23804 15654 23806 15706
rect 23806 15654 23858 15706
rect 23858 15654 23860 15706
rect 23804 15652 23860 15654
rect 23908 15706 23964 15708
rect 23908 15654 23910 15706
rect 23910 15654 23962 15706
rect 23962 15654 23964 15706
rect 23908 15652 23964 15654
rect 24012 15706 24068 15708
rect 24012 15654 24014 15706
rect 24014 15654 24066 15706
rect 24066 15654 24068 15706
rect 24012 15652 24068 15654
rect 24464 14922 24520 14924
rect 24464 14870 24466 14922
rect 24466 14870 24518 14922
rect 24518 14870 24520 14922
rect 24464 14868 24520 14870
rect 24568 14922 24624 14924
rect 24568 14870 24570 14922
rect 24570 14870 24622 14922
rect 24622 14870 24624 14922
rect 24568 14868 24624 14870
rect 24672 14922 24728 14924
rect 24672 14870 24674 14922
rect 24674 14870 24726 14922
rect 24726 14870 24728 14922
rect 24672 14868 24728 14870
rect 23804 14138 23860 14140
rect 23804 14086 23806 14138
rect 23806 14086 23858 14138
rect 23858 14086 23860 14138
rect 23804 14084 23860 14086
rect 23908 14138 23964 14140
rect 23908 14086 23910 14138
rect 23910 14086 23962 14138
rect 23962 14086 23964 14138
rect 23908 14084 23964 14086
rect 24012 14138 24068 14140
rect 24012 14086 24014 14138
rect 24014 14086 24066 14138
rect 24066 14086 24068 14138
rect 24012 14084 24068 14086
rect 23884 13580 23940 13636
rect 23884 13356 23940 13412
rect 24464 13354 24520 13356
rect 24464 13302 24466 13354
rect 24466 13302 24518 13354
rect 24518 13302 24520 13354
rect 24464 13300 24520 13302
rect 24568 13354 24624 13356
rect 24568 13302 24570 13354
rect 24570 13302 24622 13354
rect 24622 13302 24624 13354
rect 24568 13300 24624 13302
rect 24672 13354 24728 13356
rect 24672 13302 24674 13354
rect 24674 13302 24726 13354
rect 24726 13302 24728 13354
rect 24672 13300 24728 13302
rect 25564 50482 25620 50484
rect 25564 50430 25566 50482
rect 25566 50430 25618 50482
rect 25618 50430 25620 50482
rect 25564 50428 25620 50430
rect 25452 49532 25508 49588
rect 25564 48636 25620 48692
rect 27580 56028 27636 56084
rect 26236 55298 26292 55300
rect 26236 55246 26238 55298
rect 26238 55246 26290 55298
rect 26290 55246 26292 55298
rect 26236 55244 26292 55246
rect 26236 54236 26292 54292
rect 26236 53730 26292 53732
rect 26236 53678 26238 53730
rect 26238 53678 26290 53730
rect 26290 53678 26292 53730
rect 26236 53676 26292 53678
rect 27244 54012 27300 54068
rect 27020 53116 27076 53172
rect 26236 52332 26292 52388
rect 26236 52162 26292 52164
rect 26236 52110 26238 52162
rect 26238 52110 26290 52162
rect 26290 52110 26292 52162
rect 26236 52108 26292 52110
rect 27244 52220 27300 52276
rect 27356 52892 27412 52948
rect 27132 51324 27188 51380
rect 26236 51266 26292 51268
rect 26236 51214 26238 51266
rect 26238 51214 26290 51266
rect 26290 51214 26292 51266
rect 26236 51212 26292 51214
rect 26236 50706 26292 50708
rect 26236 50654 26238 50706
rect 26238 50654 26290 50706
rect 26290 50654 26292 50706
rect 26236 50652 26292 50654
rect 27244 50876 27300 50932
rect 27020 49980 27076 50036
rect 26236 49026 26292 49028
rect 26236 48974 26238 49026
rect 26238 48974 26290 49026
rect 26290 48974 26292 49026
rect 26236 48972 26292 48974
rect 26348 48748 26404 48804
rect 27244 49084 27300 49140
rect 27132 48188 27188 48244
rect 26236 48130 26292 48132
rect 26236 48078 26238 48130
rect 26238 48078 26290 48130
rect 26290 48078 26292 48130
rect 26236 48076 26292 48078
rect 25340 48018 25396 48020
rect 25340 47966 25342 48018
rect 25342 47966 25394 48018
rect 25394 47966 25396 48018
rect 25340 47964 25396 47966
rect 25676 47346 25732 47348
rect 25676 47294 25678 47346
rect 25678 47294 25730 47346
rect 25730 47294 25732 47346
rect 25676 47292 25732 47294
rect 27244 47740 27300 47796
rect 27020 46844 27076 46900
rect 26236 46732 26292 46788
rect 26236 46562 26292 46564
rect 26236 46510 26238 46562
rect 26238 46510 26290 46562
rect 26290 46510 26292 46562
rect 26236 46508 26292 46510
rect 25676 46396 25732 46452
rect 25676 45500 25732 45556
rect 25676 44210 25732 44212
rect 25676 44158 25678 44210
rect 25678 44158 25730 44210
rect 25730 44158 25732 44210
rect 25676 44156 25732 44158
rect 25676 43260 25732 43316
rect 25676 42364 25732 42420
rect 25676 41074 25732 41076
rect 25676 41022 25678 41074
rect 25678 41022 25730 41074
rect 25730 41022 25732 41074
rect 25676 41020 25732 41022
rect 25676 40124 25732 40180
rect 25676 39228 25732 39284
rect 25452 38556 25508 38612
rect 25676 37938 25732 37940
rect 25676 37886 25678 37938
rect 25678 37886 25730 37938
rect 25730 37886 25732 37938
rect 25676 37884 25732 37886
rect 25452 36988 25508 37044
rect 25788 37100 25844 37156
rect 25676 36092 25732 36148
rect 25340 35532 25396 35588
rect 25228 34860 25284 34916
rect 25676 34802 25732 34804
rect 25676 34750 25678 34802
rect 25678 34750 25730 34802
rect 25730 34750 25732 34802
rect 25676 34748 25732 34750
rect 25676 33852 25732 33908
rect 25788 33516 25844 33572
rect 25676 32956 25732 33012
rect 25228 27804 25284 27860
rect 25340 32844 25396 32900
rect 25228 26348 25284 26404
rect 25228 24668 25284 24724
rect 25564 32732 25620 32788
rect 25452 30716 25508 30772
rect 25452 29932 25508 29988
rect 25676 31666 25732 31668
rect 25676 31614 25678 31666
rect 25678 31614 25730 31666
rect 25730 31614 25732 31666
rect 25676 31612 25732 31614
rect 25676 27132 25732 27188
rect 25564 26348 25620 26404
rect 25676 26236 25732 26292
rect 25452 24780 25508 24836
rect 25564 25900 25620 25956
rect 25452 23996 25508 24052
rect 25340 20188 25396 20244
rect 25116 14700 25172 14756
rect 24892 12684 24948 12740
rect 23804 12570 23860 12572
rect 23804 12518 23806 12570
rect 23806 12518 23858 12570
rect 23858 12518 23860 12570
rect 23804 12516 23860 12518
rect 23908 12570 23964 12572
rect 23908 12518 23910 12570
rect 23910 12518 23962 12570
rect 23962 12518 23964 12570
rect 23908 12516 23964 12518
rect 24012 12570 24068 12572
rect 24012 12518 24014 12570
rect 24014 12518 24066 12570
rect 24066 12518 24068 12570
rect 24012 12516 24068 12518
rect 25676 24892 25732 24948
rect 25788 25116 25844 25172
rect 25676 23100 25732 23156
rect 25676 21756 25732 21812
rect 26236 41858 26292 41860
rect 26236 41806 26238 41858
rect 26238 41806 26290 41858
rect 26290 41806 26292 41858
rect 26236 41804 26292 41806
rect 26796 45836 26852 45892
rect 26348 41356 26404 41412
rect 26236 41186 26292 41188
rect 26236 41134 26238 41186
rect 26238 41134 26290 41186
rect 26290 41134 26292 41186
rect 26236 41132 26292 41134
rect 26236 39618 26292 39620
rect 26236 39566 26238 39618
rect 26238 39566 26290 39618
rect 26290 39566 26292 39618
rect 26236 39564 26292 39566
rect 26348 38668 26404 38724
rect 26236 38050 26292 38052
rect 26236 37998 26238 38050
rect 26238 37998 26290 38050
rect 26290 37998 26292 38050
rect 26236 37996 26292 37998
rect 26236 37154 26292 37156
rect 26236 37102 26238 37154
rect 26238 37102 26290 37154
rect 26290 37102 26292 37154
rect 26236 37100 26292 37102
rect 26124 34972 26180 35028
rect 26236 34914 26292 34916
rect 26236 34862 26238 34914
rect 26238 34862 26290 34914
rect 26290 34862 26292 34914
rect 26236 34860 26292 34862
rect 26348 34300 26404 34356
rect 26236 34018 26292 34020
rect 26236 33966 26238 34018
rect 26238 33966 26290 34018
rect 26290 33966 26292 34018
rect 26236 33964 26292 33966
rect 26460 32844 26516 32900
rect 26572 32732 26628 32788
rect 26684 33292 26740 33348
rect 26236 32620 26292 32676
rect 26124 30380 26180 30436
rect 26236 29314 26292 29316
rect 26236 29262 26238 29314
rect 26238 29262 26290 29314
rect 26290 29262 26292 29314
rect 26236 29260 26292 29262
rect 26348 28028 26404 28084
rect 26236 27580 26292 27636
rect 26236 26012 26292 26068
rect 26124 25900 26180 25956
rect 26236 25506 26292 25508
rect 26236 25454 26238 25506
rect 26238 25454 26290 25506
rect 26290 25454 26292 25506
rect 26236 25452 26292 25454
rect 26572 28700 26628 28756
rect 26460 25116 26516 25172
rect 26348 25004 26404 25060
rect 25900 22540 25956 22596
rect 26012 24780 26068 24836
rect 25900 20860 25956 20916
rect 26236 24108 26292 24164
rect 26236 23212 26292 23268
rect 26236 22482 26292 22484
rect 26236 22430 26238 22482
rect 26238 22430 26290 22482
rect 26290 22430 26292 22482
rect 26236 22428 26292 22430
rect 26124 21644 26180 21700
rect 25564 19852 25620 19908
rect 26012 20076 26068 20132
rect 25900 19292 25956 19348
rect 26236 21308 26292 21364
rect 26348 20972 26404 21028
rect 26460 22092 26516 22148
rect 26348 18396 26404 18452
rect 26124 17836 26180 17892
rect 25900 16156 25956 16212
rect 25676 13020 25732 13076
rect 25788 16044 25844 16100
rect 25452 12348 25508 12404
rect 24464 11786 24520 11788
rect 24464 11734 24466 11786
rect 24466 11734 24518 11786
rect 24518 11734 24520 11786
rect 24464 11732 24520 11734
rect 24568 11786 24624 11788
rect 24568 11734 24570 11786
rect 24570 11734 24622 11786
rect 24622 11734 24624 11786
rect 24568 11732 24624 11734
rect 24672 11786 24728 11788
rect 24672 11734 24674 11786
rect 24674 11734 24726 11786
rect 24726 11734 24728 11786
rect 24672 11732 24728 11734
rect 23804 11002 23860 11004
rect 23804 10950 23806 11002
rect 23806 10950 23858 11002
rect 23858 10950 23860 11002
rect 23804 10948 23860 10950
rect 23908 11002 23964 11004
rect 23908 10950 23910 11002
rect 23910 10950 23962 11002
rect 23962 10950 23964 11002
rect 23908 10948 23964 10950
rect 24012 11002 24068 11004
rect 24012 10950 24014 11002
rect 24014 10950 24066 11002
rect 24066 10950 24068 11002
rect 24012 10948 24068 10950
rect 24464 10218 24520 10220
rect 24464 10166 24466 10218
rect 24466 10166 24518 10218
rect 24518 10166 24520 10218
rect 24464 10164 24520 10166
rect 24568 10218 24624 10220
rect 24568 10166 24570 10218
rect 24570 10166 24622 10218
rect 24622 10166 24624 10218
rect 24568 10164 24624 10166
rect 24672 10218 24728 10220
rect 24672 10166 24674 10218
rect 24674 10166 24726 10218
rect 24726 10166 24728 10218
rect 24672 10164 24728 10166
rect 26012 15986 26068 15988
rect 26012 15934 26014 15986
rect 26014 15934 26066 15986
rect 26066 15934 26068 15986
rect 26012 15932 26068 15934
rect 26236 15260 26292 15316
rect 26012 13132 26068 13188
rect 26012 12290 26068 12292
rect 26012 12238 26014 12290
rect 26014 12238 26066 12290
rect 26066 12238 26068 12290
rect 26012 12236 26068 12238
rect 26124 11900 26180 11956
rect 26012 9996 26068 10052
rect 23804 9434 23860 9436
rect 23804 9382 23806 9434
rect 23806 9382 23858 9434
rect 23858 9382 23860 9434
rect 23804 9380 23860 9382
rect 23908 9434 23964 9436
rect 23908 9382 23910 9434
rect 23910 9382 23962 9434
rect 23962 9382 23964 9434
rect 23908 9380 23964 9382
rect 24012 9434 24068 9436
rect 24012 9382 24014 9434
rect 24014 9382 24066 9434
rect 24066 9382 24068 9434
rect 24012 9380 24068 9382
rect 25788 9212 25844 9268
rect 24464 8650 24520 8652
rect 24464 8598 24466 8650
rect 24466 8598 24518 8650
rect 24518 8598 24520 8650
rect 24464 8596 24520 8598
rect 24568 8650 24624 8652
rect 24568 8598 24570 8650
rect 24570 8598 24622 8650
rect 24622 8598 24624 8650
rect 24568 8596 24624 8598
rect 24672 8650 24728 8652
rect 24672 8598 24674 8650
rect 24674 8598 24726 8650
rect 24726 8598 24728 8650
rect 24672 8596 24728 8598
rect 23804 7866 23860 7868
rect 23804 7814 23806 7866
rect 23806 7814 23858 7866
rect 23858 7814 23860 7866
rect 23804 7812 23860 7814
rect 23908 7866 23964 7868
rect 23908 7814 23910 7866
rect 23910 7814 23962 7866
rect 23962 7814 23964 7866
rect 23908 7812 23964 7814
rect 24012 7866 24068 7868
rect 24012 7814 24014 7866
rect 24014 7814 24066 7866
rect 24066 7814 24068 7866
rect 24012 7812 24068 7814
rect 24464 7082 24520 7084
rect 24464 7030 24466 7082
rect 24466 7030 24518 7082
rect 24518 7030 24520 7082
rect 24464 7028 24520 7030
rect 24568 7082 24624 7084
rect 24568 7030 24570 7082
rect 24570 7030 24622 7082
rect 24622 7030 24624 7082
rect 24568 7028 24624 7030
rect 24672 7082 24728 7084
rect 24672 7030 24674 7082
rect 24674 7030 24726 7082
rect 24726 7030 24728 7082
rect 24672 7028 24728 7030
rect 23436 6748 23492 6804
rect 23804 6298 23860 6300
rect 23804 6246 23806 6298
rect 23806 6246 23858 6298
rect 23858 6246 23860 6298
rect 23804 6244 23860 6246
rect 23908 6298 23964 6300
rect 23908 6246 23910 6298
rect 23910 6246 23962 6298
rect 23962 6246 23964 6298
rect 23908 6244 23964 6246
rect 24012 6298 24068 6300
rect 24012 6246 24014 6298
rect 24014 6246 24066 6298
rect 24066 6246 24068 6298
rect 24012 6244 24068 6246
rect 24464 5514 24520 5516
rect 24464 5462 24466 5514
rect 24466 5462 24518 5514
rect 24518 5462 24520 5514
rect 24464 5460 24520 5462
rect 24568 5514 24624 5516
rect 24568 5462 24570 5514
rect 24570 5462 24622 5514
rect 24622 5462 24624 5514
rect 24568 5460 24624 5462
rect 24672 5514 24728 5516
rect 24672 5462 24674 5514
rect 24674 5462 24726 5514
rect 24726 5462 24728 5514
rect 24672 5460 24728 5462
rect 23804 4730 23860 4732
rect 23804 4678 23806 4730
rect 23806 4678 23858 4730
rect 23858 4678 23860 4730
rect 23804 4676 23860 4678
rect 23908 4730 23964 4732
rect 23908 4678 23910 4730
rect 23910 4678 23962 4730
rect 23962 4678 23964 4730
rect 23908 4676 23964 4678
rect 24012 4730 24068 4732
rect 24012 4678 24014 4730
rect 24014 4678 24066 4730
rect 24066 4678 24068 4730
rect 24012 4676 24068 4678
rect 24464 3946 24520 3948
rect 24464 3894 24466 3946
rect 24466 3894 24518 3946
rect 24518 3894 24520 3946
rect 24464 3892 24520 3894
rect 24568 3946 24624 3948
rect 24568 3894 24570 3946
rect 24570 3894 24622 3946
rect 24622 3894 24624 3946
rect 24568 3892 24624 3894
rect 24672 3946 24728 3948
rect 24672 3894 24674 3946
rect 24674 3894 24726 3946
rect 24726 3894 24728 3946
rect 24672 3892 24728 3894
rect 23804 3162 23860 3164
rect 23804 3110 23806 3162
rect 23806 3110 23858 3162
rect 23858 3110 23860 3162
rect 23804 3108 23860 3110
rect 23908 3162 23964 3164
rect 23908 3110 23910 3162
rect 23910 3110 23962 3162
rect 23962 3110 23964 3162
rect 23908 3108 23964 3110
rect 24012 3162 24068 3164
rect 24012 3110 24014 3162
rect 24014 3110 24066 3162
rect 24066 3110 24068 3162
rect 24012 3108 24068 3110
rect 24464 2378 24520 2380
rect 24464 2326 24466 2378
rect 24466 2326 24518 2378
rect 24518 2326 24520 2378
rect 24464 2324 24520 2326
rect 24568 2378 24624 2380
rect 24568 2326 24570 2378
rect 24570 2326 24622 2378
rect 24622 2326 24624 2378
rect 24568 2324 24624 2326
rect 24672 2378 24728 2380
rect 24672 2326 24674 2378
rect 24674 2326 24726 2378
rect 24726 2326 24728 2378
rect 24672 2324 24728 2326
rect 26348 10780 26404 10836
rect 26572 19964 26628 20020
rect 26572 18620 26628 18676
rect 26684 18396 26740 18452
rect 26684 17724 26740 17780
rect 26572 16828 26628 16884
rect 26572 15484 26628 15540
rect 26684 14588 26740 14644
rect 26572 13692 26628 13748
rect 26572 12348 26628 12404
rect 26684 11452 26740 11508
rect 26572 10556 26628 10612
rect 26572 9212 26628 9268
rect 26012 6578 26068 6580
rect 26012 6526 26014 6578
rect 26014 6526 26066 6578
rect 26066 6526 26068 6578
rect 26012 6524 26068 6526
rect 26012 5794 26068 5796
rect 26012 5742 26014 5794
rect 26014 5742 26066 5794
rect 26066 5742 26068 5794
rect 26012 5740 26068 5742
rect 26684 8316 26740 8372
rect 27244 45948 27300 46004
rect 27132 45052 27188 45108
rect 27244 44604 27300 44660
rect 27020 43708 27076 43764
rect 27244 42812 27300 42868
rect 27132 41916 27188 41972
rect 27244 41468 27300 41524
rect 27020 40572 27076 40628
rect 27244 39676 27300 39732
rect 27132 38780 27188 38836
rect 27244 38332 27300 38388
rect 27020 37436 27076 37492
rect 27244 36540 27300 36596
rect 27132 35644 27188 35700
rect 27244 35196 27300 35252
rect 27020 34300 27076 34356
rect 27244 33404 27300 33460
rect 27132 32508 27188 32564
rect 27244 32060 27300 32116
rect 27020 31164 27076 31220
rect 27244 30268 27300 30324
rect 27020 29820 27076 29876
rect 27132 29372 27188 29428
rect 27244 28924 27300 28980
rect 27244 28530 27300 28532
rect 27244 28478 27246 28530
rect 27246 28478 27298 28530
rect 27298 28478 27300 28530
rect 27244 28476 27300 28478
rect 27244 28082 27300 28084
rect 27244 28030 27246 28082
rect 27246 28030 27298 28082
rect 27298 28030 27300 28082
rect 27244 28028 27300 28030
rect 27244 27580 27300 27636
rect 26908 27244 26964 27300
rect 27244 26684 27300 26740
rect 27020 26124 27076 26180
rect 27244 25788 27300 25844
rect 27132 25340 27188 25396
rect 27244 24444 27300 24500
rect 27132 23548 27188 23604
rect 27244 22652 27300 22708
rect 27132 22204 27188 22260
rect 27020 20130 27076 20132
rect 27020 20078 27022 20130
rect 27022 20078 27074 20130
rect 27074 20078 27076 20130
rect 27020 20076 27076 20078
rect 26908 18450 26964 18452
rect 26908 18398 26910 18450
rect 26910 18398 26962 18450
rect 26962 18398 26964 18450
rect 26908 18396 26964 18398
rect 26908 17836 26964 17892
rect 27020 17500 27076 17556
rect 27132 16268 27188 16324
rect 27020 14252 27076 14308
rect 26908 13804 26964 13860
rect 26908 13634 26964 13636
rect 26908 13582 26910 13634
rect 26910 13582 26962 13634
rect 26962 13582 26964 13634
rect 26908 13580 26964 13582
rect 27244 15036 27300 15092
rect 27244 13468 27300 13524
rect 26908 12290 26964 12292
rect 26908 12238 26910 12290
rect 26910 12238 26962 12290
rect 26962 12238 26964 12290
rect 26908 12236 26964 12238
rect 27020 12012 27076 12068
rect 26908 11282 26964 11284
rect 26908 11230 26910 11282
rect 26910 11230 26962 11282
rect 26962 11230 26964 11282
rect 26908 11228 26964 11230
rect 26908 10722 26964 10724
rect 26908 10670 26910 10722
rect 26910 10670 26962 10722
rect 26962 10670 26964 10722
rect 26908 10668 26964 10670
rect 26908 9938 26964 9940
rect 26908 9886 26910 9938
rect 26910 9886 26962 9938
rect 26962 9886 26964 9938
rect 26908 9884 26964 9886
rect 27020 8876 27076 8932
rect 26908 7980 26964 8036
rect 26796 7644 26852 7700
rect 26572 7532 26628 7588
rect 26908 7474 26964 7476
rect 26908 7422 26910 7474
rect 26910 7422 26962 7474
rect 26962 7422 26964 7474
rect 26908 7420 26964 7422
rect 26236 6748 26292 6804
rect 26012 3442 26068 3444
rect 26012 3390 26014 3442
rect 26014 3390 26066 3442
rect 26066 3390 26068 3442
rect 26012 3388 26068 3390
rect 26012 2882 26068 2884
rect 26012 2830 26014 2882
rect 26014 2830 26066 2882
rect 26066 2830 26068 2882
rect 26012 2828 26068 2830
rect 22764 924 22820 980
rect 23548 1596 23604 1652
rect 23804 1594 23860 1596
rect 23804 1542 23806 1594
rect 23806 1542 23858 1594
rect 23858 1542 23860 1594
rect 23804 1540 23860 1542
rect 23908 1594 23964 1596
rect 23908 1542 23910 1594
rect 23910 1542 23962 1594
rect 23962 1542 23964 1594
rect 23908 1540 23964 1542
rect 24012 1594 24068 1596
rect 24012 1542 24014 1594
rect 24014 1542 24066 1594
rect 24066 1542 24068 1594
rect 24012 1540 24068 1542
rect 24892 1484 24948 1540
rect 24780 1202 24836 1204
rect 24780 1150 24782 1202
rect 24782 1150 24834 1202
rect 24834 1150 24836 1202
rect 24780 1148 24836 1150
rect 24464 810 24520 812
rect 24464 758 24466 810
rect 24466 758 24518 810
rect 24518 758 24520 810
rect 24464 756 24520 758
rect 24568 810 24624 812
rect 24568 758 24570 810
rect 24570 758 24622 810
rect 24622 758 24624 810
rect 24568 756 24624 758
rect 24672 810 24728 812
rect 24672 758 24674 810
rect 24674 758 24726 810
rect 24726 758 24728 810
rect 24672 756 24728 758
rect 25676 1090 25732 1092
rect 25676 1038 25678 1090
rect 25678 1038 25730 1090
rect 25730 1038 25732 1090
rect 25676 1036 25732 1038
rect 25340 700 25396 756
rect 26124 252 26180 308
rect 26572 6076 26628 6132
rect 26908 6690 26964 6692
rect 26908 6638 26910 6690
rect 26910 6638 26962 6690
rect 26962 6638 26964 6690
rect 26908 6636 26964 6638
rect 27244 12124 27300 12180
rect 27244 6636 27300 6692
rect 26684 5180 26740 5236
rect 27132 5740 27188 5796
rect 26460 4844 26516 4900
rect 26572 4284 26628 4340
rect 26796 5068 26852 5124
rect 26572 2940 26628 2996
rect 26684 2044 26740 2100
rect 26572 1596 26628 1652
rect 26908 4396 26964 4452
rect 27580 49196 27636 49252
rect 27468 21308 27524 21364
rect 27468 20412 27524 20468
rect 27468 19516 27524 19572
rect 27468 19068 27524 19124
rect 27468 17948 27524 18004
rect 27468 17276 27524 17332
rect 27468 16380 27524 16436
rect 27468 15932 27524 15988
rect 27468 14812 27524 14868
rect 28140 47964 28196 48020
rect 27916 31052 27972 31108
rect 27804 29484 27860 29540
rect 27580 14364 27636 14420
rect 27692 27804 27748 27860
rect 27916 20076 27972 20132
rect 28028 30156 28084 30212
rect 27804 18396 27860 18452
rect 28028 17836 28084 17892
rect 27916 17612 27972 17668
rect 27468 14140 27524 14196
rect 27804 14364 27860 14420
rect 27468 13244 27524 13300
rect 27468 12796 27524 12852
rect 27580 12124 27636 12180
rect 27692 13804 27748 13860
rect 27580 11900 27636 11956
rect 27468 11004 27524 11060
rect 27468 10108 27524 10164
rect 27468 9660 27524 9716
rect 27580 8764 27636 8820
rect 27468 7868 27524 7924
rect 27468 6972 27524 7028
rect 27468 6524 27524 6580
rect 27580 5628 27636 5684
rect 27468 4732 27524 4788
rect 27356 4172 27412 4228
rect 27468 3836 27524 3892
rect 26908 3442 26964 3444
rect 26908 3390 26910 3442
rect 26910 3390 26962 3442
rect 26962 3390 26964 3442
rect 26908 3388 26964 3390
rect 26908 2882 26964 2884
rect 26908 2830 26910 2882
rect 26910 2830 26962 2882
rect 26962 2830 26964 2882
rect 26908 2828 26964 2830
rect 27468 3388 27524 3444
rect 27692 3276 27748 3332
rect 27916 12236 27972 12292
rect 28028 13916 28084 13972
rect 27916 3500 27972 3556
rect 27804 2828 27860 2884
rect 27580 2492 27636 2548
rect 28252 21420 28308 21476
rect 28252 17052 28308 17108
rect 28364 14364 28420 14420
rect 28252 8876 28308 8932
rect 28140 1484 28196 1540
rect 27132 1202 27188 1204
rect 27132 1150 27134 1202
rect 27134 1150 27186 1202
rect 27186 1150 27188 1202
rect 27132 1148 27188 1150
rect 26796 140 26852 196
rect 27580 140 27636 196
<< metal3 >>
rect 4722 57260 4732 57316
rect 4788 57260 5516 57316
rect 5572 57260 5582 57316
rect 25442 57260 25452 57316
rect 25508 57260 26236 57316
rect 26292 57260 26302 57316
rect 28448 57204 28560 57232
rect 24210 57148 24220 57204
rect 24276 57148 28560 57204
rect 28448 57120 28560 57148
rect 28448 56756 28560 56784
rect 25330 56700 25340 56756
rect 25396 56700 28560 56756
rect 28448 56672 28560 56700
rect 3794 56420 3804 56476
rect 3860 56420 3908 56476
rect 3964 56420 4012 56476
rect 4068 56420 4078 56476
rect 23794 56420 23804 56476
rect 23860 56420 23908 56476
rect 23964 56420 24012 56476
rect 24068 56420 24078 56476
rect 28448 56308 28560 56336
rect 15474 56252 15484 56308
rect 15540 56252 16492 56308
rect 16548 56252 16558 56308
rect 19506 56252 19516 56308
rect 19572 56252 20636 56308
rect 20692 56252 20702 56308
rect 20850 56252 20860 56308
rect 20916 56252 21868 56308
rect 21924 56252 21934 56308
rect 23538 56252 23548 56308
rect 23604 56252 24444 56308
rect 24500 56252 24510 56308
rect 24882 56252 24892 56308
rect 24948 56252 26012 56308
rect 26068 56252 26078 56308
rect 26236 56252 28560 56308
rect 26236 56196 26292 56252
rect 28448 56224 28560 56252
rect 22530 56140 22540 56196
rect 22596 56140 26292 56196
rect 23538 56028 23548 56084
rect 23604 56028 27580 56084
rect 27636 56028 27646 56084
rect 2482 55916 2492 55972
rect 2548 55916 3052 55972
rect 3108 55916 3118 55972
rect 8082 55916 8092 55972
rect 8148 55916 21084 55972
rect 21140 55916 21150 55972
rect 21970 55916 21980 55972
rect 22036 55916 23884 55972
rect 23940 55916 23950 55972
rect 28448 55860 28560 55888
rect 21634 55804 21644 55860
rect 21700 55804 28560 55860
rect 28448 55776 28560 55804
rect 4454 55636 4464 55692
rect 4520 55636 4568 55692
rect 4624 55636 4672 55692
rect 4728 55636 4738 55692
rect 24454 55636 24464 55692
rect 24520 55636 24568 55692
rect 24624 55636 24672 55692
rect 24728 55636 24738 55692
rect 15586 55468 15596 55524
rect 15652 55468 23212 55524
rect 23268 55468 23278 55524
rect 28448 55412 28560 55440
rect 11554 55356 11564 55412
rect 11620 55356 11630 55412
rect 18834 55356 18844 55412
rect 18900 55356 20188 55412
rect 20244 55356 20254 55412
rect 24994 55356 25004 55412
rect 25060 55356 28560 55412
rect 11564 55300 11620 55356
rect 28448 55328 28560 55356
rect 11564 55244 20524 55300
rect 20580 55244 20590 55300
rect 20738 55244 20748 55300
rect 20804 55244 26236 55300
rect 26292 55244 26302 55300
rect 28448 54964 28560 54992
rect 26124 54908 28560 54964
rect 3794 54852 3804 54908
rect 3860 54852 3908 54908
rect 3964 54852 4012 54908
rect 4068 54852 4078 54908
rect 23794 54852 23804 54908
rect 23860 54852 23908 54908
rect 23964 54852 24012 54908
rect 24068 54852 24078 54908
rect 26124 54740 26180 54908
rect 28448 54880 28560 54908
rect 24098 54684 24108 54740
rect 24164 54684 26180 54740
rect 9986 54572 9996 54628
rect 10052 54572 19516 54628
rect 19572 54572 19582 54628
rect 28448 54516 28560 54544
rect 23762 54460 23772 54516
rect 23828 54460 25004 54516
rect 25060 54460 25070 54516
rect 25554 54460 25564 54516
rect 25620 54460 28560 54516
rect 28448 54432 28560 54460
rect 10882 54348 10892 54404
rect 10948 54348 23100 54404
rect 23156 54348 23166 54404
rect 13570 54236 13580 54292
rect 13636 54236 18956 54292
rect 19012 54236 19022 54292
rect 20132 54236 26236 54292
rect 26292 54236 26302 54292
rect 20132 54180 20188 54236
rect 17602 54124 17612 54180
rect 17668 54124 20188 54180
rect 4454 54068 4464 54124
rect 4520 54068 4568 54124
rect 4624 54068 4672 54124
rect 4728 54068 4738 54124
rect 24454 54068 24464 54124
rect 24520 54068 24568 54124
rect 24624 54068 24672 54124
rect 24728 54068 24738 54124
rect 28448 54068 28560 54096
rect 9202 54012 9212 54068
rect 9268 54012 20636 54068
rect 20692 54012 20702 54068
rect 27234 54012 27244 54068
rect 27300 54012 28560 54068
rect 28448 53984 28560 54012
rect 13010 53900 13020 53956
rect 13076 53900 21532 53956
rect 21588 53900 21598 53956
rect 14018 53788 14028 53844
rect 14084 53788 22204 53844
rect 22260 53788 22270 53844
rect 20514 53676 20524 53732
rect 20580 53676 21532 53732
rect 21588 53676 21598 53732
rect 26198 53676 26236 53732
rect 26292 53676 26302 53732
rect 0 53620 112 53648
rect 28448 53620 28560 53648
rect 0 53564 1036 53620
rect 1092 53564 1102 53620
rect 17490 53564 17500 53620
rect 17556 53564 21308 53620
rect 21364 53564 21374 53620
rect 25554 53564 25564 53620
rect 25620 53564 28560 53620
rect 0 53536 112 53564
rect 28448 53536 28560 53564
rect 21074 53452 21084 53508
rect 21140 53452 24668 53508
rect 24724 53452 24734 53508
rect 12898 53340 12908 53396
rect 12964 53340 23492 53396
rect 3794 53284 3804 53340
rect 3860 53284 3908 53340
rect 3964 53284 4012 53340
rect 4068 53284 4078 53340
rect 19618 53228 19628 53284
rect 19684 53228 22652 53284
rect 22708 53228 22718 53284
rect 18274 53116 18284 53172
rect 18340 53116 21756 53172
rect 21812 53116 21822 53172
rect 19618 53004 19628 53060
rect 19684 53004 21868 53060
rect 21924 53004 21934 53060
rect 23436 52948 23492 53340
rect 23794 53284 23804 53340
rect 23860 53284 23908 53340
rect 23964 53284 24012 53340
rect 24068 53284 24078 53340
rect 28448 53172 28560 53200
rect 27010 53116 27020 53172
rect 27076 53116 28560 53172
rect 28448 53088 28560 53116
rect 1362 52892 1372 52948
rect 1428 52892 15148 52948
rect 15204 52892 15214 52948
rect 23436 52892 24220 52948
rect 24276 52892 24286 52948
rect 24444 52892 27356 52948
rect 27412 52892 27422 52948
rect 24444 52836 24500 52892
rect 242 52780 252 52836
rect 308 52780 1596 52836
rect 1652 52780 1662 52836
rect 21298 52780 21308 52836
rect 21364 52780 24500 52836
rect 24658 52780 24668 52836
rect 24724 52780 25228 52836
rect 25284 52780 25294 52836
rect 28448 52724 28560 52752
rect 16706 52668 16716 52724
rect 16772 52668 22204 52724
rect 22260 52668 22270 52724
rect 25442 52668 25452 52724
rect 25508 52668 28560 52724
rect 28448 52640 28560 52668
rect 19954 52556 19964 52612
rect 20020 52556 22764 52612
rect 22820 52556 22830 52612
rect 4454 52500 4464 52556
rect 4520 52500 4568 52556
rect 4624 52500 4672 52556
rect 4728 52500 4738 52556
rect 24454 52500 24464 52556
rect 24520 52500 24568 52556
rect 24624 52500 24672 52556
rect 24728 52500 24738 52556
rect 12786 52332 12796 52388
rect 12852 52332 26236 52388
rect 26292 52332 26302 52388
rect 0 52276 112 52304
rect 28448 52276 28560 52304
rect 0 52220 1036 52276
rect 1092 52220 1102 52276
rect 6514 52220 6524 52276
rect 6580 52220 24668 52276
rect 24724 52220 24734 52276
rect 27234 52220 27244 52276
rect 27300 52220 28560 52276
rect 0 52192 112 52220
rect 28448 52192 28560 52220
rect 16034 52108 16044 52164
rect 16100 52108 26236 52164
rect 26292 52108 26302 52164
rect 23538 51996 23548 52052
rect 23604 51996 24332 52052
rect 24388 51996 24398 52052
rect 28448 51828 28560 51856
rect 25554 51772 25564 51828
rect 25620 51772 28560 51828
rect 3794 51716 3804 51772
rect 3860 51716 3908 51772
rect 3964 51716 4012 51772
rect 4068 51716 4078 51772
rect 23794 51716 23804 51772
rect 23860 51716 23908 51772
rect 23964 51716 24012 51772
rect 24068 51716 24078 51772
rect 28448 51744 28560 51772
rect 28448 51380 28560 51408
rect 6626 51324 6636 51380
rect 6692 51324 22876 51380
rect 22932 51324 22942 51380
rect 27122 51324 27132 51380
rect 27188 51324 28560 51380
rect 28448 51296 28560 51324
rect 17826 51212 17836 51268
rect 17892 51212 26236 51268
rect 26292 51212 26302 51268
rect 12562 51100 12572 51156
rect 12628 51100 23772 51156
rect 23828 51100 23838 51156
rect 0 50932 112 50960
rect 4454 50932 4464 50988
rect 4520 50932 4568 50988
rect 4624 50932 4672 50988
rect 4728 50932 4738 50988
rect 24454 50932 24464 50988
rect 24520 50932 24568 50988
rect 24624 50932 24672 50988
rect 24728 50932 24738 50988
rect 28448 50932 28560 50960
rect 0 50876 1036 50932
rect 1092 50876 1102 50932
rect 27234 50876 27244 50932
rect 27300 50876 28560 50932
rect 0 50848 112 50876
rect 28448 50848 28560 50876
rect 10994 50652 11004 50708
rect 11060 50652 26236 50708
rect 26292 50652 26302 50708
rect 28448 50484 28560 50512
rect 14242 50428 14252 50484
rect 14308 50428 24668 50484
rect 24724 50428 24734 50484
rect 25554 50428 25564 50484
rect 25620 50428 28560 50484
rect 28448 50400 28560 50428
rect 3794 50148 3804 50204
rect 3860 50148 3908 50204
rect 3964 50148 4012 50204
rect 4068 50148 4078 50204
rect 23794 50148 23804 50204
rect 23860 50148 23908 50204
rect 23964 50148 24012 50204
rect 24068 50148 24078 50204
rect 28448 50036 28560 50064
rect 27010 49980 27020 50036
rect 27076 49980 28560 50036
rect 28448 49952 28560 49980
rect 466 49868 476 49924
rect 532 49868 1596 49924
rect 1652 49868 1662 49924
rect 22978 49868 22988 49924
rect 23044 49868 24220 49924
rect 24276 49868 24286 49924
rect 1586 49644 1596 49700
rect 1652 49644 5740 49700
rect 5796 49644 5806 49700
rect 0 49588 112 49616
rect 28448 49588 28560 49616
rect 0 49532 1036 49588
rect 1092 49532 1102 49588
rect 25442 49532 25452 49588
rect 25508 49532 28560 49588
rect 0 49504 112 49532
rect 28448 49504 28560 49532
rect 4454 49364 4464 49420
rect 4520 49364 4568 49420
rect 4624 49364 4672 49420
rect 4728 49364 4738 49420
rect 24454 49364 24464 49420
rect 24520 49364 24568 49420
rect 24624 49364 24672 49420
rect 24728 49364 24738 49420
rect 23762 49196 23772 49252
rect 23828 49196 27580 49252
rect 27636 49196 27646 49252
rect 28448 49140 28560 49168
rect 27234 49084 27244 49140
rect 27300 49084 28560 49140
rect 28448 49056 28560 49084
rect 9986 48972 9996 49028
rect 10052 48972 26236 49028
rect 26292 48972 26302 49028
rect 1586 48860 1596 48916
rect 1652 48860 6076 48916
rect 6132 48860 6142 48916
rect 7410 48860 7420 48916
rect 7476 48860 24668 48916
rect 24724 48860 24734 48916
rect 11666 48748 11676 48804
rect 11732 48748 26348 48804
rect 26404 48748 26414 48804
rect 28448 48692 28560 48720
rect 20290 48636 20300 48692
rect 20356 48636 20860 48692
rect 20916 48636 20926 48692
rect 25554 48636 25564 48692
rect 25620 48636 28560 48692
rect 3794 48580 3804 48636
rect 3860 48580 3908 48636
rect 3964 48580 4012 48636
rect 4068 48580 4078 48636
rect 23794 48580 23804 48636
rect 23860 48580 23908 48636
rect 23964 48580 24012 48636
rect 24068 48580 24078 48636
rect 28448 48608 28560 48636
rect 24882 48524 24892 48580
rect 24948 48524 24958 48580
rect 0 48244 112 48272
rect 24892 48244 24948 48524
rect 28448 48244 28560 48272
rect 0 48188 1036 48244
rect 1092 48188 1102 48244
rect 7074 48188 7084 48244
rect 7140 48188 24948 48244
rect 27122 48188 27132 48244
rect 27188 48188 28560 48244
rect 0 48160 112 48188
rect 28448 48160 28560 48188
rect 15810 48076 15820 48132
rect 15876 48076 26236 48132
rect 26292 48076 26302 48132
rect 17266 47964 17276 48020
rect 17332 47964 24444 48020
rect 24500 47964 24510 48020
rect 24658 47964 24668 48020
rect 24724 47964 25004 48020
rect 25060 47964 25070 48020
rect 25330 47964 25340 48020
rect 25396 47964 28140 48020
rect 28196 47964 28206 48020
rect 4454 47796 4464 47852
rect 4520 47796 4568 47852
rect 4624 47796 4672 47852
rect 4728 47796 4738 47852
rect 24454 47796 24464 47852
rect 24520 47796 24568 47852
rect 24624 47796 24672 47852
rect 24728 47796 24738 47852
rect 28448 47796 28560 47824
rect 27234 47740 27244 47796
rect 27300 47740 28560 47796
rect 28448 47712 28560 47740
rect 28448 47348 28560 47376
rect 25666 47292 25676 47348
rect 25732 47292 28560 47348
rect 28448 47264 28560 47292
rect 3794 47012 3804 47068
rect 3860 47012 3908 47068
rect 3964 47012 4012 47068
rect 4068 47012 4078 47068
rect 23794 47012 23804 47068
rect 23860 47012 23908 47068
rect 23964 47012 24012 47068
rect 24068 47012 24078 47068
rect 0 46900 112 46928
rect 28448 46900 28560 46928
rect 0 46844 1036 46900
rect 1092 46844 1102 46900
rect 19842 46844 19852 46900
rect 19908 46844 24668 46900
rect 24724 46844 24734 46900
rect 27010 46844 27020 46900
rect 27076 46844 28560 46900
rect 0 46816 112 46844
rect 28448 46816 28560 46844
rect 16146 46732 16156 46788
rect 16212 46732 26236 46788
rect 26292 46732 26302 46788
rect 26114 46508 26124 46564
rect 26180 46508 26236 46564
rect 26292 46508 26302 46564
rect 28448 46452 28560 46480
rect 25666 46396 25676 46452
rect 25732 46396 28560 46452
rect 28448 46368 28560 46396
rect 4454 46228 4464 46284
rect 4520 46228 4568 46284
rect 4624 46228 4672 46284
rect 4728 46228 4738 46284
rect 24454 46228 24464 46284
rect 24520 46228 24568 46284
rect 24624 46228 24672 46284
rect 24728 46228 24738 46284
rect 28448 46004 28560 46032
rect 27234 45948 27244 46004
rect 27300 45948 28560 46004
rect 28448 45920 28560 45948
rect 24770 45836 24780 45892
rect 24836 45836 26796 45892
rect 26852 45836 26862 45892
rect 1446 45724 1484 45780
rect 1540 45724 1550 45780
rect 0 45556 112 45584
rect 28448 45556 28560 45584
rect 0 45500 1036 45556
rect 1092 45500 1102 45556
rect 25666 45500 25676 45556
rect 25732 45500 28560 45556
rect 0 45472 112 45500
rect 3794 45444 3804 45500
rect 3860 45444 3908 45500
rect 3964 45444 4012 45500
rect 4068 45444 4078 45500
rect 23794 45444 23804 45500
rect 23860 45444 23908 45500
rect 23964 45444 24012 45500
rect 24068 45444 24078 45500
rect 28448 45472 28560 45500
rect 19842 45388 19852 45444
rect 19908 45388 20076 45444
rect 20132 45388 20142 45444
rect 28448 45108 28560 45136
rect 27122 45052 27132 45108
rect 27188 45052 28560 45108
rect 28448 45024 28560 45052
rect 4454 44660 4464 44716
rect 4520 44660 4568 44716
rect 4624 44660 4672 44716
rect 4728 44660 4738 44716
rect 24454 44660 24464 44716
rect 24520 44660 24568 44716
rect 24624 44660 24672 44716
rect 24728 44660 24738 44716
rect 28448 44660 28560 44688
rect 27234 44604 27244 44660
rect 27300 44604 28560 44660
rect 28448 44576 28560 44604
rect 4834 44268 4844 44324
rect 4900 44268 24668 44324
rect 24724 44268 24734 44324
rect 0 44212 112 44240
rect 28448 44212 28560 44240
rect 0 44156 1036 44212
rect 1092 44156 1102 44212
rect 25666 44156 25676 44212
rect 25732 44156 28560 44212
rect 0 44128 112 44156
rect 28448 44128 28560 44156
rect 3794 43876 3804 43932
rect 3860 43876 3908 43932
rect 3964 43876 4012 43932
rect 4068 43876 4078 43932
rect 23794 43876 23804 43932
rect 23860 43876 23908 43932
rect 23964 43876 24012 43932
rect 24068 43876 24078 43932
rect 28448 43764 28560 43792
rect 1586 43708 1596 43764
rect 1652 43708 3612 43764
rect 3668 43708 3678 43764
rect 27010 43708 27020 43764
rect 27076 43708 28560 43764
rect 28448 43680 28560 43708
rect 1474 43596 1484 43652
rect 1540 43596 3388 43652
rect 3490 43596 3500 43652
rect 3556 43596 11340 43652
rect 11396 43596 11406 43652
rect 1558 43372 1596 43428
rect 1652 43372 1662 43428
rect 0 42868 112 42896
rect 3332 42868 3388 43596
rect 28448 43316 28560 43344
rect 25666 43260 25676 43316
rect 25732 43260 28560 43316
rect 28448 43232 28560 43260
rect 4454 43092 4464 43148
rect 4520 43092 4568 43148
rect 4624 43092 4672 43148
rect 4728 43092 4738 43148
rect 24454 43092 24464 43148
rect 24520 43092 24568 43148
rect 24624 43092 24672 43148
rect 24728 43092 24738 43148
rect 12226 42924 12236 42980
rect 12292 42924 24220 42980
rect 24276 42924 24286 42980
rect 28448 42868 28560 42896
rect 0 42812 924 42868
rect 980 42812 990 42868
rect 3332 42812 17948 42868
rect 18004 42812 18014 42868
rect 27234 42812 27244 42868
rect 27300 42812 28560 42868
rect 0 42784 112 42812
rect 28448 42784 28560 42812
rect 13010 42700 13020 42756
rect 13076 42700 24668 42756
rect 24724 42700 24734 42756
rect 1810 42476 1820 42532
rect 1876 42476 14476 42532
rect 14532 42476 14542 42532
rect 28448 42420 28560 42448
rect 25666 42364 25676 42420
rect 25732 42364 28560 42420
rect 3794 42308 3804 42364
rect 3860 42308 3908 42364
rect 3964 42308 4012 42364
rect 4068 42308 4078 42364
rect 23794 42308 23804 42364
rect 23860 42308 23908 42364
rect 23964 42308 24012 42364
rect 24068 42308 24078 42364
rect 28448 42336 28560 42364
rect 2146 42028 2156 42084
rect 2212 42028 11004 42084
rect 11060 42028 11070 42084
rect 28448 41972 28560 42000
rect 3332 41916 24892 41972
rect 24948 41916 24958 41972
rect 27122 41916 27132 41972
rect 27188 41916 28560 41972
rect 3332 41860 3388 41916
rect 28448 41888 28560 41916
rect 578 41804 588 41860
rect 644 41804 1596 41860
rect 1652 41804 1662 41860
rect 2594 41804 2604 41860
rect 2660 41804 3388 41860
rect 4162 41804 4172 41860
rect 4228 41804 10892 41860
rect 10948 41804 10958 41860
rect 20132 41804 26236 41860
rect 26292 41804 26302 41860
rect 20132 41748 20188 41804
rect 12002 41692 12012 41748
rect 12068 41692 20188 41748
rect 0 41524 112 41552
rect 4454 41524 4464 41580
rect 4520 41524 4568 41580
rect 4624 41524 4672 41580
rect 4728 41524 4738 41580
rect 24454 41524 24464 41580
rect 24520 41524 24568 41580
rect 24624 41524 24672 41580
rect 24728 41524 24738 41580
rect 28448 41524 28560 41552
rect 0 41468 1148 41524
rect 1204 41468 1214 41524
rect 27234 41468 27244 41524
rect 27300 41468 28560 41524
rect 0 41440 112 41468
rect 28448 41440 28560 41468
rect 2482 41356 2492 41412
rect 2548 41356 26348 41412
rect 26404 41356 26414 41412
rect 2034 41244 2044 41300
rect 2100 41244 2380 41300
rect 2436 41244 4284 41300
rect 4340 41244 4350 41300
rect 8978 41132 8988 41188
rect 9044 41132 26236 41188
rect 26292 41132 26302 41188
rect 28448 41076 28560 41104
rect 690 41020 700 41076
rect 756 41020 1484 41076
rect 1540 41020 1550 41076
rect 3490 41020 3500 41076
rect 3556 41020 10556 41076
rect 10612 41020 10622 41076
rect 25666 41020 25676 41076
rect 25732 41020 28560 41076
rect 28448 40992 28560 41020
rect 3794 40740 3804 40796
rect 3860 40740 3908 40796
rect 3964 40740 4012 40796
rect 4068 40740 4078 40796
rect 23794 40740 23804 40796
rect 23860 40740 23908 40796
rect 23964 40740 24012 40796
rect 24068 40740 24078 40796
rect 28448 40628 28560 40656
rect 6626 40572 6636 40628
rect 6692 40572 7644 40628
rect 7700 40572 7710 40628
rect 8642 40572 8652 40628
rect 8708 40572 9324 40628
rect 9380 40572 9390 40628
rect 15092 40572 24892 40628
rect 24948 40572 24958 40628
rect 27010 40572 27020 40628
rect 27076 40572 28560 40628
rect 15092 40516 15148 40572
rect 28448 40544 28560 40572
rect 6962 40460 6972 40516
rect 7028 40460 15148 40516
rect 19282 40460 19292 40516
rect 19348 40460 24668 40516
rect 24724 40460 24734 40516
rect 4274 40348 4284 40404
rect 4340 40348 8764 40404
rect 8820 40348 8830 40404
rect 9426 40348 9436 40404
rect 9492 40348 10108 40404
rect 10164 40348 10174 40404
rect 15362 40348 15372 40404
rect 15428 40348 17724 40404
rect 17780 40348 17790 40404
rect 1698 40236 1708 40292
rect 1764 40236 2268 40292
rect 2324 40236 3052 40292
rect 3108 40236 3118 40292
rect 0 40180 112 40208
rect 28448 40180 28560 40208
rect 0 40124 924 40180
rect 980 40124 990 40180
rect 25666 40124 25676 40180
rect 25732 40124 28560 40180
rect 0 40096 112 40124
rect 28448 40096 28560 40124
rect 802 40012 812 40068
rect 868 40012 1932 40068
rect 1988 40012 1998 40068
rect 4454 39956 4464 40012
rect 4520 39956 4568 40012
rect 4624 39956 4672 40012
rect 4728 39956 4738 40012
rect 24454 39956 24464 40012
rect 24520 39956 24568 40012
rect 24624 39956 24672 40012
rect 24728 39956 24738 40012
rect 5842 39900 5852 39956
rect 5908 39900 6188 39956
rect 6244 39900 6254 39956
rect 7522 39900 7532 39956
rect 7588 39900 15148 39956
rect 6188 39844 6244 39900
rect 15092 39844 15148 39900
rect 6188 39788 9884 39844
rect 9940 39788 9950 39844
rect 11778 39788 11788 39844
rect 11844 39788 12908 39844
rect 12964 39788 12974 39844
rect 15092 39788 18844 39844
rect 18900 39788 18910 39844
rect 28448 39732 28560 39760
rect 5058 39676 5068 39732
rect 5124 39676 8092 39732
rect 8148 39676 8158 39732
rect 27234 39676 27244 39732
rect 27300 39676 28560 39732
rect 28448 39648 28560 39676
rect 2034 39564 2044 39620
rect 2100 39564 2940 39620
rect 2996 39564 3006 39620
rect 8194 39564 8204 39620
rect 8260 39564 9772 39620
rect 9828 39564 9838 39620
rect 10994 39564 11004 39620
rect 11060 39564 11788 39620
rect 11844 39564 11854 39620
rect 20132 39564 26236 39620
rect 26292 39564 26302 39620
rect 20132 39508 20188 39564
rect 6290 39452 6300 39508
rect 6356 39452 6636 39508
rect 6692 39452 6702 39508
rect 11218 39452 11228 39508
rect 11284 39452 20188 39508
rect 28448 39284 28560 39312
rect 25666 39228 25676 39284
rect 25732 39228 28560 39284
rect 3794 39172 3804 39228
rect 3860 39172 3908 39228
rect 3964 39172 4012 39228
rect 4068 39172 4078 39228
rect 23794 39172 23804 39228
rect 23860 39172 23908 39228
rect 23964 39172 24012 39228
rect 24068 39172 24078 39228
rect 28448 39200 28560 39228
rect 6738 39004 6748 39060
rect 6804 39004 7196 39060
rect 7252 39004 7262 39060
rect 2930 38892 2940 38948
rect 2996 38892 5964 38948
rect 6020 38892 6030 38948
rect 0 38836 112 38864
rect 28448 38836 28560 38864
rect 0 38780 1036 38836
rect 1092 38780 1102 38836
rect 2706 38780 2716 38836
rect 2772 38780 3612 38836
rect 3668 38780 5516 38836
rect 5572 38780 5582 38836
rect 12674 38780 12684 38836
rect 12740 38780 15260 38836
rect 15316 38780 16716 38836
rect 16772 38780 16782 38836
rect 27122 38780 27132 38836
rect 27188 38780 28560 38836
rect 0 38752 112 38780
rect 28448 38752 28560 38780
rect 4274 38668 4284 38724
rect 4340 38668 8988 38724
rect 9044 38668 9054 38724
rect 13346 38668 13356 38724
rect 13412 38668 26348 38724
rect 26404 38668 26414 38724
rect 3826 38556 3836 38612
rect 3892 38556 17836 38612
rect 17892 38556 17902 38612
rect 20300 38556 25452 38612
rect 25508 38556 25518 38612
rect 20300 38500 20356 38556
rect 7746 38444 7756 38500
rect 7812 38444 20356 38500
rect 4454 38388 4464 38444
rect 4520 38388 4568 38444
rect 4624 38388 4672 38444
rect 4728 38388 4738 38444
rect 24454 38388 24464 38444
rect 24520 38388 24568 38444
rect 24624 38388 24672 38444
rect 24728 38388 24738 38444
rect 28448 38388 28560 38416
rect 12786 38332 12796 38388
rect 12852 38332 13132 38388
rect 13188 38332 13198 38388
rect 27234 38332 27244 38388
rect 27300 38332 28560 38388
rect 28448 38304 28560 38332
rect 1474 38220 1484 38276
rect 1540 38220 18172 38276
rect 18228 38220 18238 38276
rect 11778 38108 11788 38164
rect 11844 38108 13244 38164
rect 13300 38108 13310 38164
rect 9398 37996 9436 38052
rect 9492 37996 10556 38052
rect 10612 37996 10622 38052
rect 11106 37996 11116 38052
rect 11172 37996 11900 38052
rect 11956 37996 11966 38052
rect 12114 37996 12124 38052
rect 12180 37996 13132 38052
rect 13188 37996 13198 38052
rect 13458 37996 13468 38052
rect 13524 37996 17500 38052
rect 17556 37996 17566 38052
rect 21858 37996 21868 38052
rect 21924 37996 26236 38052
rect 26292 37996 26302 38052
rect 28448 37940 28560 37968
rect 1586 37884 1596 37940
rect 1652 37884 13804 37940
rect 13860 37884 13870 37940
rect 15092 37884 19740 37940
rect 19796 37884 19806 37940
rect 25666 37884 25676 37940
rect 25732 37884 28560 37940
rect 3266 37772 3276 37828
rect 3332 37772 7420 37828
rect 7476 37772 7486 37828
rect 9986 37772 9996 37828
rect 10052 37772 12348 37828
rect 12404 37772 12414 37828
rect 3794 37604 3804 37660
rect 3860 37604 3908 37660
rect 3964 37604 4012 37660
rect 4068 37604 4078 37660
rect 15092 37604 15148 37884
rect 28448 37856 28560 37884
rect 23794 37604 23804 37660
rect 23860 37604 23908 37660
rect 23964 37604 24012 37660
rect 24068 37604 24078 37660
rect 5170 37548 5180 37604
rect 5236 37548 5516 37604
rect 5572 37548 5582 37604
rect 13234 37548 13244 37604
rect 13300 37548 15148 37604
rect 0 37492 112 37520
rect 28448 37492 28560 37520
rect 0 37436 1036 37492
rect 1092 37436 1102 37492
rect 4834 37436 4844 37492
rect 4900 37436 8316 37492
rect 8372 37436 15596 37492
rect 15652 37436 17276 37492
rect 17332 37436 17342 37492
rect 27010 37436 27020 37492
rect 27076 37436 28560 37492
rect 0 37408 112 37436
rect 28448 37408 28560 37436
rect 1036 37324 1484 37380
rect 1540 37324 1550 37380
rect 2482 37324 2492 37380
rect 2548 37324 11788 37380
rect 11844 37324 11854 37380
rect 1036 37268 1092 37324
rect 1026 37212 1036 37268
rect 1092 37212 1102 37268
rect 6972 37212 12460 37268
rect 12516 37212 13356 37268
rect 13412 37212 13422 37268
rect 6972 37156 7028 37212
rect 1586 37100 1596 37156
rect 1652 37100 6524 37156
rect 6580 37100 6590 37156
rect 6962 37100 6972 37156
rect 7028 37100 7038 37156
rect 7522 37100 7532 37156
rect 7588 37100 8204 37156
rect 8260 37100 13580 37156
rect 13636 37100 13646 37156
rect 25778 37100 25788 37156
rect 25844 37100 26236 37156
rect 26292 37100 26302 37156
rect 28448 37044 28560 37072
rect 3378 36988 3388 37044
rect 3444 36988 3948 37044
rect 4004 36988 9996 37044
rect 10052 36988 10062 37044
rect 25442 36988 25452 37044
rect 25508 36988 28560 37044
rect 28448 36960 28560 36988
rect 2818 36876 2828 36932
rect 2884 36876 3612 36932
rect 3668 36876 3678 36932
rect 4454 36820 4464 36876
rect 4520 36820 4568 36876
rect 4624 36820 4672 36876
rect 4728 36820 4738 36876
rect 24454 36820 24464 36876
rect 24520 36820 24568 36876
rect 24624 36820 24672 36876
rect 24728 36820 24738 36876
rect 802 36764 812 36820
rect 868 36764 1260 36820
rect 1316 36764 2716 36820
rect 2772 36764 2782 36820
rect 2930 36764 2940 36820
rect 2996 36764 3500 36820
rect 3556 36764 3566 36820
rect 1698 36652 1708 36708
rect 1764 36652 2828 36708
rect 2884 36652 2894 36708
rect 3602 36652 3612 36708
rect 3668 36652 5068 36708
rect 5124 36652 5516 36708
rect 5572 36652 5582 36708
rect 28448 36596 28560 36624
rect 2706 36540 2716 36596
rect 2772 36540 3052 36596
rect 3108 36540 3118 36596
rect 27234 36540 27244 36596
rect 27300 36540 28560 36596
rect 28448 36512 28560 36540
rect 14354 36428 14364 36484
rect 14420 36428 14812 36484
rect 14868 36428 14878 36484
rect 17154 36428 17164 36484
rect 17220 36428 24668 36484
rect 24724 36428 24734 36484
rect 1922 36316 1932 36372
rect 1988 36316 3276 36372
rect 3332 36316 10108 36372
rect 10164 36316 10174 36372
rect 17042 36316 17052 36372
rect 17108 36316 18284 36372
rect 18340 36316 18350 36372
rect 1698 36204 1708 36260
rect 1764 36204 3388 36260
rect 3444 36204 3454 36260
rect 5058 36204 5068 36260
rect 5124 36204 5516 36260
rect 5572 36204 5582 36260
rect 13346 36204 13356 36260
rect 13412 36204 14028 36260
rect 14084 36204 14094 36260
rect 0 36148 112 36176
rect 28448 36148 28560 36176
rect 0 36092 924 36148
rect 980 36092 990 36148
rect 9174 36092 9212 36148
rect 9268 36092 9278 36148
rect 25666 36092 25676 36148
rect 25732 36092 28560 36148
rect 0 36064 112 36092
rect 3794 36036 3804 36092
rect 3860 36036 3908 36092
rect 3964 36036 4012 36092
rect 4068 36036 4078 36092
rect 23794 36036 23804 36092
rect 23860 36036 23908 36092
rect 23964 36036 24012 36092
rect 24068 36036 24078 36092
rect 28448 36064 28560 36092
rect 10658 35980 10668 36036
rect 10724 35980 11228 36036
rect 11284 35980 11294 36036
rect 3378 35868 3388 35924
rect 3444 35868 6748 35924
rect 6804 35868 11004 35924
rect 11060 35868 11070 35924
rect 5842 35756 5852 35812
rect 5908 35756 10556 35812
rect 10612 35756 17052 35812
rect 17108 35756 17118 35812
rect 28448 35700 28560 35728
rect 8082 35644 8092 35700
rect 8148 35644 8652 35700
rect 8708 35644 8718 35700
rect 8978 35644 8988 35700
rect 9044 35644 9324 35700
rect 9380 35644 9390 35700
rect 9650 35644 9660 35700
rect 9716 35644 9884 35700
rect 9940 35644 9950 35700
rect 27122 35644 27132 35700
rect 27188 35644 28560 35700
rect 28448 35616 28560 35644
rect 1586 35532 1596 35588
rect 1652 35532 3388 35588
rect 8306 35532 8316 35588
rect 8372 35532 8876 35588
rect 8932 35532 8942 35588
rect 9174 35532 9212 35588
rect 9268 35532 9278 35588
rect 16930 35532 16940 35588
rect 16996 35532 25340 35588
rect 25396 35532 25406 35588
rect 3332 35476 3388 35532
rect 3332 35420 8652 35476
rect 8708 35420 8718 35476
rect 9090 35420 9100 35476
rect 9156 35420 9436 35476
rect 9492 35420 9502 35476
rect 20962 35420 20972 35476
rect 21028 35420 25340 35476
rect 25396 35420 25406 35476
rect 3154 35308 3164 35364
rect 3220 35308 3388 35364
rect 3444 35308 3454 35364
rect 5730 35308 5740 35364
rect 5796 35308 6300 35364
rect 6356 35308 6366 35364
rect 7410 35308 7420 35364
rect 7476 35308 8204 35364
rect 8260 35308 8270 35364
rect 4454 35252 4464 35308
rect 4520 35252 4568 35308
rect 4624 35252 4672 35308
rect 4728 35252 4738 35308
rect 24454 35252 24464 35308
rect 24520 35252 24568 35308
rect 24624 35252 24672 35308
rect 24728 35252 24738 35308
rect 28448 35252 28560 35280
rect 2594 35196 2604 35252
rect 2660 35196 3500 35252
rect 3556 35196 3566 35252
rect 27234 35196 27244 35252
rect 27300 35196 28560 35252
rect 28448 35168 28560 35196
rect 4274 35084 4284 35140
rect 4340 35084 4956 35140
rect 5012 35084 5022 35140
rect 12002 35084 12012 35140
rect 12068 35084 13244 35140
rect 13300 35084 13310 35140
rect 15922 35084 15932 35140
rect 15988 35084 16828 35140
rect 16884 35084 16894 35140
rect 17938 35084 17948 35140
rect 18004 35084 19852 35140
rect 19908 35084 19918 35140
rect 6626 34972 6636 35028
rect 6692 34972 26124 35028
rect 26180 34972 26190 35028
rect 4274 34860 4284 34916
rect 4340 34860 5404 34916
rect 5460 34860 5470 34916
rect 25218 34860 25228 34916
rect 25284 34860 26236 34916
rect 26292 34860 26302 34916
rect 0 34804 112 34832
rect 28448 34804 28560 34832
rect 0 34748 1372 34804
rect 1428 34748 1438 34804
rect 5058 34748 5068 34804
rect 5124 34748 6300 34804
rect 6356 34748 6366 34804
rect 25666 34748 25676 34804
rect 25732 34748 28560 34804
rect 0 34720 112 34748
rect 28448 34720 28560 34748
rect 12114 34636 12124 34692
rect 12180 34636 12908 34692
rect 12964 34636 12974 34692
rect 3794 34468 3804 34524
rect 3860 34468 3908 34524
rect 3964 34468 4012 34524
rect 4068 34468 4078 34524
rect 23794 34468 23804 34524
rect 23860 34468 23908 34524
rect 23964 34468 24012 34524
rect 24068 34468 24078 34524
rect 5842 34412 5852 34468
rect 5908 34412 7084 34468
rect 7140 34412 15148 34468
rect 15204 34412 15214 34468
rect 28448 34356 28560 34384
rect 6626 34300 6636 34356
rect 6692 34300 26348 34356
rect 26404 34300 26414 34356
rect 27010 34300 27020 34356
rect 27076 34300 28560 34356
rect 28448 34272 28560 34300
rect 4050 34188 4060 34244
rect 4116 34188 12572 34244
rect 12628 34188 14028 34244
rect 14084 34188 14094 34244
rect 15698 34188 15708 34244
rect 15764 34188 24892 34244
rect 24948 34188 24958 34244
rect 3490 34076 3500 34132
rect 3556 34076 5180 34132
rect 5236 34076 5246 34132
rect 16594 34076 16604 34132
rect 16660 34076 18508 34132
rect 18564 34076 18574 34132
rect 12450 33964 12460 34020
rect 12516 33964 26236 34020
rect 26292 33964 26302 34020
rect 28448 33908 28560 33936
rect 3826 33852 3836 33908
rect 3892 33852 24780 33908
rect 24836 33852 24846 33908
rect 25666 33852 25676 33908
rect 25732 33852 28560 33908
rect 28448 33824 28560 33852
rect 8166 33740 8204 33796
rect 8260 33740 8270 33796
rect 17378 33740 17388 33796
rect 17444 33740 22204 33796
rect 22260 33740 22270 33796
rect 4454 33684 4464 33740
rect 4520 33684 4568 33740
rect 4624 33684 4672 33740
rect 4728 33684 4738 33740
rect 24454 33684 24464 33740
rect 24520 33684 24568 33740
rect 24624 33684 24672 33740
rect 24728 33684 24738 33740
rect 5170 33628 5180 33684
rect 5236 33628 8092 33684
rect 8148 33628 9548 33684
rect 9604 33628 9614 33684
rect 16930 33628 16940 33684
rect 16996 33628 17612 33684
rect 17668 33628 17678 33684
rect 2146 33516 2156 33572
rect 2212 33516 3276 33572
rect 3332 33516 3342 33572
rect 6066 33516 6076 33572
rect 6132 33516 6524 33572
rect 6580 33516 6590 33572
rect 8194 33516 8204 33572
rect 8260 33516 25788 33572
rect 25844 33516 25854 33572
rect 0 33460 112 33488
rect 6524 33460 6580 33516
rect 28448 33460 28560 33488
rect 0 33404 924 33460
rect 980 33404 990 33460
rect 1586 33404 1596 33460
rect 1652 33404 2716 33460
rect 2772 33404 2782 33460
rect 6524 33404 9884 33460
rect 9940 33404 14588 33460
rect 14644 33404 14654 33460
rect 15138 33404 15148 33460
rect 15204 33404 16044 33460
rect 16100 33404 16110 33460
rect 27234 33404 27244 33460
rect 27300 33404 28560 33460
rect 0 33376 112 33404
rect 14588 33348 14644 33404
rect 28448 33376 28560 33404
rect 7186 33292 7196 33348
rect 7252 33292 7262 33348
rect 14588 33292 15596 33348
rect 15652 33292 15662 33348
rect 24882 33292 24892 33348
rect 24948 33292 26684 33348
rect 26740 33292 26750 33348
rect 7196 33124 7252 33292
rect 7196 33068 7420 33124
rect 7476 33068 7486 33124
rect 19394 33068 19404 33124
rect 19460 33068 19516 33124
rect 19572 33068 19582 33124
rect 28448 33012 28560 33040
rect 690 32956 700 33012
rect 756 32956 1596 33012
rect 1652 32956 1662 33012
rect 5170 32956 5180 33012
rect 5236 32956 5628 33012
rect 5684 32956 9100 33012
rect 9156 32956 9166 33012
rect 12898 32956 12908 33012
rect 12964 32956 13356 33012
rect 13412 32956 13422 33012
rect 17378 32956 17388 33012
rect 17444 32956 23660 33012
rect 23716 32956 23726 33012
rect 25666 32956 25676 33012
rect 25732 32956 28560 33012
rect 3794 32900 3804 32956
rect 3860 32900 3908 32956
rect 3964 32900 4012 32956
rect 4068 32900 4078 32956
rect 23794 32900 23804 32956
rect 23860 32900 23908 32956
rect 23964 32900 24012 32956
rect 24068 32900 24078 32956
rect 28448 32928 28560 32956
rect 1698 32844 1708 32900
rect 1764 32844 2044 32900
rect 2100 32844 2110 32900
rect 13122 32844 13132 32900
rect 13188 32844 19908 32900
rect 25330 32844 25340 32900
rect 25396 32844 26460 32900
rect 26516 32844 26526 32900
rect 19852 32788 19908 32844
rect 8754 32732 8764 32788
rect 8820 32732 9548 32788
rect 9604 32732 9614 32788
rect 18274 32732 18284 32788
rect 18340 32732 18956 32788
rect 19012 32732 19022 32788
rect 19852 32732 24892 32788
rect 24948 32732 24958 32788
rect 25554 32732 25564 32788
rect 25620 32732 26572 32788
rect 26628 32732 26638 32788
rect 1250 32620 1260 32676
rect 1316 32620 1708 32676
rect 1764 32620 1774 32676
rect 4386 32620 4396 32676
rect 4452 32620 26236 32676
rect 26292 32620 26302 32676
rect 28448 32564 28560 32592
rect 6738 32508 6748 32564
rect 6804 32508 7196 32564
rect 7252 32508 7262 32564
rect 7410 32508 7420 32564
rect 7476 32508 8428 32564
rect 8484 32508 8494 32564
rect 9426 32508 9436 32564
rect 9492 32508 10556 32564
rect 10612 32508 11788 32564
rect 11844 32508 11854 32564
rect 13794 32508 13804 32564
rect 13860 32508 14252 32564
rect 14308 32508 14318 32564
rect 17266 32508 17276 32564
rect 17332 32508 18620 32564
rect 18676 32508 18686 32564
rect 19366 32508 19404 32564
rect 19460 32508 19470 32564
rect 27122 32508 27132 32564
rect 27188 32508 28560 32564
rect 28448 32480 28560 32508
rect 8194 32396 8204 32452
rect 8260 32396 9212 32452
rect 9268 32396 9278 32452
rect 19170 32396 19180 32452
rect 19236 32396 19852 32452
rect 19908 32396 19918 32452
rect 7074 32284 7084 32340
rect 7140 32284 7756 32340
rect 7812 32284 7822 32340
rect 12114 32284 12124 32340
rect 12180 32284 12348 32340
rect 12404 32284 12414 32340
rect 13906 32172 13916 32228
rect 13972 32172 14812 32228
rect 14868 32172 14878 32228
rect 0 32116 112 32144
rect 4454 32116 4464 32172
rect 4520 32116 4568 32172
rect 4624 32116 4672 32172
rect 4728 32116 4738 32172
rect 24454 32116 24464 32172
rect 24520 32116 24568 32172
rect 24624 32116 24672 32172
rect 24728 32116 24738 32172
rect 28448 32116 28560 32144
rect 0 32060 1036 32116
rect 1092 32060 1102 32116
rect 2258 32060 2268 32116
rect 2324 32060 2828 32116
rect 2884 32060 2894 32116
rect 17602 32060 17612 32116
rect 17668 32060 18172 32116
rect 18228 32060 18238 32116
rect 27234 32060 27244 32116
rect 27300 32060 28560 32116
rect 0 32032 112 32060
rect 28448 32032 28560 32060
rect 12786 31948 12796 32004
rect 12852 31948 13356 32004
rect 13412 31948 13422 32004
rect 2818 31836 2828 31892
rect 2884 31836 3724 31892
rect 3780 31836 3790 31892
rect 8642 31836 8652 31892
rect 8708 31836 13692 31892
rect 13748 31836 14588 31892
rect 14644 31836 14654 31892
rect 15026 31836 15036 31892
rect 15092 31836 15372 31892
rect 15428 31836 15438 31892
rect 16818 31836 16828 31892
rect 16884 31836 18172 31892
rect 18228 31836 18238 31892
rect 4050 31724 4060 31780
rect 4116 31724 4732 31780
rect 4788 31724 4798 31780
rect 7298 31724 7308 31780
rect 7364 31724 8876 31780
rect 8932 31724 8942 31780
rect 14914 31724 14924 31780
rect 14980 31724 16716 31780
rect 16772 31724 19180 31780
rect 19236 31724 19246 31780
rect 28448 31668 28560 31696
rect 1250 31612 1260 31668
rect 1316 31612 1708 31668
rect 1764 31612 4844 31668
rect 4900 31612 4910 31668
rect 16818 31612 16828 31668
rect 16884 31612 17164 31668
rect 17220 31612 17230 31668
rect 25666 31612 25676 31668
rect 25732 31612 28560 31668
rect 28448 31584 28560 31612
rect 3574 31500 3612 31556
rect 3668 31500 3678 31556
rect 5058 31500 5068 31556
rect 5124 31500 6524 31556
rect 6580 31500 7644 31556
rect 7700 31500 7710 31556
rect 15026 31500 15036 31556
rect 15092 31500 15148 31556
rect 15204 31500 15214 31556
rect 11890 31388 11900 31444
rect 11956 31388 16156 31444
rect 16212 31388 16222 31444
rect 3794 31332 3804 31388
rect 3860 31332 3908 31388
rect 3964 31332 4012 31388
rect 4068 31332 4078 31388
rect 23794 31332 23804 31388
rect 23860 31332 23908 31388
rect 23964 31332 24012 31388
rect 24068 31332 24078 31388
rect 28448 31220 28560 31248
rect 3332 31164 4844 31220
rect 4900 31164 4910 31220
rect 15810 31164 15820 31220
rect 15876 31164 17052 31220
rect 17108 31164 17118 31220
rect 27010 31164 27020 31220
rect 27076 31164 28560 31220
rect 3332 31108 3388 31164
rect 28448 31136 28560 31164
rect 2370 31052 2380 31108
rect 2436 31052 3388 31108
rect 4386 31052 4396 31108
rect 4452 31052 12012 31108
rect 12068 31052 27916 31108
rect 27972 31052 27982 31108
rect 466 30940 476 30996
rect 532 30940 1260 30996
rect 1316 30940 1326 30996
rect 2706 30940 2716 30996
rect 2772 30940 3500 30996
rect 3556 30940 4620 30996
rect 4676 30940 4686 30996
rect 7634 30940 7644 30996
rect 7700 30940 14252 30996
rect 14308 30940 15036 30996
rect 15092 30940 15102 30996
rect 1810 30828 1820 30884
rect 1876 30828 4396 30884
rect 4452 30828 4462 30884
rect 6290 30828 6300 30884
rect 6356 30828 6636 30884
rect 6692 30828 6702 30884
rect 0 30772 112 30800
rect 28448 30772 28560 30800
rect 0 30716 3500 30772
rect 3556 30716 3566 30772
rect 7074 30716 7084 30772
rect 7140 30716 7308 30772
rect 7364 30716 7644 30772
rect 7700 30716 7710 30772
rect 17266 30716 17276 30772
rect 17332 30716 17948 30772
rect 18004 30716 18014 30772
rect 19852 30716 24780 30772
rect 24836 30716 24846 30772
rect 25442 30716 25452 30772
rect 25508 30716 28560 30772
rect 0 30688 112 30716
rect 19852 30660 19908 30716
rect 28448 30688 28560 30716
rect 12674 30604 12684 30660
rect 12740 30604 19908 30660
rect 4454 30548 4464 30604
rect 4520 30548 4568 30604
rect 4624 30548 4672 30604
rect 4728 30548 4738 30604
rect 24454 30548 24464 30604
rect 24520 30548 24568 30604
rect 24624 30548 24672 30604
rect 24728 30548 24738 30604
rect 11890 30492 11900 30548
rect 11956 30492 12460 30548
rect 12516 30492 12526 30548
rect 3154 30380 3164 30436
rect 3220 30380 3388 30436
rect 3444 30380 3454 30436
rect 10770 30380 10780 30436
rect 10836 30380 26124 30436
rect 26180 30380 26190 30436
rect 28448 30324 28560 30352
rect 2818 30268 2828 30324
rect 2884 30268 3220 30324
rect 27234 30268 27244 30324
rect 27300 30268 28560 30324
rect 3164 30212 3220 30268
rect 28448 30240 28560 30268
rect 3154 30156 3164 30212
rect 3220 30156 3230 30212
rect 5842 30156 5852 30212
rect 5908 30156 7308 30212
rect 7364 30156 7374 30212
rect 8306 30156 8316 30212
rect 8372 30156 10220 30212
rect 10276 30156 28028 30212
rect 28084 30156 28094 30212
rect 802 30044 812 30100
rect 868 30044 1260 30100
rect 1316 30044 1326 30100
rect 2818 30044 2828 30100
rect 2884 30044 3948 30100
rect 4004 30044 4014 30100
rect 6626 30044 6636 30100
rect 6692 30044 7084 30100
rect 7140 30044 15148 30100
rect 19730 30044 19740 30100
rect 19796 30044 24892 30100
rect 24948 30044 24958 30100
rect 15092 29988 15148 30044
rect 2706 29932 2716 29988
rect 2772 29932 9268 29988
rect 15092 29932 16716 29988
rect 16772 29932 25452 29988
rect 25508 29932 25518 29988
rect 9212 29876 9268 29932
rect 28448 29876 28560 29904
rect 9212 29820 21868 29876
rect 21924 29820 21934 29876
rect 27010 29820 27020 29876
rect 27076 29820 28560 29876
rect 3794 29764 3804 29820
rect 3860 29764 3908 29820
rect 3964 29764 4012 29820
rect 4068 29764 4078 29820
rect 23794 29764 23804 29820
rect 23860 29764 23908 29820
rect 23964 29764 24012 29820
rect 24068 29764 24078 29820
rect 28448 29792 28560 29820
rect 11330 29596 11340 29652
rect 11396 29596 11676 29652
rect 11732 29596 11742 29652
rect 17602 29596 17612 29652
rect 17668 29596 18508 29652
rect 18564 29596 18574 29652
rect 3602 29484 3612 29540
rect 3668 29484 3724 29540
rect 3780 29484 3790 29540
rect 5058 29484 5068 29540
rect 5124 29484 9212 29540
rect 9268 29484 27804 29540
rect 27860 29484 27870 29540
rect 0 29428 112 29456
rect 28448 29428 28560 29456
rect 0 29372 1036 29428
rect 1092 29372 1102 29428
rect 9762 29372 9772 29428
rect 9828 29372 10220 29428
rect 10276 29372 10286 29428
rect 11330 29372 11340 29428
rect 11396 29372 11788 29428
rect 11844 29372 12236 29428
rect 12292 29372 12302 29428
rect 15138 29372 15148 29428
rect 15204 29372 15820 29428
rect 15876 29372 16828 29428
rect 16884 29372 16894 29428
rect 27122 29372 27132 29428
rect 27188 29372 28560 29428
rect 0 29344 112 29372
rect 28448 29344 28560 29372
rect 578 29260 588 29316
rect 644 29260 1708 29316
rect 1764 29260 1774 29316
rect 2594 29260 2604 29316
rect 2660 29260 8876 29316
rect 8932 29260 8942 29316
rect 9426 29260 9436 29316
rect 9492 29260 26236 29316
rect 26292 29260 26302 29316
rect 1708 29204 1764 29260
rect 1708 29148 8428 29204
rect 8484 29148 8494 29204
rect 14354 29148 14364 29204
rect 14420 29148 17724 29204
rect 17780 29148 17790 29204
rect 578 29036 588 29092
rect 644 29036 2604 29092
rect 2660 29036 2670 29092
rect 5058 29036 5068 29092
rect 5124 29036 5404 29092
rect 5460 29036 5470 29092
rect 16818 29036 16828 29092
rect 16884 29036 24332 29092
rect 24388 29036 24398 29092
rect 4454 28980 4464 29036
rect 4520 28980 4568 29036
rect 4624 28980 4672 29036
rect 4728 28980 4738 29036
rect 24454 28980 24464 29036
rect 24520 28980 24568 29036
rect 24624 28980 24672 29036
rect 24728 28980 24738 29036
rect 28448 28980 28560 29008
rect 18610 28924 18620 28980
rect 18676 28924 19852 28980
rect 19908 28924 19918 28980
rect 27234 28924 27244 28980
rect 27300 28924 28560 28980
rect 28448 28896 28560 28924
rect 11106 28812 11116 28868
rect 11172 28812 11340 28868
rect 11396 28812 11406 28868
rect 12898 28812 12908 28868
rect 12964 28812 13580 28868
rect 13636 28812 13804 28868
rect 13860 28812 13870 28868
rect 18946 28812 18956 28868
rect 19012 28812 20412 28868
rect 20468 28812 20478 28868
rect 130 28700 140 28756
rect 196 28700 1596 28756
rect 1652 28700 1662 28756
rect 2146 28700 2156 28756
rect 2212 28700 6972 28756
rect 7028 28700 7038 28756
rect 12124 28700 15148 28756
rect 16146 28700 16156 28756
rect 16212 28700 26572 28756
rect 26628 28700 26638 28756
rect 12124 28644 12180 28700
rect 15092 28644 15148 28700
rect 5506 28588 5516 28644
rect 5572 28588 12180 28644
rect 12450 28588 12460 28644
rect 12516 28588 14364 28644
rect 14420 28588 14430 28644
rect 15092 28588 24220 28644
rect 24276 28588 24286 28644
rect 28448 28532 28560 28560
rect 1250 28476 1260 28532
rect 1316 28476 2716 28532
rect 2772 28476 3500 28532
rect 3556 28476 4732 28532
rect 4788 28476 5180 28532
rect 5236 28476 5246 28532
rect 6626 28476 6636 28532
rect 6692 28476 7420 28532
rect 7476 28476 8540 28532
rect 8596 28476 10892 28532
rect 10948 28476 10958 28532
rect 14578 28476 14588 28532
rect 14644 28476 14924 28532
rect 14980 28476 14990 28532
rect 27234 28476 27244 28532
rect 27300 28476 28560 28532
rect 28448 28448 28560 28476
rect 6402 28364 6412 28420
rect 6468 28364 24668 28420
rect 24724 28364 24734 28420
rect 9090 28252 9100 28308
rect 9156 28252 14028 28308
rect 14084 28252 14094 28308
rect 3794 28196 3804 28252
rect 3860 28196 3908 28252
rect 3964 28196 4012 28252
rect 4068 28196 4078 28252
rect 23794 28196 23804 28252
rect 23860 28196 23908 28252
rect 23964 28196 24012 28252
rect 24068 28196 24078 28252
rect 13682 28140 13692 28196
rect 13748 28140 14364 28196
rect 14420 28140 14430 28196
rect 0 28084 112 28112
rect 28448 28084 28560 28112
rect 0 28028 3388 28084
rect 3444 28028 3454 28084
rect 8978 28028 8988 28084
rect 9044 28028 9324 28084
rect 9380 28028 18396 28084
rect 18452 28028 18462 28084
rect 20066 28028 20076 28084
rect 20132 28028 26348 28084
rect 26404 28028 26414 28084
rect 27234 28028 27244 28084
rect 27300 28028 28560 28084
rect 0 28000 112 28028
rect 28448 28000 28560 28028
rect 14466 27916 14476 27972
rect 14532 27916 16212 27972
rect 16370 27916 16380 27972
rect 16436 27916 17500 27972
rect 17556 27916 17836 27972
rect 17892 27916 17902 27972
rect 16156 27860 16212 27916
rect 4274 27804 4284 27860
rect 4340 27804 5292 27860
rect 5348 27804 5358 27860
rect 5730 27804 5740 27860
rect 5796 27804 6972 27860
rect 7028 27804 7038 27860
rect 8194 27804 8204 27860
rect 8260 27804 9324 27860
rect 9380 27804 9390 27860
rect 10966 27804 11004 27860
rect 11060 27804 11452 27860
rect 11508 27804 11518 27860
rect 14018 27804 14028 27860
rect 14084 27804 15148 27860
rect 15204 27804 15214 27860
rect 16156 27804 25228 27860
rect 25284 27804 25294 27860
rect 26852 27804 27692 27860
rect 27748 27804 27758 27860
rect 26852 27748 26908 27804
rect 3154 27692 3164 27748
rect 3220 27692 13356 27748
rect 13412 27692 13422 27748
rect 14914 27692 14924 27748
rect 14980 27692 15820 27748
rect 15876 27692 26908 27748
rect 28448 27636 28560 27664
rect 354 27580 364 27636
rect 420 27580 1036 27636
rect 1092 27580 1102 27636
rect 1810 27580 1820 27636
rect 1876 27580 3164 27636
rect 3220 27580 3230 27636
rect 14578 27580 14588 27636
rect 14644 27580 15596 27636
rect 15652 27580 15662 27636
rect 17490 27580 17500 27636
rect 17556 27580 18396 27636
rect 18452 27580 18462 27636
rect 20636 27580 26236 27636
rect 26292 27580 26302 27636
rect 27234 27580 27244 27636
rect 27300 27580 28560 27636
rect 11442 27468 11452 27524
rect 11508 27468 11564 27524
rect 11620 27468 11630 27524
rect 4454 27412 4464 27468
rect 4520 27412 4568 27468
rect 4624 27412 4672 27468
rect 4728 27412 4738 27468
rect 20636 27412 20692 27580
rect 28448 27552 28560 27580
rect 24454 27412 24464 27468
rect 24520 27412 24568 27468
rect 24624 27412 24672 27468
rect 24728 27412 24738 27468
rect 4946 27356 4956 27412
rect 5012 27356 6244 27412
rect 8642 27356 8652 27412
rect 8708 27356 20692 27412
rect 6188 27300 6244 27356
rect 5394 27244 5404 27300
rect 5460 27244 5964 27300
rect 6020 27244 6030 27300
rect 6188 27244 26908 27300
rect 26964 27244 26974 27300
rect 28448 27188 28560 27216
rect 1138 27132 1148 27188
rect 1204 27132 1708 27188
rect 1764 27132 1774 27188
rect 3042 27132 3052 27188
rect 3108 27132 4172 27188
rect 4228 27132 4238 27188
rect 5506 27132 5516 27188
rect 5572 27132 6076 27188
rect 6132 27132 6142 27188
rect 11218 27132 11228 27188
rect 11284 27132 11676 27188
rect 11732 27132 11742 27188
rect 14690 27132 14700 27188
rect 14756 27132 24668 27188
rect 24724 27132 24734 27188
rect 25666 27132 25676 27188
rect 25732 27132 28560 27188
rect 28448 27104 28560 27132
rect 354 27020 364 27076
rect 420 27020 2268 27076
rect 2324 27020 3388 27076
rect 3444 27020 3454 27076
rect 10882 27020 10892 27076
rect 10948 27020 16380 27076
rect 16436 27020 16446 27076
rect 17350 27020 17388 27076
rect 17444 27020 17454 27076
rect 18050 27020 18060 27076
rect 18116 27020 18396 27076
rect 18452 27020 18462 27076
rect 11340 26964 11396 27020
rect 1698 26908 1708 26964
rect 1764 26908 3724 26964
rect 3780 26908 3790 26964
rect 4946 26908 4956 26964
rect 5012 26908 6300 26964
rect 6356 26908 6366 26964
rect 11330 26908 11340 26964
rect 11396 26908 11406 26964
rect 16482 26908 16492 26964
rect 16548 26908 17612 26964
rect 17668 26908 17678 26964
rect 4386 26796 4396 26852
rect 4452 26796 16940 26852
rect 16996 26796 17006 26852
rect 17350 26796 17388 26852
rect 17444 26796 18284 26852
rect 18340 26796 18350 26852
rect 0 26740 112 26768
rect 28448 26740 28560 26768
rect 0 26684 1036 26740
rect 1092 26684 1102 26740
rect 5730 26684 5740 26740
rect 5796 26684 5964 26740
rect 6020 26684 6030 26740
rect 9100 26684 12796 26740
rect 12852 26684 12862 26740
rect 27234 26684 27244 26740
rect 27300 26684 28560 26740
rect 0 26656 112 26684
rect 3794 26628 3804 26684
rect 3860 26628 3908 26684
rect 3964 26628 4012 26684
rect 4068 26628 4078 26684
rect 242 26572 252 26628
rect 308 26572 700 26628
rect 756 26572 766 26628
rect 4274 26572 4284 26628
rect 4340 26572 6300 26628
rect 6356 26572 6366 26628
rect 9100 26516 9156 26684
rect 23794 26628 23804 26684
rect 23860 26628 23908 26684
rect 23964 26628 24012 26684
rect 24068 26628 24078 26684
rect 28448 26656 28560 26684
rect 2930 26460 2940 26516
rect 2996 26460 9156 26516
rect 9212 26572 16268 26628
rect 16324 26572 16940 26628
rect 16996 26572 17006 26628
rect 9212 26404 9268 26572
rect 11414 26460 11452 26516
rect 11508 26460 11518 26516
rect 13346 26460 13356 26516
rect 13412 26460 17164 26516
rect 17220 26460 17230 26516
rect 18274 26460 18284 26516
rect 18340 26460 19180 26516
rect 19236 26460 20188 26516
rect 242 26348 252 26404
rect 308 26348 9268 26404
rect 20132 26292 20188 26460
rect 25218 26348 25228 26404
rect 25284 26348 25564 26404
rect 25620 26348 25630 26404
rect 28448 26292 28560 26320
rect 2818 26236 2828 26292
rect 2884 26236 5964 26292
rect 6020 26236 6030 26292
rect 6290 26236 6300 26292
rect 6356 26236 7644 26292
rect 7700 26236 13468 26292
rect 13524 26236 13534 26292
rect 18498 26236 18508 26292
rect 18564 26236 19180 26292
rect 19236 26236 19246 26292
rect 20132 26236 25284 26292
rect 25666 26236 25676 26292
rect 25732 26236 28560 26292
rect 25228 26180 25284 26236
rect 28448 26208 28560 26236
rect 1474 26124 1484 26180
rect 1540 26124 7980 26180
rect 8036 26124 9324 26180
rect 9380 26124 9390 26180
rect 19730 26124 19740 26180
rect 19796 26124 25004 26180
rect 25060 26124 25070 26180
rect 25228 26124 27020 26180
rect 27076 26124 27086 26180
rect 2146 26012 2156 26068
rect 2212 26012 2828 26068
rect 2884 26012 2894 26068
rect 11778 26012 11788 26068
rect 11844 26012 12572 26068
rect 12628 26012 12638 26068
rect 19506 26012 19516 26068
rect 19572 26012 26236 26068
rect 26292 26012 26302 26068
rect 25554 25900 25564 25956
rect 25620 25900 26124 25956
rect 26180 25900 26190 25956
rect 4454 25844 4464 25900
rect 4520 25844 4568 25900
rect 4624 25844 4672 25900
rect 4728 25844 4738 25900
rect 24454 25844 24464 25900
rect 24520 25844 24568 25900
rect 24624 25844 24672 25900
rect 24728 25844 24738 25900
rect 28448 25844 28560 25872
rect 12898 25788 12908 25844
rect 12964 25788 20188 25844
rect 20244 25788 20254 25844
rect 27234 25788 27244 25844
rect 27300 25788 28560 25844
rect 28448 25760 28560 25788
rect 3042 25676 3052 25732
rect 3108 25676 3724 25732
rect 3780 25676 3790 25732
rect 12786 25676 12796 25732
rect 12852 25676 13132 25732
rect 13188 25676 14140 25732
rect 14196 25676 14206 25732
rect 19730 25676 19740 25732
rect 19796 25676 20412 25732
rect 20468 25676 20972 25732
rect 21028 25676 21038 25732
rect 1362 25564 1372 25620
rect 1428 25564 2044 25620
rect 2100 25564 2110 25620
rect 5954 25564 5964 25620
rect 6020 25564 6636 25620
rect 6692 25564 10332 25620
rect 10388 25564 10398 25620
rect 10770 25564 10780 25620
rect 10836 25564 24668 25620
rect 24724 25564 24734 25620
rect 3266 25452 3276 25508
rect 3332 25452 6300 25508
rect 6356 25452 6366 25508
rect 19170 25452 19180 25508
rect 19236 25452 19404 25508
rect 19460 25452 19470 25508
rect 26002 25452 26012 25508
rect 26068 25452 26236 25508
rect 26292 25452 26302 25508
rect 0 25396 112 25424
rect 28448 25396 28560 25424
rect 0 25340 1036 25396
rect 1092 25340 1102 25396
rect 1586 25340 1596 25396
rect 1652 25340 3612 25396
rect 3668 25340 3678 25396
rect 27122 25340 27132 25396
rect 27188 25340 28560 25396
rect 0 25312 112 25340
rect 28448 25312 28560 25340
rect 3042 25228 3052 25284
rect 3108 25228 3500 25284
rect 3556 25228 3566 25284
rect 12002 25228 12012 25284
rect 12068 25228 13132 25284
rect 13188 25228 13198 25284
rect 16930 25228 16940 25284
rect 16996 25228 17948 25284
rect 18004 25228 18014 25284
rect 6738 25116 6748 25172
rect 6804 25116 7420 25172
rect 7476 25116 7486 25172
rect 10546 25116 10556 25172
rect 10612 25116 12572 25172
rect 12628 25116 18060 25172
rect 18116 25116 18126 25172
rect 25778 25116 25788 25172
rect 25844 25116 26460 25172
rect 26516 25116 26526 25172
rect 3794 25060 3804 25116
rect 3860 25060 3908 25116
rect 3964 25060 4012 25116
rect 4068 25060 4078 25116
rect 23794 25060 23804 25116
rect 23860 25060 23908 25116
rect 23964 25060 24012 25116
rect 24068 25060 24078 25116
rect 2930 25004 2940 25060
rect 2996 25004 3276 25060
rect 3332 25004 3342 25060
rect 5180 25004 6860 25060
rect 6916 25004 6926 25060
rect 7074 25004 7084 25060
rect 7140 25004 7532 25060
rect 7588 25004 7598 25060
rect 10658 25004 10668 25060
rect 10724 25004 13692 25060
rect 13748 25004 13758 25060
rect 24220 25004 26348 25060
rect 26404 25004 26414 25060
rect 5180 24948 5236 25004
rect 1362 24892 1372 24948
rect 1428 24892 5236 24948
rect 5394 24892 5404 24948
rect 5460 24892 9548 24948
rect 9604 24892 9614 24948
rect 12114 24892 12124 24948
rect 12180 24892 13244 24948
rect 13300 24892 14924 24948
rect 14980 24892 14990 24948
rect 24220 24836 24276 25004
rect 28448 24948 28560 24976
rect 25666 24892 25676 24948
rect 25732 24892 28560 24948
rect 28448 24864 28560 24892
rect 1362 24780 1372 24836
rect 1428 24780 6020 24836
rect 6178 24780 6188 24836
rect 6244 24780 24276 24836
rect 25442 24780 25452 24836
rect 25508 24780 26012 24836
rect 26068 24780 26078 24836
rect 5964 24724 6020 24780
rect 2258 24668 2268 24724
rect 2324 24668 5516 24724
rect 5572 24668 5582 24724
rect 5964 24668 12684 24724
rect 12740 24668 12750 24724
rect 13346 24668 13356 24724
rect 13412 24668 16604 24724
rect 16660 24668 16670 24724
rect 18722 24668 18732 24724
rect 18788 24668 18956 24724
rect 19012 24668 19022 24724
rect 22092 24668 25228 24724
rect 25284 24668 25294 24724
rect 6178 24556 6188 24612
rect 6244 24556 10836 24612
rect 13906 24556 13916 24612
rect 13972 24556 14700 24612
rect 14756 24556 14766 24612
rect 17714 24556 17724 24612
rect 17780 24556 18060 24612
rect 18116 24556 18126 24612
rect 10780 24500 10836 24556
rect 22092 24500 22148 24668
rect 28448 24500 28560 24528
rect 4050 24444 4060 24500
rect 4116 24444 4956 24500
rect 5012 24444 5022 24500
rect 7970 24444 7980 24500
rect 8036 24444 10556 24500
rect 10612 24444 10622 24500
rect 10780 24444 22148 24500
rect 22428 24444 24668 24500
rect 24724 24444 24734 24500
rect 27234 24444 27244 24500
rect 27300 24444 28560 24500
rect 8194 24332 8204 24388
rect 8260 24332 18508 24388
rect 18564 24332 18574 24388
rect 4454 24276 4464 24332
rect 4520 24276 4568 24332
rect 4624 24276 4672 24332
rect 4728 24276 4738 24332
rect 22428 24276 22484 24444
rect 28448 24416 28560 24444
rect 24454 24276 24464 24332
rect 24520 24276 24568 24332
rect 24624 24276 24672 24332
rect 24728 24276 24738 24332
rect 8530 24220 8540 24276
rect 8596 24220 9884 24276
rect 9940 24220 9950 24276
rect 10546 24220 10556 24276
rect 10612 24220 22484 24276
rect 1362 24108 1372 24164
rect 1428 24108 8932 24164
rect 9314 24108 9324 24164
rect 9380 24108 26236 24164
rect 26292 24108 26302 24164
rect 0 24052 112 24080
rect 8876 24052 8932 24108
rect 28448 24052 28560 24080
rect 0 23996 924 24052
rect 980 23996 990 24052
rect 2370 23996 2380 24052
rect 2436 23996 4620 24052
rect 4676 23996 4686 24052
rect 8876 23996 10892 24052
rect 10948 23996 10958 24052
rect 25442 23996 25452 24052
rect 25508 23996 28560 24052
rect 0 23968 112 23996
rect 28448 23968 28560 23996
rect 4274 23884 4284 23940
rect 4340 23884 5404 23940
rect 5460 23884 5470 23940
rect 7634 23884 7644 23940
rect 7700 23884 7868 23940
rect 7924 23884 7934 23940
rect 18162 23884 18172 23940
rect 18228 23884 18396 23940
rect 18452 23884 18732 23940
rect 18788 23884 18956 23940
rect 19012 23884 19022 23940
rect 1586 23772 1596 23828
rect 1652 23772 2380 23828
rect 2436 23772 2446 23828
rect 12338 23772 12348 23828
rect 12404 23772 14252 23828
rect 14308 23772 14318 23828
rect 18498 23772 18508 23828
rect 18564 23772 20076 23828
rect 20132 23772 20142 23828
rect 6850 23660 6860 23716
rect 6916 23660 7644 23716
rect 7700 23660 7710 23716
rect 14690 23660 14700 23716
rect 14756 23660 16828 23716
rect 16884 23660 16894 23716
rect 28448 23604 28560 23632
rect 4274 23548 4284 23604
rect 4340 23548 10556 23604
rect 10612 23548 10780 23604
rect 10836 23548 10846 23604
rect 17378 23548 17388 23604
rect 17444 23548 18508 23604
rect 18564 23548 19516 23604
rect 19572 23548 19582 23604
rect 27122 23548 27132 23604
rect 27188 23548 28560 23604
rect 3794 23492 3804 23548
rect 3860 23492 3908 23548
rect 3964 23492 4012 23548
rect 4068 23492 4078 23548
rect 23794 23492 23804 23548
rect 23860 23492 23908 23548
rect 23964 23492 24012 23548
rect 24068 23492 24078 23548
rect 28448 23520 28560 23548
rect 2258 23436 2268 23492
rect 2324 23436 3612 23492
rect 3668 23436 3678 23492
rect 8082 23436 8092 23492
rect 8148 23436 9324 23492
rect 9380 23436 9390 23492
rect 1586 23324 1596 23380
rect 1652 23324 6300 23380
rect 6356 23324 6366 23380
rect 15922 23324 15932 23380
rect 15988 23324 20636 23380
rect 20692 23324 21196 23380
rect 21252 23324 21262 23380
rect 7158 23212 7196 23268
rect 7252 23212 7262 23268
rect 11974 23212 12012 23268
rect 12068 23212 12078 23268
rect 12226 23212 12236 23268
rect 12292 23212 13804 23268
rect 13860 23212 13870 23268
rect 14028 23212 26236 23268
rect 26292 23212 26302 23268
rect 14028 23156 14084 23212
rect 28448 23156 28560 23184
rect 690 23100 700 23156
rect 756 23100 2716 23156
rect 2772 23100 2782 23156
rect 6178 23100 6188 23156
rect 6244 23100 14084 23156
rect 14802 23100 14812 23156
rect 14868 23100 16044 23156
rect 16100 23100 16110 23156
rect 25666 23100 25676 23156
rect 25732 23100 28560 23156
rect 28448 23072 28560 23100
rect 7522 22988 7532 23044
rect 7588 22988 8764 23044
rect 8820 22988 8830 23044
rect 10546 22988 10556 23044
rect 10612 22988 12012 23044
rect 12068 22988 14364 23044
rect 14420 22988 14430 23044
rect 690 22876 700 22932
rect 756 22876 11676 22932
rect 11732 22876 11742 22932
rect 15138 22876 15148 22932
rect 15204 22876 16380 22932
rect 16436 22876 16446 22932
rect 0 22708 112 22736
rect 4454 22708 4464 22764
rect 4520 22708 4568 22764
rect 4624 22708 4672 22764
rect 4728 22708 4738 22764
rect 24454 22708 24464 22764
rect 24520 22708 24568 22764
rect 24624 22708 24672 22764
rect 24728 22708 24738 22764
rect 28448 22708 28560 22736
rect 0 22652 812 22708
rect 868 22652 878 22708
rect 11890 22652 11900 22708
rect 11956 22652 12236 22708
rect 12292 22652 12302 22708
rect 27234 22652 27244 22708
rect 27300 22652 28560 22708
rect 0 22624 112 22652
rect 28448 22624 28560 22652
rect 1698 22540 1708 22596
rect 1764 22540 3276 22596
rect 3332 22540 3342 22596
rect 5964 22540 25900 22596
rect 25956 22540 25966 22596
rect 5964 22484 6020 22540
rect 1138 22428 1148 22484
rect 1204 22428 6020 22484
rect 8306 22428 8316 22484
rect 8372 22428 10332 22484
rect 10388 22428 10398 22484
rect 14914 22428 14924 22484
rect 14980 22428 26236 22484
rect 26292 22428 26302 22484
rect 5394 22316 5404 22372
rect 5460 22316 5740 22372
rect 5796 22316 5806 22372
rect 6962 22316 6972 22372
rect 7028 22316 7532 22372
rect 7588 22316 7598 22372
rect 8194 22316 8204 22372
rect 8260 22316 9212 22372
rect 9268 22316 9278 22372
rect 9426 22316 9436 22372
rect 9492 22316 9660 22372
rect 9716 22316 10892 22372
rect 10948 22316 10958 22372
rect 11890 22316 11900 22372
rect 11956 22316 13692 22372
rect 13748 22316 13758 22372
rect 15810 22316 15820 22372
rect 15876 22316 17388 22372
rect 17444 22316 17454 22372
rect 28448 22260 28560 22288
rect 8082 22204 8092 22260
rect 8148 22204 13916 22260
rect 13972 22204 14476 22260
rect 14532 22204 15148 22260
rect 27122 22204 27132 22260
rect 27188 22204 28560 22260
rect 15092 22148 15148 22204
rect 28448 22176 28560 22204
rect 13010 22092 13020 22148
rect 13076 22092 13580 22148
rect 13636 22092 13646 22148
rect 15092 22092 16828 22148
rect 16884 22092 26460 22148
rect 26516 22092 26526 22148
rect 9426 21980 9436 22036
rect 9492 21980 20748 22036
rect 20804 21980 20814 22036
rect 3794 21924 3804 21980
rect 3860 21924 3908 21980
rect 3964 21924 4012 21980
rect 4068 21924 4078 21980
rect 23794 21924 23804 21980
rect 23860 21924 23908 21980
rect 23964 21924 24012 21980
rect 24068 21924 24078 21980
rect 2482 21868 2492 21924
rect 2548 21868 3052 21924
rect 3108 21868 3164 21924
rect 3220 21868 3230 21924
rect 8306 21868 8316 21924
rect 8372 21868 9660 21924
rect 9716 21868 9726 21924
rect 12002 21868 12012 21924
rect 12068 21868 12124 21924
rect 12180 21868 12190 21924
rect 13570 21868 13580 21924
rect 13636 21868 14924 21924
rect 14980 21868 14990 21924
rect 28448 21812 28560 21840
rect 2146 21756 2156 21812
rect 2212 21756 2828 21812
rect 2884 21756 2894 21812
rect 4274 21756 4284 21812
rect 4340 21756 5292 21812
rect 5348 21756 5358 21812
rect 7858 21756 7868 21812
rect 7924 21756 8092 21812
rect 8148 21756 8158 21812
rect 11330 21756 11340 21812
rect 11396 21756 11676 21812
rect 11732 21756 13132 21812
rect 13188 21756 13198 21812
rect 13356 21756 20188 21812
rect 25666 21756 25676 21812
rect 25732 21756 28560 21812
rect 13356 21700 13412 21756
rect 20132 21700 20188 21756
rect 28448 21728 28560 21756
rect 2034 21644 2044 21700
rect 2100 21644 6300 21700
rect 6356 21644 7980 21700
rect 8036 21644 9772 21700
rect 9828 21644 13412 21700
rect 13794 21644 13804 21700
rect 13860 21644 16156 21700
rect 16212 21644 16716 21700
rect 16772 21644 17892 21700
rect 20132 21644 26124 21700
rect 26180 21644 26190 21700
rect 17836 21588 17892 21644
rect 2146 21532 2156 21588
rect 2212 21532 2604 21588
rect 2660 21532 2670 21588
rect 6962 21532 6972 21588
rect 7028 21532 7084 21588
rect 7140 21532 7150 21588
rect 8978 21532 8988 21588
rect 9044 21532 10108 21588
rect 10164 21532 10174 21588
rect 16370 21532 16380 21588
rect 16436 21532 17612 21588
rect 17668 21532 17678 21588
rect 17836 21532 20188 21588
rect 20132 21476 20188 21532
rect 15250 21420 15260 21476
rect 15316 21420 17164 21476
rect 17220 21420 17230 21476
rect 19282 21420 19292 21476
rect 19348 21420 19358 21476
rect 20132 21420 28252 21476
rect 28308 21420 28318 21476
rect 0 21364 112 21392
rect 19292 21364 19348 21420
rect 28448 21364 28560 21392
rect 0 21308 1148 21364
rect 1204 21308 1214 21364
rect 5954 21308 5964 21364
rect 6020 21308 7308 21364
rect 7364 21308 7374 21364
rect 9762 21308 9772 21364
rect 9828 21308 11452 21364
rect 11508 21308 12124 21364
rect 12180 21308 12190 21364
rect 12898 21308 12908 21364
rect 12964 21308 13244 21364
rect 13300 21308 13310 21364
rect 14690 21308 14700 21364
rect 14756 21308 15708 21364
rect 15764 21308 15774 21364
rect 16930 21308 16940 21364
rect 16996 21308 18396 21364
rect 18452 21308 18462 21364
rect 19292 21308 26236 21364
rect 26292 21308 26302 21364
rect 27458 21308 27468 21364
rect 27524 21308 28560 21364
rect 0 21280 112 21308
rect 28448 21280 28560 21308
rect 12450 21196 12460 21252
rect 12516 21196 13020 21252
rect 13076 21196 13086 21252
rect 17714 21196 17724 21252
rect 17780 21196 18284 21252
rect 18340 21196 18350 21252
rect 4454 21140 4464 21196
rect 4520 21140 4568 21196
rect 4624 21140 4672 21196
rect 4728 21140 4738 21196
rect 24454 21140 24464 21196
rect 24520 21140 24568 21196
rect 24624 21140 24672 21196
rect 24728 21140 24738 21196
rect 5058 21084 5068 21140
rect 5124 21084 5292 21140
rect 5348 21084 14812 21140
rect 14868 21084 14878 21140
rect 2034 20972 2044 21028
rect 2100 20972 2268 21028
rect 2324 20972 2334 21028
rect 6290 20972 6300 21028
rect 6356 20972 26348 21028
rect 26404 20972 26414 21028
rect 28448 20916 28560 20944
rect 1334 20860 1372 20916
rect 1428 20860 1438 20916
rect 1922 20860 1932 20916
rect 1988 20860 3276 20916
rect 3332 20860 3342 20916
rect 5618 20860 5628 20916
rect 5684 20860 6636 20916
rect 6692 20860 7196 20916
rect 7252 20860 7262 20916
rect 9874 20860 9884 20916
rect 9940 20860 10444 20916
rect 10500 20860 10510 20916
rect 13234 20860 13244 20916
rect 13300 20860 17052 20916
rect 17108 20860 17118 20916
rect 17714 20860 17724 20916
rect 17780 20860 17948 20916
rect 18004 20860 18014 20916
rect 19170 20860 19180 20916
rect 19236 20860 19404 20916
rect 19460 20860 19470 20916
rect 19730 20860 19740 20916
rect 19796 20860 20412 20916
rect 20468 20860 20478 20916
rect 25890 20860 25900 20916
rect 25956 20860 28560 20916
rect 28448 20832 28560 20860
rect 2482 20748 2492 20804
rect 2548 20748 2940 20804
rect 2996 20748 3006 20804
rect 5842 20748 5852 20804
rect 5908 20748 6188 20804
rect 6244 20748 7196 20804
rect 7252 20748 7262 20804
rect 11554 20748 11564 20804
rect 11620 20748 12012 20804
rect 12068 20748 12078 20804
rect 12338 20748 12348 20804
rect 12404 20748 12684 20804
rect 12740 20748 12750 20804
rect 13346 20748 13356 20804
rect 13412 20748 15820 20804
rect 15876 20748 16716 20804
rect 16772 20748 17388 20804
rect 17444 20748 17454 20804
rect 354 20636 364 20692
rect 420 20636 1036 20692
rect 1092 20636 1102 20692
rect 3602 20636 3612 20692
rect 3668 20636 10780 20692
rect 10836 20636 10846 20692
rect 17042 20636 17052 20692
rect 17108 20636 18396 20692
rect 18452 20636 18462 20692
rect 18946 20636 18956 20692
rect 19012 20636 19180 20692
rect 19236 20636 19246 20692
rect 1586 20524 1596 20580
rect 1652 20524 15148 20580
rect 15092 20468 15148 20524
rect 28448 20468 28560 20496
rect 578 20412 588 20468
rect 644 20412 1372 20468
rect 1428 20412 1438 20468
rect 7410 20412 7420 20468
rect 7476 20412 14196 20468
rect 15092 20412 16940 20468
rect 16996 20412 17006 20468
rect 27458 20412 27468 20468
rect 27524 20412 28560 20468
rect 3794 20356 3804 20412
rect 3860 20356 3908 20412
rect 3964 20356 4012 20412
rect 4068 20356 4078 20412
rect 14140 20356 14196 20412
rect 23794 20356 23804 20412
rect 23860 20356 23908 20412
rect 23964 20356 24012 20412
rect 24068 20356 24078 20412
rect 28448 20384 28560 20412
rect 10098 20300 10108 20356
rect 10164 20300 13804 20356
rect 13860 20300 13870 20356
rect 14140 20300 20188 20356
rect 20132 20244 20188 20300
rect 1250 20188 1260 20244
rect 1316 20188 1326 20244
rect 9426 20188 9436 20244
rect 9492 20188 10556 20244
rect 10612 20188 11900 20244
rect 11956 20188 11966 20244
rect 16034 20188 16044 20244
rect 16100 20188 16716 20244
rect 16772 20188 16782 20244
rect 20132 20188 25340 20244
rect 25396 20188 25406 20244
rect 1260 20132 1316 20188
rect 1260 20076 1596 20132
rect 1652 20076 1662 20132
rect 2034 20076 2044 20132
rect 2100 20076 3836 20132
rect 3892 20076 4172 20132
rect 4228 20076 4238 20132
rect 6150 20076 6188 20132
rect 6244 20076 6254 20132
rect 6738 20076 6748 20132
rect 6804 20076 8988 20132
rect 9044 20076 9054 20132
rect 11106 20076 11116 20132
rect 11172 20076 12012 20132
rect 12068 20076 14364 20132
rect 14420 20076 14430 20132
rect 17826 20076 17836 20132
rect 17892 20076 18172 20132
rect 18228 20076 18238 20132
rect 20132 20076 26012 20132
rect 26068 20076 26078 20132
rect 27010 20076 27020 20132
rect 27076 20076 27916 20132
rect 27972 20076 27982 20132
rect 0 20020 112 20048
rect 20132 20020 20188 20076
rect 28448 20020 28560 20048
rect 0 19964 1932 20020
rect 1988 19964 1998 20020
rect 4498 19964 4508 20020
rect 4564 19964 5740 20020
rect 5796 19964 7476 20020
rect 8306 19964 8316 20020
rect 8372 19964 12180 20020
rect 0 19936 112 19964
rect 3332 19852 7196 19908
rect 7252 19852 7262 19908
rect 3332 19796 3388 19852
rect 130 19740 140 19796
rect 196 19740 3388 19796
rect 7420 19796 7476 19964
rect 12124 19908 12180 19964
rect 13244 19964 20188 20020
rect 26562 19964 26572 20020
rect 26628 19964 28560 20020
rect 8418 19852 8428 19908
rect 8484 19852 9324 19908
rect 9380 19852 9390 19908
rect 12114 19852 12124 19908
rect 12180 19852 13020 19908
rect 13076 19852 13086 19908
rect 13244 19796 13300 19964
rect 28448 19936 28560 19964
rect 14018 19852 14028 19908
rect 14084 19852 14476 19908
rect 14532 19852 14542 19908
rect 15026 19852 15036 19908
rect 15092 19852 25564 19908
rect 25620 19852 25630 19908
rect 7420 19740 13300 19796
rect 14242 19740 14252 19796
rect 14308 19740 15596 19796
rect 15652 19740 15662 19796
rect 1586 19628 1596 19684
rect 1652 19628 2716 19684
rect 2772 19628 2782 19684
rect 9538 19628 9548 19684
rect 9604 19628 12348 19684
rect 12404 19628 12572 19684
rect 12628 19628 12638 19684
rect 13234 19628 13244 19684
rect 13300 19628 13804 19684
rect 13860 19628 13870 19684
rect 14018 19628 14028 19684
rect 14084 19628 14588 19684
rect 14644 19628 16044 19684
rect 16100 19628 16110 19684
rect 4454 19572 4464 19628
rect 4520 19572 4568 19628
rect 4624 19572 4672 19628
rect 4728 19572 4738 19628
rect 24454 19572 24464 19628
rect 24520 19572 24568 19628
rect 24624 19572 24672 19628
rect 24728 19572 24738 19628
rect 28448 19572 28560 19600
rect 11666 19516 11676 19572
rect 11732 19516 13412 19572
rect 13906 19516 13916 19572
rect 13972 19516 16716 19572
rect 16772 19516 16782 19572
rect 27458 19516 27468 19572
rect 27524 19516 28560 19572
rect 13356 19460 13412 19516
rect 28448 19488 28560 19516
rect 1586 19404 1596 19460
rect 1652 19404 2604 19460
rect 2660 19404 2670 19460
rect 5730 19404 5740 19460
rect 5796 19404 6524 19460
rect 6580 19404 6590 19460
rect 9986 19404 9996 19460
rect 10052 19404 11564 19460
rect 11620 19404 11630 19460
rect 13356 19404 15484 19460
rect 15540 19404 16604 19460
rect 16660 19404 16670 19460
rect 2706 19292 2716 19348
rect 2772 19292 3388 19348
rect 3444 19292 4508 19348
rect 4564 19292 4574 19348
rect 5954 19292 5964 19348
rect 6020 19292 6636 19348
rect 6692 19292 6702 19348
rect 6962 19292 6972 19348
rect 7028 19292 7420 19348
rect 7476 19292 7486 19348
rect 10210 19292 10220 19348
rect 10276 19292 11676 19348
rect 11732 19292 12572 19348
rect 12628 19292 12638 19348
rect 13122 19292 13132 19348
rect 13188 19292 13916 19348
rect 13972 19292 13982 19348
rect 14802 19292 14812 19348
rect 14868 19292 25900 19348
rect 25956 19292 25966 19348
rect 8082 19180 8092 19236
rect 8148 19180 10332 19236
rect 10388 19180 10398 19236
rect 12226 19180 12236 19236
rect 12292 19180 13356 19236
rect 13412 19180 13422 19236
rect 15026 19180 15036 19236
rect 15092 19180 16604 19236
rect 16660 19180 16670 19236
rect 10332 19124 10388 19180
rect 28448 19124 28560 19152
rect 2258 19068 2268 19124
rect 2324 19068 3164 19124
rect 3220 19068 3612 19124
rect 3668 19068 3678 19124
rect 6626 19068 6636 19124
rect 6692 19068 6860 19124
rect 6916 19068 7420 19124
rect 7476 19068 7486 19124
rect 10332 19068 13244 19124
rect 13300 19068 13310 19124
rect 27458 19068 27468 19124
rect 27524 19068 28560 19124
rect 28448 19040 28560 19068
rect 3612 18956 3836 19012
rect 3892 18956 3902 19012
rect 3612 18900 3668 18956
rect 3602 18844 3612 18900
rect 3668 18844 3678 18900
rect 4274 18844 4284 18900
rect 4340 18844 13356 18900
rect 13412 18844 17836 18900
rect 17892 18844 17902 18900
rect 3794 18788 3804 18844
rect 3860 18788 3908 18844
rect 3964 18788 4012 18844
rect 4068 18788 4078 18844
rect 23794 18788 23804 18844
rect 23860 18788 23908 18844
rect 23964 18788 24012 18844
rect 24068 18788 24078 18844
rect 0 18676 112 18704
rect 28448 18676 28560 18704
rect 0 18620 924 18676
rect 980 18620 990 18676
rect 3490 18620 3500 18676
rect 3556 18620 4172 18676
rect 4228 18620 4238 18676
rect 13580 18620 13692 18676
rect 13748 18620 13758 18676
rect 15810 18620 15820 18676
rect 15876 18620 16828 18676
rect 16884 18620 16894 18676
rect 26562 18620 26572 18676
rect 26628 18620 28560 18676
rect 0 18592 112 18620
rect 3266 18508 3276 18564
rect 3332 18508 5180 18564
rect 5236 18508 5246 18564
rect 6626 18508 6636 18564
rect 6692 18508 8092 18564
rect 8148 18508 8158 18564
rect 8978 18508 8988 18564
rect 9044 18508 10332 18564
rect 10388 18508 10398 18564
rect 10994 18508 11004 18564
rect 11060 18508 12908 18564
rect 12964 18508 12974 18564
rect 13580 18452 13636 18620
rect 28448 18592 28560 18620
rect 13794 18508 13804 18564
rect 13860 18508 15260 18564
rect 15316 18508 15372 18564
rect 15428 18508 15438 18564
rect 16482 18508 16492 18564
rect 16548 18508 17052 18564
rect 17108 18508 17118 18564
rect 1698 18396 1708 18452
rect 1764 18396 2604 18452
rect 2660 18396 2670 18452
rect 3126 18396 3164 18452
rect 3220 18396 3230 18452
rect 4386 18396 4396 18452
rect 4452 18396 4844 18452
rect 4900 18396 4910 18452
rect 5506 18396 5516 18452
rect 5572 18396 8540 18452
rect 8596 18396 8606 18452
rect 10770 18396 10780 18452
rect 10836 18396 14420 18452
rect 14578 18396 14588 18452
rect 14644 18396 14924 18452
rect 14980 18396 15708 18452
rect 15764 18396 15774 18452
rect 15922 18396 15932 18452
rect 15988 18396 18004 18452
rect 19506 18396 19516 18452
rect 19572 18396 21084 18452
rect 21140 18396 21150 18452
rect 26338 18396 26348 18452
rect 26404 18396 26684 18452
rect 26740 18396 26750 18452
rect 26898 18396 26908 18452
rect 26964 18396 27804 18452
rect 27860 18396 27870 18452
rect 2604 18340 2660 18396
rect 14364 18340 14420 18396
rect 17948 18340 18004 18396
rect 2604 18284 10668 18340
rect 10724 18284 10734 18340
rect 11890 18284 11900 18340
rect 11956 18284 14028 18340
rect 14084 18284 14094 18340
rect 14364 18284 14812 18340
rect 14868 18284 14878 18340
rect 15362 18284 15372 18340
rect 15428 18284 15820 18340
rect 15876 18284 15886 18340
rect 16034 18284 16044 18340
rect 16100 18284 17388 18340
rect 17444 18284 17454 18340
rect 17938 18284 17948 18340
rect 18004 18284 21308 18340
rect 21364 18284 21374 18340
rect 28448 18228 28560 18256
rect 2034 18172 2044 18228
rect 2100 18172 3836 18228
rect 3892 18172 6076 18228
rect 6132 18172 6972 18228
rect 7028 18172 7038 18228
rect 14364 18172 15148 18228
rect 15204 18172 17164 18228
rect 17220 18172 17230 18228
rect 17826 18172 17836 18228
rect 17892 18172 18620 18228
rect 18676 18172 18956 18228
rect 19012 18172 19022 18228
rect 27468 18172 28560 18228
rect 14364 18116 14420 18172
rect 1698 18060 1708 18116
rect 1764 18060 2492 18116
rect 2548 18060 2558 18116
rect 14354 18060 14364 18116
rect 14420 18060 14430 18116
rect 14578 18060 14588 18116
rect 14644 18060 14682 18116
rect 4454 18004 4464 18060
rect 4520 18004 4568 18060
rect 4624 18004 4672 18060
rect 4728 18004 4738 18060
rect 24454 18004 24464 18060
rect 24520 18004 24568 18060
rect 24624 18004 24672 18060
rect 24728 18004 24738 18060
rect 27468 18004 27524 18172
rect 28448 18144 28560 18172
rect 11554 17948 11564 18004
rect 11620 17948 14700 18004
rect 14756 17948 14766 18004
rect 27458 17948 27468 18004
rect 27524 17948 27534 18004
rect 662 17836 700 17892
rect 756 17836 766 17892
rect 3714 17836 3724 17892
rect 3780 17836 4620 17892
rect 4676 17836 4686 17892
rect 4834 17836 4844 17892
rect 4900 17836 5404 17892
rect 5460 17836 9996 17892
rect 10052 17836 10062 17892
rect 14578 17836 14588 17892
rect 14644 17836 16940 17892
rect 16996 17836 17006 17892
rect 18386 17836 18396 17892
rect 18452 17836 26124 17892
rect 26180 17836 26190 17892
rect 26898 17836 26908 17892
rect 26964 17836 28028 17892
rect 28084 17836 28094 17892
rect 28448 17780 28560 17808
rect 242 17724 252 17780
rect 308 17724 1596 17780
rect 1652 17724 1662 17780
rect 2146 17724 2156 17780
rect 2212 17724 4284 17780
rect 4340 17724 4350 17780
rect 14690 17724 14700 17780
rect 14756 17724 17108 17780
rect 26674 17724 26684 17780
rect 26740 17724 28560 17780
rect 2482 17612 2492 17668
rect 2548 17612 3388 17668
rect 3602 17612 3612 17668
rect 3668 17612 6636 17668
rect 6692 17612 6702 17668
rect 3332 17556 3388 17612
rect 17052 17556 17108 17724
rect 28448 17696 28560 17724
rect 17490 17612 17500 17668
rect 17556 17612 27916 17668
rect 27972 17612 27982 17668
rect 3332 17500 10892 17556
rect 10948 17500 10958 17556
rect 11218 17500 11228 17556
rect 11284 17500 15260 17556
rect 15316 17500 16044 17556
rect 16100 17500 16828 17556
rect 16884 17500 16894 17556
rect 17052 17500 27020 17556
rect 27076 17500 27086 17556
rect 662 17388 700 17444
rect 756 17388 766 17444
rect 3332 17388 5516 17444
rect 5572 17388 5582 17444
rect 0 17332 112 17360
rect 0 17276 1932 17332
rect 1988 17276 1998 17332
rect 0 17248 112 17276
rect 3332 17108 3388 17388
rect 28448 17332 28560 17360
rect 8306 17276 8316 17332
rect 8372 17276 15708 17332
rect 15764 17276 15774 17332
rect 27458 17276 27468 17332
rect 27524 17276 28560 17332
rect 3794 17220 3804 17276
rect 3860 17220 3908 17276
rect 3964 17220 4012 17276
rect 4068 17220 4078 17276
rect 23794 17220 23804 17276
rect 23860 17220 23908 17276
rect 23964 17220 24012 17276
rect 24068 17220 24078 17276
rect 28448 17248 28560 17276
rect 11778 17164 11788 17220
rect 11844 17164 14476 17220
rect 14532 17164 14542 17220
rect 14802 17164 14812 17220
rect 14868 17164 15820 17220
rect 15876 17164 15886 17220
rect 354 17052 364 17108
rect 420 17052 3388 17108
rect 10322 17052 10332 17108
rect 10388 17052 10398 17108
rect 14018 17052 14028 17108
rect 14084 17052 16492 17108
rect 16548 17052 16558 17108
rect 21298 17052 21308 17108
rect 21364 17052 28252 17108
rect 28308 17052 28318 17108
rect 3238 16940 3276 16996
rect 3332 16940 3342 16996
rect 2930 16828 2940 16884
rect 2996 16828 3612 16884
rect 3668 16828 3678 16884
rect 3826 16828 3836 16884
rect 3892 16828 4956 16884
rect 5012 16828 5740 16884
rect 5796 16828 6636 16884
rect 6692 16828 7868 16884
rect 7924 16828 7934 16884
rect 9650 16828 9660 16884
rect 9716 16828 10164 16884
rect 10108 16772 10164 16828
rect 10332 16772 10388 17052
rect 13570 16940 13580 16996
rect 13636 16940 16380 16996
rect 16436 16940 16446 16996
rect 28448 16884 28560 16912
rect 13122 16828 13132 16884
rect 13188 16828 13356 16884
rect 13412 16828 13422 16884
rect 15026 16828 15036 16884
rect 15092 16828 15260 16884
rect 15316 16828 15326 16884
rect 15586 16828 15596 16884
rect 15652 16828 16604 16884
rect 16660 16828 16940 16884
rect 16996 16828 17006 16884
rect 26562 16828 26572 16884
rect 26628 16828 28560 16884
rect 28448 16800 28560 16828
rect 5170 16716 5180 16772
rect 5236 16716 6188 16772
rect 6244 16716 7084 16772
rect 7140 16716 7150 16772
rect 10108 16716 13748 16772
rect 14578 16716 14588 16772
rect 14644 16716 15708 16772
rect 15764 16716 15774 16772
rect 13692 16660 13748 16716
rect 1138 16604 1148 16660
rect 1204 16604 1708 16660
rect 1764 16604 1774 16660
rect 2258 16604 2268 16660
rect 2324 16604 2828 16660
rect 2884 16604 5404 16660
rect 5460 16604 5470 16660
rect 10770 16604 10780 16660
rect 10836 16604 12124 16660
rect 12180 16604 12190 16660
rect 13682 16604 13692 16660
rect 13748 16604 13758 16660
rect 13906 16604 13916 16660
rect 13972 16604 20188 16660
rect 9986 16492 9996 16548
rect 10052 16492 15764 16548
rect 4454 16436 4464 16492
rect 4520 16436 4568 16492
rect 4624 16436 4672 16492
rect 4728 16436 4738 16492
rect 9538 16380 9548 16436
rect 9604 16380 12236 16436
rect 12292 16380 12302 16436
rect 14354 16380 14364 16436
rect 14420 16380 14588 16436
rect 14644 16380 14654 16436
rect 3042 16268 3052 16324
rect 3108 16268 3388 16324
rect 4274 16268 4284 16324
rect 4340 16268 5628 16324
rect 5684 16268 7980 16324
rect 8036 16268 8046 16324
rect 8194 16268 8204 16324
rect 8260 16268 11116 16324
rect 11172 16268 11182 16324
rect 3332 16212 3388 16268
rect 15708 16212 15764 16492
rect 20132 16324 20188 16604
rect 24454 16436 24464 16492
rect 24520 16436 24568 16492
rect 24624 16436 24672 16492
rect 24728 16436 24738 16492
rect 28448 16436 28560 16464
rect 27458 16380 27468 16436
rect 27524 16380 28560 16436
rect 28448 16352 28560 16380
rect 20132 16268 27132 16324
rect 27188 16268 27198 16324
rect 3332 16156 4732 16212
rect 4788 16156 8316 16212
rect 8372 16156 8382 16212
rect 10098 16156 10108 16212
rect 10164 16156 11676 16212
rect 11732 16156 15540 16212
rect 15708 16156 25900 16212
rect 25956 16156 25966 16212
rect 15484 16100 15540 16156
rect 3014 16044 3052 16100
rect 3108 16044 3118 16100
rect 3490 16044 3500 16100
rect 3556 16044 4284 16100
rect 4340 16044 4350 16100
rect 9314 16044 9324 16100
rect 9380 16044 9996 16100
rect 10052 16044 10062 16100
rect 13906 16044 13916 16100
rect 13972 16044 15260 16100
rect 15316 16044 15326 16100
rect 15474 16044 15484 16100
rect 15540 16044 25788 16100
rect 25844 16044 25854 16100
rect 0 15988 112 16016
rect 28448 15988 28560 16016
rect 0 15932 588 15988
rect 644 15932 654 15988
rect 8082 15932 8092 15988
rect 8148 15932 9884 15988
rect 9940 15932 9950 15988
rect 10994 15932 11004 15988
rect 11060 15932 15372 15988
rect 15428 15932 17724 15988
rect 17780 15932 17790 15988
rect 18386 15932 18396 15988
rect 18452 15932 18620 15988
rect 18676 15932 19068 15988
rect 19124 15932 19134 15988
rect 20066 15932 20076 15988
rect 20132 15932 26012 15988
rect 26068 15932 26078 15988
rect 27458 15932 27468 15988
rect 27524 15932 28560 15988
rect 0 15904 112 15932
rect 28448 15904 28560 15932
rect 1922 15820 1932 15876
rect 1988 15820 2604 15876
rect 2660 15820 2670 15876
rect 16034 15820 16044 15876
rect 16100 15820 17612 15876
rect 17668 15820 17678 15876
rect 1698 15708 1708 15764
rect 1764 15708 2156 15764
rect 2212 15708 2222 15764
rect 7298 15708 7308 15764
rect 7364 15708 10220 15764
rect 10276 15708 10892 15764
rect 10948 15708 11116 15764
rect 11172 15708 11182 15764
rect 3794 15652 3804 15708
rect 3860 15652 3908 15708
rect 3964 15652 4012 15708
rect 4068 15652 4078 15708
rect 23794 15652 23804 15708
rect 23860 15652 23908 15708
rect 23964 15652 24012 15708
rect 24068 15652 24078 15708
rect 8316 15596 13356 15652
rect 13412 15596 13422 15652
rect 15250 15596 15260 15652
rect 15316 15596 15932 15652
rect 15988 15596 15998 15652
rect 8316 15540 8372 15596
rect 28448 15540 28560 15568
rect 3042 15484 3052 15540
rect 3108 15484 8372 15540
rect 9090 15484 9100 15540
rect 9156 15484 11900 15540
rect 11956 15484 11966 15540
rect 13906 15484 13916 15540
rect 13972 15484 18620 15540
rect 18676 15484 18686 15540
rect 26562 15484 26572 15540
rect 26628 15484 28560 15540
rect 28448 15456 28560 15484
rect 9538 15372 9548 15428
rect 9604 15372 11004 15428
rect 11060 15372 11070 15428
rect 15362 15372 15372 15428
rect 15428 15372 16380 15428
rect 16436 15372 16446 15428
rect 3052 15260 6860 15316
rect 6916 15260 6926 15316
rect 9650 15260 9660 15316
rect 9716 15260 10556 15316
rect 10612 15260 10622 15316
rect 11330 15260 11340 15316
rect 11396 15260 11406 15316
rect 14700 15260 26236 15316
rect 26292 15260 26302 15316
rect 3052 15204 3108 15260
rect 11340 15204 11396 15260
rect 14700 15204 14756 15260
rect 2818 15148 2828 15204
rect 2884 15148 3052 15204
rect 3108 15148 3118 15204
rect 3266 15148 3276 15204
rect 3332 15148 6188 15204
rect 6244 15148 6254 15204
rect 10098 15148 10108 15204
rect 10164 15148 11788 15204
rect 11844 15148 11854 15204
rect 12002 15148 12012 15204
rect 12068 15148 14756 15204
rect 14914 15148 14924 15204
rect 14980 15148 16044 15204
rect 16100 15148 16940 15204
rect 16996 15148 17006 15204
rect 14700 15092 14756 15148
rect 28448 15092 28560 15120
rect 1474 15036 1484 15092
rect 1540 15036 1932 15092
rect 1988 15036 1998 15092
rect 4284 15036 6972 15092
rect 7028 15036 13580 15092
rect 13636 15036 13646 15092
rect 14700 15036 15148 15092
rect 15204 15036 15214 15092
rect 20132 15036 27244 15092
rect 27300 15036 27310 15092
rect 27468 15036 28560 15092
rect 2034 14924 2044 14980
rect 2100 14924 3052 14980
rect 3108 14924 3118 14980
rect 4284 14868 4340 15036
rect 20132 14980 20188 15036
rect 5282 14924 5292 14980
rect 5348 14924 20188 14980
rect 4454 14868 4464 14924
rect 4520 14868 4568 14924
rect 4624 14868 4672 14924
rect 4728 14868 4738 14924
rect 24454 14868 24464 14924
rect 24520 14868 24568 14924
rect 24624 14868 24672 14924
rect 24728 14868 24738 14924
rect 27468 14868 27524 15036
rect 28448 15008 28560 15036
rect 1810 14812 1820 14868
rect 1876 14812 4340 14868
rect 5852 14812 20188 14868
rect 27458 14812 27468 14868
rect 27524 14812 27534 14868
rect 5852 14756 5908 14812
rect 20132 14756 20188 14812
rect 3266 14700 3276 14756
rect 3332 14700 5908 14756
rect 7634 14700 7644 14756
rect 7700 14700 9436 14756
rect 9492 14700 9502 14756
rect 14914 14700 14924 14756
rect 14980 14700 15820 14756
rect 15876 14700 15886 14756
rect 20132 14700 25116 14756
rect 25172 14700 25182 14756
rect 0 14644 112 14672
rect 28448 14644 28560 14672
rect 0 14588 1708 14644
rect 1764 14588 1774 14644
rect 2454 14588 2492 14644
rect 2548 14588 2558 14644
rect 9538 14588 9548 14644
rect 9604 14588 10108 14644
rect 10164 14588 10174 14644
rect 12002 14588 12012 14644
rect 12068 14588 13020 14644
rect 13076 14588 14812 14644
rect 14868 14588 16044 14644
rect 16100 14588 17052 14644
rect 17108 14588 17118 14644
rect 26674 14588 26684 14644
rect 26740 14588 28560 14644
rect 0 14560 112 14588
rect 28448 14560 28560 14588
rect 1250 14476 1260 14532
rect 1316 14476 1932 14532
rect 1988 14476 1998 14532
rect 9426 14476 9436 14532
rect 9492 14476 9502 14532
rect 9986 14476 9996 14532
rect 10052 14476 12684 14532
rect 12740 14476 13244 14532
rect 13300 14476 13310 14532
rect 15698 14476 15708 14532
rect 15764 14476 17164 14532
rect 17220 14476 17230 14532
rect 9436 14420 9492 14476
rect 466 14364 476 14420
rect 532 14364 1148 14420
rect 1204 14364 5292 14420
rect 5348 14364 5358 14420
rect 9436 14364 11284 14420
rect 15922 14364 15932 14420
rect 15988 14364 16492 14420
rect 16548 14364 16558 14420
rect 17042 14364 17052 14420
rect 17108 14364 17500 14420
rect 17556 14364 17566 14420
rect 27542 14364 27580 14420
rect 27636 14364 27646 14420
rect 27794 14364 27804 14420
rect 27860 14364 28364 14420
rect 28420 14364 28430 14420
rect 4844 14308 4900 14364
rect 11228 14308 11284 14364
rect 4834 14252 4844 14308
rect 4900 14252 4910 14308
rect 9426 14252 9436 14308
rect 9492 14252 11004 14308
rect 11060 14252 11070 14308
rect 11228 14252 15260 14308
rect 15316 14252 15326 14308
rect 16370 14252 16380 14308
rect 16436 14252 16940 14308
rect 16996 14252 17006 14308
rect 20132 14252 27020 14308
rect 27076 14252 27086 14308
rect 20132 14196 20188 14252
rect 28448 14196 28560 14224
rect 4162 14140 4172 14196
rect 4228 14140 4508 14196
rect 4564 14140 20188 14196
rect 27458 14140 27468 14196
rect 27524 14140 28560 14196
rect 3794 14084 3804 14140
rect 3860 14084 3908 14140
rect 3964 14084 4012 14140
rect 4068 14084 4078 14140
rect 23794 14084 23804 14140
rect 23860 14084 23908 14140
rect 23964 14084 24012 14140
rect 24068 14084 24078 14140
rect 28448 14112 28560 14140
rect 4946 14028 4956 14084
rect 5012 14028 14308 14084
rect 2482 13916 2492 13972
rect 2548 13916 4284 13972
rect 4340 13916 5628 13972
rect 5684 13916 5694 13972
rect 14252 13860 14308 14028
rect 14914 13916 14924 13972
rect 14980 13916 17052 13972
rect 17108 13916 17118 13972
rect 18386 13916 18396 13972
rect 18452 13916 28028 13972
rect 28084 13916 28094 13972
rect 1586 13804 1596 13860
rect 1652 13804 9772 13860
rect 9828 13804 9838 13860
rect 14252 13804 26908 13860
rect 26964 13804 26974 13860
rect 27570 13804 27580 13860
rect 27636 13804 27692 13860
rect 27748 13804 27758 13860
rect 28448 13748 28560 13776
rect 466 13692 476 13748
rect 532 13692 1932 13748
rect 1988 13692 1998 13748
rect 2146 13692 2156 13748
rect 2212 13692 2222 13748
rect 4274 13692 4284 13748
rect 4340 13692 6412 13748
rect 6468 13692 6478 13748
rect 16034 13692 16044 13748
rect 16100 13692 16828 13748
rect 16884 13692 16894 13748
rect 17042 13692 17052 13748
rect 17108 13692 23716 13748
rect 26562 13692 26572 13748
rect 26628 13692 28560 13748
rect 1110 13580 1148 13636
rect 1204 13580 1214 13636
rect 1026 13468 1036 13524
rect 1092 13468 1260 13524
rect 1316 13468 1326 13524
rect 0 13300 112 13328
rect 2156 13300 2212 13692
rect 3378 13580 3388 13636
rect 3444 13580 4172 13636
rect 4228 13580 4238 13636
rect 8754 13580 8764 13636
rect 8820 13580 14420 13636
rect 15250 13580 15260 13636
rect 15316 13580 15820 13636
rect 15876 13580 15886 13636
rect 14364 13524 14420 13580
rect 20132 13524 20244 13636
rect 23660 13524 23716 13692
rect 28448 13664 28560 13692
rect 23874 13580 23884 13636
rect 23940 13580 26908 13636
rect 26964 13580 26974 13636
rect 5842 13468 5852 13524
rect 5908 13468 6748 13524
rect 6804 13468 6814 13524
rect 13570 13468 13580 13524
rect 13636 13468 14140 13524
rect 14196 13468 14206 13524
rect 14364 13468 23604 13524
rect 23660 13468 27244 13524
rect 27300 13468 27310 13524
rect 23548 13412 23604 13468
rect 15222 13356 15260 13412
rect 15316 13356 15326 13412
rect 23548 13356 23884 13412
rect 23940 13356 23950 13412
rect 4454 13300 4464 13356
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4728 13300 4738 13356
rect 24454 13300 24464 13356
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24728 13300 24738 13356
rect 28448 13300 28560 13328
rect 0 13244 1148 13300
rect 1204 13244 1214 13300
rect 2146 13244 2156 13300
rect 2212 13244 3388 13300
rect 5170 13244 5180 13300
rect 5236 13244 7756 13300
rect 7812 13244 7822 13300
rect 27458 13244 27468 13300
rect 27524 13244 28560 13300
rect 0 13216 112 13244
rect 3332 13188 3388 13244
rect 5180 13188 5236 13244
rect 28448 13216 28560 13244
rect 3332 13132 5236 13188
rect 6402 13132 6412 13188
rect 6468 13132 26012 13188
rect 26068 13132 26078 13188
rect 12786 13020 12796 13076
rect 12852 13020 25676 13076
rect 25732 13020 25742 13076
rect 3714 12908 3724 12964
rect 3780 12908 4508 12964
rect 4564 12908 4574 12964
rect 7298 12908 7308 12964
rect 7364 12908 9940 12964
rect 10098 12908 10108 12964
rect 10164 12908 12236 12964
rect 12292 12908 12302 12964
rect 15474 12908 15484 12964
rect 15540 12908 16156 12964
rect 16212 12908 16222 12964
rect 8194 12796 8204 12852
rect 8260 12796 9100 12852
rect 9156 12796 9166 12852
rect 9884 12740 9940 12908
rect 28448 12852 28560 12880
rect 11890 12796 11900 12852
rect 11956 12796 26012 12852
rect 26068 12796 26078 12852
rect 27458 12796 27468 12852
rect 27524 12796 28560 12852
rect 28448 12768 28560 12796
rect 9884 12684 11788 12740
rect 11844 12684 13580 12740
rect 13636 12684 13646 12740
rect 14914 12684 14924 12740
rect 14980 12684 24892 12740
rect 24948 12684 24958 12740
rect 14578 12572 14588 12628
rect 14644 12572 14812 12628
rect 14868 12572 14878 12628
rect 3794 12516 3804 12572
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 4068 12516 4078 12572
rect 23794 12516 23804 12572
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 24068 12516 24078 12572
rect 4274 12460 4284 12516
rect 4340 12460 23380 12516
rect 23324 12404 23380 12460
rect 28448 12404 28560 12432
rect 3266 12348 3276 12404
rect 3332 12348 23100 12404
rect 23156 12348 23166 12404
rect 23324 12348 25452 12404
rect 25508 12348 25518 12404
rect 26562 12348 26572 12404
rect 26628 12348 28560 12404
rect 28448 12320 28560 12348
rect 7522 12236 7532 12292
rect 7588 12236 26012 12292
rect 26068 12236 26078 12292
rect 26898 12236 26908 12292
rect 26964 12236 27916 12292
rect 27972 12236 27982 12292
rect 1894 12124 1932 12180
rect 1988 12124 1998 12180
rect 2258 12124 2268 12180
rect 2324 12124 3724 12180
rect 3780 12124 3790 12180
rect 6626 12124 6636 12180
rect 6692 12124 6972 12180
rect 7028 12124 8204 12180
rect 8260 12124 8270 12180
rect 8530 12124 8540 12180
rect 8596 12124 9324 12180
rect 9380 12124 9390 12180
rect 15026 12124 15036 12180
rect 15092 12124 27244 12180
rect 27300 12124 27310 12180
rect 27570 12124 27580 12180
rect 27636 12124 27646 12180
rect 27580 12068 27636 12124
rect 2482 12012 2492 12068
rect 2548 12012 7084 12068
rect 7140 12012 7420 12068
rect 7476 12012 7486 12068
rect 8754 12012 8764 12068
rect 8820 12012 8988 12068
rect 9044 12012 9940 12068
rect 12114 12012 12124 12068
rect 12180 12012 14252 12068
rect 14308 12012 14318 12068
rect 27010 12012 27020 12068
rect 27076 12012 27636 12068
rect 0 11956 112 11984
rect 9884 11956 9940 12012
rect 28448 11956 28560 11984
rect 0 11900 924 11956
rect 980 11900 990 11956
rect 9874 11900 9884 11956
rect 9940 11900 26124 11956
rect 26180 11900 26190 11956
rect 27570 11900 27580 11956
rect 27636 11900 28560 11956
rect 0 11872 112 11900
rect 28448 11872 28560 11900
rect 9762 11788 9772 11844
rect 9828 11788 10108 11844
rect 10164 11788 10780 11844
rect 10836 11788 11564 11844
rect 11620 11788 11630 11844
rect 4454 11732 4464 11788
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4728 11732 4738 11788
rect 24454 11732 24464 11788
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24728 11732 24738 11788
rect 5842 11676 5852 11732
rect 5908 11676 20188 11732
rect 20132 11620 20188 11676
rect 2258 11564 2268 11620
rect 2324 11564 10556 11620
rect 10612 11564 10622 11620
rect 11666 11564 11676 11620
rect 11732 11564 12572 11620
rect 12628 11564 12638 11620
rect 13458 11564 13468 11620
rect 13524 11564 14476 11620
rect 14532 11564 14542 11620
rect 20132 11564 25340 11620
rect 25396 11564 25406 11620
rect 28448 11508 28560 11536
rect 3266 11452 3276 11508
rect 3332 11452 25228 11508
rect 25284 11452 25294 11508
rect 26674 11452 26684 11508
rect 26740 11452 28560 11508
rect 28448 11424 28560 11452
rect 1586 11340 1596 11396
rect 1652 11340 3612 11396
rect 3668 11340 4396 11396
rect 4452 11340 4462 11396
rect 8194 11340 8204 11396
rect 8260 11340 10220 11396
rect 10276 11340 10286 11396
rect 11218 11340 11228 11396
rect 11284 11340 12012 11396
rect 12068 11340 12078 11396
rect 2930 11228 2940 11284
rect 2996 11228 9436 11284
rect 9492 11228 9502 11284
rect 20132 11228 26908 11284
rect 26964 11228 26974 11284
rect 3154 11116 3164 11172
rect 3220 11116 11676 11172
rect 11732 11116 11742 11172
rect 20132 11060 20188 11228
rect 28448 11060 28560 11088
rect 9538 11004 9548 11060
rect 9604 11004 20188 11060
rect 27458 11004 27468 11060
rect 27524 11004 28560 11060
rect 3794 10948 3804 11004
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 4068 10948 4078 11004
rect 23794 10948 23804 11004
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 24068 10948 24078 11004
rect 28448 10976 28560 11004
rect 354 10780 364 10836
rect 420 10780 1596 10836
rect 1652 10780 1662 10836
rect 14018 10780 14028 10836
rect 14084 10780 26348 10836
rect 26404 10780 26414 10836
rect 578 10668 588 10724
rect 644 10668 1036 10724
rect 1092 10668 1102 10724
rect 5730 10668 5740 10724
rect 5796 10668 8204 10724
rect 8260 10668 8270 10724
rect 10994 10668 11004 10724
rect 11060 10668 26908 10724
rect 26964 10668 26974 10724
rect 0 10612 112 10640
rect 28448 10612 28560 10640
rect 0 10556 1260 10612
rect 1316 10556 1326 10612
rect 5058 10556 5068 10612
rect 5124 10556 5292 10612
rect 5348 10556 5358 10612
rect 5954 10556 5964 10612
rect 6020 10556 7084 10612
rect 7140 10556 7150 10612
rect 9650 10556 9660 10612
rect 9716 10556 10220 10612
rect 10276 10556 10892 10612
rect 10948 10556 10958 10612
rect 11218 10556 11228 10612
rect 11284 10556 13132 10612
rect 13188 10556 13198 10612
rect 13570 10556 13580 10612
rect 13636 10556 13804 10612
rect 13860 10556 13870 10612
rect 26562 10556 26572 10612
rect 26628 10556 28560 10612
rect 0 10528 112 10556
rect 28448 10528 28560 10556
rect 2146 10444 2156 10500
rect 2212 10444 13468 10500
rect 13524 10444 13534 10500
rect 4386 10332 4396 10388
rect 4452 10332 9548 10388
rect 9604 10332 10444 10388
rect 10500 10332 10510 10388
rect 4454 10164 4464 10220
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4728 10164 4738 10220
rect 24454 10164 24464 10220
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24728 10164 24738 10220
rect 28448 10164 28560 10192
rect 27458 10108 27468 10164
rect 27524 10108 28560 10164
rect 28448 10080 28560 10108
rect 3154 9996 3164 10052
rect 3220 9996 8428 10052
rect 8484 9996 8494 10052
rect 20962 9996 20972 10052
rect 21028 9996 26012 10052
rect 26068 9996 26078 10052
rect 4722 9884 4732 9940
rect 4788 9884 6300 9940
rect 6356 9884 6366 9940
rect 12002 9884 12012 9940
rect 12068 9884 12348 9940
rect 12404 9884 26908 9940
rect 26964 9884 26974 9940
rect 9874 9772 9884 9828
rect 9940 9772 13244 9828
rect 13300 9772 15148 9828
rect 15204 9772 15214 9828
rect 28448 9716 28560 9744
rect 7074 9660 7084 9716
rect 7140 9660 11228 9716
rect 11284 9660 11294 9716
rect 27458 9660 27468 9716
rect 27524 9660 28560 9716
rect 28448 9632 28560 9660
rect 1586 9548 1596 9604
rect 1652 9548 7980 9604
rect 8036 9548 10892 9604
rect 10948 9548 10958 9604
rect 3794 9380 3804 9436
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 4068 9380 4078 9436
rect 23794 9380 23804 9436
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 24068 9380 24078 9436
rect 1026 9324 1036 9380
rect 1092 9324 1484 9380
rect 1540 9324 1550 9380
rect 7410 9324 7420 9380
rect 7476 9324 9884 9380
rect 9940 9324 9950 9380
rect 0 9268 112 9296
rect 28448 9268 28560 9296
rect 0 9212 1260 9268
rect 1316 9212 1326 9268
rect 8866 9212 8876 9268
rect 8932 9212 10444 9268
rect 10500 9212 10510 9268
rect 15138 9212 15148 9268
rect 15204 9212 25788 9268
rect 25844 9212 25854 9268
rect 26562 9212 26572 9268
rect 26628 9212 28560 9268
rect 0 9184 112 9212
rect 28448 9184 28560 9212
rect 2034 9100 2044 9156
rect 2100 9100 7196 9156
rect 7252 9100 7262 9156
rect 7298 8988 7308 9044
rect 7364 8988 8092 9044
rect 8148 8988 9660 9044
rect 9716 8988 9726 9044
rect 15138 8988 15148 9044
rect 15204 8988 15372 9044
rect 15428 8988 15438 9044
rect 2482 8876 2492 8932
rect 2548 8876 26236 8932
rect 26292 8876 26302 8932
rect 27010 8876 27020 8932
rect 27076 8876 28252 8932
rect 28308 8876 28318 8932
rect 28448 8820 28560 8848
rect 27570 8764 27580 8820
rect 27636 8764 28560 8820
rect 28448 8736 28560 8764
rect 4454 8596 4464 8652
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4728 8596 4738 8652
rect 24454 8596 24464 8652
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24728 8596 24738 8652
rect 28448 8372 28560 8400
rect 26674 8316 26684 8372
rect 26740 8316 28560 8372
rect 28448 8288 28560 8316
rect 802 8204 812 8260
rect 868 8204 1596 8260
rect 1652 8204 1662 8260
rect 8306 8092 8316 8148
rect 8372 8092 26124 8148
rect 26180 8092 26190 8148
rect 13570 7980 13580 8036
rect 13636 7980 26908 8036
rect 26964 7980 26974 8036
rect 0 7924 112 7952
rect 28448 7924 28560 7952
rect 0 7868 1036 7924
rect 1092 7868 1102 7924
rect 27458 7868 27468 7924
rect 27524 7868 28560 7924
rect 0 7840 112 7868
rect 3794 7812 3804 7868
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 4068 7812 4078 7868
rect 23794 7812 23804 7868
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 24068 7812 24078 7868
rect 28448 7840 28560 7868
rect 10658 7644 10668 7700
rect 10724 7644 26796 7700
rect 26852 7644 26862 7700
rect 11554 7532 11564 7588
rect 11620 7532 19292 7588
rect 19348 7532 19358 7588
rect 26562 7532 26572 7588
rect 26628 7532 27636 7588
rect 27580 7476 27636 7532
rect 28448 7476 28560 7504
rect 12786 7420 12796 7476
rect 12852 7420 26908 7476
rect 26964 7420 26974 7476
rect 27580 7420 28560 7476
rect 28448 7392 28560 7420
rect 4454 7028 4464 7084
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4728 7028 4738 7084
rect 24454 7028 24464 7084
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 24728 7028 24738 7084
rect 28448 7028 28560 7056
rect 27458 6972 27468 7028
rect 27524 6972 28560 7028
rect 28448 6944 28560 6972
rect 23426 6748 23436 6804
rect 23492 6748 26236 6804
rect 26292 6748 26302 6804
rect 26898 6636 26908 6692
rect 26964 6636 27244 6692
rect 27300 6636 27310 6692
rect 0 6580 112 6608
rect 28448 6580 28560 6608
rect 0 6524 1260 6580
rect 1316 6524 1326 6580
rect 15810 6524 15820 6580
rect 15876 6524 26012 6580
rect 26068 6524 26078 6580
rect 27458 6524 27468 6580
rect 27524 6524 28560 6580
rect 0 6496 112 6524
rect 28448 6496 28560 6524
rect 3794 6244 3804 6300
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 4068 6244 4078 6300
rect 23794 6244 23804 6300
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 24068 6244 24078 6300
rect 28448 6132 28560 6160
rect 26562 6076 26572 6132
rect 26628 6076 28560 6132
rect 28448 6048 28560 6076
rect 14578 5964 14588 6020
rect 14644 5964 27188 6020
rect 27132 5796 27188 5964
rect 15138 5740 15148 5796
rect 15204 5740 26012 5796
rect 26068 5740 26078 5796
rect 27122 5740 27132 5796
rect 27188 5740 27198 5796
rect 28448 5684 28560 5712
rect 27570 5628 27580 5684
rect 27636 5628 28560 5684
rect 28448 5600 28560 5628
rect 4454 5460 4464 5516
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4728 5460 4738 5516
rect 24454 5460 24464 5516
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24728 5460 24738 5516
rect 0 5236 112 5264
rect 28448 5236 28560 5264
rect 0 5180 1260 5236
rect 1316 5180 1326 5236
rect 10098 5180 10108 5236
rect 10164 5180 19964 5236
rect 20020 5180 20030 5236
rect 26674 5180 26684 5236
rect 26740 5180 28560 5236
rect 0 5152 112 5180
rect 28448 5152 28560 5180
rect 12786 5068 12796 5124
rect 12852 5068 19628 5124
rect 19684 5068 19694 5124
rect 21522 5068 21532 5124
rect 21588 5068 26796 5124
rect 26852 5068 26862 5124
rect 20738 4844 20748 4900
rect 20804 4844 26460 4900
rect 26516 4844 26526 4900
rect 28448 4788 28560 4816
rect 27458 4732 27468 4788
rect 27524 4732 28560 4788
rect 3794 4676 3804 4732
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 4068 4676 4078 4732
rect 23794 4676 23804 4732
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 24068 4676 24078 4732
rect 28448 4704 28560 4732
rect 466 4396 476 4452
rect 532 4396 1484 4452
rect 1540 4396 1550 4452
rect 14690 4396 14700 4452
rect 14756 4396 26908 4452
rect 26964 4396 26974 4452
rect 28448 4340 28560 4368
rect 26562 4284 26572 4340
rect 26628 4284 28560 4340
rect 28448 4256 28560 4284
rect 16818 4172 16828 4228
rect 16884 4172 27356 4228
rect 27412 4172 27422 4228
rect 0 3892 112 3920
rect 4454 3892 4464 3948
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4728 3892 4738 3948
rect 24454 3892 24464 3948
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24728 3892 24738 3948
rect 28448 3892 28560 3920
rect 0 3836 1036 3892
rect 1092 3836 1102 3892
rect 27458 3836 27468 3892
rect 27524 3836 28560 3892
rect 0 3808 112 3836
rect 28448 3808 28560 3836
rect 26908 3500 27916 3556
rect 27972 3500 27982 3556
rect 26908 3444 26964 3500
rect 28448 3444 28560 3472
rect 13346 3388 13356 3444
rect 13412 3388 26012 3444
rect 26068 3388 26078 3444
rect 26898 3388 26908 3444
rect 26964 3388 26974 3444
rect 27458 3388 27468 3444
rect 27524 3388 28560 3444
rect 28448 3360 28560 3388
rect 20850 3276 20860 3332
rect 20916 3276 27692 3332
rect 27748 3276 27758 3332
rect 3794 3108 3804 3164
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 4068 3108 4078 3164
rect 23794 3108 23804 3164
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 24068 3108 24078 3164
rect 28448 2996 28560 3024
rect 26562 2940 26572 2996
rect 26628 2940 28560 2996
rect 28448 2912 28560 2940
rect 21186 2828 21196 2884
rect 21252 2828 26012 2884
rect 26068 2828 26078 2884
rect 26898 2828 26908 2884
rect 26964 2828 27804 2884
rect 27860 2828 27870 2884
rect 1138 2716 1148 2772
rect 1204 2716 3388 2772
rect 3444 2716 3454 2772
rect 28448 2548 28560 2576
rect 27570 2492 27580 2548
rect 27636 2492 28560 2548
rect 28448 2464 28560 2492
rect 4454 2324 4464 2380
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4728 2324 4738 2380
rect 24454 2324 24464 2380
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24728 2324 24738 2380
rect 28448 2100 28560 2128
rect 26674 2044 26684 2100
rect 26740 2044 28560 2100
rect 28448 2016 28560 2044
rect 28448 1652 28560 1680
rect 7410 1596 7420 1652
rect 7476 1596 8988 1652
rect 9044 1596 9054 1652
rect 22418 1596 22428 1652
rect 22484 1596 23548 1652
rect 23604 1596 23614 1652
rect 26562 1596 26572 1652
rect 26628 1596 28560 1652
rect 3794 1540 3804 1596
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 4068 1540 4078 1596
rect 23794 1540 23804 1596
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 24068 1540 24078 1596
rect 28448 1568 28560 1596
rect 24882 1484 24892 1540
rect 24948 1484 28140 1540
rect 28196 1484 28206 1540
rect 2034 1372 2044 1428
rect 2100 1372 7084 1428
rect 7140 1372 7150 1428
rect 28448 1204 28560 1232
rect 15474 1148 15484 1204
rect 15540 1148 24780 1204
rect 24836 1148 24846 1204
rect 27122 1148 27132 1204
rect 27188 1148 28560 1204
rect 28448 1120 28560 1148
rect 6850 1036 6860 1092
rect 6916 1036 17164 1092
rect 17220 1036 17230 1092
rect 18610 1036 18620 1092
rect 18676 1036 25676 1092
rect 25732 1036 25742 1092
rect 14130 924 14140 980
rect 14196 924 22764 980
rect 22820 924 22830 980
rect 4454 756 4464 812
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4728 756 4738 812
rect 24454 756 24464 812
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24728 756 24738 812
rect 28448 756 28560 784
rect 25330 700 25340 756
rect 25396 700 28560 756
rect 28448 672 28560 700
rect 15474 588 15484 644
rect 15540 588 20300 644
rect 20356 588 20366 644
rect 28448 308 28560 336
rect 26114 252 26124 308
rect 26180 252 28560 308
rect 28448 224 28560 252
rect 4722 140 4732 196
rect 4788 140 4956 196
rect 5012 140 5022 196
rect 26786 140 26796 196
rect 26852 140 27580 196
rect 27636 140 27646 196
<< via3 >>
rect 3804 56420 3860 56476
rect 3908 56420 3964 56476
rect 4012 56420 4068 56476
rect 23804 56420 23860 56476
rect 23908 56420 23964 56476
rect 24012 56420 24068 56476
rect 2492 55916 2548 55972
rect 4464 55636 4520 55692
rect 4568 55636 4624 55692
rect 4672 55636 4728 55692
rect 24464 55636 24520 55692
rect 24568 55636 24624 55692
rect 24672 55636 24728 55692
rect 3804 54852 3860 54908
rect 3908 54852 3964 54908
rect 4012 54852 4068 54908
rect 23804 54852 23860 54908
rect 23908 54852 23964 54908
rect 24012 54852 24068 54908
rect 4464 54068 4520 54124
rect 4568 54068 4624 54124
rect 4672 54068 4728 54124
rect 24464 54068 24520 54124
rect 24568 54068 24624 54124
rect 24672 54068 24728 54124
rect 26236 53676 26292 53732
rect 3804 53284 3860 53340
rect 3908 53284 3964 53340
rect 4012 53284 4068 53340
rect 23804 53284 23860 53340
rect 23908 53284 23964 53340
rect 24012 53284 24068 53340
rect 25228 52780 25284 52836
rect 4464 52500 4520 52556
rect 4568 52500 4624 52556
rect 4672 52500 4728 52556
rect 24464 52500 24520 52556
rect 24568 52500 24624 52556
rect 24672 52500 24728 52556
rect 3804 51716 3860 51772
rect 3908 51716 3964 51772
rect 4012 51716 4068 51772
rect 23804 51716 23860 51772
rect 23908 51716 23964 51772
rect 24012 51716 24068 51772
rect 12572 51100 12628 51156
rect 4464 50932 4520 50988
rect 4568 50932 4624 50988
rect 4672 50932 4728 50988
rect 24464 50932 24520 50988
rect 24568 50932 24624 50988
rect 24672 50932 24728 50988
rect 3804 50148 3860 50204
rect 3908 50148 3964 50204
rect 4012 50148 4068 50204
rect 23804 50148 23860 50204
rect 23908 50148 23964 50204
rect 24012 50148 24068 50204
rect 4464 49364 4520 49420
rect 4568 49364 4624 49420
rect 4672 49364 4728 49420
rect 24464 49364 24520 49420
rect 24568 49364 24624 49420
rect 24672 49364 24728 49420
rect 11676 48748 11732 48804
rect 3804 48580 3860 48636
rect 3908 48580 3964 48636
rect 4012 48580 4068 48636
rect 23804 48580 23860 48636
rect 23908 48580 23964 48636
rect 24012 48580 24068 48636
rect 4464 47796 4520 47852
rect 4568 47796 4624 47852
rect 4672 47796 4728 47852
rect 24464 47796 24520 47852
rect 24568 47796 24624 47852
rect 24672 47796 24728 47852
rect 3804 47012 3860 47068
rect 3908 47012 3964 47068
rect 4012 47012 4068 47068
rect 23804 47012 23860 47068
rect 23908 47012 23964 47068
rect 24012 47012 24068 47068
rect 26124 46508 26180 46564
rect 4464 46228 4520 46284
rect 4568 46228 4624 46284
rect 4672 46228 4728 46284
rect 24464 46228 24520 46284
rect 24568 46228 24624 46284
rect 24672 46228 24728 46284
rect 1484 45724 1540 45780
rect 3804 45444 3860 45500
rect 3908 45444 3964 45500
rect 4012 45444 4068 45500
rect 23804 45444 23860 45500
rect 23908 45444 23964 45500
rect 24012 45444 24068 45500
rect 4464 44660 4520 44716
rect 4568 44660 4624 44716
rect 4672 44660 4728 44716
rect 24464 44660 24520 44716
rect 24568 44660 24624 44716
rect 24672 44660 24728 44716
rect 4844 44268 4900 44324
rect 3804 43876 3860 43932
rect 3908 43876 3964 43932
rect 4012 43876 4068 43932
rect 23804 43876 23860 43932
rect 23908 43876 23964 43932
rect 24012 43876 24068 43932
rect 1596 43372 1652 43428
rect 4464 43092 4520 43148
rect 4568 43092 4624 43148
rect 4672 43092 4728 43148
rect 24464 43092 24520 43148
rect 24568 43092 24624 43148
rect 24672 43092 24728 43148
rect 3804 42308 3860 42364
rect 3908 42308 3964 42364
rect 4012 42308 4068 42364
rect 23804 42308 23860 42364
rect 23908 42308 23964 42364
rect 24012 42308 24068 42364
rect 4464 41524 4520 41580
rect 4568 41524 4624 41580
rect 4672 41524 4728 41580
rect 24464 41524 24520 41580
rect 24568 41524 24624 41580
rect 24672 41524 24728 41580
rect 3804 40740 3860 40796
rect 3908 40740 3964 40796
rect 4012 40740 4068 40796
rect 23804 40740 23860 40796
rect 23908 40740 23964 40796
rect 24012 40740 24068 40796
rect 4464 39956 4520 40012
rect 4568 39956 4624 40012
rect 4672 39956 4728 40012
rect 24464 39956 24520 40012
rect 24568 39956 24624 40012
rect 24672 39956 24728 40012
rect 11228 39452 11284 39508
rect 3804 39172 3860 39228
rect 3908 39172 3964 39228
rect 4012 39172 4068 39228
rect 23804 39172 23860 39228
rect 23908 39172 23964 39228
rect 24012 39172 24068 39228
rect 4464 38388 4520 38444
rect 4568 38388 4624 38444
rect 4672 38388 4728 38444
rect 24464 38388 24520 38444
rect 24568 38388 24624 38444
rect 24672 38388 24728 38444
rect 1484 38220 1540 38276
rect 9436 37996 9492 38052
rect 1596 37884 1652 37940
rect 3804 37604 3860 37660
rect 3908 37604 3964 37660
rect 4012 37604 4068 37660
rect 23804 37604 23860 37660
rect 23908 37604 23964 37660
rect 24012 37604 24068 37660
rect 4464 36820 4520 36876
rect 4568 36820 4624 36876
rect 4672 36820 4728 36876
rect 24464 36820 24520 36876
rect 24568 36820 24624 36876
rect 24672 36820 24728 36876
rect 9212 36092 9268 36148
rect 3804 36036 3860 36092
rect 3908 36036 3964 36092
rect 4012 36036 4068 36092
rect 23804 36036 23860 36092
rect 23908 36036 23964 36092
rect 24012 36036 24068 36092
rect 9212 35532 9268 35588
rect 9436 35420 9492 35476
rect 25340 35420 25396 35476
rect 4464 35252 4520 35308
rect 4568 35252 4624 35308
rect 4672 35252 4728 35308
rect 24464 35252 24520 35308
rect 24568 35252 24624 35308
rect 24672 35252 24728 35308
rect 3804 34468 3860 34524
rect 3908 34468 3964 34524
rect 4012 34468 4068 34524
rect 23804 34468 23860 34524
rect 23908 34468 23964 34524
rect 24012 34468 24068 34524
rect 8204 33740 8260 33796
rect 4464 33684 4520 33740
rect 4568 33684 4624 33740
rect 4672 33684 4728 33740
rect 24464 33684 24520 33740
rect 24568 33684 24624 33740
rect 24672 33684 24728 33740
rect 19404 33068 19460 33124
rect 3804 32900 3860 32956
rect 3908 32900 3964 32956
rect 4012 32900 4068 32956
rect 23804 32900 23860 32956
rect 23908 32900 23964 32956
rect 24012 32900 24068 32956
rect 19404 32508 19460 32564
rect 8204 32396 8260 32452
rect 4464 32116 4520 32172
rect 4568 32116 4624 32172
rect 4672 32116 4728 32172
rect 24464 32116 24520 32172
rect 24568 32116 24624 32172
rect 24672 32116 24728 32172
rect 3612 31500 3668 31556
rect 3804 31332 3860 31388
rect 3908 31332 3964 31388
rect 4012 31332 4068 31388
rect 23804 31332 23860 31388
rect 23908 31332 23964 31388
rect 24012 31332 24068 31388
rect 7084 30716 7140 30772
rect 4464 30548 4520 30604
rect 4568 30548 4624 30604
rect 4672 30548 4728 30604
rect 24464 30548 24520 30604
rect 24568 30548 24624 30604
rect 24672 30548 24728 30604
rect 3804 29764 3860 29820
rect 3908 29764 3964 29820
rect 4012 29764 4068 29820
rect 23804 29764 23860 29820
rect 23908 29764 23964 29820
rect 24012 29764 24068 29820
rect 3612 29484 3668 29540
rect 4464 28980 4520 29036
rect 4568 28980 4624 29036
rect 4672 28980 4728 29036
rect 24464 28980 24520 29036
rect 24568 28980 24624 29036
rect 24672 28980 24728 29036
rect 3804 28196 3860 28252
rect 3908 28196 3964 28252
rect 4012 28196 4068 28252
rect 23804 28196 23860 28252
rect 23908 28196 23964 28252
rect 24012 28196 24068 28252
rect 18396 28028 18452 28084
rect 11004 27804 11060 27860
rect 3164 27692 3220 27748
rect 11452 27468 11508 27524
rect 4464 27412 4520 27468
rect 4568 27412 4624 27468
rect 4672 27412 4728 27468
rect 24464 27412 24520 27468
rect 24568 27412 24624 27468
rect 24672 27412 24728 27468
rect 17388 27020 17444 27076
rect 17388 26796 17444 26852
rect 3804 26628 3860 26684
rect 3908 26628 3964 26684
rect 4012 26628 4068 26684
rect 23804 26628 23860 26684
rect 23908 26628 23964 26684
rect 24012 26628 24068 26684
rect 11452 26460 11508 26516
rect 4464 25844 4520 25900
rect 4568 25844 4624 25900
rect 4672 25844 4728 25900
rect 24464 25844 24520 25900
rect 24568 25844 24624 25900
rect 24672 25844 24728 25900
rect 26012 25452 26068 25508
rect 3804 25060 3860 25116
rect 3908 25060 3964 25116
rect 4012 25060 4068 25116
rect 23804 25060 23860 25116
rect 23908 25060 23964 25116
rect 24012 25060 24068 25116
rect 1372 24780 1428 24836
rect 6188 24556 6244 24612
rect 10556 24444 10612 24500
rect 4464 24276 4520 24332
rect 4568 24276 4624 24332
rect 4672 24276 4728 24332
rect 24464 24276 24520 24332
rect 24568 24276 24624 24332
rect 24672 24276 24728 24332
rect 10556 24220 10612 24276
rect 3804 23492 3860 23548
rect 3908 23492 3964 23548
rect 4012 23492 4068 23548
rect 23804 23492 23860 23548
rect 23908 23492 23964 23548
rect 24012 23492 24068 23548
rect 7196 23212 7252 23268
rect 12012 23212 12068 23268
rect 4464 22708 4520 22764
rect 4568 22708 4624 22764
rect 4672 22708 4728 22764
rect 24464 22708 24520 22764
rect 24568 22708 24624 22764
rect 24672 22708 24728 22764
rect 3804 21924 3860 21980
rect 3908 21924 3964 21980
rect 4012 21924 4068 21980
rect 23804 21924 23860 21980
rect 23908 21924 23964 21980
rect 24012 21924 24068 21980
rect 3052 21868 3108 21924
rect 12012 21868 12068 21924
rect 6972 21532 7028 21588
rect 4464 21140 4520 21196
rect 4568 21140 4624 21196
rect 4672 21140 4728 21196
rect 24464 21140 24520 21196
rect 24568 21140 24624 21196
rect 24672 21140 24728 21196
rect 1372 20860 1428 20916
rect 7196 20748 7252 20804
rect 3612 20636 3668 20692
rect 3804 20356 3860 20412
rect 3908 20356 3964 20412
rect 4012 20356 4068 20412
rect 23804 20356 23860 20412
rect 23908 20356 23964 20412
rect 24012 20356 24068 20412
rect 6188 20076 6244 20132
rect 4464 19572 4520 19628
rect 4568 19572 4624 19628
rect 4672 19572 4728 19628
rect 24464 19572 24520 19628
rect 24568 19572 24624 19628
rect 24672 19572 24728 19628
rect 3804 18788 3860 18844
rect 3908 18788 3964 18844
rect 4012 18788 4068 18844
rect 23804 18788 23860 18844
rect 23908 18788 23964 18844
rect 24012 18788 24068 18844
rect 3276 18508 3332 18564
rect 15260 18508 15316 18564
rect 3164 18396 3220 18452
rect 4844 18396 4900 18452
rect 14588 18060 14644 18116
rect 4464 18004 4520 18060
rect 4568 18004 4624 18060
rect 4672 18004 4728 18060
rect 24464 18004 24520 18060
rect 24568 18004 24624 18060
rect 24672 18004 24728 18060
rect 14700 17948 14756 18004
rect 700 17836 756 17892
rect 18396 17836 18452 17892
rect 14700 17724 14756 17780
rect 700 17388 756 17444
rect 1932 17276 1988 17332
rect 3804 17220 3860 17276
rect 3908 17220 3964 17276
rect 4012 17220 4068 17276
rect 23804 17220 23860 17276
rect 23908 17220 23964 17276
rect 24012 17220 24068 17276
rect 11788 17164 11844 17220
rect 3276 16940 3332 16996
rect 3612 16828 3668 16884
rect 4464 16436 4520 16492
rect 4568 16436 4624 16492
rect 4672 16436 4728 16492
rect 14588 16380 14644 16436
rect 24464 16436 24520 16492
rect 24568 16436 24624 16492
rect 24672 16436 24728 16492
rect 3052 16044 3108 16100
rect 3804 15652 3860 15708
rect 3908 15652 3964 15708
rect 4012 15652 4068 15708
rect 23804 15652 23860 15708
rect 23908 15652 23964 15708
rect 24012 15652 24068 15708
rect 3052 15484 3108 15540
rect 6972 15036 7028 15092
rect 3052 14924 3108 14980
rect 4464 14868 4520 14924
rect 4568 14868 4624 14924
rect 4672 14868 4728 14924
rect 24464 14868 24520 14924
rect 24568 14868 24624 14924
rect 24672 14868 24728 14924
rect 2492 14588 2548 14644
rect 17052 14588 17108 14644
rect 1148 14364 1204 14420
rect 27580 14364 27636 14420
rect 15260 14252 15316 14308
rect 3804 14084 3860 14140
rect 3908 14084 3964 14140
rect 4012 14084 4068 14140
rect 23804 14084 23860 14140
rect 23908 14084 23964 14140
rect 24012 14084 24068 14140
rect 27580 13804 27636 13860
rect 17052 13692 17108 13748
rect 1148 13580 1204 13636
rect 15260 13356 15316 13412
rect 4464 13300 4520 13356
rect 4568 13300 4624 13356
rect 4672 13300 4728 13356
rect 24464 13300 24520 13356
rect 24568 13300 24624 13356
rect 24672 13300 24728 13356
rect 26012 12796 26068 12852
rect 11788 12684 11844 12740
rect 3804 12516 3860 12572
rect 3908 12516 3964 12572
rect 4012 12516 4068 12572
rect 23804 12516 23860 12572
rect 23908 12516 23964 12572
rect 24012 12516 24068 12572
rect 1932 12124 1988 12180
rect 4464 11732 4520 11788
rect 4568 11732 4624 11788
rect 4672 11732 4728 11788
rect 24464 11732 24520 11788
rect 24568 11732 24624 11788
rect 24672 11732 24728 11788
rect 12572 11564 12628 11620
rect 25340 11564 25396 11620
rect 25228 11452 25284 11508
rect 11676 11116 11732 11172
rect 3804 10948 3860 11004
rect 3908 10948 3964 11004
rect 4012 10948 4068 11004
rect 23804 10948 23860 11004
rect 23908 10948 23964 11004
rect 24012 10948 24068 11004
rect 11004 10668 11060 10724
rect 4464 10164 4520 10220
rect 4568 10164 4624 10220
rect 4672 10164 4728 10220
rect 24464 10164 24520 10220
rect 24568 10164 24624 10220
rect 24672 10164 24728 10220
rect 11228 9660 11284 9716
rect 3804 9380 3860 9436
rect 3908 9380 3964 9436
rect 4012 9380 4068 9436
rect 23804 9380 23860 9436
rect 23908 9380 23964 9436
rect 24012 9380 24068 9436
rect 26236 8876 26292 8932
rect 4464 8596 4520 8652
rect 4568 8596 4624 8652
rect 4672 8596 4728 8652
rect 24464 8596 24520 8652
rect 24568 8596 24624 8652
rect 24672 8596 24728 8652
rect 26124 8092 26180 8148
rect 3804 7812 3860 7868
rect 3908 7812 3964 7868
rect 4012 7812 4068 7868
rect 23804 7812 23860 7868
rect 23908 7812 23964 7868
rect 24012 7812 24068 7868
rect 4464 7028 4520 7084
rect 4568 7028 4624 7084
rect 4672 7028 4728 7084
rect 24464 7028 24520 7084
rect 24568 7028 24624 7084
rect 24672 7028 24728 7084
rect 3804 6244 3860 6300
rect 3908 6244 3964 6300
rect 4012 6244 4068 6300
rect 23804 6244 23860 6300
rect 23908 6244 23964 6300
rect 24012 6244 24068 6300
rect 4464 5460 4520 5516
rect 4568 5460 4624 5516
rect 4672 5460 4728 5516
rect 24464 5460 24520 5516
rect 24568 5460 24624 5516
rect 24672 5460 24728 5516
rect 3804 4676 3860 4732
rect 3908 4676 3964 4732
rect 4012 4676 4068 4732
rect 23804 4676 23860 4732
rect 23908 4676 23964 4732
rect 24012 4676 24068 4732
rect 4464 3892 4520 3948
rect 4568 3892 4624 3948
rect 4672 3892 4728 3948
rect 24464 3892 24520 3948
rect 24568 3892 24624 3948
rect 24672 3892 24728 3948
rect 3804 3108 3860 3164
rect 3908 3108 3964 3164
rect 4012 3108 4068 3164
rect 23804 3108 23860 3164
rect 23908 3108 23964 3164
rect 24012 3108 24068 3164
rect 4464 2324 4520 2380
rect 4568 2324 4624 2380
rect 4672 2324 4728 2380
rect 24464 2324 24520 2380
rect 24568 2324 24624 2380
rect 24672 2324 24728 2380
rect 3804 1540 3860 1596
rect 3908 1540 3964 1596
rect 4012 1540 4068 1596
rect 23804 1540 23860 1596
rect 23908 1540 23964 1596
rect 24012 1540 24068 1596
rect 7084 1372 7140 1428
rect 4464 756 4520 812
rect 4568 756 4624 812
rect 4672 756 4728 812
rect 24464 756 24520 812
rect 24568 756 24624 812
rect 24672 756 24728 812
<< metal4 >>
rect 3776 56476 4096 57456
rect 3776 56420 3804 56476
rect 3860 56420 3908 56476
rect 3964 56420 4012 56476
rect 4068 56420 4096 56476
rect 2492 55972 2548 55982
rect 1484 45780 1540 45790
rect 1484 38276 1540 45724
rect 1484 38210 1540 38220
rect 1596 43428 1652 43438
rect 1596 37940 1652 43372
rect 1596 37874 1652 37884
rect 1372 24836 1428 24846
rect 1372 20916 1428 24780
rect 1372 20850 1428 20860
rect 700 17892 756 17902
rect 700 17444 756 17836
rect 700 17378 756 17388
rect 1932 17332 1988 17342
rect 1148 14420 1204 14430
rect 1148 13636 1204 14364
rect 1148 13570 1204 13580
rect 1932 12180 1988 17276
rect 2492 14644 2548 55916
rect 3776 54908 4096 56420
rect 3776 54852 3804 54908
rect 3860 54852 3908 54908
rect 3964 54852 4012 54908
rect 4068 54852 4096 54908
rect 3776 53340 4096 54852
rect 3776 53284 3804 53340
rect 3860 53284 3908 53340
rect 3964 53284 4012 53340
rect 4068 53284 4096 53340
rect 3776 51772 4096 53284
rect 3776 51716 3804 51772
rect 3860 51716 3908 51772
rect 3964 51716 4012 51772
rect 4068 51716 4096 51772
rect 3776 50204 4096 51716
rect 3776 50148 3804 50204
rect 3860 50148 3908 50204
rect 3964 50148 4012 50204
rect 4068 50148 4096 50204
rect 3776 48636 4096 50148
rect 3776 48580 3804 48636
rect 3860 48580 3908 48636
rect 3964 48580 4012 48636
rect 4068 48580 4096 48636
rect 3776 47068 4096 48580
rect 3776 47012 3804 47068
rect 3860 47012 3908 47068
rect 3964 47012 4012 47068
rect 4068 47012 4096 47068
rect 3776 45500 4096 47012
rect 3776 45444 3804 45500
rect 3860 45444 3908 45500
rect 3964 45444 4012 45500
rect 4068 45444 4096 45500
rect 3776 43932 4096 45444
rect 3776 43876 3804 43932
rect 3860 43876 3908 43932
rect 3964 43876 4012 43932
rect 4068 43876 4096 43932
rect 3776 42364 4096 43876
rect 3776 42308 3804 42364
rect 3860 42308 3908 42364
rect 3964 42308 4012 42364
rect 4068 42308 4096 42364
rect 3776 40796 4096 42308
rect 3776 40740 3804 40796
rect 3860 40740 3908 40796
rect 3964 40740 4012 40796
rect 4068 40740 4096 40796
rect 3776 39228 4096 40740
rect 3776 39172 3804 39228
rect 3860 39172 3908 39228
rect 3964 39172 4012 39228
rect 4068 39172 4096 39228
rect 3776 37660 4096 39172
rect 3776 37604 3804 37660
rect 3860 37604 3908 37660
rect 3964 37604 4012 37660
rect 4068 37604 4096 37660
rect 3776 36092 4096 37604
rect 3776 36036 3804 36092
rect 3860 36036 3908 36092
rect 3964 36036 4012 36092
rect 4068 36036 4096 36092
rect 3776 34524 4096 36036
rect 3776 34468 3804 34524
rect 3860 34468 3908 34524
rect 3964 34468 4012 34524
rect 4068 34468 4096 34524
rect 3776 32956 4096 34468
rect 3776 32900 3804 32956
rect 3860 32900 3908 32956
rect 3964 32900 4012 32956
rect 4068 32900 4096 32956
rect 3612 31556 3668 31566
rect 3612 29540 3668 31500
rect 3612 29474 3668 29484
rect 3776 31388 4096 32900
rect 3776 31332 3804 31388
rect 3860 31332 3908 31388
rect 3964 31332 4012 31388
rect 4068 31332 4096 31388
rect 3776 29820 4096 31332
rect 3776 29764 3804 29820
rect 3860 29764 3908 29820
rect 3964 29764 4012 29820
rect 4068 29764 4096 29820
rect 3776 28252 4096 29764
rect 3776 28196 3804 28252
rect 3860 28196 3908 28252
rect 3964 28196 4012 28252
rect 4068 28196 4096 28252
rect 3164 27748 3220 27758
rect 3052 21924 3108 21934
rect 3052 16100 3108 21868
rect 3164 18452 3220 27692
rect 3776 26684 4096 28196
rect 3776 26628 3804 26684
rect 3860 26628 3908 26684
rect 3964 26628 4012 26684
rect 4068 26628 4096 26684
rect 3776 25116 4096 26628
rect 3776 25060 3804 25116
rect 3860 25060 3908 25116
rect 3964 25060 4012 25116
rect 4068 25060 4096 25116
rect 3776 23548 4096 25060
rect 3776 23492 3804 23548
rect 3860 23492 3908 23548
rect 3964 23492 4012 23548
rect 4068 23492 4096 23548
rect 3776 21980 4096 23492
rect 3776 21924 3804 21980
rect 3860 21924 3908 21980
rect 3964 21924 4012 21980
rect 4068 21924 4096 21980
rect 3612 20692 3668 20702
rect 3164 18386 3220 18396
rect 3276 18564 3332 18574
rect 3276 16996 3332 18508
rect 3276 16930 3332 16940
rect 3612 16884 3668 20636
rect 3612 16818 3668 16828
rect 3776 20412 4096 21924
rect 3776 20356 3804 20412
rect 3860 20356 3908 20412
rect 3964 20356 4012 20412
rect 4068 20356 4096 20412
rect 3776 18844 4096 20356
rect 3776 18788 3804 18844
rect 3860 18788 3908 18844
rect 3964 18788 4012 18844
rect 4068 18788 4096 18844
rect 3776 17276 4096 18788
rect 3776 17220 3804 17276
rect 3860 17220 3908 17276
rect 3964 17220 4012 17276
rect 4068 17220 4096 17276
rect 3052 16034 3108 16044
rect 3776 15708 4096 17220
rect 3776 15652 3804 15708
rect 3860 15652 3908 15708
rect 3964 15652 4012 15708
rect 4068 15652 4096 15708
rect 3052 15540 3108 15550
rect 3052 14980 3108 15484
rect 3052 14914 3108 14924
rect 2492 14578 2548 14588
rect 1932 12114 1988 12124
rect 3776 14140 4096 15652
rect 3776 14084 3804 14140
rect 3860 14084 3908 14140
rect 3964 14084 4012 14140
rect 4068 14084 4096 14140
rect 3776 12572 4096 14084
rect 3776 12516 3804 12572
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 4068 12516 4096 12572
rect 3776 11004 4096 12516
rect 3776 10948 3804 11004
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 4068 10948 4096 11004
rect 3776 9436 4096 10948
rect 3776 9380 3804 9436
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 4068 9380 4096 9436
rect 3776 7868 4096 9380
rect 3776 7812 3804 7868
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 4068 7812 4096 7868
rect 3776 6300 4096 7812
rect 3776 6244 3804 6300
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 4068 6244 4096 6300
rect 3776 4732 4096 6244
rect 3776 4676 3804 4732
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 4068 4676 4096 4732
rect 3776 3164 4096 4676
rect 3776 3108 3804 3164
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 4068 3108 4096 3164
rect 3776 1596 4096 3108
rect 3776 1540 3804 1596
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 4068 1540 4096 1596
rect 3776 0 4096 1540
rect 4436 55692 4756 57456
rect 4436 55636 4464 55692
rect 4520 55636 4568 55692
rect 4624 55636 4672 55692
rect 4728 55636 4756 55692
rect 4436 54124 4756 55636
rect 4436 54068 4464 54124
rect 4520 54068 4568 54124
rect 4624 54068 4672 54124
rect 4728 54068 4756 54124
rect 4436 52556 4756 54068
rect 4436 52500 4464 52556
rect 4520 52500 4568 52556
rect 4624 52500 4672 52556
rect 4728 52500 4756 52556
rect 4436 50988 4756 52500
rect 23776 56476 24096 57456
rect 23776 56420 23804 56476
rect 23860 56420 23908 56476
rect 23964 56420 24012 56476
rect 24068 56420 24096 56476
rect 23776 54908 24096 56420
rect 23776 54852 23804 54908
rect 23860 54852 23908 54908
rect 23964 54852 24012 54908
rect 24068 54852 24096 54908
rect 23776 53340 24096 54852
rect 23776 53284 23804 53340
rect 23860 53284 23908 53340
rect 23964 53284 24012 53340
rect 24068 53284 24096 53340
rect 23776 51772 24096 53284
rect 23776 51716 23804 51772
rect 23860 51716 23908 51772
rect 23964 51716 24012 51772
rect 24068 51716 24096 51772
rect 4436 50932 4464 50988
rect 4520 50932 4568 50988
rect 4624 50932 4672 50988
rect 4728 50932 4756 50988
rect 4436 49420 4756 50932
rect 4436 49364 4464 49420
rect 4520 49364 4568 49420
rect 4624 49364 4672 49420
rect 4728 49364 4756 49420
rect 4436 47852 4756 49364
rect 12572 51156 12628 51166
rect 4436 47796 4464 47852
rect 4520 47796 4568 47852
rect 4624 47796 4672 47852
rect 4728 47796 4756 47852
rect 4436 46284 4756 47796
rect 4436 46228 4464 46284
rect 4520 46228 4568 46284
rect 4624 46228 4672 46284
rect 4728 46228 4756 46284
rect 4436 44716 4756 46228
rect 4436 44660 4464 44716
rect 4520 44660 4568 44716
rect 4624 44660 4672 44716
rect 4728 44660 4756 44716
rect 4436 43148 4756 44660
rect 11676 48804 11732 48814
rect 4436 43092 4464 43148
rect 4520 43092 4568 43148
rect 4624 43092 4672 43148
rect 4728 43092 4756 43148
rect 4436 41580 4756 43092
rect 4436 41524 4464 41580
rect 4520 41524 4568 41580
rect 4624 41524 4672 41580
rect 4728 41524 4756 41580
rect 4436 40012 4756 41524
rect 4436 39956 4464 40012
rect 4520 39956 4568 40012
rect 4624 39956 4672 40012
rect 4728 39956 4756 40012
rect 4436 38444 4756 39956
rect 4436 38388 4464 38444
rect 4520 38388 4568 38444
rect 4624 38388 4672 38444
rect 4728 38388 4756 38444
rect 4436 36876 4756 38388
rect 4436 36820 4464 36876
rect 4520 36820 4568 36876
rect 4624 36820 4672 36876
rect 4728 36820 4756 36876
rect 4436 35308 4756 36820
rect 4436 35252 4464 35308
rect 4520 35252 4568 35308
rect 4624 35252 4672 35308
rect 4728 35252 4756 35308
rect 4436 33740 4756 35252
rect 4436 33684 4464 33740
rect 4520 33684 4568 33740
rect 4624 33684 4672 33740
rect 4728 33684 4756 33740
rect 4436 32172 4756 33684
rect 4436 32116 4464 32172
rect 4520 32116 4568 32172
rect 4624 32116 4672 32172
rect 4728 32116 4756 32172
rect 4436 30604 4756 32116
rect 4436 30548 4464 30604
rect 4520 30548 4568 30604
rect 4624 30548 4672 30604
rect 4728 30548 4756 30604
rect 4436 29036 4756 30548
rect 4436 28980 4464 29036
rect 4520 28980 4568 29036
rect 4624 28980 4672 29036
rect 4728 28980 4756 29036
rect 4436 27468 4756 28980
rect 4436 27412 4464 27468
rect 4520 27412 4568 27468
rect 4624 27412 4672 27468
rect 4728 27412 4756 27468
rect 4436 25900 4756 27412
rect 4436 25844 4464 25900
rect 4520 25844 4568 25900
rect 4624 25844 4672 25900
rect 4728 25844 4756 25900
rect 4436 24332 4756 25844
rect 4436 24276 4464 24332
rect 4520 24276 4568 24332
rect 4624 24276 4672 24332
rect 4728 24276 4756 24332
rect 4436 22764 4756 24276
rect 4436 22708 4464 22764
rect 4520 22708 4568 22764
rect 4624 22708 4672 22764
rect 4728 22708 4756 22764
rect 4436 21196 4756 22708
rect 4436 21140 4464 21196
rect 4520 21140 4568 21196
rect 4624 21140 4672 21196
rect 4728 21140 4756 21196
rect 4436 19628 4756 21140
rect 4436 19572 4464 19628
rect 4520 19572 4568 19628
rect 4624 19572 4672 19628
rect 4728 19572 4756 19628
rect 4436 18060 4756 19572
rect 4844 44324 4900 44334
rect 4844 18452 4900 44268
rect 11228 39508 11284 39518
rect 9436 38052 9492 38062
rect 9212 36148 9268 36158
rect 9212 35588 9268 36092
rect 9212 35522 9268 35532
rect 9436 35476 9492 37996
rect 9436 35410 9492 35420
rect 8204 33796 8260 33806
rect 8204 32452 8260 33740
rect 8204 32386 8260 32396
rect 7084 30772 7140 30782
rect 6188 24612 6244 24622
rect 6188 20132 6244 24556
rect 6188 20066 6244 20076
rect 6972 21588 7028 21598
rect 4844 18386 4900 18396
rect 4436 18004 4464 18060
rect 4520 18004 4568 18060
rect 4624 18004 4672 18060
rect 4728 18004 4756 18060
rect 4436 16492 4756 18004
rect 4436 16436 4464 16492
rect 4520 16436 4568 16492
rect 4624 16436 4672 16492
rect 4728 16436 4756 16492
rect 4436 14924 4756 16436
rect 6972 15092 7028 21532
rect 6972 15026 7028 15036
rect 4436 14868 4464 14924
rect 4520 14868 4568 14924
rect 4624 14868 4672 14924
rect 4728 14868 4756 14924
rect 4436 13356 4756 14868
rect 4436 13300 4464 13356
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4728 13300 4756 13356
rect 4436 11788 4756 13300
rect 4436 11732 4464 11788
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4728 11732 4756 11788
rect 4436 10220 4756 11732
rect 4436 10164 4464 10220
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4728 10164 4756 10220
rect 4436 8652 4756 10164
rect 4436 8596 4464 8652
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4728 8596 4756 8652
rect 4436 7084 4756 8596
rect 4436 7028 4464 7084
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4728 7028 4756 7084
rect 4436 5516 4756 7028
rect 4436 5460 4464 5516
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4728 5460 4756 5516
rect 4436 3948 4756 5460
rect 4436 3892 4464 3948
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4728 3892 4756 3948
rect 4436 2380 4756 3892
rect 4436 2324 4464 2380
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4728 2324 4756 2380
rect 4436 812 4756 2324
rect 7084 1428 7140 30716
rect 11004 27860 11060 27870
rect 10556 24500 10612 24510
rect 10556 24276 10612 24444
rect 10556 24210 10612 24220
rect 7196 23268 7252 23278
rect 7196 20804 7252 23212
rect 7196 20738 7252 20748
rect 11004 10724 11060 27804
rect 11004 10658 11060 10668
rect 11228 9716 11284 39452
rect 11452 27524 11508 27534
rect 11452 26516 11508 27468
rect 11452 26450 11508 26460
rect 11676 11172 11732 48748
rect 12012 23268 12068 23278
rect 12012 21924 12068 23212
rect 12012 21858 12068 21868
rect 11788 17220 11844 17230
rect 11788 12740 11844 17164
rect 11788 12674 11844 12684
rect 12572 11620 12628 51100
rect 23776 50204 24096 51716
rect 23776 50148 23804 50204
rect 23860 50148 23908 50204
rect 23964 50148 24012 50204
rect 24068 50148 24096 50204
rect 23776 48636 24096 50148
rect 23776 48580 23804 48636
rect 23860 48580 23908 48636
rect 23964 48580 24012 48636
rect 24068 48580 24096 48636
rect 23776 47068 24096 48580
rect 23776 47012 23804 47068
rect 23860 47012 23908 47068
rect 23964 47012 24012 47068
rect 24068 47012 24096 47068
rect 23776 45500 24096 47012
rect 23776 45444 23804 45500
rect 23860 45444 23908 45500
rect 23964 45444 24012 45500
rect 24068 45444 24096 45500
rect 23776 43932 24096 45444
rect 23776 43876 23804 43932
rect 23860 43876 23908 43932
rect 23964 43876 24012 43932
rect 24068 43876 24096 43932
rect 23776 42364 24096 43876
rect 23776 42308 23804 42364
rect 23860 42308 23908 42364
rect 23964 42308 24012 42364
rect 24068 42308 24096 42364
rect 23776 40796 24096 42308
rect 23776 40740 23804 40796
rect 23860 40740 23908 40796
rect 23964 40740 24012 40796
rect 24068 40740 24096 40796
rect 23776 39228 24096 40740
rect 23776 39172 23804 39228
rect 23860 39172 23908 39228
rect 23964 39172 24012 39228
rect 24068 39172 24096 39228
rect 23776 37660 24096 39172
rect 23776 37604 23804 37660
rect 23860 37604 23908 37660
rect 23964 37604 24012 37660
rect 24068 37604 24096 37660
rect 23776 36092 24096 37604
rect 23776 36036 23804 36092
rect 23860 36036 23908 36092
rect 23964 36036 24012 36092
rect 24068 36036 24096 36092
rect 23776 34524 24096 36036
rect 23776 34468 23804 34524
rect 23860 34468 23908 34524
rect 23964 34468 24012 34524
rect 24068 34468 24096 34524
rect 19404 33124 19460 33134
rect 19404 32564 19460 33068
rect 19404 32498 19460 32508
rect 23776 32956 24096 34468
rect 23776 32900 23804 32956
rect 23860 32900 23908 32956
rect 23964 32900 24012 32956
rect 24068 32900 24096 32956
rect 23776 31388 24096 32900
rect 23776 31332 23804 31388
rect 23860 31332 23908 31388
rect 23964 31332 24012 31388
rect 24068 31332 24096 31388
rect 23776 29820 24096 31332
rect 23776 29764 23804 29820
rect 23860 29764 23908 29820
rect 23964 29764 24012 29820
rect 24068 29764 24096 29820
rect 23776 28252 24096 29764
rect 23776 28196 23804 28252
rect 23860 28196 23908 28252
rect 23964 28196 24012 28252
rect 24068 28196 24096 28252
rect 18396 28084 18452 28094
rect 17388 27076 17444 27086
rect 17388 26852 17444 27020
rect 17388 26786 17444 26796
rect 15260 18564 15316 18574
rect 14588 18116 14644 18126
rect 14588 16436 14644 18060
rect 14700 18004 14756 18014
rect 14700 17780 14756 17948
rect 14700 17714 14756 17724
rect 14588 16370 14644 16380
rect 15260 14308 15316 18508
rect 18396 17892 18452 28028
rect 18396 17826 18452 17836
rect 23776 26684 24096 28196
rect 23776 26628 23804 26684
rect 23860 26628 23908 26684
rect 23964 26628 24012 26684
rect 24068 26628 24096 26684
rect 23776 25116 24096 26628
rect 23776 25060 23804 25116
rect 23860 25060 23908 25116
rect 23964 25060 24012 25116
rect 24068 25060 24096 25116
rect 23776 23548 24096 25060
rect 23776 23492 23804 23548
rect 23860 23492 23908 23548
rect 23964 23492 24012 23548
rect 24068 23492 24096 23548
rect 23776 21980 24096 23492
rect 23776 21924 23804 21980
rect 23860 21924 23908 21980
rect 23964 21924 24012 21980
rect 24068 21924 24096 21980
rect 23776 20412 24096 21924
rect 23776 20356 23804 20412
rect 23860 20356 23908 20412
rect 23964 20356 24012 20412
rect 24068 20356 24096 20412
rect 23776 18844 24096 20356
rect 23776 18788 23804 18844
rect 23860 18788 23908 18844
rect 23964 18788 24012 18844
rect 24068 18788 24096 18844
rect 23776 17276 24096 18788
rect 23776 17220 23804 17276
rect 23860 17220 23908 17276
rect 23964 17220 24012 17276
rect 24068 17220 24096 17276
rect 23776 15708 24096 17220
rect 23776 15652 23804 15708
rect 23860 15652 23908 15708
rect 23964 15652 24012 15708
rect 24068 15652 24096 15708
rect 15260 13412 15316 14252
rect 17052 14644 17108 14654
rect 17052 13748 17108 14588
rect 17052 13682 17108 13692
rect 23776 14140 24096 15652
rect 23776 14084 23804 14140
rect 23860 14084 23908 14140
rect 23964 14084 24012 14140
rect 24068 14084 24096 14140
rect 15260 13346 15316 13356
rect 12572 11554 12628 11564
rect 23776 12572 24096 14084
rect 23776 12516 23804 12572
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 24068 12516 24096 12572
rect 11676 11106 11732 11116
rect 11228 9650 11284 9660
rect 23776 11004 24096 12516
rect 23776 10948 23804 11004
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 24068 10948 24096 11004
rect 7084 1362 7140 1372
rect 23776 9436 24096 10948
rect 23776 9380 23804 9436
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 24068 9380 24096 9436
rect 23776 7868 24096 9380
rect 23776 7812 23804 7868
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 24068 7812 24096 7868
rect 23776 6300 24096 7812
rect 23776 6244 23804 6300
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 24068 6244 24096 6300
rect 23776 4732 24096 6244
rect 23776 4676 23804 4732
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 24068 4676 24096 4732
rect 23776 3164 24096 4676
rect 23776 3108 23804 3164
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 24068 3108 24096 3164
rect 23776 1596 24096 3108
rect 23776 1540 23804 1596
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 24068 1540 24096 1596
rect 4436 756 4464 812
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4728 756 4756 812
rect 4436 0 4756 756
rect 23776 0 24096 1540
rect 24436 55692 24756 57456
rect 24436 55636 24464 55692
rect 24520 55636 24568 55692
rect 24624 55636 24672 55692
rect 24728 55636 24756 55692
rect 24436 54124 24756 55636
rect 24436 54068 24464 54124
rect 24520 54068 24568 54124
rect 24624 54068 24672 54124
rect 24728 54068 24756 54124
rect 24436 52556 24756 54068
rect 26236 53732 26292 53742
rect 24436 52500 24464 52556
rect 24520 52500 24568 52556
rect 24624 52500 24672 52556
rect 24728 52500 24756 52556
rect 24436 50988 24756 52500
rect 24436 50932 24464 50988
rect 24520 50932 24568 50988
rect 24624 50932 24672 50988
rect 24728 50932 24756 50988
rect 24436 49420 24756 50932
rect 24436 49364 24464 49420
rect 24520 49364 24568 49420
rect 24624 49364 24672 49420
rect 24728 49364 24756 49420
rect 24436 47852 24756 49364
rect 24436 47796 24464 47852
rect 24520 47796 24568 47852
rect 24624 47796 24672 47852
rect 24728 47796 24756 47852
rect 24436 46284 24756 47796
rect 24436 46228 24464 46284
rect 24520 46228 24568 46284
rect 24624 46228 24672 46284
rect 24728 46228 24756 46284
rect 24436 44716 24756 46228
rect 24436 44660 24464 44716
rect 24520 44660 24568 44716
rect 24624 44660 24672 44716
rect 24728 44660 24756 44716
rect 24436 43148 24756 44660
rect 24436 43092 24464 43148
rect 24520 43092 24568 43148
rect 24624 43092 24672 43148
rect 24728 43092 24756 43148
rect 24436 41580 24756 43092
rect 24436 41524 24464 41580
rect 24520 41524 24568 41580
rect 24624 41524 24672 41580
rect 24728 41524 24756 41580
rect 24436 40012 24756 41524
rect 24436 39956 24464 40012
rect 24520 39956 24568 40012
rect 24624 39956 24672 40012
rect 24728 39956 24756 40012
rect 24436 38444 24756 39956
rect 24436 38388 24464 38444
rect 24520 38388 24568 38444
rect 24624 38388 24672 38444
rect 24728 38388 24756 38444
rect 24436 36876 24756 38388
rect 24436 36820 24464 36876
rect 24520 36820 24568 36876
rect 24624 36820 24672 36876
rect 24728 36820 24756 36876
rect 24436 35308 24756 36820
rect 24436 35252 24464 35308
rect 24520 35252 24568 35308
rect 24624 35252 24672 35308
rect 24728 35252 24756 35308
rect 24436 33740 24756 35252
rect 24436 33684 24464 33740
rect 24520 33684 24568 33740
rect 24624 33684 24672 33740
rect 24728 33684 24756 33740
rect 24436 32172 24756 33684
rect 24436 32116 24464 32172
rect 24520 32116 24568 32172
rect 24624 32116 24672 32172
rect 24728 32116 24756 32172
rect 24436 30604 24756 32116
rect 24436 30548 24464 30604
rect 24520 30548 24568 30604
rect 24624 30548 24672 30604
rect 24728 30548 24756 30604
rect 24436 29036 24756 30548
rect 24436 28980 24464 29036
rect 24520 28980 24568 29036
rect 24624 28980 24672 29036
rect 24728 28980 24756 29036
rect 24436 27468 24756 28980
rect 24436 27412 24464 27468
rect 24520 27412 24568 27468
rect 24624 27412 24672 27468
rect 24728 27412 24756 27468
rect 24436 25900 24756 27412
rect 24436 25844 24464 25900
rect 24520 25844 24568 25900
rect 24624 25844 24672 25900
rect 24728 25844 24756 25900
rect 24436 24332 24756 25844
rect 24436 24276 24464 24332
rect 24520 24276 24568 24332
rect 24624 24276 24672 24332
rect 24728 24276 24756 24332
rect 24436 22764 24756 24276
rect 24436 22708 24464 22764
rect 24520 22708 24568 22764
rect 24624 22708 24672 22764
rect 24728 22708 24756 22764
rect 24436 21196 24756 22708
rect 24436 21140 24464 21196
rect 24520 21140 24568 21196
rect 24624 21140 24672 21196
rect 24728 21140 24756 21196
rect 24436 19628 24756 21140
rect 24436 19572 24464 19628
rect 24520 19572 24568 19628
rect 24624 19572 24672 19628
rect 24728 19572 24756 19628
rect 24436 18060 24756 19572
rect 24436 18004 24464 18060
rect 24520 18004 24568 18060
rect 24624 18004 24672 18060
rect 24728 18004 24756 18060
rect 24436 16492 24756 18004
rect 24436 16436 24464 16492
rect 24520 16436 24568 16492
rect 24624 16436 24672 16492
rect 24728 16436 24756 16492
rect 24436 14924 24756 16436
rect 24436 14868 24464 14924
rect 24520 14868 24568 14924
rect 24624 14868 24672 14924
rect 24728 14868 24756 14924
rect 24436 13356 24756 14868
rect 24436 13300 24464 13356
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24728 13300 24756 13356
rect 24436 11788 24756 13300
rect 24436 11732 24464 11788
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24728 11732 24756 11788
rect 24436 10220 24756 11732
rect 25228 52836 25284 52846
rect 25228 11508 25284 52780
rect 26124 46564 26180 46574
rect 25340 35476 25396 35486
rect 25340 11620 25396 35420
rect 26012 25508 26068 25518
rect 26012 12852 26068 25452
rect 26012 12786 26068 12796
rect 25340 11554 25396 11564
rect 25228 11442 25284 11452
rect 24436 10164 24464 10220
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24728 10164 24756 10220
rect 24436 8652 24756 10164
rect 24436 8596 24464 8652
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24728 8596 24756 8652
rect 24436 7084 24756 8596
rect 26124 8148 26180 46508
rect 26236 8932 26292 53676
rect 27580 14420 27636 14430
rect 27580 13860 27636 14364
rect 27580 13794 27636 13804
rect 26236 8866 26292 8876
rect 26124 8082 26180 8092
rect 24436 7028 24464 7084
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 24728 7028 24756 7084
rect 24436 5516 24756 7028
rect 24436 5460 24464 5516
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24728 5460 24756 5516
rect 24436 3948 24756 5460
rect 24436 3892 24464 3948
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24728 3892 24756 3948
rect 24436 2380 24756 3892
rect 24436 2324 24464 2380
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24728 2324 24756 2380
rect 24436 812 24756 2324
rect 24436 756 24464 812
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24728 756 24756 812
rect 24436 0 24756 756
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _042_
timestamp 1486834041
transform -1 0 17024 0 -1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _043_
timestamp 1486834041
transform -1 0 15456 0 1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _044_
timestamp 1486834041
transform 1 0 15120 0 -1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _045_
timestamp 1486834041
transform 1 0 15120 0 1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _046_
timestamp 1486834041
transform -1 0 12432 0 1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _047_
timestamp 1486834041
transform -1 0 16352 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _048_
timestamp 1486834041
transform -1 0 10304 0 1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _049_
timestamp 1486834041
transform 1 0 14784 0 1 16464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _050_
timestamp 1486834041
transform 1 0 15680 0 -1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _051_
timestamp 1486834041
transform -1 0 15680 0 -1 18032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _052_
timestamp 1486834041
transform 1 0 16800 0 1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _053_
timestamp 1486834041
transform 1 0 12768 0 -1 21168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _054_
timestamp 1486834041
transform 1 0 16576 0 -1 19600
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _055_
timestamp 1486834041
transform 1 0 13216 0 1 18032
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _056_
timestamp 1486834041
transform -1 0 17248 0 -1 21168
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _057_
timestamp 1486834041
transform 1 0 15344 0 1 19600
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _058_
timestamp 1486834041
transform 1 0 13664 0 1 16464
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _059_
timestamp 1486834041
transform 1 0 15456 0 1 18032
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _060_
timestamp 1486834041
transform 1 0 12768 0 -1 19600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _061_
timestamp 1486834041
transform -1 0 13328 0 1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _062_
timestamp 1486834041
transform -1 0 12768 0 -1 19600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _063_
timestamp 1486834041
transform -1 0 10192 0 -1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _064_
timestamp 1486834041
transform 1 0 12656 0 1 22736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _065_
timestamp 1486834041
transform -1 0 12432 0 1 24304
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _066_
timestamp 1486834041
transform 1 0 12656 0 1 19600
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _067_
timestamp 1486834041
transform -1 0 13328 0 1 21168
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _068_
timestamp 1486834041
transform 1 0 11312 0 1 19600
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _069_
timestamp 1486834041
transform -1 0 12432 0 1 22736
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _070_
timestamp 1486834041
transform -1 0 12768 0 -1 21168
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _071_
timestamp 1486834041
transform 1 0 16576 0 -1 32144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _072_
timestamp 1486834041
transform 1 0 12432 0 -1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _073_
timestamp 1486834041
transform 1 0 7392 0 1 36848
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _074_
timestamp 1486834041
transform -1 0 4592 0 1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _075_
timestamp 1486834041
transform 1 0 16576 0 1 30576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _076_
timestamp 1486834041
transform 1 0 11872 0 -1 32144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _077_
timestamp 1486834041
transform 1 0 9968 0 -1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _078_
timestamp 1486834041
transform 1 0 6160 0 1 21168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _079_
timestamp 1486834041
transform 1 0 4928 0 -1 39984
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _080_
timestamp 1486834041
transform 1 0 1008 0 1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _081_
timestamp 1486834041
transform 1 0 6608 0 1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _082_
timestamp 1486834041
transform 1 0 4816 0 1 27440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _083_
timestamp 1486834041
transform -1 0 16912 0 1 21168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _084_
timestamp 1486834041
transform 1 0 12768 0 1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _085_
timestamp 1486834041
transform -1 0 4592 0 1 30576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _086_
timestamp 1486834041
transform 1 0 1904 0 -1 25872
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _087_
timestamp 1486834041
transform 1 0 6160 0 1 32144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _088_
timestamp 1486834041
transform 1 0 11424 0 -1 38416
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _089_
timestamp 1486834041
transform 1 0 1008 0 1 33712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _090_
timestamp 1486834041
transform 1 0 4928 0 -1 30576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _091_
timestamp 1486834041
transform -1 0 16352 0 -1 22736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _092_
timestamp 1486834041
transform 1 0 12656 0 -1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _093_
timestamp 1486834041
transform 1 0 12656 0 1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _094_
timestamp 1486834041
transform 1 0 10640 0 -1 16464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _095_
timestamp 1486834041
transform 1 0 1680 0 -1 32144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _096_
timestamp 1486834041
transform 1 0 2128 0 -1 21168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _097_
timestamp 1486834041
transform 1 0 4928 0 -1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _098_
timestamp 1486834041
transform 1 0 11312 0 -1 39984
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _099_
timestamp 1486834041
transform 1 0 18256 0 -1 29008
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _100_
timestamp 1486834041
transform 1 0 13440 0 1 27440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _101_
timestamp 1486834041
transform 1 0 8848 0 1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _102_
timestamp 1486834041
transform 1 0 7392 0 1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _103_
timestamp 1486834041
transform 1 0 9296 0 -1 30576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _104_
timestamp 1486834041
transform 1 0 4480 0 -1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _105_
timestamp 1486834041
transform 1 0 7168 0 1 39984
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _106_
timestamp 1486834041
transform 1 0 4032 0 -1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _107_
timestamp 1486834041
transform 1 0 17360 0 -1 25872
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _108_
timestamp 1486834041
transform 1 0 12768 0 -1 29008
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _109_
timestamp 1486834041
transform 1 0 9744 0 -1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _110_
timestamp 1486834041
transform 1 0 8736 0 -1 22736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _111_
timestamp 1486834041
transform 1 0 8848 0 1 27440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _112_
timestamp 1486834041
transform 1 0 4816 0 -1 22736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _113_
timestamp 1486834041
transform 1 0 7728 0 1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _114_
timestamp 1486834041
transform 1 0 4368 0 -1 14896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _115_
timestamp 1486834041
transform 1 0 18032 0 1 32144
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _116_
timestamp 1486834041
transform 1 0 14560 0 -1 36848
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _117_
timestamp 1486834041
transform 1 0 19600 0 -1 21168
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _118_
timestamp 1486834041
transform 1 0 13888 0 -1 11760
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _119_
timestamp 1486834041
transform -1 0 15680 0 -1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _120_
timestamp 1486834041
transform -1 0 16688 0 1 13328
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _121_
timestamp 1486834041
transform 1 0 15568 0 1 14896
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _122_
timestamp 1486834041
transform 1 0 16688 0 1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _123_
timestamp 1486834041
transform -1 0 15568 0 1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _124_
timestamp 1486834041
transform 1 0 15792 0 -1 14896
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _125_
timestamp 1486834041
transform -1 0 16352 0 -1 16464
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _126_
timestamp 1486834041
transform 1 0 16576 0 -1 14896
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _127_
timestamp 1486834041
transform 1 0 9744 0 1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _128_
timestamp 1486834041
transform -1 0 11536 0 1 16464
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _129_
timestamp 1486834041
transform 1 0 9744 0 -1 14896
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _130_
timestamp 1486834041
transform -1 0 9744 0 -1 14896
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _131_
timestamp 1486834041
transform 1 0 10864 0 -1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _132_
timestamp 1486834041
transform 1 0 9744 0 -1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _133_
timestamp 1486834041
transform 1 0 11648 0 1 14896
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _134_
timestamp 1486834041
transform 1 0 8960 0 -1 16464
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _135_
timestamp 1486834041
transform -1 0 11648 0 1 14896
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _136_
timestamp 1486834041
transform 1 0 12880 0 1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _137_
timestamp 1486834041
transform 1 0 17808 0 1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _138_
timestamp 1486834041
transform -1 0 18816 0 -1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _139_
timestamp 1486834041
transform 1 0 17584 0 -1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _140_
timestamp 1486834041
transform 1 0 1792 0 -1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _141_
timestamp 1486834041
transform 1 0 4032 0 -1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _142_
timestamp 1486834041
transform 1 0 5488 0 1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _143_
timestamp 1486834041
transform -1 0 10976 0 -1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _144_
timestamp 1486834041
transform 1 0 2352 0 1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _145_
timestamp 1486834041
transform 1 0 3808 0 -1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _146_
timestamp 1486834041
transform 1 0 6272 0 -1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _147_
timestamp 1486834041
transform 1 0 8176 0 1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _148_
timestamp 1486834041
transform 1 0 6272 0 -1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _149_
timestamp 1486834041
transform 1 0 6384 0 1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _150_
timestamp 1486834041
transform 1 0 6272 0 -1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _151_
timestamp 1486834041
transform 1 0 9072 0 1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _152_
timestamp 1486834041
transform 1 0 10976 0 -1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _153_
timestamp 1486834041
transform 1 0 10528 0 -1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _154_
timestamp 1486834041
transform 1 0 16128 0 1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _155_
timestamp 1486834041
transform 1 0 17472 0 -1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _156_
timestamp 1486834041
transform 1 0 1792 0 -1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _157_
timestamp 1486834041
transform 1 0 4816 0 1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _158_
timestamp 1486834041
transform 1 0 4368 0 -1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _159_
timestamp 1486834041
transform 1 0 2352 0 1 39984
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _160_
timestamp 1486834041
transform 1 0 2352 0 1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _161_
timestamp 1486834041
transform 1 0 3136 0 -1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _162_
timestamp 1486834041
transform 1 0 7840 0 1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _163_
timestamp 1486834041
transform 1 0 9184 0 -1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _164_
timestamp 1486834041
transform 1 0 5936 0 -1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _165_
timestamp 1486834041
transform 1 0 7280 0 1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _166_
timestamp 1486834041
transform 1 0 6608 0 1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _167_
timestamp 1486834041
transform 1 0 8736 0 -1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _168_
timestamp 1486834041
transform 1 0 13216 0 -1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _169_
timestamp 1486834041
transform 1 0 13328 0 1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _170_
timestamp 1486834041
transform 1 0 17136 0 1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _171_
timestamp 1486834041
transform 1 0 17808 0 1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _172_
timestamp 1486834041
transform 1 0 9856 0 -1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _173_
timestamp 1486834041
transform 1 0 9072 0 -1 39984
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _174_
timestamp 1486834041
transform 1 0 4816 0 1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _175_
timestamp 1486834041
transform 1 0 2352 0 -1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _176_
timestamp 1486834041
transform 1 0 1904 0 -1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _177_
timestamp 1486834041
transform -1 0 3584 0 -1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _178_
timestamp 1486834041
transform 1 0 1344 0 1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _179_
timestamp 1486834041
transform 1 0 896 0 -1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _180_
timestamp 1486834041
transform 1 0 6272 0 -1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _181_
timestamp 1486834041
transform 1 0 7728 0 1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _182_
timestamp 1486834041
transform 1 0 9184 0 1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _183_
timestamp 1486834041
transform 1 0 10192 0 1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _184_
timestamp 1486834041
transform 1 0 10416 0 -1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _185_
timestamp 1486834041
transform 1 0 10080 0 -1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _186_
timestamp 1486834041
transform -1 0 18816 0 -1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _187_
timestamp 1486834041
transform -1 0 19376 0 1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _188_
timestamp 1486834041
transform 1 0 4816 0 1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _189_
timestamp 1486834041
transform 1 0 3136 0 -1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _190_
timestamp 1486834041
transform 1 0 896 0 -1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _191_
timestamp 1486834041
transform -1 0 3136 0 -1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _192_
timestamp 1486834041
transform 1 0 10192 0 1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _193_
timestamp 1486834041
transform 1 0 9184 0 -1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _194_
timestamp 1486834041
transform -1 0 9520 0 1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _195_
timestamp 1486834041
transform 1 0 5264 0 -1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _196_
timestamp 1486834041
transform 1 0 1344 0 1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _197_
timestamp 1486834041
transform 1 0 896 0 -1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _198_
timestamp 1486834041
transform 1 0 896 0 -1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _199_
timestamp 1486834041
transform 1 0 896 0 1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _200_
timestamp 1486834041
transform 1 0 12320 0 -1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _201_
timestamp 1486834041
transform -1 0 18592 0 1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _202_
timestamp 1486834041
transform -1 0 19152 0 1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _203_
timestamp 1486834041
transform -1 0 19600 0 -1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _204_
timestamp 1486834041
transform 1 0 2352 0 1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _205_
timestamp 1486834041
transform 1 0 4592 0 -1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _206_
timestamp 1486834041
transform 1 0 4032 0 -1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _207_
timestamp 1486834041
transform 1 0 3920 0 -1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _208_
timestamp 1486834041
transform -1 0 3920 0 1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _209_
timestamp 1486834041
transform -1 0 3920 0 -1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _210_
timestamp 1486834041
transform 1 0 3584 0 -1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _211_
timestamp 1486834041
transform 1 0 5264 0 1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _212_
timestamp 1486834041
transform 1 0 5264 0 1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _213_
timestamp 1486834041
transform 1 0 5936 0 -1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _214_
timestamp 1486834041
transform 1 0 6944 0 1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _215_
timestamp 1486834041
transform 1 0 9408 0 -1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _216_
timestamp 1486834041
transform 1 0 10192 0 1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _217_
timestamp 1486834041
transform 1 0 11536 0 -1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _218_
timestamp 1486834041
transform 1 0 15568 0 1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _219_
timestamp 1486834041
transform 1 0 16576 0 -1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _220_
timestamp 1486834041
transform 1 0 1904 0 1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _221_
timestamp 1486834041
transform -1 0 4480 0 -1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _222_
timestamp 1486834041
transform 1 0 4816 0 1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _223_
timestamp 1486834041
transform 1 0 2352 0 1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _224_
timestamp 1486834041
transform 1 0 10192 0 -1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _225_
timestamp 1486834041
transform 1 0 11424 0 -1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _226_
timestamp 1486834041
transform 1 0 13888 0 1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _227_
timestamp 1486834041
transform 1 0 14896 0 1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _228_
timestamp 1486834041
transform 1 0 9744 0 1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _229_
timestamp 1486834041
transform 1 0 8624 0 1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _230_
timestamp 1486834041
transform 1 0 6384 0 1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _231_
timestamp 1486834041
transform 1 0 8624 0 1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _232_
timestamp 1486834041
transform 1 0 13552 0 -1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _233_
timestamp 1486834041
transform -1 0 18816 0 -1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _234_
timestamp 1486834041
transform -1 0 18928 0 1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _235_
timestamp 1486834041
transform -1 0 19376 0 -1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _236_
timestamp 1486834041
transform 1 0 9968 0 1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _237_
timestamp 1486834041
transform 1 0 9296 0 -1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _238_
timestamp 1486834041
transform 1 0 6384 0 1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _239_
timestamp 1486834041
transform 1 0 7616 0 1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _240_
timestamp 1486834041
transform 1 0 6160 0 -1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _241_
timestamp 1486834041
transform 1 0 5376 0 1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_4  _242_
timestamp 1486834041
transform 1 0 16576 0 -1 38416
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_4  _243_
timestamp 1486834041
transform -1 0 18704 0 1 39984
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _244_
timestamp 1486834041
transform -1 0 2128 0 -1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _245_
timestamp 1486834041
transform 1 0 3584 0 1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _246_
timestamp 1486834041
transform 1 0 11536 0 1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _247_
timestamp 1486834041
transform 1 0 13328 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _248_
timestamp 1486834041
transform 1 0 13888 0 1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _249_
timestamp 1486834041
transform 1 0 16240 0 1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _250_
timestamp 1486834041
transform 1 0 6048 0 1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _251_
timestamp 1486834041
transform 1 0 3136 0 -1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _252_
timestamp 1486834041
transform 1 0 12768 0 1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _253_
timestamp 1486834041
transform 1 0 7504 0 -1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _254_
timestamp 1486834041
transform 1 0 3584 0 1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _255_
timestamp 1486834041
transform -1 0 3360 0 -1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _256_
timestamp 1486834041
transform 1 0 14560 0 -1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _257_
timestamp 1486834041
transform 1 0 14448 0 1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _258_
timestamp 1486834041
transform 1 0 1904 0 -1 41552
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _259_
timestamp 1486834041
transform 1 0 1792 0 -1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _260_
timestamp 1486834041
transform 1 0 3696 0 1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _261_
timestamp 1486834041
transform 1 0 5488 0 1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _262_
timestamp 1486834041
transform 1 0 7616 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _263_
timestamp 1486834041
transform 1 0 9968 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _264_
timestamp 1486834041
transform 1 0 11200 0 1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _265_
timestamp 1486834041
transform 1 0 11536 0 1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _266_
timestamp 1486834041
transform 1 0 15456 0 -1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _267_
timestamp 1486834041
transform 1 0 19264 0 -1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _268_
timestamp 1486834041
transform 1 0 2464 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _269_
timestamp 1486834041
transform 1 0 2464 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _270_
timestamp 1486834041
transform 1 0 2688 0 1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _271_
timestamp 1486834041
transform 1 0 1456 0 1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _272_
timestamp 1486834041
transform 1 0 6608 0 -1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _273_
timestamp 1486834041
transform 1 0 3136 0 -1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _274_
timestamp 1486834041
transform 1 0 13664 0 1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _275_
timestamp 1486834041
transform 1 0 14448 0 -1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _276_
timestamp 1486834041
transform 1 0 2464 0 1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _277_
timestamp 1486834041
transform 1 0 1008 0 1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _278_
timestamp 1486834041
transform 1 0 1792 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _279_
timestamp 1486834041
transform 1 0 2688 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _280_
timestamp 1486834041
transform 1 0 12656 0 1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _281_
timestamp 1486834041
transform 1 0 18816 0 1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _282_
timestamp 1486834041
transform 1 0 19712 0 -1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _283_
timestamp 1486834041
transform 1 0 19040 0 1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _284_
timestamp 1486834041
transform 1 0 3472 0 1 41552
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _285_
timestamp 1486834041
transform 1 0 5936 0 -1 41552
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _286_
timestamp 1486834041
transform 1 0 5152 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _287_
timestamp 1486834041
transform 1 0 1792 0 1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _288_
timestamp 1486834041
transform 1 0 2688 0 -1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _289_
timestamp 1486834041
transform 1 0 2688 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _290_
timestamp 1486834041
transform -1 0 12208 0 1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _291_
timestamp 1486834041
transform 1 0 1792 0 -1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _292_
timestamp 1486834041
transform 1 0 2688 0 1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _293_
timestamp 1486834041
transform 1 0 18144 0 -1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _294_
timestamp 1486834041
transform 1 0 20496 0 1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _295_
timestamp 1486834041
transform 1 0 18816 0 1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _296_
timestamp 1486834041
transform 1 0 19824 0 -1 55664
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _297_
timestamp 1486834041
transform 1 0 23632 0 1 50960
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _298_
timestamp 1486834041
transform 1 0 21616 0 -1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _299_
timestamp 1486834041
transform 1 0 22624 0 1 50960
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _300_
timestamp 1486834041
transform 1 0 20720 0 -1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _301_
timestamp 1486834041
transform 1 0 21168 0 1 52528
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _302_
timestamp 1486834041
transform 1 0 22064 0 1 52528
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _303_
timestamp 1486834041
transform -1 0 19600 0 -1 55664
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _304_
timestamp 1486834041
transform 1 0 23632 0 1 49392
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _305_
timestamp 1486834041
transform 1 0 24304 0 1 47824
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _306_
timestamp 1486834041
transform -1 0 22624 0 -1 52528
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _307_
timestamp 1486834041
transform 1 0 25200 0 1 47824
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _308_
timestamp 1486834041
transform -1 0 24192 0 -1 50960
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _309_
timestamp 1486834041
transform -1 0 20720 0 -1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _310_
timestamp 1486834041
transform -1 0 15680 0 -1 38416
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _311_
timestamp 1486834041
transform 1 0 14224 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _312_
timestamp 1486834041
transform -1 0 20048 0 1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _313_
timestamp 1486834041
transform -1 0 14560 0 -1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _314_
timestamp 1486834041
transform 1 0 18816 0 -1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _315_
timestamp 1486834041
transform 1 0 5264 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _316_
timestamp 1486834041
transform -1 0 8512 0 -1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _317_
timestamp 1486834041
transform 1 0 5488 0 1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _318_
timestamp 1486834041
transform 1 0 10080 0 -1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _319_
timestamp 1486834041
transform -1 0 10080 0 -1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _320_
timestamp 1486834041
transform 1 0 11200 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _321_
timestamp 1486834041
transform 1 0 14000 0 -1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _322_
timestamp 1486834041
transform 1 0 18816 0 1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _323_
timestamp 1486834041
transform -1 0 5488 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _324_
timestamp 1486834041
transform 1 0 8736 0 -1 41552
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _325_
timestamp 1486834041
transform 1 0 5488 0 1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _326_
timestamp 1486834041
transform 1 0 10192 0 1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _327_
timestamp 1486834041
transform 1 0 8736 0 -1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _328_
timestamp 1486834041
transform 1 0 12096 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _329_
timestamp 1486834041
transform 1 0 15456 0 -1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _330_
timestamp 1486834041
transform 1 0 19376 0 1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _331_
timestamp 1486834041
transform -1 0 6272 0 -1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _332_
timestamp 1486834041
transform -1 0 7728 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _333_
timestamp 1486834041
transform 1 0 3584 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _334_
timestamp 1486834041
transform 1 0 6272 0 1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _335_
timestamp 1486834041
transform -1 0 6160 0 1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _336_
timestamp 1486834041
transform 1 0 10864 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _337_
timestamp 1486834041
transform 1 0 12768 0 1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _338_
timestamp 1486834041
transform -1 0 18032 0 1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _339_
timestamp 1486834041
transform -1 0 1904 0 -1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _340_
timestamp 1486834041
transform -1 0 8512 0 -1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _341_
timestamp 1486834041
transform -1 0 13552 0 1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _342_
timestamp 1486834041
transform -1 0 17584 0 -1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _343_
timestamp 1486834041
transform 1 0 12768 0 1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _344_
timestamp 1486834041
transform 1 0 6048 0 -1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_UserCLK
timestamp 1486834041
transform 1 0 16576 0 -1 39984
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_UserCLK_regs
timestamp 1486834041
transform -1 0 20272 0 1 36848
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_UserCLK
timestamp 1486834041
transform -1 0 19152 0 1 35280
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_UserCLK_regs
timestamp 1486834041
transform -1 0 20160 0 1 33712
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_UserCLK_regs
timestamp 1486834041
transform 1 0 14672 0 1 41552
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_regs_0_UserCLK
timestamp 1486834041
transform 1 0 14672 0 1 38416
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout27
timestamp 1486834041
transform -1 0 18144 0 -1 36848
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout28
timestamp 1486834041
transform -1 0 8624 0 1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout29
timestamp 1486834041
transform 1 0 7616 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout30
timestamp 1486834041
transform -1 0 2464 0 1 18032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout31
timestamp 1486834041
transform -1 0 4032 0 1 19600
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout32
timestamp 1486834041
transform 1 0 896 0 1 19600
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout33
timestamp 1486834041
transform 1 0 896 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout34
timestamp 1486834041
transform -1 0 2464 0 -1 30576
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout35
timestamp 1486834041
transform 1 0 3136 0 -1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout36
timestamp 1486834041
transform -1 0 1792 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout37
timestamp 1486834041
transform 1 0 4816 0 1 16464
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout38
timestamp 1486834041
transform -1 0 4592 0 1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout39
timestamp 1486834041
transform -1 0 7840 0 1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout40
timestamp 1486834041
transform 1 0 6944 0 -1 32144
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout41
timestamp 1486834041
transform 1 0 8736 0 -1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2
timestamp 1486834041
transform 1 0 896 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36
timestamp 1486834041
transform 1 0 4704 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45
timestamp 1486834041
transform 1 0 5712 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57
timestamp 1486834041
transform 1 0 7056 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65
timestamp 1486834041
transform 1 0 7952 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67
timestamp 1486834041
transform 1 0 8176 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_70
timestamp 1486834041
transform 1 0 8512 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_104
timestamp 1486834041
transform 1 0 12320 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_138
timestamp 1486834041
transform 1 0 16128 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_172
timestamp 1486834041
transform 1 0 19936 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_206
timestamp 1486834041
transform 1 0 23744 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_240
timestamp 1486834041
transform 1 0 27552 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_2
timestamp 1486834041
transform 1 0 896 0 -1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_66
timestamp 1486834041
transform 1 0 8064 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_72
timestamp 1486834041
transform 1 0 8736 0 -1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_136
timestamp 1486834041
transform 1 0 15904 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_142
timestamp 1486834041
transform 1 0 16576 0 -1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_206
timestamp 1486834041
transform 1 0 23744 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_212
timestamp 1486834041
transform 1 0 24416 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_220
timestamp 1486834041
transform 1 0 25312 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_224
timestamp 1486834041
transform 1 0 25760 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_2
timestamp 1486834041
transform 1 0 896 0 1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1486834041
transform 1 0 4480 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_37
timestamp 1486834041
transform 1 0 4816 0 1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_101
timestamp 1486834041
transform 1 0 11984 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_107
timestamp 1486834041
transform 1 0 12656 0 1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_171
timestamp 1486834041
transform 1 0 19824 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_177
timestamp 1486834041
transform 1 0 20496 0 1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_209
timestamp 1486834041
transform 1 0 24080 0 1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_2
timestamp 1486834041
transform 1 0 896 0 -1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_66
timestamp 1486834041
transform 1 0 8064 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_72
timestamp 1486834041
transform 1 0 8736 0 -1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_136
timestamp 1486834041
transform 1 0 15904 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_142
timestamp 1486834041
transform 1 0 16576 0 -1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_206
timestamp 1486834041
transform 1 0 23744 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_212
timestamp 1486834041
transform 1 0 24416 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_220
timestamp 1486834041
transform 1 0 25312 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_224
timestamp 1486834041
transform 1 0 25760 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_10
timestamp 1486834041
transform 1 0 1792 0 1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_26
timestamp 1486834041
transform 1 0 3584 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1486834041
transform 1 0 4480 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_37
timestamp 1486834041
transform 1 0 4816 0 1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_101
timestamp 1486834041
transform 1 0 11984 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_107
timestamp 1486834041
transform 1 0 12656 0 1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_171
timestamp 1486834041
transform 1 0 19824 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_177
timestamp 1486834041
transform 1 0 20496 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_209
timestamp 1486834041
transform 1 0 24080 0 1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_225
timestamp 1486834041
transform 1 0 25872 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_2
timestamp 1486834041
transform 1 0 896 0 -1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_66
timestamp 1486834041
transform 1 0 8064 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_72
timestamp 1486834041
transform 1 0 8736 0 -1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_136
timestamp 1486834041
transform 1 0 15904 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_142
timestamp 1486834041
transform 1 0 16576 0 -1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_206
timestamp 1486834041
transform 1 0 23744 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_212
timestamp 1486834041
transform 1 0 24416 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_220
timestamp 1486834041
transform 1 0 25312 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_224
timestamp 1486834041
transform 1 0 25760 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_16
timestamp 1486834041
transform 1 0 2464 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_32
timestamp 1486834041
transform 1 0 4256 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1486834041
transform 1 0 4480 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_37
timestamp 1486834041
transform 1 0 4816 0 1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_101
timestamp 1486834041
transform 1 0 11984 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_107
timestamp 1486834041
transform 1 0 12656 0 1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_171
timestamp 1486834041
transform 1 0 19824 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_177
timestamp 1486834041
transform 1 0 20496 0 1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_209
timestamp 1486834041
transform 1 0 24080 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_16
timestamp 1486834041
transform 1 0 2464 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_48
timestamp 1486834041
transform 1 0 6048 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_64
timestamp 1486834041
transform 1 0 7840 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_68
timestamp 1486834041
transform 1 0 8288 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_72
timestamp 1486834041
transform 1 0 8736 0 -1 7056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_136
timestamp 1486834041
transform 1 0 15904 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_142
timestamp 1486834041
transform 1 0 16576 0 -1 7056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_206
timestamp 1486834041
transform 1 0 23744 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_212
timestamp 1486834041
transform 1 0 24416 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_220
timestamp 1486834041
transform 1 0 25312 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_224
timestamp 1486834041
transform 1 0 25760 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_10
timestamp 1486834041
transform 1 0 1792 0 1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_26
timestamp 1486834041
transform 1 0 3584 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1486834041
transform 1 0 4480 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_37
timestamp 1486834041
transform 1 0 4816 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_69
timestamp 1486834041
transform 1 0 8400 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_77
timestamp 1486834041
transform 1 0 9296 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_81
timestamp 1486834041
transform 1 0 9744 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_99
timestamp 1486834041
transform 1 0 11760 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_103
timestamp 1486834041
transform 1 0 12208 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_107
timestamp 1486834041
transform 1 0 12656 0 1 7056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_171
timestamp 1486834041
transform 1 0 19824 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_177
timestamp 1486834041
transform 1 0 20496 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_209
timestamp 1486834041
transform 1 0 24080 0 1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_225
timestamp 1486834041
transform 1 0 25872 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_10
timestamp 1486834041
transform 1 0 1792 0 -1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_42
timestamp 1486834041
transform 1 0 5376 0 -1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_58
timestamp 1486834041
transform 1 0 7168 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_72
timestamp 1486834041
transform 1 0 8736 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_76
timestamp 1486834041
transform 1 0 9184 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_98
timestamp 1486834041
transform 1 0 11648 0 -1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_130
timestamp 1486834041
transform 1 0 15232 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_138
timestamp 1486834041
transform 1 0 16128 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_142
timestamp 1486834041
transform 1 0 16576 0 -1 8624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_206
timestamp 1486834041
transform 1 0 23744 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_212
timestamp 1486834041
transform 1 0 24416 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_220
timestamp 1486834041
transform 1 0 25312 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_224
timestamp 1486834041
transform 1 0 25760 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_18
timestamp 1486834041
transform 1 0 2688 0 1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1486834041
transform 1 0 4480 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_37
timestamp 1486834041
transform 1 0 4816 0 1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_53
timestamp 1486834041
transform 1 0 6608 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_55
timestamp 1486834041
transform 1 0 6832 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_96
timestamp 1486834041
transform 1 0 11424 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_104
timestamp 1486834041
transform 1 0 12320 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_107
timestamp 1486834041
transform 1 0 12656 0 1 8624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_171
timestamp 1486834041
transform 1 0 19824 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_177
timestamp 1486834041
transform 1 0 20496 0 1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_209
timestamp 1486834041
transform 1 0 24080 0 1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_24
timestamp 1486834041
transform 1 0 3360 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_32
timestamp 1486834041
transform 1 0 4256 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_34
timestamp 1486834041
transform 1 0 4480 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_43
timestamp 1486834041
transform 1 0 5488 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_51
timestamp 1486834041
transform 1 0 6384 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_63
timestamp 1486834041
transform 1 0 7728 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_67
timestamp 1486834041
transform 1 0 8176 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_69
timestamp 1486834041
transform 1 0 8400 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_72
timestamp 1486834041
transform 1 0 8736 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_80
timestamp 1486834041
transform 1 0 9632 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_82
timestamp 1486834041
transform 1 0 9856 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_115
timestamp 1486834041
transform 1 0 13552 0 -1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_131
timestamp 1486834041
transform 1 0 15344 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_139
timestamp 1486834041
transform 1 0 16240 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_142
timestamp 1486834041
transform 1 0 16576 0 -1 10192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_206
timestamp 1486834041
transform 1 0 23744 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_212
timestamp 1486834041
transform 1 0 24416 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_220
timestamp 1486834041
transform 1 0 25312 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_224
timestamp 1486834041
transform 1 0 25760 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_26
timestamp 1486834041
transform 1 0 3584 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1486834041
transform 1 0 4480 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_37
timestamp 1486834041
transform 1 0 4816 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_39
timestamp 1486834041
transform 1 0 5040 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_48
timestamp 1486834041
transform 1 0 6048 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_52
timestamp 1486834041
transform 1 0 6496 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_107
timestamp 1486834041
transform 1 0 12656 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_111
timestamp 1486834041
transform 1 0 13104 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_129
timestamp 1486834041
transform 1 0 15120 0 1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_161
timestamp 1486834041
transform 1 0 18704 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_169
timestamp 1486834041
transform 1 0 19600 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_173
timestamp 1486834041
transform 1 0 20048 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_177
timestamp 1486834041
transform 1 0 20496 0 1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_209
timestamp 1486834041
transform 1 0 24080 0 1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_225
timestamp 1486834041
transform 1 0 25872 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_24
timestamp 1486834041
transform 1 0 3360 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_28
timestamp 1486834041
transform 1 0 3808 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_72
timestamp 1486834041
transform 1 0 8736 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_80
timestamp 1486834041
transform 1 0 9632 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_113
timestamp 1486834041
transform 1 0 13328 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_117
timestamp 1486834041
transform 1 0 13776 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_133
timestamp 1486834041
transform 1 0 15568 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_137
timestamp 1486834041
transform 1 0 16016 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_139
timestamp 1486834041
transform 1 0 16240 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_142
timestamp 1486834041
transform 1 0 16576 0 -1 11760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_206
timestamp 1486834041
transform 1 0 23744 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_212
timestamp 1486834041
transform 1 0 24416 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_220
timestamp 1486834041
transform 1 0 25312 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_224
timestamp 1486834041
transform 1 0 25760 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1486834041
transform 1 0 4480 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_37
timestamp 1486834041
transform 1 0 4816 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_49
timestamp 1486834041
transform 1 0 6160 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_139
timestamp 1486834041
transform 1 0 16240 0 1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_171
timestamp 1486834041
transform 1 0 19824 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_177
timestamp 1486834041
transform 1 0 20496 0 1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_209
timestamp 1486834041
transform 1 0 24080 0 1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_92
timestamp 1486834041
transform 1 0 10976 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_110
timestamp 1486834041
transform 1 0 12992 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_118
timestamp 1486834041
transform 1 0 13888 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_134
timestamp 1486834041
transform 1 0 15680 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_142
timestamp 1486834041
transform 1 0 16576 0 -1 13328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_206
timestamp 1486834041
transform 1 0 23744 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_212
timestamp 1486834041
transform 1 0 24416 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_220
timestamp 1486834041
transform 1 0 25312 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_224
timestamp 1486834041
transform 1 0 25760 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_2
timestamp 1486834041
transform 1 0 896 0 1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_71
timestamp 1486834041
transform 1 0 8624 0 1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_95
timestamp 1486834041
transform 1 0 11312 0 1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_103
timestamp 1486834041
transform 1 0 12208 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_107
timestamp 1486834041
transform 1 0 12656 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_151
timestamp 1486834041
transform 1 0 17584 0 1 13328
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_167
timestamp 1486834041
transform 1 0 19376 0 1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_177
timestamp 1486834041
transform 1 0 20496 0 1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_209
timestamp 1486834041
transform 1 0 24080 0 1 13328
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_225
timestamp 1486834041
transform 1 0 25872 0 1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_26
timestamp 1486834041
transform 1 0 3584 0 -1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_30
timestamp 1486834041
transform 1 0 4032 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_32
timestamp 1486834041
transform 1 0 4256 0 -1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_65
timestamp 1486834041
transform 1 0 7952 0 -1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_69
timestamp 1486834041
transform 1 0 8400 0 -1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_72
timestamp 1486834041
transform 1 0 8736 0 -1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_97
timestamp 1486834041
transform 1 0 11536 0 -1 14896
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_113
timestamp 1486834041
transform 1 0 13328 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_17_154
timestamp 1486834041
transform 1 0 17920 0 -1 14896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_186
timestamp 1486834041
transform 1 0 21504 0 -1 14896
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_202
timestamp 1486834041
transform 1 0 23296 0 -1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_212
timestamp 1486834041
transform 1 0 24416 0 -1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_220
timestamp 1486834041
transform 1 0 25312 0 -1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_224
timestamp 1486834041
transform 1 0 25760 0 -1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_2
timestamp 1486834041
transform 1 0 896 0 1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_6
timestamp 1486834041
transform 1 0 1344 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_8
timestamp 1486834041
transform 1 0 1568 0 1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_29
timestamp 1486834041
transform 1 0 3920 0 1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_33
timestamp 1486834041
transform 1 0 4368 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_37
timestamp 1486834041
transform 1 0 4816 0 1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_41
timestamp 1486834041
transform 1 0 5264 0 1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_103
timestamp 1486834041
transform 1 0 12208 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_107
timestamp 1486834041
transform 1 0 12656 0 1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_111
timestamp 1486834041
transform 1 0 13104 0 1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_118
timestamp 1486834041
transform 1 0 13888 0 1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_122
timestamp 1486834041
transform 1 0 14336 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_124
timestamp 1486834041
transform 1 0 14560 0 1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_163
timestamp 1486834041
transform 1 0 18928 0 1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_171
timestamp 1486834041
transform 1 0 19824 0 1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_177
timestamp 1486834041
transform 1 0 20496 0 1 14896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_209
timestamp 1486834041
transform 1 0 24080 0 1 14896
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_2
timestamp 1486834041
transform 1 0 896 0 -1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_6
timestamp 1486834041
transform 1 0 1344 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_8
timestamp 1486834041
transform 1 0 1568 0 -1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_69
timestamp 1486834041
transform 1 0 8400 0 -1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_72
timestamp 1486834041
transform 1 0 8736 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_121
timestamp 1486834041
transform 1 0 14224 0 -1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_19_162
timestamp 1486834041
transform 1 0 18816 0 -1 16464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_194
timestamp 1486834041
transform 1 0 22400 0 -1 16464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_212
timestamp 1486834041
transform 1 0 24416 0 -1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_220
timestamp 1486834041
transform 1 0 25312 0 -1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_224
timestamp 1486834041
transform 1 0 25760 0 -1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_26
timestamp 1486834041
transform 1 0 3584 0 1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_71
timestamp 1486834041
transform 1 0 8624 0 1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_79
timestamp 1486834041
transform 1 0 9520 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_113
timestamp 1486834041
transform 1 0 13328 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_115
timestamp 1486834041
transform 1 0 13552 0 1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_158
timestamp 1486834041
transform 1 0 18368 0 1 16464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_174
timestamp 1486834041
transform 1 0 20160 0 1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_177
timestamp 1486834041
transform 1 0 20496 0 1 16464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_209
timestamp 1486834041
transform 1 0 24080 0 1 16464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_225
timestamp 1486834041
transform 1 0 25872 0 1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_72
timestamp 1486834041
transform 1 0 8736 0 -1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_76
timestamp 1486834041
transform 1 0 9184 0 -1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_97
timestamp 1486834041
transform 1 0 11536 0 -1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_101
timestamp 1486834041
transform 1 0 11984 0 -1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_142
timestamp 1486834041
transform 1 0 16576 0 -1 18032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_206
timestamp 1486834041
transform 1 0 23744 0 -1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_212
timestamp 1486834041
transform 1 0 24416 0 -1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_220
timestamp 1486834041
transform 1 0 25312 0 -1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_224
timestamp 1486834041
transform 1 0 25760 0 -1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_24
timestamp 1486834041
transform 1 0 3360 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_26
timestamp 1486834041
transform 1 0 3584 0 1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_37
timestamp 1486834041
transform 1 0 4816 0 1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_61
timestamp 1486834041
transform 1 0 7504 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_103
timestamp 1486834041
transform 1 0 12208 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_107
timestamp 1486834041
transform 1 0 12656 0 1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_111
timestamp 1486834041
transform 1 0 13104 0 1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_127
timestamp 1486834041
transform 1 0 14896 0 1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_152
timestamp 1486834041
transform 1 0 17696 0 1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_160
timestamp 1486834041
transform 1 0 18592 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_170
timestamp 1486834041
transform 1 0 19712 0 1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_174
timestamp 1486834041
transform 1 0 20160 0 1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_177
timestamp 1486834041
transform 1 0 20496 0 1 18032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_209
timestamp 1486834041
transform 1 0 24080 0 1 18032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_2
timestamp 1486834041
transform 1 0 896 0 -1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_26
timestamp 1486834041
transform 1 0 3584 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_48
timestamp 1486834041
transform 1 0 6048 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_72
timestamp 1486834041
transform 1 0 8736 0 -1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_23_148
timestamp 1486834041
transform 1 0 17248 0 -1 19600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_180
timestamp 1486834041
transform 1 0 20832 0 -1 19600
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_196
timestamp 1486834041
transform 1 0 22624 0 -1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_204
timestamp 1486834041
transform 1 0 23520 0 -1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_208
timestamp 1486834041
transform 1 0 23968 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_212
timestamp 1486834041
transform 1 0 24416 0 -1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_220
timestamp 1486834041
transform 1 0 25312 0 -1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_224
timestamp 1486834041
transform 1 0 25760 0 -1 19600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_30
timestamp 1486834041
transform 1 0 4032 0 1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_34
timestamp 1486834041
transform 1 0 4480 0 1 19600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_37
timestamp 1486834041
transform 1 0 4816 0 1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_41
timestamp 1486834041
transform 1 0 5264 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_91
timestamp 1486834041
transform 1 0 10864 0 1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_122
timestamp 1486834041
transform 1 0 14336 0 1 19600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_141
timestamp 1486834041
transform 1 0 16464 0 1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_149
timestamp 1486834041
transform 1 0 17360 0 1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_173
timestamp 1486834041
transform 1 0 20048 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_177
timestamp 1486834041
transform 1 0 20496 0 1 19600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_209
timestamp 1486834041
transform 1 0 24080 0 1 19600
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_225
timestamp 1486834041
transform 1 0 25872 0 1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_2
timestamp 1486834041
transform 1 0 896 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_4
timestamp 1486834041
transform 1 0 1120 0 -1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_45
timestamp 1486834041
transform 1 0 5712 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_67
timestamp 1486834041
transform 1 0 8176 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_69
timestamp 1486834041
transform 1 0 8400 0 -1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_72
timestamp 1486834041
transform 1 0 8736 0 -1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_76
timestamp 1486834041
transform 1 0 9184 0 -1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_148
timestamp 1486834041
transform 1 0 17248 0 -1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_184
timestamp 1486834041
transform 1 0 21280 0 -1 21168
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_200
timestamp 1486834041
transform 1 0 23072 0 -1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_208
timestamp 1486834041
transform 1 0 23968 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_212
timestamp 1486834041
transform 1 0 24416 0 -1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_220
timestamp 1486834041
transform 1 0 25312 0 -1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_224
timestamp 1486834041
transform 1 0 25760 0 -1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_10
timestamp 1486834041
transform 1 0 1792 0 1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_14
timestamp 1486834041
transform 1 0 2240 0 1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_37
timestamp 1486834041
transform 1 0 4816 0 1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_173
timestamp 1486834041
transform 1 0 20048 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_177
timestamp 1486834041
transform 1 0 20496 0 1 21168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_209
timestamp 1486834041
transform 1 0 24080 0 1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_217
timestamp 1486834041
transform 1 0 24976 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_2
timestamp 1486834041
transform 1 0 896 0 -1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_31
timestamp 1486834041
transform 1 0 4144 0 -1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_35
timestamp 1486834041
transform 1 0 4592 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_69
timestamp 1486834041
transform 1 0 8400 0 -1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_104
timestamp 1486834041
transform 1 0 12320 0 -1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_146
timestamp 1486834041
transform 1 0 17024 0 -1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_27_167
timestamp 1486834041
transform 1 0 19376 0 -1 22736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_199
timestamp 1486834041
transform 1 0 22960 0 -1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_207
timestamp 1486834041
transform 1 0 23856 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_209
timestamp 1486834041
transform 1 0 24080 0 -1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_212
timestamp 1486834041
transform 1 0 24416 0 -1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_2
timestamp 1486834041
transform 1 0 896 0 1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_31
timestamp 1486834041
transform 1 0 4144 0 1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_37
timestamp 1486834041
transform 1 0 4816 0 1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_41
timestamp 1486834041
transform 1 0 5264 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_91
timestamp 1486834041
transform 1 0 10864 0 1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_167
timestamp 1486834041
transform 1 0 19376 0 1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_177
timestamp 1486834041
transform 1 0 20496 0 1 22736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_209
timestamp 1486834041
transform 1 0 24080 0 1 22736
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_225
timestamp 1486834041
transform 1 0 25872 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_10
timestamp 1486834041
transform 1 0 1792 0 -1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_66
timestamp 1486834041
transform 1 0 8064 0 -1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_72
timestamp 1486834041
transform 1 0 8736 0 -1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_84
timestamp 1486834041
transform 1 0 10080 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_86
timestamp 1486834041
transform 1 0 10304 0 -1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_139
timestamp 1486834041
transform 1 0 16240 0 -1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_162
timestamp 1486834041
transform 1 0 18816 0 -1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_29_174
timestamp 1486834041
transform 1 0 20160 0 -1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_206
timestamp 1486834041
transform 1 0 23744 0 -1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_212
timestamp 1486834041
transform 1 0 24416 0 -1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_2
timestamp 1486834041
transform 1 0 896 0 1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_37
timestamp 1486834041
transform 1 0 4816 0 1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_41
timestamp 1486834041
transform 1 0 5264 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_51
timestamp 1486834041
transform 1 0 6384 0 1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_59
timestamp 1486834041
transform 1 0 7280 0 1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_92
timestamp 1486834041
transform 1 0 10976 0 1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_96
timestamp 1486834041
transform 1 0 11424 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_98
timestamp 1486834041
transform 1 0 11648 0 1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_107
timestamp 1486834041
transform 1 0 12656 0 1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_160
timestamp 1486834041
transform 1 0 18592 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_170
timestamp 1486834041
transform 1 0 19712 0 1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_174
timestamp 1486834041
transform 1 0 20160 0 1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_177
timestamp 1486834041
transform 1 0 20496 0 1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_209
timestamp 1486834041
transform 1 0 24080 0 1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_10
timestamp 1486834041
transform 1 0 1792 0 -1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_43
timestamp 1486834041
transform 1 0 5488 0 -1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_67
timestamp 1486834041
transform 1 0 8176 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_69
timestamp 1486834041
transform 1 0 8400 0 -1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_80
timestamp 1486834041
transform 1 0 9632 0 -1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_132
timestamp 1486834041
transform 1 0 15456 0 -1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_142
timestamp 1486834041
transform 1 0 16576 0 -1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_146
timestamp 1486834041
transform 1 0 17024 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_148
timestamp 1486834041
transform 1 0 17248 0 -1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_181
timestamp 1486834041
transform 1 0 20944 0 -1 25872
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_197
timestamp 1486834041
transform 1 0 22736 0 -1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_205
timestamp 1486834041
transform 1 0 23632 0 -1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_209
timestamp 1486834041
transform 1 0 24080 0 -1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_212
timestamp 1486834041
transform 1 0 24416 0 -1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_2
timestamp 1486834041
transform 1 0 896 0 1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_34
timestamp 1486834041
transform 1 0 4480 0 1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_37
timestamp 1486834041
transform 1 0 4816 0 1 25872
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_53
timestamp 1486834041
transform 1 0 6608 0 1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_57
timestamp 1486834041
transform 1 0 7056 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_79
timestamp 1486834041
transform 1 0 9520 0 1 25872
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_95
timestamp 1486834041
transform 1 0 11312 0 1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_103
timestamp 1486834041
transform 1 0 12208 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_115
timestamp 1486834041
transform 1 0 13552 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_117
timestamp 1486834041
transform 1 0 13776 0 1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_126
timestamp 1486834041
transform 1 0 14784 0 1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_134
timestamp 1486834041
transform 1 0 15680 0 1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_158
timestamp 1486834041
transform 1 0 18368 0 1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_162
timestamp 1486834041
transform 1 0 18816 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_172
timestamp 1486834041
transform 1 0 19936 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_174
timestamp 1486834041
transform 1 0 20160 0 1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_177
timestamp 1486834041
transform 1 0 20496 0 1 25872
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_209
timestamp 1486834041
transform 1 0 24080 0 1 25872
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_225
timestamp 1486834041
transform 1 0 25872 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_30
timestamp 1486834041
transform 1 0 4032 0 -1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_34
timestamp 1486834041
transform 1 0 4480 0 -1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_55
timestamp 1486834041
transform 1 0 6832 0 -1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_63
timestamp 1486834041
transform 1 0 7728 0 -1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_67
timestamp 1486834041
transform 1 0 8176 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_69
timestamp 1486834041
transform 1 0 8400 0 -1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_72
timestamp 1486834041
transform 1 0 8736 0 -1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_80
timestamp 1486834041
transform 1 0 9632 0 -1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_142
timestamp 1486834041
transform 1 0 16576 0 -1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_33_170
timestamp 1486834041
transform 1 0 19712 0 -1 27440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_202
timestamp 1486834041
transform 1 0 23296 0 -1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_212
timestamp 1486834041
transform 1 0 24416 0 -1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_10
timestamp 1486834041
transform 1 0 1792 0 1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_14
timestamp 1486834041
transform 1 0 2240 0 1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_69
timestamp 1486834041
transform 1 0 8400 0 1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_107
timestamp 1486834041
transform 1 0 12656 0 1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_111
timestamp 1486834041
transform 1 0 13104 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_113
timestamp 1486834041
transform 1 0 13328 0 1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_146
timestamp 1486834041
transform 1 0 17024 0 1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_177
timestamp 1486834041
transform 1 0 20496 0 1 27440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_209
timestamp 1486834041
transform 1 0 24080 0 1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_72
timestamp 1486834041
transform 1 0 8736 0 -1 29008
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_142
timestamp 1486834041
transform 1 0 16576 0 -1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_150
timestamp 1486834041
transform 1 0 17472 0 -1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_154
timestamp 1486834041
transform 1 0 17920 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_156
timestamp 1486834041
transform 1 0 18144 0 -1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_189
timestamp 1486834041
transform 1 0 21840 0 -1 29008
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_205
timestamp 1486834041
transform 1 0 23632 0 -1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_209
timestamp 1486834041
transform 1 0 24080 0 -1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_212
timestamp 1486834041
transform 1 0 24416 0 -1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_220
timestamp 1486834041
transform 1 0 25312 0 -1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_224
timestamp 1486834041
transform 1 0 25760 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_226
timestamp 1486834041
transform 1 0 25984 0 -1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_30
timestamp 1486834041
transform 1 0 4032 0 1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_34
timestamp 1486834041
transform 1 0 4480 0 1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_57
timestamp 1486834041
transform 1 0 7056 0 1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_65
timestamp 1486834041
transform 1 0 7952 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_87
timestamp 1486834041
transform 1 0 10416 0 1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_95
timestamp 1486834041
transform 1 0 11312 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_107
timestamp 1486834041
transform 1 0 12656 0 1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_111
timestamp 1486834041
transform 1 0 13104 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_173
timestamp 1486834041
transform 1 0 20048 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_177
timestamp 1486834041
transform 1 0 20496 0 1 29008
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_209
timestamp 1486834041
transform 1 0 24080 0 1 29008
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_225
timestamp 1486834041
transform 1 0 25872 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_32
timestamp 1486834041
transform 1 0 4256 0 -1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_36
timestamp 1486834041
transform 1 0 4704 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_72
timestamp 1486834041
transform 1 0 8736 0 -1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_76
timestamp 1486834041
transform 1 0 9184 0 -1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_109
timestamp 1486834041
transform 1 0 12880 0 -1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_117
timestamp 1486834041
transform 1 0 13776 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_127
timestamp 1486834041
transform 1 0 14896 0 -1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_131
timestamp 1486834041
transform 1 0 15344 0 -1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_162
timestamp 1486834041
transform 1 0 18816 0 -1 30576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_194
timestamp 1486834041
transform 1 0 22400 0 -1 30576
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_212
timestamp 1486834041
transform 1 0 24416 0 -1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_220
timestamp 1486834041
transform 1 0 25312 0 -1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_224
timestamp 1486834041
transform 1 0 25760 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_226
timestamp 1486834041
transform 1 0 25984 0 -1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_2
timestamp 1486834041
transform 1 0 896 0 1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_37
timestamp 1486834041
transform 1 0 4816 0 1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_45
timestamp 1486834041
transform 1 0 5712 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_47
timestamp 1486834041
transform 1 0 5936 0 1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_84
timestamp 1486834041
transform 1 0 10080 0 1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_93
timestamp 1486834041
transform 1 0 11088 0 1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_102
timestamp 1486834041
transform 1 0 12096 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_104
timestamp 1486834041
transform 1 0 12320 0 1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_107
timestamp 1486834041
transform 1 0 12656 0 1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_115
timestamp 1486834041
transform 1 0 13552 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_117
timestamp 1486834041
transform 1 0 13776 0 1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_138
timestamp 1486834041
transform 1 0 16128 0 1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_174
timestamp 1486834041
transform 1 0 20160 0 1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_177
timestamp 1486834041
transform 1 0 20496 0 1 30576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_209
timestamp 1486834041
transform 1 0 24080 0 1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_2
timestamp 1486834041
transform 1 0 896 0 -1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_6
timestamp 1486834041
transform 1 0 1344 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_8
timestamp 1486834041
transform 1 0 1568 0 -1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_41
timestamp 1486834041
transform 1 0 5264 0 -1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_49
timestamp 1486834041
transform 1 0 6160 0 -1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_53
timestamp 1486834041
transform 1 0 6608 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_55
timestamp 1486834041
transform 1 0 6832 0 -1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_80
timestamp 1486834041
transform 1 0 9632 0 -1 32144
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_96
timestamp 1486834041
transform 1 0 11424 0 -1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_132
timestamp 1486834041
transform 1 0 15456 0 -1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_39_174
timestamp 1486834041
transform 1 0 20160 0 -1 32144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_206
timestamp 1486834041
transform 1 0 23744 0 -1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_212
timestamp 1486834041
transform 1 0 24416 0 -1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_2
timestamp 1486834041
transform 1 0 896 0 1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_34
timestamp 1486834041
transform 1 0 4480 0 1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_37
timestamp 1486834041
transform 1 0 4816 0 1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_45
timestamp 1486834041
transform 1 0 5712 0 1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_81
timestamp 1486834041
transform 1 0 9744 0 1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_107
timestamp 1486834041
transform 1 0 12656 0 1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_124
timestamp 1486834041
transform 1 0 14560 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_126
timestamp 1486834041
transform 1 0 14784 0 1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_170
timestamp 1486834041
transform 1 0 19712 0 1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_174
timestamp 1486834041
transform 1 0 20160 0 1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_177
timestamp 1486834041
transform 1 0 20496 0 1 32144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_209
timestamp 1486834041
transform 1 0 24080 0 1 32144
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_225
timestamp 1486834041
transform 1 0 25872 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_30
timestamp 1486834041
transform 1 0 4032 0 -1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_38
timestamp 1486834041
transform 1 0 4928 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_40
timestamp 1486834041
transform 1 0 5152 0 -1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_69
timestamp 1486834041
transform 1 0 8400 0 -1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_72
timestamp 1486834041
transform 1 0 8736 0 -1 33712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_96
timestamp 1486834041
transform 1 0 11424 0 -1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_117
timestamp 1486834041
transform 1 0 13776 0 -1 33712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_121
timestamp 1486834041
transform 1 0 14224 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_131
timestamp 1486834041
transform 1 0 15344 0 -1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_139
timestamp 1486834041
transform 1 0 16240 0 -1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_142
timestamp 1486834041
transform 1 0 16576 0 -1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_41_171
timestamp 1486834041
transform 1 0 19824 0 -1 33712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_203
timestamp 1486834041
transform 1 0 23408 0 -1 33712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_207
timestamp 1486834041
transform 1 0 23856 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_209
timestamp 1486834041
transform 1 0 24080 0 -1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_212
timestamp 1486834041
transform 1 0 24416 0 -1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_2
timestamp 1486834041
transform 1 0 896 0 1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_57
timestamp 1486834041
transform 1 0 7056 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_79
timestamp 1486834041
transform 1 0 9520 0 1 33712
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_95
timestamp 1486834041
transform 1 0 11312 0 1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_103
timestamp 1486834041
transform 1 0 12208 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_107
timestamp 1486834041
transform 1 0 12656 0 1 33712
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_123
timestamp 1486834041
transform 1 0 14448 0 1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_174
timestamp 1486834041
transform 1 0 20160 0 1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_177
timestamp 1486834041
transform 1 0 20496 0 1 33712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_209
timestamp 1486834041
transform 1 0 24080 0 1 33712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_10
timestamp 1486834041
transform 1 0 1792 0 -1 35280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_14
timestamp 1486834041
transform 1 0 2240 0 -1 35280
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_35
timestamp 1486834041
transform 1 0 4592 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_37
timestamp 1486834041
transform 1 0 4816 0 -1 35280
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_72
timestamp 1486834041
transform 1 0 8736 0 -1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_80
timestamp 1486834041
transform 1 0 9632 0 -1 35280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_84
timestamp 1486834041
transform 1 0 10080 0 -1 35280
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_137
timestamp 1486834041
transform 1 0 16016 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_139
timestamp 1486834041
transform 1 0 16240 0 -1 35280
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_43_178
timestamp 1486834041
transform 1 0 20608 0 -1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_212
timestamp 1486834041
transform 1 0 24416 0 -1 35280
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_10
timestamp 1486834041
transform 1 0 1792 0 1 35280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_14
timestamp 1486834041
transform 1 0 2240 0 1 35280
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_37
timestamp 1486834041
transform 1 0 4816 0 1 35280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_41
timestamp 1486834041
transform 1 0 5264 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_103
timestamp 1486834041
transform 1 0 12208 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_165
timestamp 1486834041
transform 1 0 19152 0 1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_173
timestamp 1486834041
transform 1 0 20048 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_177
timestamp 1486834041
transform 1 0 20496 0 1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_209
timestamp 1486834041
transform 1 0 24080 0 1 35280
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_225
timestamp 1486834041
transform 1 0 25872 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_42
timestamp 1486834041
transform 1 0 5376 0 -1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_46
timestamp 1486834041
transform 1 0 5824 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_56
timestamp 1486834041
transform 1 0 6944 0 -1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_60
timestamp 1486834041
transform 1 0 7392 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_92
timestamp 1486834041
transform 1 0 10976 0 -1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_139
timestamp 1486834041
transform 1 0 16240 0 -1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_45_164
timestamp 1486834041
transform 1 0 19040 0 -1 36848
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_196
timestamp 1486834041
transform 1 0 22624 0 -1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_204
timestamp 1486834041
transform 1 0 23520 0 -1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_208
timestamp 1486834041
transform 1 0 23968 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_212
timestamp 1486834041
transform 1 0 24416 0 -1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_26
timestamp 1486834041
transform 1 0 3584 0 1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_34
timestamp 1486834041
transform 1 0 4480 0 1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_57
timestamp 1486834041
transform 1 0 7056 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_59
timestamp 1486834041
transform 1 0 7280 0 1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_92
timestamp 1486834041
transform 1 0 10976 0 1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_100
timestamp 1486834041
transform 1 0 11872 0 1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_104
timestamp 1486834041
transform 1 0 12320 0 1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_107
timestamp 1486834041
transform 1 0 12656 0 1 36848
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_123
timestamp 1486834041
transform 1 0 14448 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_46_177
timestamp 1486834041
transform 1 0 20496 0 1 36848
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_209
timestamp 1486834041
transform 1 0 24080 0 1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_30
timestamp 1486834041
transform 1 0 4032 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_32
timestamp 1486834041
transform 1 0 4256 0 -1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_61
timestamp 1486834041
transform 1 0 7504 0 -1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_72
timestamp 1486834041
transform 1 0 8736 0 -1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_134
timestamp 1486834041
transform 1 0 15680 0 -1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_138
timestamp 1486834041
transform 1 0 16128 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_178
timestamp 1486834041
transform 1 0 20608 0 -1 38416
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_212
timestamp 1486834041
transform 1 0 24416 0 -1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_10
timestamp 1486834041
transform 1 0 1792 0 1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_14
timestamp 1486834041
transform 1 0 2240 0 1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_37
timestamp 1486834041
transform 1 0 4816 0 1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_61
timestamp 1486834041
transform 1 0 7504 0 1 38416
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_77
timestamp 1486834041
transform 1 0 9296 0 1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_107
timestamp 1486834041
transform 1 0 12656 0 1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_116
timestamp 1486834041
transform 1 0 13664 0 1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_124
timestamp 1486834041
transform 1 0 14560 0 1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_48_177
timestamp 1486834041
transform 1 0 20496 0 1 38416
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_209
timestamp 1486834041
transform 1 0 24080 0 1 38416
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_225
timestamp 1486834041
transform 1 0 25872 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_18
timestamp 1486834041
transform 1 0 2688 0 -1 39984
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_34
timestamp 1486834041
transform 1 0 4480 0 -1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_72
timestamp 1486834041
transform 1 0 8736 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_74
timestamp 1486834041
transform 1 0 8960 0 -1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_127
timestamp 1486834041
transform 1 0 14896 0 -1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_135
timestamp 1486834041
transform 1 0 15792 0 -1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_139
timestamp 1486834041
transform 1 0 16240 0 -1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_192
timestamp 1486834041
transform 1 0 22176 0 -1 39984
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_208
timestamp 1486834041
transform 1 0 23968 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_212
timestamp 1486834041
transform 1 0 24416 0 -1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_2
timestamp 1486834041
transform 1 0 896 0 1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_6
timestamp 1486834041
transform 1 0 1344 0 1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_37
timestamp 1486834041
transform 1 0 4816 0 1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_45
timestamp 1486834041
transform 1 0 5712 0 1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_49
timestamp 1486834041
transform 1 0 6160 0 1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_90
timestamp 1486834041
transform 1 0 10752 0 1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_98
timestamp 1486834041
transform 1 0 11648 0 1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_102
timestamp 1486834041
transform 1 0 12096 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_104
timestamp 1486834041
transform 1 0 12320 0 1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_107
timestamp 1486834041
transform 1 0 12656 0 1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_116
timestamp 1486834041
transform 1 0 13664 0 1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_124
timestamp 1486834041
transform 1 0 14560 0 1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_161
timestamp 1486834041
transform 1 0 18704 0 1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_169
timestamp 1486834041
transform 1 0 19600 0 1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_173
timestamp 1486834041
transform 1 0 20048 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_177
timestamp 1486834041
transform 1 0 20496 0 1 39984
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_209
timestamp 1486834041
transform 1 0 24080 0 1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_10
timestamp 1486834041
transform 1 0 1792 0 -1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_19
timestamp 1486834041
transform 1 0 2800 0 -1 41552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_23
timestamp 1486834041
transform 1 0 3248 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_25
timestamp 1486834041
transform 1 0 3472 0 -1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_46
timestamp 1486834041
transform 1 0 5824 0 -1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_55
timestamp 1486834041
transform 1 0 6832 0 -1 41552
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_63
timestamp 1486834041
transform 1 0 7728 0 -1 41552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_67
timestamp 1486834041
transform 1 0 8176 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_69
timestamp 1486834041
transform 1 0 8400 0 -1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_80
timestamp 1486834041
transform 1 0 9632 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_51_102
timestamp 1486834041
transform 1 0 12096 0 -1 41552
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_134
timestamp 1486834041
transform 1 0 15680 0 -1 41552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_138
timestamp 1486834041
transform 1 0 16128 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_142
timestamp 1486834041
transform 1 0 16576 0 -1 41552
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_206
timestamp 1486834041
transform 1 0 23744 0 -1 41552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_212
timestamp 1486834041
transform 1 0 24416 0 -1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_10
timestamp 1486834041
transform 1 0 1792 0 1 41552
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_18
timestamp 1486834041
transform 1 0 2688 0 1 41552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_22
timestamp 1486834041
transform 1 0 3136 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_24
timestamp 1486834041
transform 1 0 3360 0 1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_33
timestamp 1486834041
transform 1 0 4368 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_37
timestamp 1486834041
transform 1 0 4816 0 1 41552
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_101
timestamp 1486834041
transform 1 0 11984 0 1 41552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_107
timestamp 1486834041
transform 1 0 12656 0 1 41552
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_123
timestamp 1486834041
transform 1 0 14448 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_52_177
timestamp 1486834041
transform 1 0 20496 0 1 41552
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_209
timestamp 1486834041
transform 1 0 24080 0 1 41552
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_225
timestamp 1486834041
transform 1 0 25872 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_53_10
timestamp 1486834041
transform 1 0 1792 0 -1 43120
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_42
timestamp 1486834041
transform 1 0 5376 0 -1 43120
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_58
timestamp 1486834041
transform 1 0 7168 0 -1 43120
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_66
timestamp 1486834041
transform 1 0 8064 0 -1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_72
timestamp 1486834041
transform 1 0 8736 0 -1 43120
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_136
timestamp 1486834041
transform 1 0 15904 0 -1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_142
timestamp 1486834041
transform 1 0 16576 0 -1 43120
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_206
timestamp 1486834041
transform 1 0 23744 0 -1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_212
timestamp 1486834041
transform 1 0 24416 0 -1 43120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_10
timestamp 1486834041
transform 1 0 1792 0 1 43120
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_26
timestamp 1486834041
transform 1 0 3584 0 1 43120
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_34
timestamp 1486834041
transform 1 0 4480 0 1 43120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_37
timestamp 1486834041
transform 1 0 4816 0 1 43120
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_101
timestamp 1486834041
transform 1 0 11984 0 1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_107
timestamp 1486834041
transform 1 0 12656 0 1 43120
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_171
timestamp 1486834041
transform 1 0 19824 0 1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_177
timestamp 1486834041
transform 1 0 20496 0 1 43120
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_209
timestamp 1486834041
transform 1 0 24080 0 1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_55_10
timestamp 1486834041
transform 1 0 1792 0 -1 44688
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_42
timestamp 1486834041
transform 1 0 5376 0 -1 44688
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_58
timestamp 1486834041
transform 1 0 7168 0 -1 44688
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_66
timestamp 1486834041
transform 1 0 8064 0 -1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_72
timestamp 1486834041
transform 1 0 8736 0 -1 44688
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_136
timestamp 1486834041
transform 1 0 15904 0 -1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_142
timestamp 1486834041
transform 1 0 16576 0 -1 44688
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_206
timestamp 1486834041
transform 1 0 23744 0 -1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_212
timestamp 1486834041
transform 1 0 24416 0 -1 44688
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_56_2
timestamp 1486834041
transform 1 0 896 0 1 44688
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_34
timestamp 1486834041
transform 1 0 4480 0 1 44688
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_37
timestamp 1486834041
transform 1 0 4816 0 1 44688
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_101
timestamp 1486834041
transform 1 0 11984 0 1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_107
timestamp 1486834041
transform 1 0 12656 0 1 44688
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_171
timestamp 1486834041
transform 1 0 19824 0 1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_56_177
timestamp 1486834041
transform 1 0 20496 0 1 44688
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_56_209
timestamp 1486834041
transform 1 0 24080 0 1 44688
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_225
timestamp 1486834041
transform 1 0 25872 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_57_10
timestamp 1486834041
transform 1 0 1792 0 -1 46256
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_57_42
timestamp 1486834041
transform 1 0 5376 0 -1 46256
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_57_58
timestamp 1486834041
transform 1 0 7168 0 -1 46256
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_66
timestamp 1486834041
transform 1 0 8064 0 -1 46256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_72
timestamp 1486834041
transform 1 0 8736 0 -1 46256
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_136
timestamp 1486834041
transform 1 0 15904 0 -1 46256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_142
timestamp 1486834041
transform 1 0 16576 0 -1 46256
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_206
timestamp 1486834041
transform 1 0 23744 0 -1 46256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_212
timestamp 1486834041
transform 1 0 24416 0 -1 46256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_58_2
timestamp 1486834041
transform 1 0 896 0 1 46256
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_34
timestamp 1486834041
transform 1 0 4480 0 1 46256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_37
timestamp 1486834041
transform 1 0 4816 0 1 46256
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_101
timestamp 1486834041
transform 1 0 11984 0 1 46256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_107
timestamp 1486834041
transform 1 0 12656 0 1 46256
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_171
timestamp 1486834041
transform 1 0 19824 0 1 46256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_58_177
timestamp 1486834041
transform 1 0 20496 0 1 46256
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_209
timestamp 1486834041
transform 1 0 24080 0 1 46256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_59_10
timestamp 1486834041
transform 1 0 1792 0 -1 47824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_59_42
timestamp 1486834041
transform 1 0 5376 0 -1 47824
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_59_58
timestamp 1486834041
transform 1 0 7168 0 -1 47824
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_66
timestamp 1486834041
transform 1 0 8064 0 -1 47824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_72
timestamp 1486834041
transform 1 0 8736 0 -1 47824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_136
timestamp 1486834041
transform 1 0 15904 0 -1 47824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_142
timestamp 1486834041
transform 1 0 16576 0 -1 47824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_206
timestamp 1486834041
transform 1 0 23744 0 -1 47824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_212
timestamp 1486834041
transform 1 0 24416 0 -1 47824
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_2
timestamp 1486834041
transform 1 0 896 0 1 47824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_34
timestamp 1486834041
transform 1 0 4480 0 1 47824
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_37
timestamp 1486834041
transform 1 0 4816 0 1 47824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_101
timestamp 1486834041
transform 1 0 11984 0 1 47824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_107
timestamp 1486834041
transform 1 0 12656 0 1 47824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_171
timestamp 1486834041
transform 1 0 19824 0 1 47824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_177
timestamp 1486834041
transform 1 0 20496 0 1 47824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_209
timestamp 1486834041
transform 1 0 24080 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_61_10
timestamp 1486834041
transform 1 0 1792 0 -1 49392
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_61_42
timestamp 1486834041
transform 1 0 5376 0 -1 49392
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_58
timestamp 1486834041
transform 1 0 7168 0 -1 49392
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_66
timestamp 1486834041
transform 1 0 8064 0 -1 49392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_72
timestamp 1486834041
transform 1 0 8736 0 -1 49392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_136
timestamp 1486834041
transform 1 0 15904 0 -1 49392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_142
timestamp 1486834041
transform 1 0 16576 0 -1 49392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_206
timestamp 1486834041
transform 1 0 23744 0 -1 49392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_212
timestamp 1486834041
transform 1 0 24416 0 -1 49392
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_62_10
timestamp 1486834041
transform 1 0 1792 0 1 49392
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_26
timestamp 1486834041
transform 1 0 3584 0 1 49392
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_34
timestamp 1486834041
transform 1 0 4480 0 1 49392
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_37
timestamp 1486834041
transform 1 0 4816 0 1 49392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_101
timestamp 1486834041
transform 1 0 11984 0 1 49392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_107
timestamp 1486834041
transform 1 0 12656 0 1 49392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_171
timestamp 1486834041
transform 1 0 19824 0 1 49392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_62_177
timestamp 1486834041
transform 1 0 20496 0 1 49392
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_193
timestamp 1486834041
transform 1 0 22288 0 1 49392
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_201
timestamp 1486834041
transform 1 0 23184 0 1 49392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_2
timestamp 1486834041
transform 1 0 896 0 -1 50960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_66
timestamp 1486834041
transform 1 0 8064 0 -1 50960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_72
timestamp 1486834041
transform 1 0 8736 0 -1 50960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_136
timestamp 1486834041
transform 1 0 15904 0 -1 50960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_63_142
timestamp 1486834041
transform 1 0 16576 0 -1 50960
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_63_174
timestamp 1486834041
transform 1 0 20160 0 -1 50960
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_190
timestamp 1486834041
transform 1 0 21952 0 -1 50960
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_198
timestamp 1486834041
transform 1 0 22848 0 -1 50960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_212
timestamp 1486834041
transform 1 0 24416 0 -1 50960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_64_10
timestamp 1486834041
transform 1 0 1792 0 1 50960
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_26
timestamp 1486834041
transform 1 0 3584 0 1 50960
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_34
timestamp 1486834041
transform 1 0 4480 0 1 50960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_37
timestamp 1486834041
transform 1 0 4816 0 1 50960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_101
timestamp 1486834041
transform 1 0 11984 0 1 50960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_107
timestamp 1486834041
transform 1 0 12656 0 1 50960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_171
timestamp 1486834041
transform 1 0 19824 0 1 50960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_64_177
timestamp 1486834041
transform 1 0 20496 0 1 50960
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_193
timestamp 1486834041
transform 1 0 22288 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_195
timestamp 1486834041
transform 1 0 22512 0 1 50960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_204
timestamp 1486834041
transform 1 0 23520 0 1 50960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_2
timestamp 1486834041
transform 1 0 896 0 -1 52528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_66
timestamp 1486834041
transform 1 0 8064 0 -1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_72
timestamp 1486834041
transform 1 0 8736 0 -1 52528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_136
timestamp 1486834041
transform 1 0 15904 0 -1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_65_142
timestamp 1486834041
transform 1 0 16576 0 -1 52528
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_174
timestamp 1486834041
transform 1 0 20160 0 -1 52528
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_182
timestamp 1486834041
transform 1 0 21056 0 -1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_186
timestamp 1486834041
transform 1 0 21504 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_212
timestamp 1486834041
transform 1 0 24416 0 -1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_10
timestamp 1486834041
transform 1 0 1792 0 1 52528
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_26
timestamp 1486834041
transform 1 0 3584 0 1 52528
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_34
timestamp 1486834041
transform 1 0 4480 0 1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_37
timestamp 1486834041
transform 1 0 4816 0 1 52528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_101
timestamp 1486834041
transform 1 0 11984 0 1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_107
timestamp 1486834041
transform 1 0 12656 0 1 52528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_171
timestamp 1486834041
transform 1 0 19824 0 1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_177
timestamp 1486834041
transform 1 0 20496 0 1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_181
timestamp 1486834041
transform 1 0 20944 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_10
timestamp 1486834041
transform 1 0 1792 0 -1 54096
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_42
timestamp 1486834041
transform 1 0 5376 0 -1 54096
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_58
timestamp 1486834041
transform 1 0 7168 0 -1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_66
timestamp 1486834041
transform 1 0 8064 0 -1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_72
timestamp 1486834041
transform 1 0 8736 0 -1 54096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_136
timestamp 1486834041
transform 1 0 15904 0 -1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_142
timestamp 1486834041
transform 1 0 16576 0 -1 54096
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_158
timestamp 1486834041
transform 1 0 18368 0 -1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_166
timestamp 1486834041
transform 1 0 19264 0 -1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_170
timestamp 1486834041
transform 1 0 19712 0 -1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_195
timestamp 1486834041
transform 1 0 22512 0 -1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_212
timestamp 1486834041
transform 1 0 24416 0 -1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_68_2
timestamp 1486834041
transform 1 0 896 0 1 54096
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_34
timestamp 1486834041
transform 1 0 4480 0 1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_37
timestamp 1486834041
transform 1 0 4816 0 1 54096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_101
timestamp 1486834041
transform 1 0 11984 0 1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_68_107
timestamp 1486834041
transform 1 0 12656 0 1 54096
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_68_139
timestamp 1486834041
transform 1 0 16240 0 1 54096
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_155
timestamp 1486834041
transform 1 0 18032 0 1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_159
timestamp 1486834041
transform 1 0 18480 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_161
timestamp 1486834041
transform 1 0 18704 0 1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_170
timestamp 1486834041
transform 1 0 19712 0 1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_174
timestamp 1486834041
transform 1 0 20160 0 1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_69_2
timestamp 1486834041
transform 1 0 896 0 -1 55664
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_10
timestamp 1486834041
transform 1 0 1792 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_12
timestamp 1486834041
transform 1 0 2016 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_69_27
timestamp 1486834041
transform 1 0 3696 0 -1 55664
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_43
timestamp 1486834041
transform 1 0 5488 0 -1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_47
timestamp 1486834041
transform 1 0 5936 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_63
timestamp 1486834041
transform 1 0 7728 0 -1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_67
timestamp 1486834041
transform 1 0 8176 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_69
timestamp 1486834041
transform 1 0 8400 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_69_72
timestamp 1486834041
transform 1 0 8736 0 -1 55664
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_69_88
timestamp 1486834041
transform 1 0 10528 0 -1 55664
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_96
timestamp 1486834041
transform 1 0 11424 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_69_111
timestamp 1486834041
transform 1 0 13104 0 -1 55664
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_69_127
timestamp 1486834041
transform 1 0 14896 0 -1 55664
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_135
timestamp 1486834041
transform 1 0 15792 0 -1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_139
timestamp 1486834041
transform 1 0 16240 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_142
timestamp 1486834041
transform 1 0 16576 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_144
timestamp 1486834041
transform 1 0 16800 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_159
timestamp 1486834041
transform 1 0 18480 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_169
timestamp 1486834041
transform 1 0 19600 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_207
timestamp 1486834041
transform 1 0 23856 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_209
timestamp 1486834041
transform 1 0 24080 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_212
timestamp 1486834041
transform 1 0 24416 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_70_8
timestamp 1486834041
transform 1 0 1568 0 1 55664
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_16
timestamp 1486834041
transform 1 0 2464 0 1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_36
timestamp 1486834041
transform 1 0 4704 0 1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_51
timestamp 1486834041
transform 1 0 6384 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_53
timestamp 1486834041
transform 1 0 6608 0 1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_70
timestamp 1486834041
transform 1 0 8512 0 1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_99
timestamp 1486834041
transform 1 0 11760 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_101
timestamp 1486834041
transform 1 0 11984 0 1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_104
timestamp 1486834041
transform 1 0 12320 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_106
timestamp 1486834041
transform 1 0 12544 0 1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_135
timestamp 1486834041
transform 1 0 15792 0 1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_152
timestamp 1486834041
transform 1 0 17696 0 1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_200
timestamp 1486834041
transform 1 0 23072 0 1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_234
timestamp 1486834041
transform 1 0 26880 0 1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_240
timestamp 1486834041
transform 1 0 27552 0 1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input1
timestamp 1486834041
transform 1 0 896 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input2
timestamp 1486834041
transform 1 0 896 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input3
timestamp 1486834041
transform 1 0 896 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input4
timestamp 1486834041
transform 1 0 896 0 -1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input5
timestamp 1486834041
transform 1 0 896 0 -1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input6
timestamp 1486834041
transform 1 0 3136 0 1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input7
timestamp 1486834041
transform 1 0 896 0 1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input8
timestamp 1486834041
transform 1 0 3360 0 -1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input9
timestamp 1486834041
transform 1 0 896 0 -1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input10
timestamp 1486834041
transform 1 0 896 0 1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input11
timestamp 1486834041
transform 1 0 896 0 1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input12
timestamp 1486834041
transform 1 0 896 0 1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input13
timestamp 1486834041
transform 1 0 896 0 -1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input14
timestamp 1486834041
transform 1 0 896 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input15
timestamp 1486834041
transform 1 0 896 0 -1 41552
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input16
timestamp 1486834041
transform 1 0 896 0 1 41552
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input17
timestamp 1486834041
transform 1 0 896 0 -1 43120
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input18
timestamp 1486834041
transform 1 0 896 0 1 43120
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input19
timestamp 1486834041
transform 1 0 896 0 -1 44688
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input20
timestamp 1486834041
transform 1 0 896 0 -1 46256
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input21
timestamp 1486834041
transform 1 0 896 0 -1 47824
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input22
timestamp 1486834041
transform 1 0 896 0 -1 49392
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input23
timestamp 1486834041
transform 1 0 896 0 1 49392
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input24
timestamp 1486834041
transform 1 0 896 0 1 50960
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input25
timestamp 1486834041
transform 1 0 1792 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input26
timestamp 1486834041
transform 1 0 896 0 1 52528
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input27
timestamp 1486834041
transform 1 0 896 0 -1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input28
timestamp 1486834041
transform 1 0 896 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input29
timestamp 1486834041
transform 1 0 1792 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input30
timestamp 1486834041
transform 1 0 896 0 -1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input31
timestamp 1486834041
transform 1 0 1792 0 1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input32
timestamp 1486834041
transform 1 0 896 0 1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input33
timestamp 1486834041
transform 1 0 896 0 -1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input34
timestamp 1486834041
transform 1 0 896 0 1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input35
timestamp 1486834041
transform 1 0 4816 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input36
timestamp 1486834041
transform 1 0 6160 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input37
timestamp 1486834041
transform -1 0 26432 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input38
timestamp 1486834041
transform -1 0 25536 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input39
timestamp 1486834041
transform -1 0 27328 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input40
timestamp 1486834041
transform -1 0 26768 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input41
timestamp 1486834041
transform -1 0 27664 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input42
timestamp 1486834041
transform -1 0 26768 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input43
timestamp 1486834041
transform -1 0 27664 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input44
timestamp 1486834041
transform -1 0 27664 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input45
timestamp 1486834041
transform -1 0 26768 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input46
timestamp 1486834041
transform -1 0 27664 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input47
timestamp 1486834041
transform -1 0 26768 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input48
timestamp 1486834041
transform -1 0 27664 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input49
timestamp 1486834041
transform -1 0 26768 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input50
timestamp 1486834041
transform -1 0 27664 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input51
timestamp 1486834041
transform -1 0 26768 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input52
timestamp 1486834041
transform -1 0 27664 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input53
timestamp 1486834041
transform -1 0 27664 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input54
timestamp 1486834041
transform -1 0 26768 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input55
timestamp 1486834041
transform -1 0 27664 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input56
timestamp 1486834041
transform -1 0 26768 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input57
timestamp 1486834041
transform -1 0 27664 0 -1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input58
timestamp 1486834041
transform -1 0 26096 0 1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input59
timestamp 1486834041
transform -1 0 27664 0 -1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input60
timestamp 1486834041
transform -1 0 26768 0 -1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input61
timestamp 1486834041
transform -1 0 27664 0 1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input62
timestamp 1486834041
transform -1 0 26768 0 1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input63
timestamp 1486834041
transform -1 0 27664 0 -1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input64
timestamp 1486834041
transform -1 0 26768 0 -1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input65
timestamp 1486834041
transform -1 0 27664 0 1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input66
timestamp 1486834041
transform -1 0 27664 0 -1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input67
timestamp 1486834041
transform -1 0 26768 0 -1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input68
timestamp 1486834041
transform -1 0 27664 0 1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input69
timestamp 1486834041
transform -1 0 26768 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input70
timestamp 1486834041
transform -1 0 26768 0 -1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input71
timestamp 1486834041
transform -1 0 27664 0 1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input72
timestamp 1486834041
transform -1 0 26768 0 1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input73
timestamp 1486834041
transform -1 0 27664 0 -1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input74
timestamp 1486834041
transform -1 0 26768 0 -1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input75
timestamp 1486834041
transform -1 0 27664 0 1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input76
timestamp 1486834041
transform -1 0 27664 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input77
timestamp 1486834041
transform -1 0 27664 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input78
timestamp 1486834041
transform -1 0 26768 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input79
timestamp 1486834041
transform -1 0 27664 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input80
timestamp 1486834041
transform -1 0 26768 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input81
timestamp 1486834041
transform -1 0 27664 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input82
timestamp 1486834041
transform -1 0 26768 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input83
timestamp 1486834041
transform -1 0 27664 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input84
timestamp 1486834041
transform -1 0 27664 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output85
timestamp 1486834041
transform -1 0 2464 0 1 5488
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output86
timestamp 1486834041
transform -1 0 2464 0 -1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output87
timestamp 1486834041
transform -1 0 2464 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output88
timestamp 1486834041
transform -1 0 2464 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output89
timestamp 1486834041
transform 1 0 24528 0 -1 22736
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output90
timestamp 1486834041
transform 1 0 26096 0 1 21168
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output91
timestamp 1486834041
transform 1 0 26096 0 -1 22736
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output92
timestamp 1486834041
transform 1 0 24528 0 -1 24304
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output93
timestamp 1486834041
transform 1 0 26096 0 1 22736
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output94
timestamp 1486834041
transform 1 0 24528 0 1 24304
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output95
timestamp 1486834041
transform 1 0 26096 0 -1 24304
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output96
timestamp 1486834041
transform 1 0 24528 0 -1 25872
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output97
timestamp 1486834041
transform 1 0 26096 0 1 24304
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output98
timestamp 1486834041
transform 1 0 26096 0 -1 25872
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output99
timestamp 1486834041
transform 1 0 24528 0 -1 27440
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output100
timestamp 1486834041
transform 1 0 26096 0 1 25872
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output101
timestamp 1486834041
transform 1 0 24528 0 1 27440
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output102
timestamp 1486834041
transform 1 0 26096 0 -1 27440
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output103
timestamp 1486834041
transform 1 0 26096 0 1 27440
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output104
timestamp 1486834041
transform 1 0 26096 0 -1 29008
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output105
timestamp 1486834041
transform 1 0 26096 0 1 29008
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output106
timestamp 1486834041
transform 1 0 26096 0 -1 30576
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output107
timestamp 1486834041
transform 1 0 26096 0 1 30576
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output108
timestamp 1486834041
transform 1 0 26096 0 -1 32144
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output109
timestamp 1486834041
transform 1 0 24528 0 -1 38416
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output110
timestamp 1486834041
transform 1 0 24528 0 -1 43120
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output111
timestamp 1486834041
transform 1 0 26096 0 -1 44688
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output112
timestamp 1486834041
transform 1 0 26096 0 -1 39984
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output113
timestamp 1486834041
transform 1 0 26096 0 1 39984
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output114
timestamp 1486834041
transform 1 0 24528 0 -1 39984
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output115
timestamp 1486834041
transform 1 0 26096 0 -1 41552
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output116
timestamp 1486834041
transform 1 0 24528 0 1 39984
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output117
timestamp 1486834041
transform 1 0 26096 0 1 41552
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output118
timestamp 1486834041
transform 1 0 24528 0 -1 41552
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output119
timestamp 1486834041
transform 1 0 26096 0 -1 43120
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output120
timestamp 1486834041
transform 1 0 26096 0 1 43120
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output121
timestamp 1486834041
transform 1 0 24528 0 1 30576
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output122
timestamp 1486834041
transform 1 0 26096 0 -1 36848
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output123
timestamp 1486834041
transform 1 0 26096 0 1 36848
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output124
timestamp 1486834041
transform 1 0 24528 0 -1 36848
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output125
timestamp 1486834041
transform 1 0 26096 0 -1 38416
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output126
timestamp 1486834041
transform 1 0 24528 0 1 36848
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output127
timestamp 1486834041
transform 1 0 26096 0 1 38416
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output128
timestamp 1486834041
transform 1 0 26096 0 1 32144
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output129
timestamp 1486834041
transform 1 0 24528 0 -1 32144
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output130
timestamp 1486834041
transform 1 0 26096 0 -1 33712
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output131
timestamp 1486834041
transform 1 0 26096 0 1 33712
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output132
timestamp 1486834041
transform 1 0 24528 0 -1 33712
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output133
timestamp 1486834041
transform 1 0 26096 0 -1 35280
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output134
timestamp 1486834041
transform 1 0 24528 0 1 33712
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output135
timestamp 1486834041
transform 1 0 26096 0 1 35280
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output136
timestamp 1486834041
transform 1 0 24528 0 -1 35280
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output137
timestamp 1486834041
transform 1 0 24528 0 1 43120
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output138
timestamp 1486834041
transform 1 0 26096 0 -1 49392
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output139
timestamp 1486834041
transform 1 0 26096 0 1 49392
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output140
timestamp 1486834041
transform 1 0 24528 0 -1 49392
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output141
timestamp 1486834041
transform 1 0 26096 0 -1 50960
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output142
timestamp 1486834041
transform 1 0 24528 0 1 49392
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output143
timestamp 1486834041
transform 1 0 26096 0 1 50960
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output144
timestamp 1486834041
transform 1 0 24528 0 -1 50960
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output145
timestamp 1486834041
transform 1 0 26096 0 -1 52528
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output146
timestamp 1486834041
transform 1 0 26096 0 1 52528
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output147
timestamp 1486834041
transform 1 0 24528 0 -1 52528
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output148
timestamp 1486834041
transform 1 0 26096 0 1 44688
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output149
timestamp 1486834041
transform 1 0 26096 0 -1 54096
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output150
timestamp 1486834041
transform 1 0 24528 0 1 52528
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output151
timestamp 1486834041
transform 1 0 26096 0 1 54096
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output152
timestamp 1486834041
transform 1 0 24528 0 -1 54096
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output153
timestamp 1486834041
transform 1 0 26096 0 -1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output154
timestamp 1486834041
transform 1 0 24528 0 -1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output155
timestamp 1486834041
transform 1 0 22960 0 1 54096
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output156
timestamp 1486834041
transform 1 0 22624 0 -1 54096
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output157
timestamp 1486834041
transform 1 0 20720 0 -1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output158
timestamp 1486834041
transform 1 0 21392 0 1 54096
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output159
timestamp 1486834041
transform 1 0 24528 0 -1 44688
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output160
timestamp 1486834041
transform 1 0 24528 0 1 50960
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output161
timestamp 1486834041
transform 1 0 22960 0 1 52528
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output162
timestamp 1486834041
transform 1 0 26096 0 -1 46256
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output163
timestamp 1486834041
transform 1 0 26096 0 1 46256
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output164
timestamp 1486834041
transform 1 0 24528 0 -1 46256
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output165
timestamp 1486834041
transform 1 0 26096 0 -1 47824
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output166
timestamp 1486834041
transform 1 0 24528 0 1 46256
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output167
timestamp 1486834041
transform 1 0 26096 0 1 47824
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output168
timestamp 1486834041
transform 1 0 24528 0 -1 47824
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output169
timestamp 1486834041
transform -1 0 3696 0 -1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output170
timestamp 1486834041
transform -1 0 17696 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output171
timestamp 1486834041
transform -1 0 18480 0 -1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output172
timestamp 1486834041
transform -1 0 19712 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output173
timestamp 1486834041
transform 1 0 19936 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output174
timestamp 1486834041
transform -1 0 23072 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output175
timestamp 1486834041
transform -1 0 23856 0 -1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output176
timestamp 1486834041
transform 1 0 23744 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output177
timestamp 1486834041
transform 1 0 25312 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output178
timestamp 1486834041
transform 1 0 24528 0 1 54096
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output179
timestamp 1486834041
transform 1 0 22624 0 -1 52528
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output180
timestamp 1486834041
transform 1 0 2912 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output181
timestamp 1486834041
transform 1 0 4816 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output182
timestamp 1486834041
transform -1 0 7728 0 -1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output183
timestamp 1486834041
transform -1 0 8288 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output184
timestamp 1486834041
transform -1 0 10192 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output185
timestamp 1486834041
transform -1 0 11760 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output186
timestamp 1486834041
transform -1 0 13104 0 -1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output187
timestamp 1486834041
transform -1 0 14224 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output188
timestamp 1486834041
transform -1 0 15792 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output189
timestamp 1486834041
transform -1 0 1568 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_71
timestamp 1486834041
transform 1 0 672 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1486834041
transform -1 0 27888 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_72
timestamp 1486834041
transform 1 0 672 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1486834041
transform -1 0 27888 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_73
timestamp 1486834041
transform 1 0 672 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1486834041
transform -1 0 27888 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_74
timestamp 1486834041
transform 1 0 672 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1486834041
transform -1 0 27888 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_75
timestamp 1486834041
transform 1 0 672 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1486834041
transform -1 0 27888 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_76
timestamp 1486834041
transform 1 0 672 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1486834041
transform -1 0 27888 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_77
timestamp 1486834041
transform 1 0 672 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1486834041
transform -1 0 27888 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_78
timestamp 1486834041
transform 1 0 672 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1486834041
transform -1 0 27888 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_79
timestamp 1486834041
transform 1 0 672 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1486834041
transform -1 0 27888 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_80
timestamp 1486834041
transform 1 0 672 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1486834041
transform -1 0 27888 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_81
timestamp 1486834041
transform 1 0 672 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1486834041
transform -1 0 27888 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_82
timestamp 1486834041
transform 1 0 672 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1486834041
transform -1 0 27888 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_83
timestamp 1486834041
transform 1 0 672 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1486834041
transform -1 0 27888 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_84
timestamp 1486834041
transform 1 0 672 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1486834041
transform -1 0 27888 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_85
timestamp 1486834041
transform 1 0 672 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1486834041
transform -1 0 27888 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_86
timestamp 1486834041
transform 1 0 672 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1486834041
transform -1 0 27888 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_87
timestamp 1486834041
transform 1 0 672 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1486834041
transform -1 0 27888 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_88
timestamp 1486834041
transform 1 0 672 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1486834041
transform -1 0 27888 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_89
timestamp 1486834041
transform 1 0 672 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1486834041
transform -1 0 27888 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_90
timestamp 1486834041
transform 1 0 672 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1486834041
transform -1 0 27888 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_91
timestamp 1486834041
transform 1 0 672 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1486834041
transform -1 0 27888 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_92
timestamp 1486834041
transform 1 0 672 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1486834041
transform -1 0 27888 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_93
timestamp 1486834041
transform 1 0 672 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1486834041
transform -1 0 27888 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_94
timestamp 1486834041
transform 1 0 672 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1486834041
transform -1 0 27888 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_95
timestamp 1486834041
transform 1 0 672 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1486834041
transform -1 0 27888 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_96
timestamp 1486834041
transform 1 0 672 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1486834041
transform -1 0 27888 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_97
timestamp 1486834041
transform 1 0 672 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1486834041
transform -1 0 27888 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_98
timestamp 1486834041
transform 1 0 672 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1486834041
transform -1 0 27888 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_99
timestamp 1486834041
transform 1 0 672 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1486834041
transform -1 0 27888 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_100
timestamp 1486834041
transform 1 0 672 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1486834041
transform -1 0 27888 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_101
timestamp 1486834041
transform 1 0 672 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1486834041
transform -1 0 27888 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_102
timestamp 1486834041
transform 1 0 672 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1486834041
transform -1 0 27888 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_103
timestamp 1486834041
transform 1 0 672 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1486834041
transform -1 0 27888 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_104
timestamp 1486834041
transform 1 0 672 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1486834041
transform -1 0 27888 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_105
timestamp 1486834041
transform 1 0 672 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1486834041
transform -1 0 27888 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_106
timestamp 1486834041
transform 1 0 672 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1486834041
transform -1 0 27888 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_107
timestamp 1486834041
transform 1 0 672 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1486834041
transform -1 0 27888 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_108
timestamp 1486834041
transform 1 0 672 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1486834041
transform -1 0 27888 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_109
timestamp 1486834041
transform 1 0 672 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1486834041
transform -1 0 27888 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_110
timestamp 1486834041
transform 1 0 672 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1486834041
transform -1 0 27888 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_111
timestamp 1486834041
transform 1 0 672 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1486834041
transform -1 0 27888 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_112
timestamp 1486834041
transform 1 0 672 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1486834041
transform -1 0 27888 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_113
timestamp 1486834041
transform 1 0 672 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1486834041
transform -1 0 27888 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_114
timestamp 1486834041
transform 1 0 672 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1486834041
transform -1 0 27888 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_115
timestamp 1486834041
transform 1 0 672 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1486834041
transform -1 0 27888 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_116
timestamp 1486834041
transform 1 0 672 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1486834041
transform -1 0 27888 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_117
timestamp 1486834041
transform 1 0 672 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1486834041
transform -1 0 27888 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_118
timestamp 1486834041
transform 1 0 672 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1486834041
transform -1 0 27888 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_119
timestamp 1486834041
transform 1 0 672 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1486834041
transform -1 0 27888 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_120
timestamp 1486834041
transform 1 0 672 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1486834041
transform -1 0 27888 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_121
timestamp 1486834041
transform 1 0 672 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1486834041
transform -1 0 27888 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_122
timestamp 1486834041
transform 1 0 672 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1486834041
transform -1 0 27888 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_123
timestamp 1486834041
transform 1 0 672 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1486834041
transform -1 0 27888 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_124
timestamp 1486834041
transform 1 0 672 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1486834041
transform -1 0 27888 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_125
timestamp 1486834041
transform 1 0 672 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1486834041
transform -1 0 27888 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_126
timestamp 1486834041
transform 1 0 672 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1486834041
transform -1 0 27888 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_127
timestamp 1486834041
transform 1 0 672 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1486834041
transform -1 0 27888 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_128
timestamp 1486834041
transform 1 0 672 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1486834041
transform -1 0 27888 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_129
timestamp 1486834041
transform 1 0 672 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1486834041
transform -1 0 27888 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_130
timestamp 1486834041
transform 1 0 672 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1486834041
transform -1 0 27888 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_131
timestamp 1486834041
transform 1 0 672 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1486834041
transform -1 0 27888 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_132
timestamp 1486834041
transform 1 0 672 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1486834041
transform -1 0 27888 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Left_133
timestamp 1486834041
transform 1 0 672 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Right_62
timestamp 1486834041
transform -1 0 27888 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Left_134
timestamp 1486834041
transform 1 0 672 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Right_63
timestamp 1486834041
transform -1 0 27888 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Left_135
timestamp 1486834041
transform 1 0 672 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Right_64
timestamp 1486834041
transform -1 0 27888 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Left_136
timestamp 1486834041
transform 1 0 672 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Right_65
timestamp 1486834041
transform -1 0 27888 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Left_137
timestamp 1486834041
transform 1 0 672 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Right_66
timestamp 1486834041
transform -1 0 27888 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Left_138
timestamp 1486834041
transform 1 0 672 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Right_67
timestamp 1486834041
transform -1 0 27888 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Left_139
timestamp 1486834041
transform 1 0 672 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Right_68
timestamp 1486834041
transform -1 0 27888 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Left_140
timestamp 1486834041
transform 1 0 672 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Right_69
timestamp 1486834041
transform -1 0 27888 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Left_141
timestamp 1486834041
transform 1 0 672 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Right_70
timestamp 1486834041
transform -1 0 27888 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_142
timestamp 1486834041
transform 1 0 4480 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_143
timestamp 1486834041
transform 1 0 8288 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_144
timestamp 1486834041
transform 1 0 12096 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_145
timestamp 1486834041
transform 1 0 15904 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_146
timestamp 1486834041
transform 1 0 19712 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_147
timestamp 1486834041
transform 1 0 23520 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_148
timestamp 1486834041
transform 1 0 27328 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_149
timestamp 1486834041
transform 1 0 8512 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_150
timestamp 1486834041
transform 1 0 16352 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_151
timestamp 1486834041
transform 1 0 24192 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_152
timestamp 1486834041
transform 1 0 4592 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_153
timestamp 1486834041
transform 1 0 12432 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_154
timestamp 1486834041
transform 1 0 20272 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_155
timestamp 1486834041
transform 1 0 8512 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_156
timestamp 1486834041
transform 1 0 16352 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_157
timestamp 1486834041
transform 1 0 24192 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_158
timestamp 1486834041
transform 1 0 4592 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_159
timestamp 1486834041
transform 1 0 12432 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_160
timestamp 1486834041
transform 1 0 20272 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_161
timestamp 1486834041
transform 1 0 8512 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_162
timestamp 1486834041
transform 1 0 16352 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_163
timestamp 1486834041
transform 1 0 24192 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_164
timestamp 1486834041
transform 1 0 4592 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_165
timestamp 1486834041
transform 1 0 12432 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_166
timestamp 1486834041
transform 1 0 20272 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_167
timestamp 1486834041
transform 1 0 8512 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_168
timestamp 1486834041
transform 1 0 16352 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_169
timestamp 1486834041
transform 1 0 24192 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_170
timestamp 1486834041
transform 1 0 4592 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_171
timestamp 1486834041
transform 1 0 12432 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_172
timestamp 1486834041
transform 1 0 20272 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_173
timestamp 1486834041
transform 1 0 8512 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_174
timestamp 1486834041
transform 1 0 16352 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_175
timestamp 1486834041
transform 1 0 24192 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_176
timestamp 1486834041
transform 1 0 4592 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_177
timestamp 1486834041
transform 1 0 12432 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_178
timestamp 1486834041
transform 1 0 20272 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_179
timestamp 1486834041
transform 1 0 8512 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_180
timestamp 1486834041
transform 1 0 16352 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_181
timestamp 1486834041
transform 1 0 24192 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_182
timestamp 1486834041
transform 1 0 4592 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_183
timestamp 1486834041
transform 1 0 12432 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_184
timestamp 1486834041
transform 1 0 20272 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_185
timestamp 1486834041
transform 1 0 8512 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_186
timestamp 1486834041
transform 1 0 16352 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_187
timestamp 1486834041
transform 1 0 24192 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_188
timestamp 1486834041
transform 1 0 4592 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_189
timestamp 1486834041
transform 1 0 12432 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_190
timestamp 1486834041
transform 1 0 20272 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_191
timestamp 1486834041
transform 1 0 8512 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_192
timestamp 1486834041
transform 1 0 16352 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_193
timestamp 1486834041
transform 1 0 24192 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_194
timestamp 1486834041
transform 1 0 4592 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_195
timestamp 1486834041
transform 1 0 12432 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_196
timestamp 1486834041
transform 1 0 20272 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_197
timestamp 1486834041
transform 1 0 8512 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_198
timestamp 1486834041
transform 1 0 16352 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_199
timestamp 1486834041
transform 1 0 24192 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_200
timestamp 1486834041
transform 1 0 4592 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_201
timestamp 1486834041
transform 1 0 12432 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_202
timestamp 1486834041
transform 1 0 20272 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_203
timestamp 1486834041
transform 1 0 8512 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_204
timestamp 1486834041
transform 1 0 16352 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_205
timestamp 1486834041
transform 1 0 24192 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_206
timestamp 1486834041
transform 1 0 4592 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_207
timestamp 1486834041
transform 1 0 12432 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_208
timestamp 1486834041
transform 1 0 20272 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_209
timestamp 1486834041
transform 1 0 8512 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_210
timestamp 1486834041
transform 1 0 16352 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_211
timestamp 1486834041
transform 1 0 24192 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_212
timestamp 1486834041
transform 1 0 4592 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_213
timestamp 1486834041
transform 1 0 12432 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_214
timestamp 1486834041
transform 1 0 20272 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_215
timestamp 1486834041
transform 1 0 8512 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_216
timestamp 1486834041
transform 1 0 16352 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_217
timestamp 1486834041
transform 1 0 24192 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_218
timestamp 1486834041
transform 1 0 4592 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_219
timestamp 1486834041
transform 1 0 12432 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_220
timestamp 1486834041
transform 1 0 20272 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_221
timestamp 1486834041
transform 1 0 8512 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_222
timestamp 1486834041
transform 1 0 16352 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_223
timestamp 1486834041
transform 1 0 24192 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_224
timestamp 1486834041
transform 1 0 4592 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_225
timestamp 1486834041
transform 1 0 12432 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_226
timestamp 1486834041
transform 1 0 20272 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_227
timestamp 1486834041
transform 1 0 8512 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_228
timestamp 1486834041
transform 1 0 16352 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_229
timestamp 1486834041
transform 1 0 24192 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_230
timestamp 1486834041
transform 1 0 4592 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_231
timestamp 1486834041
transform 1 0 12432 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_232
timestamp 1486834041
transform 1 0 20272 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_233
timestamp 1486834041
transform 1 0 8512 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_234
timestamp 1486834041
transform 1 0 16352 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_235
timestamp 1486834041
transform 1 0 24192 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_236
timestamp 1486834041
transform 1 0 4592 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_237
timestamp 1486834041
transform 1 0 12432 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_238
timestamp 1486834041
transform 1 0 20272 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_239
timestamp 1486834041
transform 1 0 8512 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_240
timestamp 1486834041
transform 1 0 16352 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_241
timestamp 1486834041
transform 1 0 24192 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1486834041
transform 1 0 4592 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1486834041
transform 1 0 12432 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_244
timestamp 1486834041
transform 1 0 20272 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1486834041
transform 1 0 8512 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1486834041
transform 1 0 16352 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1486834041
transform 1 0 24192 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1486834041
transform 1 0 4592 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1486834041
transform 1 0 12432 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1486834041
transform 1 0 20272 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_251
timestamp 1486834041
transform 1 0 8512 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_252
timestamp 1486834041
transform 1 0 16352 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1486834041
transform 1 0 24192 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_254
timestamp 1486834041
transform 1 0 4592 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_255
timestamp 1486834041
transform 1 0 12432 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_256
timestamp 1486834041
transform 1 0 20272 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_257
timestamp 1486834041
transform 1 0 8512 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_258
timestamp 1486834041
transform 1 0 16352 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_259
timestamp 1486834041
transform 1 0 24192 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_260
timestamp 1486834041
transform 1 0 4592 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_261
timestamp 1486834041
transform 1 0 12432 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_262
timestamp 1486834041
transform 1 0 20272 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_263
timestamp 1486834041
transform 1 0 8512 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_264
timestamp 1486834041
transform 1 0 16352 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_265
timestamp 1486834041
transform 1 0 24192 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_266
timestamp 1486834041
transform 1 0 4592 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_267
timestamp 1486834041
transform 1 0 12432 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_268
timestamp 1486834041
transform 1 0 20272 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_269
timestamp 1486834041
transform 1 0 8512 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_270
timestamp 1486834041
transform 1 0 16352 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_271
timestamp 1486834041
transform 1 0 24192 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_272
timestamp 1486834041
transform 1 0 4592 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_273
timestamp 1486834041
transform 1 0 12432 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_274
timestamp 1486834041
transform 1 0 20272 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_275
timestamp 1486834041
transform 1 0 8512 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_276
timestamp 1486834041
transform 1 0 16352 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_277
timestamp 1486834041
transform 1 0 24192 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_278
timestamp 1486834041
transform 1 0 4592 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_279
timestamp 1486834041
transform 1 0 12432 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_280
timestamp 1486834041
transform 1 0 20272 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_281
timestamp 1486834041
transform 1 0 8512 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_282
timestamp 1486834041
transform 1 0 16352 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_283
timestamp 1486834041
transform 1 0 24192 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_284
timestamp 1486834041
transform 1 0 4592 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_285
timestamp 1486834041
transform 1 0 12432 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_286
timestamp 1486834041
transform 1 0 20272 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_287
timestamp 1486834041
transform 1 0 8512 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_288
timestamp 1486834041
transform 1 0 16352 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_289
timestamp 1486834041
transform 1 0 24192 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_290
timestamp 1486834041
transform 1 0 4592 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_291
timestamp 1486834041
transform 1 0 12432 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_292
timestamp 1486834041
transform 1 0 20272 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_293
timestamp 1486834041
transform 1 0 8512 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_294
timestamp 1486834041
transform 1 0 16352 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_295
timestamp 1486834041
transform 1 0 24192 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_296
timestamp 1486834041
transform 1 0 4592 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_297
timestamp 1486834041
transform 1 0 12432 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_298
timestamp 1486834041
transform 1 0 20272 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_299
timestamp 1486834041
transform 1 0 8512 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_300
timestamp 1486834041
transform 1 0 16352 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_301
timestamp 1486834041
transform 1 0 24192 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_302
timestamp 1486834041
transform 1 0 4592 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_303
timestamp 1486834041
transform 1 0 12432 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_304
timestamp 1486834041
transform 1 0 20272 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_305
timestamp 1486834041
transform 1 0 8512 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_306
timestamp 1486834041
transform 1 0 16352 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_307
timestamp 1486834041
transform 1 0 24192 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_308
timestamp 1486834041
transform 1 0 4592 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_309
timestamp 1486834041
transform 1 0 12432 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_310
timestamp 1486834041
transform 1 0 20272 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_311
timestamp 1486834041
transform 1 0 8512 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_312
timestamp 1486834041
transform 1 0 16352 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_313
timestamp 1486834041
transform 1 0 24192 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_314
timestamp 1486834041
transform 1 0 4592 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_315
timestamp 1486834041
transform 1 0 12432 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_316
timestamp 1486834041
transform 1 0 20272 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_317
timestamp 1486834041
transform 1 0 8512 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_318
timestamp 1486834041
transform 1 0 16352 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_319
timestamp 1486834041
transform 1 0 24192 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_320
timestamp 1486834041
transform 1 0 4592 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_321
timestamp 1486834041
transform 1 0 12432 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_322
timestamp 1486834041
transform 1 0 20272 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_323
timestamp 1486834041
transform 1 0 8512 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_324
timestamp 1486834041
transform 1 0 16352 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_325
timestamp 1486834041
transform 1 0 24192 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_326
timestamp 1486834041
transform 1 0 4592 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_327
timestamp 1486834041
transform 1 0 12432 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_328
timestamp 1486834041
transform 1 0 20272 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_329
timestamp 1486834041
transform 1 0 8512 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_330
timestamp 1486834041
transform 1 0 16352 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_331
timestamp 1486834041
transform 1 0 24192 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_332
timestamp 1486834041
transform 1 0 4592 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_333
timestamp 1486834041
transform 1 0 12432 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_334
timestamp 1486834041
transform 1 0 20272 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_335
timestamp 1486834041
transform 1 0 8512 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_336
timestamp 1486834041
transform 1 0 16352 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_337
timestamp 1486834041
transform 1 0 24192 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_338
timestamp 1486834041
transform 1 0 4592 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_339
timestamp 1486834041
transform 1 0 12432 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_340
timestamp 1486834041
transform 1 0 20272 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_341
timestamp 1486834041
transform 1 0 8512 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_342
timestamp 1486834041
transform 1 0 16352 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_343
timestamp 1486834041
transform 1 0 24192 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_344
timestamp 1486834041
transform 1 0 4592 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_345
timestamp 1486834041
transform 1 0 12432 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_346
timestamp 1486834041
transform 1 0 20272 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_347
timestamp 1486834041
transform 1 0 8512 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_348
timestamp 1486834041
transform 1 0 16352 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_349
timestamp 1486834041
transform 1 0 24192 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_350
timestamp 1486834041
transform 1 0 4592 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_351
timestamp 1486834041
transform 1 0 12432 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_352
timestamp 1486834041
transform 1 0 20272 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_353
timestamp 1486834041
transform 1 0 8512 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_354
timestamp 1486834041
transform 1 0 16352 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_355
timestamp 1486834041
transform 1 0 24192 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_356
timestamp 1486834041
transform 1 0 4480 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_357
timestamp 1486834041
transform 1 0 8288 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_358
timestamp 1486834041
transform 1 0 12096 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_359
timestamp 1486834041
transform 1 0 15904 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_360
timestamp 1486834041
transform 1 0 19712 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_361
timestamp 1486834041
transform 1 0 23520 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_362
timestamp 1486834041
transform 1 0 27328 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  wire190
timestamp 1486834041
transform -1 0 13888 0 1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  wire191
timestamp 1486834041
transform -1 0 15008 0 -1 13328
box -86 -86 758 870
<< labels >>
flabel metal3 s 0 5152 112 5264 0 FreeSans 448 0 0 0 A_I_top
port 0 nsew signal output
flabel metal3 s 0 3808 112 3920 0 FreeSans 448 0 0 0 A_O_top
port 1 nsew signal input
flabel metal3 s 0 6496 112 6608 0 FreeSans 448 0 0 0 A_T_top
port 2 nsew signal output
flabel metal3 s 0 9184 112 9296 0 FreeSans 448 0 0 0 B_I_top
port 3 nsew signal output
flabel metal3 s 0 7840 112 7952 0 FreeSans 448 0 0 0 B_O_top
port 4 nsew signal input
flabel metal3 s 0 10528 112 10640 0 FreeSans 448 0 0 0 B_T_top
port 5 nsew signal output
flabel metal3 s 28448 21728 28560 21840 0 FreeSans 448 0 0 0 E1BEG[0]
port 6 nsew signal output
flabel metal3 s 28448 22176 28560 22288 0 FreeSans 448 0 0 0 E1BEG[1]
port 7 nsew signal output
flabel metal3 s 28448 22624 28560 22736 0 FreeSans 448 0 0 0 E1BEG[2]
port 8 nsew signal output
flabel metal3 s 28448 23072 28560 23184 0 FreeSans 448 0 0 0 E1BEG[3]
port 9 nsew signal output
flabel metal3 s 28448 23520 28560 23632 0 FreeSans 448 0 0 0 E2BEG[0]
port 10 nsew signal output
flabel metal3 s 28448 23968 28560 24080 0 FreeSans 448 0 0 0 E2BEG[1]
port 11 nsew signal output
flabel metal3 s 28448 24416 28560 24528 0 FreeSans 448 0 0 0 E2BEG[2]
port 12 nsew signal output
flabel metal3 s 28448 24864 28560 24976 0 FreeSans 448 0 0 0 E2BEG[3]
port 13 nsew signal output
flabel metal3 s 28448 25312 28560 25424 0 FreeSans 448 0 0 0 E2BEG[4]
port 14 nsew signal output
flabel metal3 s 28448 25760 28560 25872 0 FreeSans 448 0 0 0 E2BEG[5]
port 15 nsew signal output
flabel metal3 s 28448 26208 28560 26320 0 FreeSans 448 0 0 0 E2BEG[6]
port 16 nsew signal output
flabel metal3 s 28448 26656 28560 26768 0 FreeSans 448 0 0 0 E2BEG[7]
port 17 nsew signal output
flabel metal3 s 28448 27104 28560 27216 0 FreeSans 448 0 0 0 E2BEGb[0]
port 18 nsew signal output
flabel metal3 s 28448 27552 28560 27664 0 FreeSans 448 0 0 0 E2BEGb[1]
port 19 nsew signal output
flabel metal3 s 28448 28000 28560 28112 0 FreeSans 448 0 0 0 E2BEGb[2]
port 20 nsew signal output
flabel metal3 s 28448 28448 28560 28560 0 FreeSans 448 0 0 0 E2BEGb[3]
port 21 nsew signal output
flabel metal3 s 28448 28896 28560 29008 0 FreeSans 448 0 0 0 E2BEGb[4]
port 22 nsew signal output
flabel metal3 s 28448 29344 28560 29456 0 FreeSans 448 0 0 0 E2BEGb[5]
port 23 nsew signal output
flabel metal3 s 28448 29792 28560 29904 0 FreeSans 448 0 0 0 E2BEGb[6]
port 24 nsew signal output
flabel metal3 s 28448 30240 28560 30352 0 FreeSans 448 0 0 0 E2BEGb[7]
port 25 nsew signal output
flabel metal3 s 28448 37856 28560 37968 0 FreeSans 448 0 0 0 E6BEG[0]
port 26 nsew signal output
flabel metal3 s 28448 42336 28560 42448 0 FreeSans 448 0 0 0 E6BEG[10]
port 27 nsew signal output
flabel metal3 s 28448 42784 28560 42896 0 FreeSans 448 0 0 0 E6BEG[11]
port 28 nsew signal output
flabel metal3 s 28448 38304 28560 38416 0 FreeSans 448 0 0 0 E6BEG[1]
port 29 nsew signal output
flabel metal3 s 28448 38752 28560 38864 0 FreeSans 448 0 0 0 E6BEG[2]
port 30 nsew signal output
flabel metal3 s 28448 39200 28560 39312 0 FreeSans 448 0 0 0 E6BEG[3]
port 31 nsew signal output
flabel metal3 s 28448 39648 28560 39760 0 FreeSans 448 0 0 0 E6BEG[4]
port 32 nsew signal output
flabel metal3 s 28448 40096 28560 40208 0 FreeSans 448 0 0 0 E6BEG[5]
port 33 nsew signal output
flabel metal3 s 28448 40544 28560 40656 0 FreeSans 448 0 0 0 E6BEG[6]
port 34 nsew signal output
flabel metal3 s 28448 40992 28560 41104 0 FreeSans 448 0 0 0 E6BEG[7]
port 35 nsew signal output
flabel metal3 s 28448 41440 28560 41552 0 FreeSans 448 0 0 0 E6BEG[8]
port 36 nsew signal output
flabel metal3 s 28448 41888 28560 42000 0 FreeSans 448 0 0 0 E6BEG[9]
port 37 nsew signal output
flabel metal3 s 28448 30688 28560 30800 0 FreeSans 448 0 0 0 EE4BEG[0]
port 38 nsew signal output
flabel metal3 s 28448 35168 28560 35280 0 FreeSans 448 0 0 0 EE4BEG[10]
port 39 nsew signal output
flabel metal3 s 28448 35616 28560 35728 0 FreeSans 448 0 0 0 EE4BEG[11]
port 40 nsew signal output
flabel metal3 s 28448 36064 28560 36176 0 FreeSans 448 0 0 0 EE4BEG[12]
port 41 nsew signal output
flabel metal3 s 28448 36512 28560 36624 0 FreeSans 448 0 0 0 EE4BEG[13]
port 42 nsew signal output
flabel metal3 s 28448 36960 28560 37072 0 FreeSans 448 0 0 0 EE4BEG[14]
port 43 nsew signal output
flabel metal3 s 28448 37408 28560 37520 0 FreeSans 448 0 0 0 EE4BEG[15]
port 44 nsew signal output
flabel metal3 s 28448 31136 28560 31248 0 FreeSans 448 0 0 0 EE4BEG[1]
port 45 nsew signal output
flabel metal3 s 28448 31584 28560 31696 0 FreeSans 448 0 0 0 EE4BEG[2]
port 46 nsew signal output
flabel metal3 s 28448 32032 28560 32144 0 FreeSans 448 0 0 0 EE4BEG[3]
port 47 nsew signal output
flabel metal3 s 28448 32480 28560 32592 0 FreeSans 448 0 0 0 EE4BEG[4]
port 48 nsew signal output
flabel metal3 s 28448 32928 28560 33040 0 FreeSans 448 0 0 0 EE4BEG[5]
port 49 nsew signal output
flabel metal3 s 28448 33376 28560 33488 0 FreeSans 448 0 0 0 EE4BEG[6]
port 50 nsew signal output
flabel metal3 s 28448 33824 28560 33936 0 FreeSans 448 0 0 0 EE4BEG[7]
port 51 nsew signal output
flabel metal3 s 28448 34272 28560 34384 0 FreeSans 448 0 0 0 EE4BEG[8]
port 52 nsew signal output
flabel metal3 s 28448 34720 28560 34832 0 FreeSans 448 0 0 0 EE4BEG[9]
port 53 nsew signal output
flabel metal3 s 0 11872 112 11984 0 FreeSans 448 0 0 0 FrameData[0]
port 54 nsew signal input
flabel metal3 s 0 25312 112 25424 0 FreeSans 448 0 0 0 FrameData[10]
port 55 nsew signal input
flabel metal3 s 0 26656 112 26768 0 FreeSans 448 0 0 0 FrameData[11]
port 56 nsew signal input
flabel metal3 s 0 28000 112 28112 0 FreeSans 448 0 0 0 FrameData[12]
port 57 nsew signal input
flabel metal3 s 0 29344 112 29456 0 FreeSans 448 0 0 0 FrameData[13]
port 58 nsew signal input
flabel metal3 s 0 30688 112 30800 0 FreeSans 448 0 0 0 FrameData[14]
port 59 nsew signal input
flabel metal3 s 0 32032 112 32144 0 FreeSans 448 0 0 0 FrameData[15]
port 60 nsew signal input
flabel metal3 s 0 33376 112 33488 0 FreeSans 448 0 0 0 FrameData[16]
port 61 nsew signal input
flabel metal3 s 0 34720 112 34832 0 FreeSans 448 0 0 0 FrameData[17]
port 62 nsew signal input
flabel metal3 s 0 36064 112 36176 0 FreeSans 448 0 0 0 FrameData[18]
port 63 nsew signal input
flabel metal3 s 0 37408 112 37520 0 FreeSans 448 0 0 0 FrameData[19]
port 64 nsew signal input
flabel metal3 s 0 13216 112 13328 0 FreeSans 448 0 0 0 FrameData[1]
port 65 nsew signal input
flabel metal3 s 0 38752 112 38864 0 FreeSans 448 0 0 0 FrameData[20]
port 66 nsew signal input
flabel metal3 s 0 40096 112 40208 0 FreeSans 448 0 0 0 FrameData[21]
port 67 nsew signal input
flabel metal3 s 0 41440 112 41552 0 FreeSans 448 0 0 0 FrameData[22]
port 68 nsew signal input
flabel metal3 s 0 42784 112 42896 0 FreeSans 448 0 0 0 FrameData[23]
port 69 nsew signal input
flabel metal3 s 0 44128 112 44240 0 FreeSans 448 0 0 0 FrameData[24]
port 70 nsew signal input
flabel metal3 s 0 45472 112 45584 0 FreeSans 448 0 0 0 FrameData[25]
port 71 nsew signal input
flabel metal3 s 0 46816 112 46928 0 FreeSans 448 0 0 0 FrameData[26]
port 72 nsew signal input
flabel metal3 s 0 48160 112 48272 0 FreeSans 448 0 0 0 FrameData[27]
port 73 nsew signal input
flabel metal3 s 0 49504 112 49616 0 FreeSans 448 0 0 0 FrameData[28]
port 74 nsew signal input
flabel metal3 s 0 50848 112 50960 0 FreeSans 448 0 0 0 FrameData[29]
port 75 nsew signal input
flabel metal3 s 0 14560 112 14672 0 FreeSans 448 0 0 0 FrameData[2]
port 76 nsew signal input
flabel metal3 s 0 52192 112 52304 0 FreeSans 448 0 0 0 FrameData[30]
port 77 nsew signal input
flabel metal3 s 0 53536 112 53648 0 FreeSans 448 0 0 0 FrameData[31]
port 78 nsew signal input
flabel metal3 s 0 15904 112 16016 0 FreeSans 448 0 0 0 FrameData[3]
port 79 nsew signal input
flabel metal3 s 0 17248 112 17360 0 FreeSans 448 0 0 0 FrameData[4]
port 80 nsew signal input
flabel metal3 s 0 18592 112 18704 0 FreeSans 448 0 0 0 FrameData[5]
port 81 nsew signal input
flabel metal3 s 0 19936 112 20048 0 FreeSans 448 0 0 0 FrameData[6]
port 82 nsew signal input
flabel metal3 s 0 21280 112 21392 0 FreeSans 448 0 0 0 FrameData[7]
port 83 nsew signal input
flabel metal3 s 0 22624 112 22736 0 FreeSans 448 0 0 0 FrameData[8]
port 84 nsew signal input
flabel metal3 s 0 23968 112 24080 0 FreeSans 448 0 0 0 FrameData[9]
port 85 nsew signal input
flabel metal3 s 28448 43232 28560 43344 0 FreeSans 448 0 0 0 FrameData_O[0]
port 86 nsew signal output
flabel metal3 s 28448 47712 28560 47824 0 FreeSans 448 0 0 0 FrameData_O[10]
port 87 nsew signal output
flabel metal3 s 28448 48160 28560 48272 0 FreeSans 448 0 0 0 FrameData_O[11]
port 88 nsew signal output
flabel metal3 s 28448 48608 28560 48720 0 FreeSans 448 0 0 0 FrameData_O[12]
port 89 nsew signal output
flabel metal3 s 28448 49056 28560 49168 0 FreeSans 448 0 0 0 FrameData_O[13]
port 90 nsew signal output
flabel metal3 s 28448 49504 28560 49616 0 FreeSans 448 0 0 0 FrameData_O[14]
port 91 nsew signal output
flabel metal3 s 28448 49952 28560 50064 0 FreeSans 448 0 0 0 FrameData_O[15]
port 92 nsew signal output
flabel metal3 s 28448 50400 28560 50512 0 FreeSans 448 0 0 0 FrameData_O[16]
port 93 nsew signal output
flabel metal3 s 28448 50848 28560 50960 0 FreeSans 448 0 0 0 FrameData_O[17]
port 94 nsew signal output
flabel metal3 s 28448 51296 28560 51408 0 FreeSans 448 0 0 0 FrameData_O[18]
port 95 nsew signal output
flabel metal3 s 28448 51744 28560 51856 0 FreeSans 448 0 0 0 FrameData_O[19]
port 96 nsew signal output
flabel metal3 s 28448 43680 28560 43792 0 FreeSans 448 0 0 0 FrameData_O[1]
port 97 nsew signal output
flabel metal3 s 28448 52192 28560 52304 0 FreeSans 448 0 0 0 FrameData_O[20]
port 98 nsew signal output
flabel metal3 s 28448 52640 28560 52752 0 FreeSans 448 0 0 0 FrameData_O[21]
port 99 nsew signal output
flabel metal3 s 28448 53088 28560 53200 0 FreeSans 448 0 0 0 FrameData_O[22]
port 100 nsew signal output
flabel metal3 s 28448 53536 28560 53648 0 FreeSans 448 0 0 0 FrameData_O[23]
port 101 nsew signal output
flabel metal3 s 28448 53984 28560 54096 0 FreeSans 448 0 0 0 FrameData_O[24]
port 102 nsew signal output
flabel metal3 s 28448 54432 28560 54544 0 FreeSans 448 0 0 0 FrameData_O[25]
port 103 nsew signal output
flabel metal3 s 28448 54880 28560 54992 0 FreeSans 448 0 0 0 FrameData_O[26]
port 104 nsew signal output
flabel metal3 s 28448 55328 28560 55440 0 FreeSans 448 0 0 0 FrameData_O[27]
port 105 nsew signal output
flabel metal3 s 28448 55776 28560 55888 0 FreeSans 448 0 0 0 FrameData_O[28]
port 106 nsew signal output
flabel metal3 s 28448 56224 28560 56336 0 FreeSans 448 0 0 0 FrameData_O[29]
port 107 nsew signal output
flabel metal3 s 28448 44128 28560 44240 0 FreeSans 448 0 0 0 FrameData_O[2]
port 108 nsew signal output
flabel metal3 s 28448 56672 28560 56784 0 FreeSans 448 0 0 0 FrameData_O[30]
port 109 nsew signal output
flabel metal3 s 28448 57120 28560 57232 0 FreeSans 448 0 0 0 FrameData_O[31]
port 110 nsew signal output
flabel metal3 s 28448 44576 28560 44688 0 FreeSans 448 0 0 0 FrameData_O[3]
port 111 nsew signal output
flabel metal3 s 28448 45024 28560 45136 0 FreeSans 448 0 0 0 FrameData_O[4]
port 112 nsew signal output
flabel metal3 s 28448 45472 28560 45584 0 FreeSans 448 0 0 0 FrameData_O[5]
port 113 nsew signal output
flabel metal3 s 28448 45920 28560 46032 0 FreeSans 448 0 0 0 FrameData_O[6]
port 114 nsew signal output
flabel metal3 s 28448 46368 28560 46480 0 FreeSans 448 0 0 0 FrameData_O[7]
port 115 nsew signal output
flabel metal3 s 28448 46816 28560 46928 0 FreeSans 448 0 0 0 FrameData_O[8]
port 116 nsew signal output
flabel metal3 s 28448 47264 28560 47376 0 FreeSans 448 0 0 0 FrameData_O[9]
port 117 nsew signal output
flabel metal2 s 2016 0 2128 112 0 FreeSans 448 0 0 0 FrameStrobe[0]
port 118 nsew signal input
flabel metal2 s 15456 0 15568 112 0 FreeSans 448 0 0 0 FrameStrobe[10]
port 119 nsew signal input
flabel metal2 s 16800 0 16912 112 0 FreeSans 448 0 0 0 FrameStrobe[11]
port 120 nsew signal input
flabel metal2 s 18144 0 18256 112 0 FreeSans 448 0 0 0 FrameStrobe[12]
port 121 nsew signal input
flabel metal2 s 19488 0 19600 112 0 FreeSans 448 0 0 0 FrameStrobe[13]
port 122 nsew signal input
flabel metal2 s 20832 0 20944 112 0 FreeSans 448 0 0 0 FrameStrobe[14]
port 123 nsew signal input
flabel metal2 s 22176 0 22288 112 0 FreeSans 448 0 0 0 FrameStrobe[15]
port 124 nsew signal input
flabel metal2 s 23520 0 23632 112 0 FreeSans 448 0 0 0 FrameStrobe[16]
port 125 nsew signal input
flabel metal2 s 24864 0 24976 112 0 FreeSans 448 0 0 0 FrameStrobe[17]
port 126 nsew signal input
flabel metal2 s 26208 0 26320 112 0 FreeSans 448 0 0 0 FrameStrobe[18]
port 127 nsew signal input
flabel metal2 s 27552 0 27664 112 0 FreeSans 448 0 0 0 FrameStrobe[19]
port 128 nsew signal input
flabel metal2 s 3360 0 3472 112 0 FreeSans 448 0 0 0 FrameStrobe[1]
port 129 nsew signal input
flabel metal2 s 4704 0 4816 112 0 FreeSans 448 0 0 0 FrameStrobe[2]
port 130 nsew signal input
flabel metal2 s 6048 0 6160 112 0 FreeSans 448 0 0 0 FrameStrobe[3]
port 131 nsew signal input
flabel metal2 s 7392 0 7504 112 0 FreeSans 448 0 0 0 FrameStrobe[4]
port 132 nsew signal input
flabel metal2 s 8736 0 8848 112 0 FreeSans 448 0 0 0 FrameStrobe[5]
port 133 nsew signal input
flabel metal2 s 10080 0 10192 112 0 FreeSans 448 0 0 0 FrameStrobe[6]
port 134 nsew signal input
flabel metal2 s 11424 0 11536 112 0 FreeSans 448 0 0 0 FrameStrobe[7]
port 135 nsew signal input
flabel metal2 s 12768 0 12880 112 0 FreeSans 448 0 0 0 FrameStrobe[8]
port 136 nsew signal input
flabel metal2 s 14112 0 14224 112 0 FreeSans 448 0 0 0 FrameStrobe[9]
port 137 nsew signal input
flabel metal2 s 2016 57344 2128 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[0]
port 138 nsew signal output
flabel metal2 s 15456 57344 15568 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[10]
port 139 nsew signal output
flabel metal2 s 16800 57344 16912 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[11]
port 140 nsew signal output
flabel metal2 s 18144 57344 18256 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[12]
port 141 nsew signal output
flabel metal2 s 19488 57344 19600 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[13]
port 142 nsew signal output
flabel metal2 s 20832 57344 20944 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[14]
port 143 nsew signal output
flabel metal2 s 22176 57344 22288 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[15]
port 144 nsew signal output
flabel metal2 s 23520 57344 23632 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[16]
port 145 nsew signal output
flabel metal2 s 24864 57344 24976 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[17]
port 146 nsew signal output
flabel metal2 s 26208 57344 26320 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[18]
port 147 nsew signal output
flabel metal2 s 27552 57344 27664 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[19]
port 148 nsew signal output
flabel metal2 s 3360 57344 3472 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[1]
port 149 nsew signal output
flabel metal2 s 4704 57344 4816 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[2]
port 150 nsew signal output
flabel metal2 s 6048 57344 6160 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[3]
port 151 nsew signal output
flabel metal2 s 7392 57344 7504 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[4]
port 152 nsew signal output
flabel metal2 s 8736 57344 8848 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[5]
port 153 nsew signal output
flabel metal2 s 10080 57344 10192 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[6]
port 154 nsew signal output
flabel metal2 s 11424 57344 11536 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[7]
port 155 nsew signal output
flabel metal2 s 12768 57344 12880 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[8]
port 156 nsew signal output
flabel metal2 s 14112 57344 14224 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[9]
port 157 nsew signal output
flabel metal2 s 672 0 784 112 0 FreeSans 448 0 0 0 UserCLK
port 158 nsew signal input
flabel metal2 s 672 57344 784 57456 0 FreeSans 448 0 0 0 UserCLKo
port 159 nsew signal output
flabel metal4 s 3776 0 4096 57456 0 FreeSans 1472 90 0 0 VDD
port 160 nsew power bidirectional
flabel metal4 s 3776 0 4096 56 0 FreeSans 368 0 0 0 VDD
port 160 nsew power bidirectional
flabel metal4 s 3776 57400 4096 57456 0 FreeSans 368 0 0 0 VDD
port 160 nsew power bidirectional
flabel metal4 s 23776 0 24096 57456 0 FreeSans 1472 90 0 0 VDD
port 160 nsew power bidirectional
flabel metal4 s 23776 0 24096 56 0 FreeSans 368 0 0 0 VDD
port 160 nsew power bidirectional
flabel metal4 s 23776 57400 24096 57456 0 FreeSans 368 0 0 0 VDD
port 160 nsew power bidirectional
flabel metal4 s 4436 0 4756 57456 0 FreeSans 1472 90 0 0 VSS
port 161 nsew ground bidirectional
flabel metal4 s 4436 0 4756 56 0 FreeSans 368 0 0 0 VSS
port 161 nsew ground bidirectional
flabel metal4 s 4436 57400 4756 57456 0 FreeSans 368 0 0 0 VSS
port 161 nsew ground bidirectional
flabel metal4 s 24436 0 24756 57456 0 FreeSans 1472 90 0 0 VSS
port 161 nsew ground bidirectional
flabel metal4 s 24436 0 24756 56 0 FreeSans 368 0 0 0 VSS
port 161 nsew ground bidirectional
flabel metal4 s 24436 57400 24756 57456 0 FreeSans 368 0 0 0 VSS
port 161 nsew ground bidirectional
flabel metal3 s 28448 224 28560 336 0 FreeSans 448 0 0 0 W1END[0]
port 162 nsew signal input
flabel metal3 s 28448 672 28560 784 0 FreeSans 448 0 0 0 W1END[1]
port 163 nsew signal input
flabel metal3 s 28448 1120 28560 1232 0 FreeSans 448 0 0 0 W1END[2]
port 164 nsew signal input
flabel metal3 s 28448 1568 28560 1680 0 FreeSans 448 0 0 0 W1END[3]
port 165 nsew signal input
flabel metal3 s 28448 5600 28560 5712 0 FreeSans 448 0 0 0 W2END[0]
port 166 nsew signal input
flabel metal3 s 28448 6048 28560 6160 0 FreeSans 448 0 0 0 W2END[1]
port 167 nsew signal input
flabel metal3 s 28448 6496 28560 6608 0 FreeSans 448 0 0 0 W2END[2]
port 168 nsew signal input
flabel metal3 s 28448 6944 28560 7056 0 FreeSans 448 0 0 0 W2END[3]
port 169 nsew signal input
flabel metal3 s 28448 7392 28560 7504 0 FreeSans 448 0 0 0 W2END[4]
port 170 nsew signal input
flabel metal3 s 28448 7840 28560 7952 0 FreeSans 448 0 0 0 W2END[5]
port 171 nsew signal input
flabel metal3 s 28448 8288 28560 8400 0 FreeSans 448 0 0 0 W2END[6]
port 172 nsew signal input
flabel metal3 s 28448 8736 28560 8848 0 FreeSans 448 0 0 0 W2END[7]
port 173 nsew signal input
flabel metal3 s 28448 2016 28560 2128 0 FreeSans 448 0 0 0 W2MID[0]
port 174 nsew signal input
flabel metal3 s 28448 2464 28560 2576 0 FreeSans 448 0 0 0 W2MID[1]
port 175 nsew signal input
flabel metal3 s 28448 2912 28560 3024 0 FreeSans 448 0 0 0 W2MID[2]
port 176 nsew signal input
flabel metal3 s 28448 3360 28560 3472 0 FreeSans 448 0 0 0 W2MID[3]
port 177 nsew signal input
flabel metal3 s 28448 3808 28560 3920 0 FreeSans 448 0 0 0 W2MID[4]
port 178 nsew signal input
flabel metal3 s 28448 4256 28560 4368 0 FreeSans 448 0 0 0 W2MID[5]
port 179 nsew signal input
flabel metal3 s 28448 4704 28560 4816 0 FreeSans 448 0 0 0 W2MID[6]
port 180 nsew signal input
flabel metal3 s 28448 5152 28560 5264 0 FreeSans 448 0 0 0 W2MID[7]
port 181 nsew signal input
flabel metal3 s 28448 16352 28560 16464 0 FreeSans 448 0 0 0 W6END[0]
port 182 nsew signal input
flabel metal3 s 28448 20832 28560 20944 0 FreeSans 448 0 0 0 W6END[10]
port 183 nsew signal input
flabel metal3 s 28448 21280 28560 21392 0 FreeSans 448 0 0 0 W6END[11]
port 184 nsew signal input
flabel metal3 s 28448 16800 28560 16912 0 FreeSans 448 0 0 0 W6END[1]
port 185 nsew signal input
flabel metal3 s 28448 17248 28560 17360 0 FreeSans 448 0 0 0 W6END[2]
port 186 nsew signal input
flabel metal3 s 28448 17696 28560 17808 0 FreeSans 448 0 0 0 W6END[3]
port 187 nsew signal input
flabel metal3 s 28448 18144 28560 18256 0 FreeSans 448 0 0 0 W6END[4]
port 188 nsew signal input
flabel metal3 s 28448 18592 28560 18704 0 FreeSans 448 0 0 0 W6END[5]
port 189 nsew signal input
flabel metal3 s 28448 19040 28560 19152 0 FreeSans 448 0 0 0 W6END[6]
port 190 nsew signal input
flabel metal3 s 28448 19488 28560 19600 0 FreeSans 448 0 0 0 W6END[7]
port 191 nsew signal input
flabel metal3 s 28448 19936 28560 20048 0 FreeSans 448 0 0 0 W6END[8]
port 192 nsew signal input
flabel metal3 s 28448 20384 28560 20496 0 FreeSans 448 0 0 0 W6END[9]
port 193 nsew signal input
flabel metal3 s 28448 9184 28560 9296 0 FreeSans 448 0 0 0 WW4END[0]
port 194 nsew signal input
flabel metal3 s 28448 13664 28560 13776 0 FreeSans 448 0 0 0 WW4END[10]
port 195 nsew signal input
flabel metal3 s 28448 14112 28560 14224 0 FreeSans 448 0 0 0 WW4END[11]
port 196 nsew signal input
flabel metal3 s 28448 14560 28560 14672 0 FreeSans 448 0 0 0 WW4END[12]
port 197 nsew signal input
flabel metal3 s 28448 15008 28560 15120 0 FreeSans 448 0 0 0 WW4END[13]
port 198 nsew signal input
flabel metal3 s 28448 15456 28560 15568 0 FreeSans 448 0 0 0 WW4END[14]
port 199 nsew signal input
flabel metal3 s 28448 15904 28560 16016 0 FreeSans 448 0 0 0 WW4END[15]
port 200 nsew signal input
flabel metal3 s 28448 9632 28560 9744 0 FreeSans 448 0 0 0 WW4END[1]
port 201 nsew signal input
flabel metal3 s 28448 10080 28560 10192 0 FreeSans 448 0 0 0 WW4END[2]
port 202 nsew signal input
flabel metal3 s 28448 10528 28560 10640 0 FreeSans 448 0 0 0 WW4END[3]
port 203 nsew signal input
flabel metal3 s 28448 10976 28560 11088 0 FreeSans 448 0 0 0 WW4END[4]
port 204 nsew signal input
flabel metal3 s 28448 11424 28560 11536 0 FreeSans 448 0 0 0 WW4END[5]
port 205 nsew signal input
flabel metal3 s 28448 11872 28560 11984 0 FreeSans 448 0 0 0 WW4END[6]
port 206 nsew signal input
flabel metal3 s 28448 12320 28560 12432 0 FreeSans 448 0 0 0 WW4END[7]
port 207 nsew signal input
flabel metal3 s 28448 12768 28560 12880 0 FreeSans 448 0 0 0 WW4END[8]
port 208 nsew signal input
flabel metal3 s 28448 13216 28560 13328 0 FreeSans 448 0 0 0 WW4END[9]
port 209 nsew signal input
rlabel metal1 14280 56448 14280 56448 0 VDD
rlabel metal1 14280 55664 14280 55664 0 VSS
rlabel metal3 686 5208 686 5208 0 A_I_top
rlabel metal3 574 3864 574 3864 0 A_O_top
rlabel metal3 686 6552 686 6552 0 A_T_top
rlabel metal3 686 9240 686 9240 0 B_I_top
rlabel metal2 1064 7672 1064 7672 0 B_O_top
rlabel metal3 686 10584 686 10584 0 B_T_top
rlabel metal2 25704 21952 25704 21952 0 E1BEG[0]
rlabel metal2 27160 21952 27160 21952 0 E1BEG[1]
rlabel metal3 27874 22680 27874 22680 0 E1BEG[2]
rlabel metal2 25704 23408 25704 23408 0 E1BEG[3]
rlabel metal2 27160 23408 27160 23408 0 E2BEG[0]
rlabel metal2 25480 24304 25480 24304 0 E2BEG[1]
rlabel metal3 27874 24472 27874 24472 0 E2BEG[2]
rlabel metal2 25704 25088 25704 25088 0 E2BEG[3]
rlabel metal2 27160 25088 27160 25088 0 E2BEG[4]
rlabel metal3 27874 25816 27874 25816 0 E2BEG[5]
rlabel metal2 25704 26544 25704 26544 0 E2BEG[6]
rlabel metal2 27272 26600 27272 26600 0 E2BEG[7]
rlabel metal2 25704 27552 25704 27552 0 E2BEGb[0]
rlabel metal2 27272 27272 27272 27272 0 E2BEGb[1]
rlabel metal3 27874 28056 27874 28056 0 E2BEGb[2]
rlabel metal3 27874 28504 27874 28504 0 E2BEGb[3]
rlabel metal3 27874 28952 27874 28952 0 E2BEGb[4]
rlabel metal3 27818 29400 27818 29400 0 E2BEGb[5]
rlabel metal3 27762 29848 27762 29848 0 E2BEGb[6]
rlabel metal3 27874 30296 27874 30296 0 E2BEGb[7]
rlabel metal3 27090 37912 27090 37912 0 E6BEG[0]
rlabel metal3 27090 42392 27090 42392 0 E6BEG[10]
rlabel metal3 27874 42840 27874 42840 0 E6BEG[11]
rlabel metal3 27874 38360 27874 38360 0 E6BEG[1]
rlabel metal3 27818 38808 27818 38808 0 E6BEG[2]
rlabel metal3 27090 39256 27090 39256 0 E6BEG[3]
rlabel metal3 27874 39704 27874 39704 0 E6BEG[4]
rlabel metal3 27090 40152 27090 40152 0 E6BEG[5]
rlabel metal3 27762 40600 27762 40600 0 E6BEG[6]
rlabel metal3 27090 41048 27090 41048 0 E6BEG[7]
rlabel metal3 27874 41496 27874 41496 0 E6BEG[8]
rlabel metal3 27818 41944 27818 41944 0 E6BEG[9]
rlabel metal2 25480 30800 25480 30800 0 EE4BEG[0]
rlabel metal3 27874 35224 27874 35224 0 EE4BEG[10]
rlabel metal3 27818 35672 27818 35672 0 EE4BEG[11]
rlabel metal2 25704 36176 25704 36176 0 EE4BEG[12]
rlabel metal3 27874 36568 27874 36568 0 EE4BEG[13]
rlabel metal2 25480 37072 25480 37072 0 EE4BEG[14]
rlabel metal3 27762 37464 27762 37464 0 EE4BEG[15]
rlabel metal3 27762 31192 27762 31192 0 EE4BEG[1]
rlabel metal3 27090 31640 27090 31640 0 EE4BEG[2]
rlabel metal3 27874 32088 27874 32088 0 EE4BEG[3]
rlabel metal3 27818 32536 27818 32536 0 EE4BEG[4]
rlabel metal2 25704 33040 25704 33040 0 EE4BEG[5]
rlabel metal3 27874 33432 27874 33432 0 EE4BEG[6]
rlabel metal2 25704 34048 25704 34048 0 EE4BEG[7]
rlabel metal3 27762 34328 27762 34328 0 EE4BEG[8]
rlabel metal3 27090 34776 27090 34776 0 EE4BEG[9]
rlabel metal3 518 11928 518 11928 0 FrameData[0]
rlabel metal3 574 25368 574 25368 0 FrameData[10]
rlabel metal3 574 26712 574 26712 0 FrameData[11]
rlabel metal2 3416 28728 3416 28728 0 FrameData[12]
rlabel metal2 1064 28616 1064 28616 0 FrameData[13]
rlabel metal2 3528 30576 3528 30576 0 FrameData[14]
rlabel metal3 574 32088 574 32088 0 FrameData[15]
rlabel metal3 518 33432 518 33432 0 FrameData[16]
rlabel metal3 742 34776 742 34776 0 FrameData[17]
rlabel metal2 1008 38584 1008 38584 0 FrameData[18]
rlabel metal3 574 37464 574 37464 0 FrameData[19]
rlabel metal2 1176 11144 1176 11144 0 FrameData[1]
rlabel metal3 574 38808 574 38808 0 FrameData[20]
rlabel metal3 518 40152 518 40152 0 FrameData[21]
rlabel metal3 630 41496 630 41496 0 FrameData[22]
rlabel metal3 518 42840 518 42840 0 FrameData[23]
rlabel metal3 574 44184 574 44184 0 FrameData[24]
rlabel metal3 574 45528 574 45528 0 FrameData[25]
rlabel metal3 574 46872 574 46872 0 FrameData[26]
rlabel metal3 574 48216 574 48216 0 FrameData[27]
rlabel metal3 574 49560 574 49560 0 FrameData[28]
rlabel metal3 574 50904 574 50904 0 FrameData[29]
rlabel metal2 1960 11256 1960 11256 0 FrameData[2]
rlabel metal3 574 52248 574 52248 0 FrameData[30]
rlabel metal3 574 53592 574 53592 0 FrameData[31]
rlabel metal3 350 15960 350 15960 0 FrameData[3]
rlabel metal4 1960 14728 1960 14728 0 FrameData[4]
rlabel metal3 518 18648 518 18648 0 FrameData[5]
rlabel metal2 1960 18424 1960 18424 0 FrameData[6]
rlabel metal2 1176 19096 1176 19096 0 FrameData[7]
rlabel metal3 462 22680 462 22680 0 FrameData[8]
rlabel metal2 1008 21560 1008 21560 0 FrameData[9]
rlabel metal3 27090 43288 27090 43288 0 FrameData_O[0]
rlabel metal3 27874 47768 27874 47768 0 FrameData_O[10]
rlabel metal3 27818 48216 27818 48216 0 FrameData_O[11]
rlabel metal3 27034 48664 27034 48664 0 FrameData_O[12]
rlabel metal3 27874 49112 27874 49112 0 FrameData_O[13]
rlabel metal3 26978 49560 26978 49560 0 FrameData_O[14]
rlabel metal3 27762 50008 27762 50008 0 FrameData_O[15]
rlabel metal3 27034 50456 27034 50456 0 FrameData_O[16]
rlabel metal3 27874 50904 27874 50904 0 FrameData_O[17]
rlabel metal3 27818 51352 27818 51352 0 FrameData_O[18]
rlabel metal3 27034 51800 27034 51800 0 FrameData_O[19]
rlabel metal3 27762 43736 27762 43736 0 FrameData_O[1]
rlabel metal3 27874 52248 27874 52248 0 FrameData_O[20]
rlabel metal3 26978 52696 26978 52696 0 FrameData_O[21]
rlabel metal3 27762 53144 27762 53144 0 FrameData_O[22]
rlabel metal3 27034 53592 27034 53592 0 FrameData_O[23]
rlabel metal3 27874 54040 27874 54040 0 FrameData_O[24]
rlabel metal3 27034 54488 27034 54488 0 FrameData_O[25]
rlabel metal3 25144 54712 25144 54712 0 FrameData_O[26]
rlabel metal2 23800 54040 23800 54040 0 FrameData_O[27]
rlabel metal3 25074 55832 25074 55832 0 FrameData_O[28]
rlabel metal3 27370 56280 27370 56280 0 FrameData_O[29]
rlabel metal3 27090 44184 27090 44184 0 FrameData_O[2]
rlabel metal3 26922 56728 26922 56728 0 FrameData_O[30]
rlabel metal2 24192 53144 24192 53144 0 FrameData_O[31]
rlabel metal3 27874 44632 27874 44632 0 FrameData_O[3]
rlabel metal3 27818 45080 27818 45080 0 FrameData_O[4]
rlabel metal3 27090 45528 27090 45528 0 FrameData_O[5]
rlabel metal3 27874 45976 27874 45976 0 FrameData_O[6]
rlabel metal3 27090 46424 27090 46424 0 FrameData_O[7]
rlabel metal3 27762 46872 27762 46872 0 FrameData_O[8]
rlabel metal3 27090 47320 27090 47320 0 FrameData_O[9]
rlabel metal2 2072 742 2072 742 0 FrameStrobe[0]
rlabel metal3 20608 48664 20608 48664 0 FrameStrobe[10]
rlabel metal3 25928 52920 25928 52920 0 FrameStrobe[11]
rlabel metal2 17696 24248 17696 24248 0 FrameStrobe[12]
rlabel metal2 18928 26040 18928 26040 0 FrameStrobe[13]
rlabel metal2 20888 1694 20888 1694 0 FrameStrobe[14]
rlabel metal3 20888 47992 20888 47992 0 FrameStrobe[15]
rlabel metal2 23576 854 23576 854 0 FrameStrobe[16]
rlabel metal2 24920 798 24920 798 0 FrameStrobe[17]
rlabel metal2 26264 3430 26264 3430 0 FrameStrobe[18]
rlabel metal2 27608 126 27608 126 0 FrameStrobe[19]
rlabel metal2 3416 1414 3416 1414 0 FrameStrobe[1]
rlabel metal2 4760 126 4760 126 0 FrameStrobe[2]
rlabel metal2 6104 518 6104 518 0 FrameStrobe[3]
rlabel metal2 7448 854 7448 854 0 FrameStrobe[4]
rlabel metal3 16296 54264 16296 54264 0 FrameStrobe[5]
rlabel metal2 10136 2646 10136 2646 0 FrameStrobe[6]
rlabel metal3 18200 51128 18200 51128 0 FrameStrobe[7]
rlabel metal2 21896 53368 21896 53368 0 FrameStrobe[8]
rlabel metal2 14168 518 14168 518 0 FrameStrobe[9]
rlabel metal2 2520 55300 2520 55300 0 FrameStrobe_O[0]
rlabel metal3 16016 56280 16016 56280 0 FrameStrobe_O[10]
rlabel metal2 17304 55300 17304 55300 0 FrameStrobe_O[11]
rlabel metal2 18368 56280 18368 56280 0 FrameStrobe_O[12]
rlabel metal2 19544 56826 19544 56826 0 FrameStrobe_O[13]
rlabel metal3 21392 56280 21392 56280 0 FrameStrobe_O[14]
rlabel metal2 22232 57274 22232 57274 0 FrameStrobe_O[15]
rlabel metal2 23576 56826 23576 56826 0 FrameStrobe_O[16]
rlabel metal2 24920 56826 24920 56826 0 FrameStrobe_O[17]
rlabel metal2 26264 57330 26264 57330 0 FrameStrobe_O[18]
rlabel metal2 27608 56714 27608 56714 0 FrameStrobe_O[19]
rlabel metal2 3416 56826 3416 56826 0 FrameStrobe_O[1]
rlabel metal2 4760 57330 4760 57330 0 FrameStrobe_O[2]
rlabel metal2 6552 55300 6552 55300 0 FrameStrobe_O[3]
rlabel metal2 7448 56770 7448 56770 0 FrameStrobe_O[4]
rlabel metal2 9016 56448 9016 56448 0 FrameStrobe_O[5]
rlabel metal2 10584 56504 10584 56504 0 FrameStrobe_O[6]
rlabel metal2 11704 55160 11704 55160 0 FrameStrobe_O[7]
rlabel metal2 13048 56448 13048 56448 0 FrameStrobe_O[8]
rlabel metal2 14616 56504 14616 56504 0 FrameStrobe_O[9]
rlabel metal2 20216 23296 20216 23296 0 Inst_A_IO_1_bidirectional_frame_config_pass.Q
rlabel metal2 2744 31360 2744 31360 0 Inst_B_IO_1_bidirectional_frame_config_pass.Q
rlabel metal2 5544 40264 5544 40264 0 Inst_W_IO_ConfigMem.Inst_frame0_bit0.Q
rlabel metal3 7000 39032 7000 39032 0 Inst_W_IO_ConfigMem.Inst_frame0_bit1.Q
rlabel metal2 4032 23352 4032 23352 0 Inst_W_IO_ConfigMem.Inst_frame0_bit10.Q
rlabel metal2 2520 24416 2520 24416 0 Inst_W_IO_ConfigMem.Inst_frame0_bit11.Q
rlabel metal2 7896 37352 7896 37352 0 Inst_W_IO_ConfigMem.Inst_frame0_bit12.Q
rlabel metal3 6664 38696 6664 38696 0 Inst_W_IO_ConfigMem.Inst_frame0_bit13.Q
rlabel metal3 12544 34664 12544 34664 0 Inst_W_IO_ConfigMem.Inst_frame0_bit14.Q
rlabel metal2 14056 35616 14056 35616 0 Inst_W_IO_ConfigMem.Inst_frame0_bit15.Q
rlabel metal3 16464 31192 16464 31192 0 Inst_W_IO_ConfigMem.Inst_frame0_bit16.Q
rlabel metal3 17528 31864 17528 31864 0 Inst_W_IO_ConfigMem.Inst_frame0_bit17.Q
rlabel metal2 13160 22456 13160 22456 0 Inst_W_IO_ConfigMem.Inst_frame0_bit18.Q
rlabel metal2 12040 20160 12040 20160 0 Inst_W_IO_ConfigMem.Inst_frame0_bit19.Q
rlabel metal2 7224 18984 7224 18984 0 Inst_W_IO_ConfigMem.Inst_frame0_bit2.Q
rlabel metal2 12264 21000 12264 21000 0 Inst_W_IO_ConfigMem.Inst_frame0_bit20.Q
rlabel metal2 10584 20160 10584 20160 0 Inst_W_IO_ConfigMem.Inst_frame0_bit21.Q
rlabel metal2 15512 14840 15512 14840 0 Inst_W_IO_ConfigMem.Inst_frame0_bit22.Q
rlabel metal2 16520 14280 16520 14280 0 Inst_W_IO_ConfigMem.Inst_frame0_bit23.Q
rlabel metal3 16520 15176 16520 15176 0 Inst_W_IO_ConfigMem.Inst_frame0_bit24.Q
rlabel metal3 17080 20776 17080 20776 0 Inst_W_IO_ConfigMem.Inst_frame0_bit25.Q
rlabel metal2 16072 19824 16072 19824 0 Inst_W_IO_ConfigMem.Inst_frame0_bit26.Q
rlabel metal2 15288 17920 15288 17920 0 Inst_W_IO_ConfigMem.Inst_frame0_bit27.Q
rlabel metal2 16072 18256 16072 18256 0 Inst_W_IO_ConfigMem.Inst_frame0_bit28.Q
rlabel metal3 10304 15400 10304 15400 0 Inst_W_IO_ConfigMem.Inst_frame0_bit29.Q
rlabel metal2 7896 21280 7896 21280 0 Inst_W_IO_ConfigMem.Inst_frame0_bit3.Q
rlabel metal3 10976 15176 10976 15176 0 Inst_W_IO_ConfigMem.Inst_frame0_bit30.Q
rlabel metal3 8792 15736 8792 15736 0 Inst_W_IO_ConfigMem.Inst_frame0_bit31.Q
rlabel metal3 9688 9240 9688 9240 0 Inst_W_IO_ConfigMem.Inst_frame0_bit4.Q
rlabel metal2 11592 9464 11592 9464 0 Inst_W_IO_ConfigMem.Inst_frame0_bit5.Q
rlabel metal2 12376 32032 12376 32032 0 Inst_W_IO_ConfigMem.Inst_frame0_bit6.Q
rlabel metal2 13496 32480 13496 32480 0 Inst_W_IO_ConfigMem.Inst_frame0_bit7.Q
rlabel metal2 17528 30072 17528 30072 0 Inst_W_IO_ConfigMem.Inst_frame0_bit8.Q
rlabel metal2 18536 30576 18536 30576 0 Inst_W_IO_ConfigMem.Inst_frame0_bit9.Q
rlabel metal2 3304 32088 3304 32088 0 Inst_W_IO_ConfigMem.Inst_frame1_bit0.Q
rlabel metal2 2296 31920 2296 31920 0 Inst_W_IO_ConfigMem.Inst_frame1_bit1.Q
rlabel metal2 6776 29904 6776 29904 0 Inst_W_IO_ConfigMem.Inst_frame1_bit10.Q
rlabel metal2 5096 28952 5096 28952 0 Inst_W_IO_ConfigMem.Inst_frame1_bit11.Q
rlabel metal2 2856 35168 2856 35168 0 Inst_W_IO_ConfigMem.Inst_frame1_bit12.Q
rlabel metal2 1512 35560 1512 35560 0 Inst_W_IO_ConfigMem.Inst_frame1_bit13.Q
rlabel metal3 12656 38024 12656 38024 0 Inst_W_IO_ConfigMem.Inst_frame1_bit14.Q
rlabel metal3 11536 38024 11536 38024 0 Inst_W_IO_ConfigMem.Inst_frame1_bit15.Q
rlabel metal2 7784 33208 7784 33208 0 Inst_W_IO_ConfigMem.Inst_frame1_bit16.Q
rlabel metal3 7000 32536 7000 32536 0 Inst_W_IO_ConfigMem.Inst_frame1_bit17.Q
rlabel metal2 3528 25816 3528 25816 0 Inst_W_IO_ConfigMem.Inst_frame1_bit18.Q
rlabel metal2 2688 26824 2688 26824 0 Inst_W_IO_ConfigMem.Inst_frame1_bit19.Q
rlabel metal2 11144 16184 11144 16184 0 Inst_W_IO_ConfigMem.Inst_frame1_bit2.Q
rlabel metal2 2912 28840 2912 28840 0 Inst_W_IO_ConfigMem.Inst_frame1_bit20.Q
rlabel metal2 2856 29848 2856 29848 0 Inst_W_IO_ConfigMem.Inst_frame1_bit21.Q
rlabel metal2 14336 24696 14336 24696 0 Inst_W_IO_ConfigMem.Inst_frame1_bit22.Q
rlabel metal3 15008 24696 15008 24696 0 Inst_W_IO_ConfigMem.Inst_frame1_bit23.Q
rlabel metal3 16240 21448 16240 21448 0 Inst_W_IO_ConfigMem.Inst_frame1_bit24.Q
rlabel metal2 17640 21280 17640 21280 0 Inst_W_IO_ConfigMem.Inst_frame1_bit25.Q
rlabel metal3 4816 27832 4816 27832 0 Inst_W_IO_ConfigMem.Inst_frame1_bit26.Q
rlabel metal2 6552 27552 6552 27552 0 Inst_W_IO_ConfigMem.Inst_frame1_bit27.Q
rlabel metal3 6552 10584 6552 10584 0 Inst_W_IO_ConfigMem.Inst_frame1_bit28.Q
rlabel metal2 8232 10640 8232 10640 0 Inst_W_IO_ConfigMem.Inst_frame1_bit29.Q
rlabel metal2 12264 16296 12264 16296 0 Inst_W_IO_ConfigMem.Inst_frame1_bit3.Q
rlabel metal3 1736 15064 1736 15064 0 Inst_W_IO_ConfigMem.Inst_frame1_bit30.Q
rlabel metal3 2296 15848 2296 15848 0 Inst_W_IO_ConfigMem.Inst_frame1_bit31.Q
rlabel metal2 11200 9240 11200 9240 0 Inst_W_IO_ConfigMem.Inst_frame1_bit4.Q
rlabel metal2 12152 11424 12152 11424 0 Inst_W_IO_ConfigMem.Inst_frame1_bit5.Q
rlabel metal2 14280 23856 14280 23856 0 Inst_W_IO_ConfigMem.Inst_frame1_bit6.Q
rlabel metal2 13160 24584 13160 24584 0 Inst_W_IO_ConfigMem.Inst_frame1_bit7.Q
rlabel metal2 14728 23072 14728 23072 0 Inst_W_IO_ConfigMem.Inst_frame1_bit8.Q
rlabel metal3 16632 22344 16632 22344 0 Inst_W_IO_ConfigMem.Inst_frame1_bit9.Q
rlabel metal3 8792 27832 8792 27832 0 Inst_W_IO_ConfigMem.Inst_frame2_bit0.Q
rlabel metal2 10472 28504 10472 28504 0 Inst_W_IO_ConfigMem.Inst_frame2_bit1.Q
rlabel metal3 4144 12936 4144 12936 0 Inst_W_IO_ConfigMem.Inst_frame2_bit10.Q
rlabel metal2 5880 13216 5880 13216 0 Inst_W_IO_ConfigMem.Inst_frame2_bit11.Q
rlabel metal3 6496 39480 6496 39480 0 Inst_W_IO_ConfigMem.Inst_frame2_bit12.Q
rlabel metal3 6552 40376 6552 40376 0 Inst_W_IO_ConfigMem.Inst_frame2_bit13.Q
rlabel metal2 5152 23912 5152 23912 0 Inst_W_IO_ConfigMem.Inst_frame2_bit14.Q
rlabel metal3 5824 27160 5824 27160 0 Inst_W_IO_ConfigMem.Inst_frame2_bit15.Q
rlabel metal2 9800 30464 9800 30464 0 Inst_W_IO_ConfigMem.Inst_frame2_bit16.Q
rlabel metal2 11032 30576 11032 30576 0 Inst_W_IO_ConfigMem.Inst_frame2_bit17.Q
rlabel metal2 7896 24976 7896 24976 0 Inst_W_IO_ConfigMem.Inst_frame2_bit18.Q
rlabel metal2 9240 25368 9240 25368 0 Inst_W_IO_ConfigMem.Inst_frame2_bit19.Q
rlabel metal2 8232 20888 8232 20888 0 Inst_W_IO_ConfigMem.Inst_frame2_bit2.Q
rlabel metal3 8960 12152 8960 12152 0 Inst_W_IO_ConfigMem.Inst_frame2_bit20.Q
rlabel metal2 10696 12432 10696 12432 0 Inst_W_IO_ConfigMem.Inst_frame2_bit21.Q
rlabel metal2 15176 27552 15176 27552 0 Inst_W_IO_ConfigMem.Inst_frame2_bit22.Q
rlabel metal2 15288 28504 15288 28504 0 Inst_W_IO_ConfigMem.Inst_frame2_bit23.Q
rlabel metal2 19096 28336 19096 28336 0 Inst_W_IO_ConfigMem.Inst_frame2_bit24.Q
rlabel metal2 19824 28728 19824 28728 0 Inst_W_IO_ConfigMem.Inst_frame2_bit25.Q
rlabel metal2 12936 39760 12936 39760 0 Inst_W_IO_ConfigMem.Inst_frame2_bit26.Q
rlabel metal3 11424 39592 11424 39592 0 Inst_W_IO_ConfigMem.Inst_frame2_bit27.Q
rlabel metal2 6776 34608 6776 34608 0 Inst_W_IO_ConfigMem.Inst_frame2_bit28.Q
rlabel metal3 4872 34888 4872 34888 0 Inst_W_IO_ConfigMem.Inst_frame2_bit29.Q
rlabel metal3 9352 22456 9352 22456 0 Inst_W_IO_ConfigMem.Inst_frame2_bit3.Q
rlabel metal2 3696 20888 3696 20888 0 Inst_W_IO_ConfigMem.Inst_frame2_bit30.Q
rlabel metal3 2128 19432 2128 19432 0 Inst_W_IO_ConfigMem.Inst_frame2_bit31.Q
rlabel metal3 9240 11368 9240 11368 0 Inst_W_IO_ConfigMem.Inst_frame2_bit4.Q
rlabel metal2 11480 12432 11480 12432 0 Inst_W_IO_ConfigMem.Inst_frame2_bit5.Q
rlabel metal2 12992 27272 12992 27272 0 Inst_W_IO_ConfigMem.Inst_frame2_bit6.Q
rlabel metal3 13440 28616 13440 28616 0 Inst_W_IO_ConfigMem.Inst_frame2_bit7.Q
rlabel metal2 18032 25480 18032 25480 0 Inst_W_IO_ConfigMem.Inst_frame2_bit8.Q
rlabel metal3 19320 25480 19320 25480 0 Inst_W_IO_ConfigMem.Inst_frame2_bit9.Q
rlabel metal2 14728 12488 14728 12488 0 Inst_W_IO_ConfigMem.Inst_frame3_bit22.Q
rlabel metal3 20104 20888 20104 20888 0 Inst_W_IO_ConfigMem.Inst_frame3_bit23.Q
rlabel metal3 16408 35112 16408 35112 0 Inst_W_IO_ConfigMem.Inst_frame3_bit24.Q
rlabel metal4 19432 32816 19432 32816 0 Inst_W_IO_ConfigMem.Inst_frame3_bit25.Q
rlabel metal2 4760 16632 4760 16632 0 Inst_W_IO_ConfigMem.Inst_frame3_bit26.Q
rlabel metal2 5992 16016 5992 16016 0 Inst_W_IO_ConfigMem.Inst_frame3_bit27.Q
rlabel metal2 8232 35504 8232 35504 0 Inst_W_IO_ConfigMem.Inst_frame3_bit28.Q
rlabel metal3 9184 35672 9184 35672 0 Inst_W_IO_ConfigMem.Inst_frame3_bit29.Q
rlabel metal3 4816 21784 4816 21784 0 Inst_W_IO_ConfigMem.Inst_frame3_bit30.Q
rlabel metal2 6552 20888 6552 20888 0 Inst_W_IO_ConfigMem.Inst_frame3_bit31.Q
rlabel metal2 14392 10864 14392 10864 0 Inst_W_IO_switch_matrix.E1BEG0
rlabel metal2 19880 21168 19880 21168 0 Inst_W_IO_switch_matrix.E1BEG1
rlabel metal3 14616 36456 14616 36456 0 Inst_W_IO_switch_matrix.E1BEG2
rlabel metal3 18648 32760 18648 32760 0 Inst_W_IO_switch_matrix.E1BEG3
rlabel metal2 5544 13384 5544 13384 0 Inst_W_IO_switch_matrix.E2BEG0
rlabel metal3 8624 35560 8624 35560 0 Inst_W_IO_switch_matrix.E2BEG1
rlabel metal2 5992 22848 5992 22848 0 Inst_W_IO_switch_matrix.E2BEG2
rlabel metal2 10080 27608 10080 27608 0 Inst_W_IO_switch_matrix.E2BEG3
rlabel metal2 9912 23240 9912 23240 0 Inst_W_IO_switch_matrix.E2BEG4
rlabel metal2 10920 12264 10920 12264 0 Inst_W_IO_switch_matrix.E2BEG5
rlabel metal2 13944 29512 13944 29512 0 Inst_W_IO_switch_matrix.E2BEG6
rlabel metal3 18872 24696 18872 24696 0 Inst_W_IO_switch_matrix.E2BEG7
rlabel metal2 5208 11424 5208 11424 0 Inst_W_IO_switch_matrix.E2BEGb0
rlabel metal2 8400 40264 8400 40264 0 Inst_W_IO_switch_matrix.E2BEGb1
rlabel metal2 5656 24304 5656 24304 0 Inst_W_IO_switch_matrix.E2BEGb2
rlabel metal2 10472 30688 10472 30688 0 Inst_W_IO_switch_matrix.E2BEGb3
rlabel metal2 8568 25032 8568 25032 0 Inst_W_IO_switch_matrix.E2BEGb4
rlabel metal2 10080 12040 10080 12040 0 Inst_W_IO_switch_matrix.E2BEGb5
rlabel metal2 15624 27440 15624 27440 0 Inst_W_IO_switch_matrix.E2BEGb6
rlabel metal2 19488 27832 19488 27832 0 Inst_W_IO_switch_matrix.E2BEGb7
rlabel metal2 5992 28168 5992 28168 0 Inst_W_IO_switch_matrix.E6BEG0
rlabel metal2 7784 10192 7784 10192 0 Inst_W_IO_switch_matrix.E6BEG1
rlabel metal2 13608 35336 13608 35336 0 Inst_W_IO_switch_matrix.E6BEG10
rlabel metal2 17752 32648 17752 32648 0 Inst_W_IO_switch_matrix.E6BEG11
rlabel metal2 2296 12824 2296 12824 0 Inst_W_IO_switch_matrix.E6BEG2
rlabel metal2 6104 39984 6104 39984 0 Inst_W_IO_switch_matrix.E6BEG3
rlabel metal3 6664 21336 6664 21336 0 Inst_W_IO_switch_matrix.E6BEG4
rlabel metal2 11088 9912 11088 9912 0 Inst_W_IO_switch_matrix.E6BEG5
rlabel metal2 13048 32256 13048 32256 0 Inst_W_IO_switch_matrix.E6BEG6
rlabel metal2 17808 30856 17808 30856 0 Inst_W_IO_switch_matrix.E6BEG7
rlabel metal2 3304 23520 3304 23520 0 Inst_W_IO_switch_matrix.E6BEG8
rlabel metal2 8568 37576 8568 37576 0 Inst_W_IO_switch_matrix.E6BEG9
rlabel metal2 12488 39984 12488 39984 0 Inst_W_IO_switch_matrix.EE4BEG0
rlabel metal2 6160 35112 6160 35112 0 Inst_W_IO_switch_matrix.EE4BEG1
rlabel metal2 12768 39032 12768 39032 0 Inst_W_IO_switch_matrix.EE4BEG10
rlabel metal2 7336 32872 7336 32872 0 Inst_W_IO_switch_matrix.EE4BEG11
rlabel metal2 3752 25872 3752 25872 0 Inst_W_IO_switch_matrix.EE4BEG12
rlabel metal2 3416 30576 3416 30576 0 Inst_W_IO_switch_matrix.EE4BEG13
rlabel metal3 14336 24584 14336 24584 0 Inst_W_IO_switch_matrix.EE4BEG14
rlabel metal2 14728 20664 14728 20664 0 Inst_W_IO_switch_matrix.EE4BEG15
rlabel metal3 2632 20888 2632 20888 0 Inst_W_IO_switch_matrix.EE4BEG2
rlabel metal2 3752 32088 3752 32088 0 Inst_W_IO_switch_matrix.EE4BEG3
rlabel metal2 11816 16576 11816 16576 0 Inst_W_IO_switch_matrix.EE4BEG4
rlabel metal3 13720 10584 13720 10584 0 Inst_W_IO_switch_matrix.EE4BEG5
rlabel metal2 13944 24136 13944 24136 0 Inst_W_IO_switch_matrix.EE4BEG6
rlabel metal2 15176 22736 15176 22736 0 Inst_W_IO_switch_matrix.EE4BEG7
rlabel metal2 6160 30408 6160 30408 0 Inst_W_IO_switch_matrix.EE4BEG8
rlabel metal3 2744 33544 2744 33544 0 Inst_W_IO_switch_matrix.EE4BEG9
rlabel metal2 16744 39200 16744 39200 0 UserCLK
rlabel metal2 18648 37968 18648 37968 0 UserCLK_regs
rlabel metal2 896 55944 896 55944 0 UserCLKo
rlabel metal3 27314 280 27314 280 0 W1END[0]
rlabel metal3 26922 728 26922 728 0 W1END[1]
rlabel metal3 27818 1176 27818 1176 0 W1END[2]
rlabel metal3 27538 1624 27538 1624 0 W1END[3]
rlabel metal3 28042 5656 28042 5656 0 W2END[0]
rlabel metal3 27538 6104 27538 6104 0 W2END[1]
rlabel metal2 27496 6216 27496 6216 0 W2END[2]
rlabel metal3 27986 7000 27986 7000 0 W2END[3]
rlabel metal3 28042 7448 28042 7448 0 W2END[4]
rlabel metal2 27496 7672 27496 7672 0 W2END[5]
rlabel metal3 27594 8344 27594 8344 0 W2END[6]
rlabel metal2 27552 8456 27552 8456 0 W2END[7]
rlabel metal3 27594 2072 27594 2072 0 W2MID[0]
rlabel metal3 28042 2520 28042 2520 0 W2MID[1]
rlabel metal3 27538 2968 27538 2968 0 W2MID[2]
rlabel metal2 27496 3080 27496 3080 0 W2MID[3]
rlabel metal3 27986 3864 27986 3864 0 W2MID[4]
rlabel metal3 27538 4312 27538 4312 0 W2MID[5]
rlabel metal2 27496 4536 27496 4536 0 W2MID[6]
rlabel metal3 27594 5208 27594 5208 0 W2MID[7]
rlabel metal3 27986 16408 27986 16408 0 W6END[0]
rlabel metal2 25928 21112 25928 21112 0 W6END[10]
rlabel metal3 27986 21336 27986 21336 0 W6END[11]
rlabel metal2 26600 17248 26600 17248 0 W6END[1]
rlabel metal2 27496 17080 27496 17080 0 W6END[2]
rlabel metal2 26712 17976 26712 17976 0 W6END[3]
rlabel metal3 27986 18200 27986 18200 0 W6END[4]
rlabel metal2 26600 18928 26600 18928 0 W6END[5]
rlabel metal2 27496 18760 27496 18760 0 W6END[6]
rlabel metal3 27986 19544 27986 19544 0 W6END[7]
rlabel metal2 26600 20384 26600 20384 0 W6END[8]
rlabel metal2 27496 20216 27496 20216 0 W6END[9]
rlabel metal3 27538 9240 27538 9240 0 WW4END[0]
rlabel metal3 27538 13720 27538 13720 0 WW4END[10]
rlabel metal2 27496 13944 27496 13944 0 WW4END[11]
rlabel metal3 27594 14616 27594 14616 0 WW4END[12]
rlabel metal3 27986 15064 27986 15064 0 WW4END[13]
rlabel metal2 26600 15792 26600 15792 0 WW4END[14]
rlabel metal2 27496 15624 27496 15624 0 WW4END[15]
rlabel metal2 27496 9352 27496 9352 0 WW4END[1]
rlabel metal3 27986 10136 27986 10136 0 WW4END[2]
rlabel metal3 27538 10584 27538 10584 0 WW4END[3]
rlabel metal2 27496 10808 27496 10808 0 WW4END[4]
rlabel metal3 27594 11480 27594 11480 0 WW4END[5]
rlabel metal3 28042 11928 28042 11928 0 WW4END[6]
rlabel metal3 27538 12376 27538 12376 0 WW4END[7]
rlabel metal2 27496 12488 27496 12488 0 WW4END[8]
rlabel metal3 27986 13272 27986 13272 0 WW4END[9]
rlabel metal2 16688 22120 16688 22120 0 _000_
rlabel metal3 16184 18200 16184 18200 0 _001_
rlabel metal2 17416 13720 17416 13720 0 _002_
rlabel metal2 16184 13832 16184 13832 0 _003_
rlabel metal3 10976 21336 10976 21336 0 _004_
rlabel metal2 16184 13160 16184 13160 0 _005_
rlabel metal2 10136 14672 10136 14672 0 _006_
rlabel metal2 15960 17080 15960 17080 0 _007_
rlabel metal2 16184 17864 16184 17864 0 _008_
rlabel metal2 14560 17752 14560 17752 0 _009_
rlabel metal2 16520 18480 16520 18480 0 _010_
rlabel metal2 16744 19432 16744 19432 0 _011_
rlabel metal3 16352 18648 16352 18648 0 _012_
rlabel metal2 13776 16856 13776 16856 0 _013_
rlabel metal3 16408 20216 16408 20216 0 _014_
rlabel metal2 14280 18424 14280 18424 0 _015_
rlabel metal2 14616 16688 14616 16688 0 _016_
rlabel metal2 13160 18200 13160 18200 0 _017_
rlabel metal2 12936 17752 12936 17752 0 _018_
rlabel metal3 10808 19432 10808 19432 0 _019_
rlabel metal3 10192 20888 10192 20888 0 _020_
rlabel metal2 13832 23128 13832 23128 0 _021_
rlabel metal3 11816 20776 11816 20776 0 _022_
rlabel metal2 12992 20104 12992 20104 0 _023_
rlabel metal2 12320 19992 12320 19992 0 _024_
rlabel metal2 11648 23352 11648 23352 0 _025_
rlabel metal2 11816 21784 11816 21784 0 _026_
rlabel metal2 15400 13440 15400 13440 0 _027_
rlabel metal3 16688 14280 16688 14280 0 _028_
rlabel metal2 16744 14784 16744 14784 0 _029_
rlabel metal2 17416 14224 17416 14224 0 _030_
rlabel metal2 15288 15512 15288 15512 0 _031_
rlabel metal2 16296 15400 16296 15400 0 _032_
rlabel metal2 17640 15288 17640 15288 0 _033_
rlabel metal2 10248 16912 10248 16912 0 _034_
rlabel metal2 11256 16072 11256 16072 0 _035_
rlabel metal2 10920 14504 10920 14504 0 _036_
rlabel metal3 10248 14280 10248 14280 0 _037_
rlabel metal2 11144 14896 11144 14896 0 _038_
rlabel metal3 9688 16072 9688 16072 0 _039_
rlabel metal3 10528 15512 10528 15512 0 _040_
rlabel metal3 10136 15288 10136 15288 0 _041_
rlabel metal2 18592 39480 18592 39480 0 clknet_0_UserCLK
rlabel metal2 16632 35616 16632 35616 0 clknet_0_UserCLK_regs
rlabel metal2 15512 36904 15512 36904 0 clknet_1_0__leaf_UserCLK
rlabel metal2 16744 36120 16744 36120 0 clknet_1_0__leaf_UserCLK_regs
rlabel metal2 18424 41104 18424 41104 0 clknet_1_1__leaf_UserCLK_regs
rlabel metal2 14504 11200 14504 11200 0 net1
rlabel metal3 2492 35560 2492 35560 0 net10
rlabel metal2 2912 12376 2912 12376 0 net100
rlabel metal2 14896 13048 14896 13048 0 net101
rlabel metal2 16408 17584 16408 17584 0 net102
rlabel metal2 10584 13328 10584 13328 0 net103
rlabel metal2 24920 17528 24920 17528 0 net104
rlabel metal2 26264 21392 26264 21392 0 net105
rlabel metal2 14896 24472 14896 24472 0 net106
rlabel metal3 22344 30072 22344 30072 0 net107
rlabel metal2 26376 22064 26376 22064 0 net108
rlabel metal3 22456 24360 22456 24360 0 net109
rlabel metal2 15624 32872 15624 32872 0 net11
rlabel metal2 26264 23576 26264 23576 0 net110
rlabel metal3 17752 25592 17752 25592 0 net111
rlabel metal2 26264 24360 26264 24360 0 net112
rlabel metal3 26152 25480 26152 25480 0 net113
rlabel metal2 14728 28616 14728 28616 0 net114
rlabel metal2 26264 26096 26264 26096 0 net115
rlabel metal3 5544 9912 5544 9912 0 net116
rlabel metal3 20664 27496 20664 27496 0 net117
rlabel metal3 24248 24920 24248 24920 0 net118
rlabel metal2 26152 29568 26152 29568 0 net119
rlabel metal3 2520 26040 2520 26040 0 net12
rlabel metal2 9464 27440 9464 27440 0 net120
rlabel metal3 26152 25144 26152 25144 0 net121
rlabel metal2 16184 27944 16184 27944 0 net122
rlabel metal2 20104 28000 20104 28000 0 net123
rlabel metal2 24248 33320 24248 33320 0 net124
rlabel metal3 18872 42728 18872 42728 0 net125
rlabel metal2 25704 43960 25704 43960 0 net126
rlabel metal3 9184 9688 9184 9688 0 net127
rlabel metal2 25424 23800 25424 23800 0 net128
rlabel metal2 24920 40096 24920 40096 0 net129
rlabel metal2 1400 25368 1400 25368 0 net13
rlabel metal2 5544 22904 5544 22904 0 net130
rlabel metal2 24696 40432 24696 40432 0 net131
rlabel metal3 23212 41832 23212 41832 0 net132
rlabel metal2 24192 41160 24192 41160 0 net133
rlabel metal2 26096 42728 26096 42728 0 net134
rlabel metal2 25872 43064 25872 43064 0 net135
rlabel metal3 19880 32816 19880 32816 0 net136
rlabel metal2 26376 37576 26376 37576 0 net137
rlabel metal2 25816 35336 25816 35336 0 net138
rlabel metal2 16912 30632 16912 30632 0 net139
rlabel metal3 1008 20440 1008 20440 0 net14
rlabel metal2 2744 30016 2744 30016 0 net140
rlabel metal2 15512 25592 15512 25592 0 net141
rlabel metal3 25872 25928 25872 25928 0 net142
rlabel metal2 26152 33712 26152 33712 0 net143
rlabel metal4 1400 22848 1400 22848 0 net144
rlabel metal2 26264 32984 26264 32984 0 net145
rlabel metal2 12376 16968 12376 16968 0 net146
rlabel metal2 26376 14616 26376 14616 0 net147
rlabel metal3 16184 27888 16184 27888 0 net148
rlabel metal2 16968 23576 16968 23576 0 net149
rlabel metal2 7280 12040 7280 12040 0 net15
rlabel metal2 26376 35000 26376 35000 0 net150
rlabel metal2 24808 34384 24808 34384 0 net151
rlabel metal2 24920 42728 24920 42728 0 net152
rlabel metal2 3192 9968 3192 9968 0 net153
rlabel metal2 26376 49280 26376 49280 0 net154
rlabel metal2 24696 48944 24696 48944 0 net155
rlabel metal3 18648 50680 18648 50680 0 net156
rlabel metal3 24920 48384 24920 48384 0 net157
rlabel metal3 22064 51240 22064 51240 0 net158
rlabel metal2 24696 50512 24696 50512 0 net159
rlabel metal2 9464 12152 9464 12152 0 net16
rlabel metal3 21168 52136 21168 52136 0 net160
rlabel metal2 26264 52584 26264 52584 0 net161
rlabel metal3 15624 52248 15624 52248 0 net162
rlabel metal2 26376 43232 26376 43232 0 net163
rlabel metal3 14392 8904 14392 8904 0 net164
rlabel metal3 24976 52808 24976 52808 0 net165
rlabel metal2 26264 54320 26264 54320 0 net166
rlabel metal3 22904 53480 22904 53480 0 net167
rlabel metal3 23520 55272 23520 55272 0 net168
rlabel metal2 24864 47992 24864 47992 0 net169
rlabel metal2 14224 14616 14224 14616 0 net17
rlabel metal3 17024 54376 17024 54376 0 net170
rlabel metal2 22904 52528 22904 52528 0 net171
rlabel metal2 5880 11200 5880 11200 0 net172
rlabel metal2 21560 54152 21560 54152 0 net173
rlabel metal3 4648 18424 4648 18424 0 net174
rlabel metal2 25032 51352 25032 51352 0 net175
rlabel metal2 3304 12320 3304 12320 0 net176
rlabel metal3 22120 24584 22120 24584 0 net177
rlabel metal3 26208 46536 26208 46536 0 net178
rlabel metal3 25816 45864 25816 45864 0 net179
rlabel metal3 17920 24584 17920 24584 0 net18
rlabel metal2 26264 47096 26264 47096 0 net180
rlabel metal2 24472 46536 24472 46536 0 net181
rlabel metal3 21056 48104 21056 48104 0 net182
rlabel metal2 24696 47152 24696 47152 0 net183
rlabel metal3 7448 43624 7448 43624 0 net184
rlabel metal3 19432 53592 19432 53592 0 net185
rlabel metal2 21784 53088 21784 53088 0 net186
rlabel metal2 22680 53144 22680 53144 0 net187
rlabel metal2 20216 55720 20216 55720 0 net188
rlabel metal3 23632 49896 23632 49896 0 net189
rlabel metal2 18312 23352 18312 23352 0 net19
rlabel metal2 25032 48048 25032 48048 0 net190
rlabel metal2 21952 52248 21952 52248 0 net191
rlabel metal2 25760 48328 25760 48328 0 net192
rlabel metal2 23520 50680 23520 50680 0 net193
rlabel metal2 22792 52416 22792 52416 0 net194
rlabel metal3 2800 55944 2800 55944 0 net195
rlabel metal2 5264 55440 5264 55440 0 net196
rlabel metal2 18872 38192 18872 38192 0 net197
rlabel metal2 21112 55272 21112 55272 0 net198
rlabel metal3 14784 54600 14784 54600 0 net199
rlabel metal2 7672 12040 7672 12040 0 net2
rlabel metal3 18872 26264 18872 26264 0 net20
rlabel metal3 11592 55328 11592 55328 0 net200
rlabel metal2 24360 51632 24360 51632 0 net201
rlabel metal2 22232 53704 22232 53704 0 net202
rlabel metal2 23240 53480 23240 53480 0 net203
rlabel metal2 1400 54376 1400 54376 0 net204
rlabel metal3 2576 14952 2576 14952 0 net205
rlabel metal2 13496 11032 13496 11032 0 net206
rlabel metal2 2632 18088 2632 18088 0 net21
rlabel metal3 5152 17864 5152 17864 0 net22
rlabel metal2 4984 11592 4984 11592 0 net23
rlabel metal2 1176 51464 1176 51464 0 net24
rlabel metal2 2240 16296 2240 16296 0 net25
rlabel metal3 952 52808 952 52808 0 net26
rlabel metal2 17976 26264 17976 26264 0 net27
rlabel metal2 17528 28672 17528 28672 0 net28
rlabel metal3 6832 12152 6832 12152 0 net29
rlabel metal3 1456 16632 1456 16632 0 net3
rlabel metal2 5208 13496 5208 13496 0 net30
rlabel metal2 2184 23632 2184 23632 0 net31
rlabel metal2 18144 24808 18144 24808 0 net32
rlabel metal2 4424 10808 4424 10808 0 net33
rlabel metal3 1064 30072 1064 30072 0 net34
rlabel metal3 1512 32648 1512 32648 0 net35
rlabel metal2 1064 20328 1064 20328 0 net36
rlabel metal3 18536 15960 18536 15960 0 net37
rlabel metal3 4424 16856 4424 16856 0 net38
rlabel metal3 8512 9016 8512 9016 0 net39
rlabel metal2 2520 23016 2520 23016 0 net4
rlabel metal2 2296 23352 2296 23352 0 net40
rlabel metal3 10024 32536 10024 32536 0 net41
rlabel metal2 1568 51688 1568 51688 0 net42
rlabel metal2 1624 10752 1624 10752 0 net43
rlabel metal2 7112 11816 7112 11816 0 net44
rlabel metal2 10136 7896 10136 7896 0 net45
rlabel metal2 2520 17304 2520 17304 0 net46
rlabel metal2 1512 19040 1512 19040 0 net47
rlabel metal2 16968 26376 16968 26376 0 net48
rlabel metal2 18480 22904 18480 22904 0 net49
rlabel metal2 5656 13776 5656 13776 0 net5
rlabel metal2 5544 4844 5544 4844 0 net50
rlabel metal3 12040 1064 12040 1064 0 net51
rlabel metal3 22176 1064 22176 1064 0 net52
rlabel metal3 20160 1176 20160 1176 0 net53
rlabel metal2 26544 1288 26544 1288 0 net54
rlabel metal2 25928 2072 25928 2072 0 net55
rlabel metal2 26936 5488 26936 5488 0 net56
rlabel metal3 20944 6552 20944 6552 0 net57
rlabel metal2 26936 6160 26936 6160 0 net58
rlabel metal3 27104 6664 27104 6664 0 net59
rlabel metal2 2856 36848 2856 36848 0 net6
rlabel metal2 26264 12096 26264 12096 0 net60
rlabel metal3 19880 7448 19880 7448 0 net61
rlabel metal2 26040 9408 26040 9408 0 net62
rlabel metal2 26936 8064 26936 8064 0 net63
rlabel metal3 23632 2856 23632 2856 0 net64
rlabel metal2 26936 4032 26936 4032 0 net65
rlabel metal3 19712 3416 19712 3416 0 net66
rlabel metal3 27384 2856 27384 2856 0 net67
rlabel metal3 26936 3472 26936 3472 0 net68
rlabel metal2 26096 5208 26096 5208 0 net69
rlabel metal3 2408 40264 2408 40264 0 net7
rlabel metal2 27104 4424 27104 4424 0 net70
rlabel metal2 7672 14616 7672 14616 0 net71
rlabel metal3 25256 26208 25256 26208 0 net72
rlabel metal2 25368 20832 25368 20832 0 net73
rlabel metal2 2408 31024 2408 31024 0 net74
rlabel metal2 25928 18536 25928 18536 0 net75
rlabel metal3 17080 17640 17080 17640 0 net76
rlabel metal2 26152 20104 26152 20104 0 net77
rlabel metal2 26936 17808 26936 17808 0 net78
rlabel metal2 26040 19712 26040 19712 0 net79
rlabel metal2 3192 35392 3192 35392 0 net8
rlabel metal2 8120 40040 8120 40040 0 net80
rlabel metal2 5320 14448 5320 14448 0 net81
rlabel metal3 25760 24808 25760 24808 0 net82
rlabel metal2 1848 31248 1848 31248 0 net83
rlabel metal3 23520 10024 23520 10024 0 net84
rlabel metal2 26152 13160 26152 13160 0 net85
rlabel metal3 20216 13552 20216 13552 0 net86
rlabel metal2 26152 16632 26152 16632 0 net87
rlabel metal2 26936 14112 26936 14112 0 net88
rlabel metal2 18536 24080 18536 24080 0 net89
rlabel metal2 1736 35784 1736 35784 0 net9
rlabel metal2 4536 14280 4536 14280 0 net90
rlabel metal2 27048 10584 27048 10584 0 net91
rlabel metal2 12376 9856 12376 9856 0 net92
rlabel metal2 25928 13832 25928 13832 0 net93
rlabel metal3 18984 10696 18984 10696 0 net94
rlabel metal3 16800 12264 16800 12264 0 net95
rlabel metal3 23548 11256 23548 11256 0 net96
rlabel metal2 6440 13048 6440 13048 0 net97
rlabel metal3 27440 12264 27440 12264 0 net98
rlabel metal2 27104 12824 27104 12824 0 net99
<< properties >>
string FIXED_BBOX 0 0 28560 57456
<< end >>
