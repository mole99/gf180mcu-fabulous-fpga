module RegFile (UserCLK,
    UserCLKo,
    E1BEG,
    E1END,
    E2BEG,
    E2BEGb,
    E2END,
    E2MID,
    E6BEG,
    E6END,
    EE4BEG,
    EE4END,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N1END,
    N2BEG,
    N2BEGb,
    N2END,
    N2MID,
    N4BEG,
    N4END,
    NN4BEG,
    NN4END,
    S1BEG,
    S1END,
    S2BEG,
    S2BEGb,
    S2END,
    S2MID,
    S4BEG,
    S4END,
    SS4BEG,
    SS4END,
    W1BEG,
    W1END,
    W2BEG,
    W2BEGb,
    W2END,
    W2MID,
    W6BEG,
    W6END,
    WW4BEG,
    WW4END);
 input UserCLK;
 output UserCLKo;
 output [3:0] E1BEG;
 input [3:0] E1END;
 output [7:0] E2BEG;
 output [7:0] E2BEGb;
 input [7:0] E2END;
 input [7:0] E2MID;
 output [11:0] E6BEG;
 input [11:0] E6END;
 output [15:0] EE4BEG;
 input [15:0] EE4END;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 input [3:0] N1END;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 input [7:0] N2END;
 input [7:0] N2MID;
 output [15:0] N4BEG;
 input [15:0] N4END;
 output [15:0] NN4BEG;
 input [15:0] NN4END;
 output [3:0] S1BEG;
 input [3:0] S1END;
 output [7:0] S2BEG;
 output [7:0] S2BEGb;
 input [7:0] S2END;
 input [7:0] S2MID;
 output [15:0] S4BEG;
 input [15:0] S4END;
 output [15:0] SS4BEG;
 input [15:0] SS4END;
 output [3:0] W1BEG;
 input [3:0] W1END;
 output [7:0] W2BEG;
 output [7:0] W2BEGb;
 input [7:0] W2END;
 input [7:0] W2MID;
 output [11:0] W6BEG;
 input [11:0] W6END;
 output [15:0] WW4BEG;
 input [15:0] WW4END;

 wire AD0;
 wire AD1;
 wire AD2;
 wire AD3;
 wire A_ADR0;
 wire BD0;
 wire BD1;
 wire BD2;
 wire BD3;
 wire B_ADR0;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire \Inst_RegFile_32x4.AD_comb[0] ;
 wire \Inst_RegFile_32x4.AD_comb[1] ;
 wire \Inst_RegFile_32x4.AD_comb[2] ;
 wire \Inst_RegFile_32x4.AD_comb[3] ;
 wire \Inst_RegFile_32x4.AD_reg[0] ;
 wire \Inst_RegFile_32x4.AD_reg[1] ;
 wire \Inst_RegFile_32x4.AD_reg[2] ;
 wire \Inst_RegFile_32x4.AD_reg[3] ;
 wire \Inst_RegFile_32x4.BD_comb[0] ;
 wire \Inst_RegFile_32x4.BD_comb[1] ;
 wire \Inst_RegFile_32x4.BD_comb[2] ;
 wire \Inst_RegFile_32x4.BD_comb[3] ;
 wire \Inst_RegFile_32x4.BD_reg[0] ;
 wire \Inst_RegFile_32x4.BD_reg[1] ;
 wire \Inst_RegFile_32x4.BD_reg[2] ;
 wire \Inst_RegFile_32x4.BD_reg[3] ;
 wire \Inst_RegFile_32x4.mem[0][0] ;
 wire \Inst_RegFile_32x4.mem[0][1] ;
 wire \Inst_RegFile_32x4.mem[0][2] ;
 wire \Inst_RegFile_32x4.mem[0][3] ;
 wire \Inst_RegFile_32x4.mem[10][0] ;
 wire \Inst_RegFile_32x4.mem[10][1] ;
 wire \Inst_RegFile_32x4.mem[10][2] ;
 wire \Inst_RegFile_32x4.mem[10][3] ;
 wire \Inst_RegFile_32x4.mem[11][0] ;
 wire \Inst_RegFile_32x4.mem[11][1] ;
 wire \Inst_RegFile_32x4.mem[11][2] ;
 wire \Inst_RegFile_32x4.mem[11][3] ;
 wire \Inst_RegFile_32x4.mem[12][0] ;
 wire \Inst_RegFile_32x4.mem[12][1] ;
 wire \Inst_RegFile_32x4.mem[12][2] ;
 wire \Inst_RegFile_32x4.mem[12][3] ;
 wire \Inst_RegFile_32x4.mem[13][0] ;
 wire \Inst_RegFile_32x4.mem[13][1] ;
 wire \Inst_RegFile_32x4.mem[13][2] ;
 wire \Inst_RegFile_32x4.mem[13][3] ;
 wire \Inst_RegFile_32x4.mem[14][0] ;
 wire \Inst_RegFile_32x4.mem[14][1] ;
 wire \Inst_RegFile_32x4.mem[14][2] ;
 wire \Inst_RegFile_32x4.mem[14][3] ;
 wire \Inst_RegFile_32x4.mem[15][0] ;
 wire \Inst_RegFile_32x4.mem[15][1] ;
 wire \Inst_RegFile_32x4.mem[15][2] ;
 wire \Inst_RegFile_32x4.mem[15][3] ;
 wire \Inst_RegFile_32x4.mem[16][0] ;
 wire \Inst_RegFile_32x4.mem[16][1] ;
 wire \Inst_RegFile_32x4.mem[16][2] ;
 wire \Inst_RegFile_32x4.mem[16][3] ;
 wire \Inst_RegFile_32x4.mem[17][0] ;
 wire \Inst_RegFile_32x4.mem[17][1] ;
 wire \Inst_RegFile_32x4.mem[17][2] ;
 wire \Inst_RegFile_32x4.mem[17][3] ;
 wire \Inst_RegFile_32x4.mem[18][0] ;
 wire \Inst_RegFile_32x4.mem[18][1] ;
 wire \Inst_RegFile_32x4.mem[18][2] ;
 wire \Inst_RegFile_32x4.mem[18][3] ;
 wire \Inst_RegFile_32x4.mem[19][0] ;
 wire \Inst_RegFile_32x4.mem[19][1] ;
 wire \Inst_RegFile_32x4.mem[19][2] ;
 wire \Inst_RegFile_32x4.mem[19][3] ;
 wire \Inst_RegFile_32x4.mem[1][0] ;
 wire \Inst_RegFile_32x4.mem[1][1] ;
 wire \Inst_RegFile_32x4.mem[1][2] ;
 wire \Inst_RegFile_32x4.mem[1][3] ;
 wire \Inst_RegFile_32x4.mem[20][0] ;
 wire \Inst_RegFile_32x4.mem[20][1] ;
 wire \Inst_RegFile_32x4.mem[20][2] ;
 wire \Inst_RegFile_32x4.mem[20][3] ;
 wire \Inst_RegFile_32x4.mem[21][0] ;
 wire \Inst_RegFile_32x4.mem[21][1] ;
 wire \Inst_RegFile_32x4.mem[21][2] ;
 wire \Inst_RegFile_32x4.mem[21][3] ;
 wire \Inst_RegFile_32x4.mem[22][0] ;
 wire \Inst_RegFile_32x4.mem[22][1] ;
 wire \Inst_RegFile_32x4.mem[22][2] ;
 wire \Inst_RegFile_32x4.mem[22][3] ;
 wire \Inst_RegFile_32x4.mem[23][0] ;
 wire \Inst_RegFile_32x4.mem[23][1] ;
 wire \Inst_RegFile_32x4.mem[23][2] ;
 wire \Inst_RegFile_32x4.mem[23][3] ;
 wire \Inst_RegFile_32x4.mem[24][0] ;
 wire \Inst_RegFile_32x4.mem[24][1] ;
 wire \Inst_RegFile_32x4.mem[24][2] ;
 wire \Inst_RegFile_32x4.mem[24][3] ;
 wire \Inst_RegFile_32x4.mem[25][0] ;
 wire \Inst_RegFile_32x4.mem[25][1] ;
 wire \Inst_RegFile_32x4.mem[25][2] ;
 wire \Inst_RegFile_32x4.mem[25][3] ;
 wire \Inst_RegFile_32x4.mem[26][0] ;
 wire \Inst_RegFile_32x4.mem[26][1] ;
 wire \Inst_RegFile_32x4.mem[26][2] ;
 wire \Inst_RegFile_32x4.mem[26][3] ;
 wire \Inst_RegFile_32x4.mem[27][0] ;
 wire \Inst_RegFile_32x4.mem[27][1] ;
 wire \Inst_RegFile_32x4.mem[27][2] ;
 wire \Inst_RegFile_32x4.mem[27][3] ;
 wire \Inst_RegFile_32x4.mem[28][0] ;
 wire \Inst_RegFile_32x4.mem[28][1] ;
 wire \Inst_RegFile_32x4.mem[28][2] ;
 wire \Inst_RegFile_32x4.mem[28][3] ;
 wire \Inst_RegFile_32x4.mem[29][0] ;
 wire \Inst_RegFile_32x4.mem[29][1] ;
 wire \Inst_RegFile_32x4.mem[29][2] ;
 wire \Inst_RegFile_32x4.mem[29][3] ;
 wire \Inst_RegFile_32x4.mem[2][0] ;
 wire \Inst_RegFile_32x4.mem[2][1] ;
 wire \Inst_RegFile_32x4.mem[2][2] ;
 wire \Inst_RegFile_32x4.mem[2][3] ;
 wire \Inst_RegFile_32x4.mem[30][0] ;
 wire \Inst_RegFile_32x4.mem[30][1] ;
 wire \Inst_RegFile_32x4.mem[30][2] ;
 wire \Inst_RegFile_32x4.mem[30][3] ;
 wire \Inst_RegFile_32x4.mem[31][0] ;
 wire \Inst_RegFile_32x4.mem[31][1] ;
 wire \Inst_RegFile_32x4.mem[31][2] ;
 wire \Inst_RegFile_32x4.mem[31][3] ;
 wire \Inst_RegFile_32x4.mem[3][0] ;
 wire \Inst_RegFile_32x4.mem[3][1] ;
 wire \Inst_RegFile_32x4.mem[3][2] ;
 wire \Inst_RegFile_32x4.mem[3][3] ;
 wire \Inst_RegFile_32x4.mem[4][0] ;
 wire \Inst_RegFile_32x4.mem[4][1] ;
 wire \Inst_RegFile_32x4.mem[4][2] ;
 wire \Inst_RegFile_32x4.mem[4][3] ;
 wire \Inst_RegFile_32x4.mem[5][0] ;
 wire \Inst_RegFile_32x4.mem[5][1] ;
 wire \Inst_RegFile_32x4.mem[5][2] ;
 wire \Inst_RegFile_32x4.mem[5][3] ;
 wire \Inst_RegFile_32x4.mem[6][0] ;
 wire \Inst_RegFile_32x4.mem[6][1] ;
 wire \Inst_RegFile_32x4.mem[6][2] ;
 wire \Inst_RegFile_32x4.mem[6][3] ;
 wire \Inst_RegFile_32x4.mem[7][0] ;
 wire \Inst_RegFile_32x4.mem[7][1] ;
 wire \Inst_RegFile_32x4.mem[7][2] ;
 wire \Inst_RegFile_32x4.mem[7][3] ;
 wire \Inst_RegFile_32x4.mem[8][0] ;
 wire \Inst_RegFile_32x4.mem[8][1] ;
 wire \Inst_RegFile_32x4.mem[8][2] ;
 wire \Inst_RegFile_32x4.mem[8][3] ;
 wire \Inst_RegFile_32x4.mem[9][0] ;
 wire \Inst_RegFile_32x4.mem[9][1] ;
 wire \Inst_RegFile_32x4.mem[9][2] ;
 wire \Inst_RegFile_32x4.mem[9][3] ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame10_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame11_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame12_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame5_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame6_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame7_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame8_bit9.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit0.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit1.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit10.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit11.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit14.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit15.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit18.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit19.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit2.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit20.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit21.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit22.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit23.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit24.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit25.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit27.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit29.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit3.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit30.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit4.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit5.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit7.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit8.Q ;
 wire \Inst_RegFile_ConfigMem.Inst_frame9_bit9.Q ;
 wire \Inst_RegFile_switch_matrix.E1BEG0 ;
 wire \Inst_RegFile_switch_matrix.E1BEG1 ;
 wire \Inst_RegFile_switch_matrix.E1BEG2 ;
 wire \Inst_RegFile_switch_matrix.E1BEG3 ;
 wire \Inst_RegFile_switch_matrix.E2BEG0 ;
 wire \Inst_RegFile_switch_matrix.E2BEG1 ;
 wire \Inst_RegFile_switch_matrix.E2BEG2 ;
 wire \Inst_RegFile_switch_matrix.E2BEG3 ;
 wire \Inst_RegFile_switch_matrix.E2BEG4 ;
 wire \Inst_RegFile_switch_matrix.E2BEG5 ;
 wire \Inst_RegFile_switch_matrix.E2BEG6 ;
 wire \Inst_RegFile_switch_matrix.E2BEG7 ;
 wire \Inst_RegFile_switch_matrix.E6BEG0 ;
 wire \Inst_RegFile_switch_matrix.E6BEG1 ;
 wire \Inst_RegFile_switch_matrix.EE4BEG0 ;
 wire \Inst_RegFile_switch_matrix.EE4BEG1 ;
 wire \Inst_RegFile_switch_matrix.EE4BEG2 ;
 wire \Inst_RegFile_switch_matrix.EE4BEG3 ;
 wire \Inst_RegFile_switch_matrix.JN2BEG0 ;
 wire \Inst_RegFile_switch_matrix.JN2BEG1 ;
 wire \Inst_RegFile_switch_matrix.JN2BEG2 ;
 wire \Inst_RegFile_switch_matrix.JN2BEG3 ;
 wire \Inst_RegFile_switch_matrix.JN2BEG4 ;
 wire \Inst_RegFile_switch_matrix.JN2BEG5 ;
 wire \Inst_RegFile_switch_matrix.JN2BEG6 ;
 wire \Inst_RegFile_switch_matrix.JN2BEG7 ;
 wire \Inst_RegFile_switch_matrix.JS2BEG0 ;
 wire \Inst_RegFile_switch_matrix.JS2BEG1 ;
 wire \Inst_RegFile_switch_matrix.JS2BEG2 ;
 wire \Inst_RegFile_switch_matrix.JS2BEG3 ;
 wire \Inst_RegFile_switch_matrix.JS2BEG4 ;
 wire \Inst_RegFile_switch_matrix.JS2BEG5 ;
 wire \Inst_RegFile_switch_matrix.JS2BEG6 ;
 wire \Inst_RegFile_switch_matrix.JS2BEG7 ;
 wire \Inst_RegFile_switch_matrix.JW2BEG0 ;
 wire \Inst_RegFile_switch_matrix.JW2BEG1 ;
 wire \Inst_RegFile_switch_matrix.JW2BEG2 ;
 wire \Inst_RegFile_switch_matrix.JW2BEG3 ;
 wire \Inst_RegFile_switch_matrix.JW2BEG4 ;
 wire \Inst_RegFile_switch_matrix.JW2BEG5 ;
 wire \Inst_RegFile_switch_matrix.JW2BEG6 ;
 wire \Inst_RegFile_switch_matrix.JW2BEG7 ;
 wire \Inst_RegFile_switch_matrix.N1BEG0 ;
 wire \Inst_RegFile_switch_matrix.N1BEG1 ;
 wire \Inst_RegFile_switch_matrix.N1BEG2 ;
 wire \Inst_RegFile_switch_matrix.N1BEG3 ;
 wire \Inst_RegFile_switch_matrix.N4BEG0 ;
 wire \Inst_RegFile_switch_matrix.N4BEG1 ;
 wire \Inst_RegFile_switch_matrix.N4BEG2 ;
 wire \Inst_RegFile_switch_matrix.N4BEG3 ;
 wire \Inst_RegFile_switch_matrix.NN4BEG0 ;
 wire \Inst_RegFile_switch_matrix.NN4BEG1 ;
 wire \Inst_RegFile_switch_matrix.NN4BEG2 ;
 wire \Inst_RegFile_switch_matrix.NN4BEG3 ;
 wire \Inst_RegFile_switch_matrix.S1BEG0 ;
 wire \Inst_RegFile_switch_matrix.S1BEG1 ;
 wire \Inst_RegFile_switch_matrix.S1BEG2 ;
 wire \Inst_RegFile_switch_matrix.S1BEG3 ;
 wire \Inst_RegFile_switch_matrix.S4BEG0 ;
 wire \Inst_RegFile_switch_matrix.S4BEG1 ;
 wire \Inst_RegFile_switch_matrix.S4BEG2 ;
 wire \Inst_RegFile_switch_matrix.S4BEG3 ;
 wire \Inst_RegFile_switch_matrix.SS4BEG0 ;
 wire \Inst_RegFile_switch_matrix.SS4BEG1 ;
 wire \Inst_RegFile_switch_matrix.SS4BEG2 ;
 wire \Inst_RegFile_switch_matrix.SS4BEG3 ;
 wire \Inst_RegFile_switch_matrix.W1BEG0 ;
 wire \Inst_RegFile_switch_matrix.W1BEG1 ;
 wire \Inst_RegFile_switch_matrix.W1BEG2 ;
 wire \Inst_RegFile_switch_matrix.W1BEG3 ;
 wire \Inst_RegFile_switch_matrix.W6BEG0 ;
 wire \Inst_RegFile_switch_matrix.W6BEG1 ;
 wire \Inst_RegFile_switch_matrix.WW4BEG0 ;
 wire \Inst_RegFile_switch_matrix.WW4BEG1 ;
 wire \Inst_RegFile_switch_matrix.WW4BEG2 ;
 wire \Inst_RegFile_switch_matrix.WW4BEG3 ;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire UserCLK_regs;
 wire clknet_0_UserCLK;
 wire clknet_1_0__leaf_UserCLK;
 wire clknet_0_UserCLK_regs;
 wire clknet_4_0_0_UserCLK_regs;
 wire clknet_4_1_0_UserCLK_regs;
 wire clknet_4_2_0_UserCLK_regs;
 wire clknet_4_3_0_UserCLK_regs;
 wire clknet_4_4_0_UserCLK_regs;
 wire clknet_4_5_0_UserCLK_regs;
 wire clknet_4_6_0_UserCLK_regs;
 wire clknet_4_7_0_UserCLK_regs;
 wire clknet_4_8_0_UserCLK_regs;
 wire clknet_4_9_0_UserCLK_regs;
 wire clknet_4_10_0_UserCLK_regs;
 wire clknet_4_11_0_UserCLK_regs;
 wire clknet_4_12_0_UserCLK_regs;
 wire clknet_4_13_0_UserCLK_regs;
 wire clknet_4_14_0_UserCLK_regs;
 wire clknet_4_15_0_UserCLK_regs;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1356_ (.I(E2MID[6]),
    .ZN(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1357_ (.I(S2MID[7]),
    .ZN(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1358_ (.I(\Inst_RegFile_ConfigMem.Inst_frame8_bit21.Q ),
    .ZN(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1359_ (.I(WW4END[0]),
    .ZN(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1360_ (.I(EE4END[0]),
    .ZN(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1361_ (.I(\Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q ),
    .ZN(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1362_ (.I(\Inst_RegFile_32x4.mem[1][0] ),
    .ZN(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1363_ (.I(S2MID[2]),
    .ZN(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1364_ (.I(EE4END[1]),
    .ZN(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1365_ (.I(\Inst_RegFile_ConfigMem.Inst_frame3_bit26.Q ),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1366_ (.I(\Inst_RegFile_ConfigMem.Inst_frame3_bit27.Q ),
    .ZN(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1367_ (.I(\Inst_RegFile_ConfigMem.Inst_frame7_bit27.Q ),
    .ZN(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1368_ (.I(S2MID[3]),
    .ZN(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1369_ (.I(\Inst_RegFile_ConfigMem.Inst_frame8_bit23.Q ),
    .ZN(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1370_ (.I(SS4END[2]),
    .ZN(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1371_ (.I(\Inst_RegFile_ConfigMem.Inst_frame3_bit18.Q ),
    .ZN(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1372_ (.I(\Inst_RegFile_ConfigMem.Inst_frame3_bit19.Q ),
    .ZN(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1373_ (.I(\Inst_RegFile_32x4.mem[2][0] ),
    .ZN(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1374_ (.I(\Inst_RegFile_ConfigMem.Inst_frame8_bit25.Q ),
    .ZN(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1375_ (.I(\Inst_RegFile_ConfigMem.Inst_frame2_bit26.Q ),
    .ZN(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1376_ (.I(W2MID[4]),
    .ZN(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1377_ (.I(WW4END[3]),
    .ZN(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1378_ (.I(SS4END[3]),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1379_ (.I(\Inst_RegFile_ConfigMem.Inst_frame2_bit18.Q ),
    .ZN(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1380_ (.I(\Inst_RegFile_ConfigMem.Inst_frame8_bit26.Q ),
    .ZN(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1381_ (.I(\Inst_RegFile_32x4.mem[6][0] ),
    .ZN(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1382_ (.I(\Inst_RegFile_ConfigMem.Inst_frame8_bit27.Q ),
    .ZN(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1383_ (.I(E2MID[0]),
    .ZN(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1384_ (.I(\Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q ),
    .ZN(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1385_ (.I(WW4END[1]),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1386_ (.I(\Inst_RegFile_ConfigMem.Inst_frame1_bit27.Q ),
    .ZN(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1387_ (.I(S2MID[1]),
    .ZN(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1388_ (.I(S2END[1]),
    .ZN(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1389_ (.I(E6END[0]),
    .ZN(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1390_ (.I(\Inst_RegFile_ConfigMem.Inst_frame1_bit18.Q ),
    .ZN(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1391_ (.I(\Inst_RegFile_ConfigMem.Inst_frame8_bit28.Q ),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1392_ (.I(\Inst_RegFile_32x4.mem[9][0] ),
    .ZN(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1393_ (.I(\Inst_RegFile_32x4.mem[11][0] ),
    .ZN(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1394_ (.I(\Inst_RegFile_32x4.mem[13][0] ),
    .ZN(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1395_ (.I(\Inst_RegFile_32x4.mem[15][0] ),
    .ZN(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1396_ (.I(\Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q ),
    .ZN(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1397_ (.I(W2END[4]),
    .ZN(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1398_ (.I(\Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q ),
    .ZN(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1399_ (.I(W6END[0]),
    .ZN(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1400_ (.I(\Inst_RegFile_ConfigMem.Inst_frame3_bit15.Q ),
    .ZN(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1401_ (.I(\Inst_RegFile_32x4.mem[17][0] ),
    .ZN(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1402_ (.I(\Inst_RegFile_32x4.mem[18][0] ),
    .ZN(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1403_ (.I(\Inst_RegFile_32x4.mem[21][0] ),
    .ZN(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1404_ (.I(\Inst_RegFile_32x4.mem[22][0] ),
    .ZN(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1405_ (.I(\Inst_RegFile_32x4.mem[25][0] ),
    .ZN(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1406_ (.I(\Inst_RegFile_32x4.mem[27][0] ),
    .ZN(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1407_ (.I(\Inst_RegFile_32x4.mem[29][0] ),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1408_ (.I(\Inst_RegFile_32x4.mem[31][0] ),
    .ZN(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1409_ (.I(\Inst_RegFile_32x4.mem[2][1] ),
    .ZN(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1410_ (.I(\Inst_RegFile_32x4.mem[5][1] ),
    .ZN(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1411_ (.I(\Inst_RegFile_32x4.mem[6][1] ),
    .ZN(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1412_ (.I(\Inst_RegFile_32x4.mem[13][1] ),
    .ZN(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1413_ (.I(\Inst_RegFile_32x4.mem[16][1] ),
    .ZN(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1414_ (.I(\Inst_RegFile_32x4.mem[18][1] ),
    .ZN(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1415_ (.I(\Inst_RegFile_32x4.mem[21][1] ),
    .ZN(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1416_ (.I(\Inst_RegFile_32x4.mem[24][1] ),
    .ZN(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1417_ (.I(\Inst_RegFile_32x4.mem[26][1] ),
    .ZN(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1418_ (.I(\Inst_RegFile_32x4.mem[28][1] ),
    .ZN(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1419_ (.I(\Inst_RegFile_32x4.mem[31][1] ),
    .ZN(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1420_ (.I(\Inst_RegFile_32x4.mem[1][2] ),
    .ZN(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1421_ (.I(\Inst_RegFile_32x4.mem[2][2] ),
    .ZN(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1422_ (.I(\Inst_RegFile_32x4.mem[6][2] ),
    .ZN(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1423_ (.I(\Inst_RegFile_32x4.mem[9][2] ),
    .ZN(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1424_ (.I(\Inst_RegFile_32x4.mem[11][2] ),
    .ZN(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1425_ (.I(\Inst_RegFile_32x4.mem[13][2] ),
    .ZN(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1426_ (.I(\Inst_RegFile_32x4.mem[15][2] ),
    .ZN(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1427_ (.I(\Inst_RegFile_32x4.mem[17][2] ),
    .ZN(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1428_ (.I(\Inst_RegFile_32x4.mem[18][2] ),
    .ZN(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1429_ (.I(\Inst_RegFile_32x4.mem[21][2] ),
    .ZN(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1430_ (.I(\Inst_RegFile_32x4.mem[22][2] ),
    .ZN(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1431_ (.I(\Inst_RegFile_32x4.mem[25][2] ),
    .ZN(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1432_ (.I(\Inst_RegFile_32x4.mem[27][2] ),
    .ZN(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1433_ (.I(\Inst_RegFile_32x4.mem[29][2] ),
    .ZN(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1434_ (.I(\Inst_RegFile_32x4.mem[31][2] ),
    .ZN(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1435_ (.I(\Inst_RegFile_32x4.mem[2][3] ),
    .ZN(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1436_ (.I(\Inst_RegFile_32x4.mem[5][3] ),
    .ZN(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1437_ (.I(\Inst_RegFile_32x4.mem[6][3] ),
    .ZN(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1438_ (.I(\Inst_RegFile_32x4.mem[9][3] ),
    .ZN(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1439_ (.I(\Inst_RegFile_32x4.mem[11][3] ),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1440_ (.I(\Inst_RegFile_32x4.mem[13][3] ),
    .ZN(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1441_ (.I(\Inst_RegFile_32x4.mem[15][3] ),
    .ZN(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1442_ (.I(\Inst_RegFile_32x4.mem[17][3] ),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1443_ (.I(\Inst_RegFile_32x4.mem[18][3] ),
    .ZN(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1444_ (.I(\Inst_RegFile_32x4.mem[21][3] ),
    .ZN(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1445_ (.I(\Inst_RegFile_32x4.mem[22][3] ),
    .ZN(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1446_ (.I(\Inst_RegFile_32x4.mem[25][3] ),
    .ZN(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1447_ (.I(\Inst_RegFile_32x4.mem[27][3] ),
    .ZN(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1448_ (.I(\Inst_RegFile_32x4.mem[29][3] ),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1449_ (.I(\Inst_RegFile_32x4.mem[31][3] ),
    .ZN(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1450_ (.I(\Inst_RegFile_ConfigMem.Inst_frame4_bit22.Q ),
    .ZN(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1451_ (.I(W2END[7]),
    .ZN(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1452_ (.I(\Inst_RegFile_ConfigMem.Inst_frame3_bit22.Q ),
    .ZN(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1453_ (.I(E2END[2]),
    .ZN(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1454_ (.I(\Inst_RegFile_ConfigMem.Inst_frame8_bit14.Q ),
    .ZN(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1455_ (.I(\Inst_RegFile_ConfigMem.Inst_frame2_bit22.Q ),
    .ZN(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1456_ (.I(\Inst_RegFile_ConfigMem.Inst_frame2_bit14.Q ),
    .ZN(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1457_ (.I(\Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q ),
    .ZN(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1458_ (.I(\Inst_RegFile_ConfigMem.Inst_frame1_bit23.Q ),
    .ZN(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1459_ (.I(\Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q ),
    .ZN(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1460_ (.I(\Inst_RegFile_ConfigMem.Inst_frame1_bit14.Q ),
    .ZN(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1461_ (.I(\Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q ),
    .ZN(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1462_ (.I(S2END[0]),
    .ZN(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1463_ (.I(\Inst_RegFile_ConfigMem.Inst_frame1_bit10.Q ),
    .ZN(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1464_ (.I(\Inst_RegFile_ConfigMem.Inst_frame3_bit10.Q ),
    .ZN(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1465_ (.I(\Inst_RegFile_ConfigMem.Inst_frame4_bit10.Q ),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1466_ (.I(\Inst_RegFile_ConfigMem.Inst_frame4_bit11.Q ),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1467_ (.I(\Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q ),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1468_ (.I(\Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q ),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1469_ (.I(\Inst_RegFile_ConfigMem.Inst_frame3_bit6.Q ),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1470_ (.I(\Inst_RegFile_ConfigMem.Inst_frame1_bit30.Q ),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1471_ (.I(\Inst_RegFile_ConfigMem.Inst_frame2_bit2.Q ),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1472_ (.I(\Inst_RegFile_ConfigMem.Inst_frame3_bit2.Q ),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1473_ (.I(\Inst_RegFile_ConfigMem.Inst_frame9_bit18.Q ),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1474_ (.I(\Inst_RegFile_ConfigMem.Inst_frame11_bit26.Q ),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1475_ (.I(\Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q ),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1476_ (.I(\Inst_RegFile_ConfigMem.Inst_frame10_bit3.Q ),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1477_ (.I(\Inst_RegFile_ConfigMem.Inst_frame7_bit8.Q ),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1478_ (.I(\Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q ),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1479_ (.I(\Inst_RegFile_ConfigMem.Inst_frame8_bit0.Q ),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1480_ (.I(\Inst_RegFile_ConfigMem.Inst_frame0_bit12.Q ),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1481_ (.I(\Inst_RegFile_ConfigMem.Inst_frame8_bit2.Q ),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1482_ (.I(\Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q ),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1483_ (.I(\Inst_RegFile_ConfigMem.Inst_frame8_bit8.Q ),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1484_ (.I(A_ADR0),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1485_ (.I0(AD3),
    .I1(BD0),
    .I2(BD2),
    .I3(BD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q ),
    .Z(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1486_ (.A1(_1343_),
    .A2(_0148_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1487_ (.I0(W1END[2]),
    .I1(AD0),
    .I2(AD1),
    .I3(AD2),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q ),
    .Z(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1488_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit22.Q ),
    .A2(_0150_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame3_bit23.Q ),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1489_ (.I0(EE4END[2]),
    .I1(S1END[0]),
    .I2(S1END[2]),
    .I3(S2END[6]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q ),
    .Z(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1490_ (.A1(_1343_),
    .A2(_0152_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1491_ (.I0(N1END[2]),
    .I1(N2END[6]),
    .I2(E1END[2]),
    .I3(E2END[6]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q ),
    .Z(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1492_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit22.Q ),
    .A2(_0154_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1493_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit23.Q ),
    .A2(_0153_),
    .A3(_0155_),
    .B1(_0149_),
    .B2(_0151_),
    .ZN(\Inst_RegFile_switch_matrix.E2BEG5 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1494_ (.I0(N2MID[2]),
    .I1(S2MID[2]),
    .I2(E2MID[2]),
    .I3(\Inst_RegFile_switch_matrix.E2BEG5 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit19.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit18.Q ),
    .Z(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1495_ (.I0(N2MID[3]),
    .I1(E2MID[3]),
    .S(\Inst_RegFile_ConfigMem.Inst_frame6_bit18.Q ),
    .Z(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1496_ (.A1(W2MID[3]),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame6_bit18.Q ),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1497_ (.A1(_1259_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame6_bit18.Q ),
    .B(\Inst_RegFile_ConfigMem.Inst_frame6_bit19.Q ),
    .C(_0158_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1498_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame6_bit19.Q ),
    .A2(_0157_),
    .B(_0159_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1499_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit12.Q ),
    .A2(_0160_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame8_bit13.Q ),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1500_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit12.Q ),
    .A2(_0156_),
    .B(_0161_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1501_ (.I0(W6END[0]),
    .I1(AD0),
    .I2(AD1),
    .I3(AD2),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q ),
    .Z(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1502_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q ),
    .A2(_0163_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1503_ (.I0(BD0),
    .I1(BD2),
    .I2(BD1),
    .I3(BD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q ),
    .Z(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1504_ (.A1(_1289_),
    .A2(_0165_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame3_bit15.Q ),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1505_ (.I0(N1END[2]),
    .I1(N2END[4]),
    .I2(N4END[0]),
    .I3(E2END[4]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q ),
    .Z(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1506_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q ),
    .A2(_0167_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1507_ (.I0(E6END[0]),
    .I1(S2END[4]),
    .I2(SS4END[3]),
    .I3(W2END[4]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q ),
    .Z(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1508_ (.A1(_1289_),
    .A2(_0169_),
    .B(_1291_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1509_ (.A1(_0164_),
    .A2(_0166_),
    .B1(_0168_),
    .B2(_0170_),
    .ZN(\Inst_RegFile_switch_matrix.E2BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1510_ (.A1(_0164_),
    .A2(_0166_),
    .B1(_0168_),
    .B2(_0170_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q ),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1511_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q ),
    .A2(S4END[2]),
    .Z(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1512_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit19.Q ),
    .A2(_0171_),
    .A3(_0172_),
    .Z(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1513_ (.A1(_1344_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q ),
    .B(\Inst_RegFile_ConfigMem.Inst_frame0_bit19.Q ),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1514_ (.A1(NN4END[2]),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q ),
    .B(_0174_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1515_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit12.Q ),
    .A2(_0175_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1516_ (.I0(N2END[3]),
    .I1(E2END[3]),
    .I2(S2END[3]),
    .I3(WW4END[1]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit18.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit19.Q ),
    .Z(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1517_ (.I(_0177_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1518_ (.A1(_0173_),
    .A2(_0176_),
    .B1(_0177_),
    .B2(\Inst_RegFile_ConfigMem.Inst_frame8_bit12.Q ),
    .C(\Inst_RegFile_ConfigMem.Inst_frame8_bit13.Q ),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1519_ (.A1(_0162_),
    .A2(_0179_),
    .Z(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1520_ (.A1(_0162_),
    .A2(_0179_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1521_ (.A1(\Inst_RegFile_32x4.mem[26][0] ),
    .A2(_0147_),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1522_ (.A1(_1297_),
    .A2(_0147_),
    .B(_0181_),
    .C(_0182_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1523_ (.I0(W6END[0]),
    .I1(AD0),
    .I2(AD1),
    .I3(AD2),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q ),
    .Z(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1524_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit14.Q ),
    .A2(_0184_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1525_ (.I0(BD0),
    .I1(BD2),
    .I2(BD1),
    .I3(BD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q ),
    .Z(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1526_ (.A1(_1347_),
    .A2(_0186_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame2_bit15.Q ),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1527_ (.I0(E6END[0]),
    .I1(S2END[4]),
    .I2(S4END[0]),
    .I3(W2END[4]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q ),
    .Z(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1528_ (.A1(_1347_),
    .A2(_0188_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1529_ (.I0(N2END[4]),
    .I1(E2END[4]),
    .I2(E1END[2]),
    .I3(EE4END[3]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q ),
    .Z(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1530_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit14.Q ),
    .A2(_0190_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1531_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit15.Q ),
    .A2(_0189_),
    .A3(_0191_),
    .B1(_0185_),
    .B2(_0187_),
    .ZN(\Inst_RegFile_switch_matrix.JS2BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1532_ (.I0(N4END[1]),
    .I1(SS4END[1]),
    .S(\Inst_RegFile_ConfigMem.Inst_frame0_bit20.Q ),
    .Z(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1533_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit20.Q ),
    .A2(\Inst_RegFile_switch_matrix.JS2BEG3 ),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1534_ (.A1(_1288_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame0_bit20.Q ),
    .B(\Inst_RegFile_ConfigMem.Inst_frame0_bit21.Q ),
    .C(_0193_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1535_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit21.Q ),
    .A2(_0192_),
    .B(_0194_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1536_ (.I0(N4END[1]),
    .I1(W2END[4]),
    .I2(SS4END[1]),
    .I3(\Inst_RegFile_switch_matrix.JS2BEG3 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame0_bit21.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame0_bit20.Q ),
    .Z(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1537_ (.I0(N2END[5]),
    .I1(E2END[5]),
    .I2(SS4END[1]),
    .I3(W2END[5]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit21.Q ),
    .Z(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1538_ (.I(_0197_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1539_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit14.Q ),
    .A2(_0198_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame8_bit15.Q ),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1540_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit14.Q ),
    .A2(_0196_),
    .B(_0199_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1541_ (.I0(W1END[2]),
    .I1(AD0),
    .I2(AD1),
    .I3(AD2),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q ),
    .Z(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1542_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit22.Q ),
    .A2(_0201_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1543_ (.I0(AD3),
    .I1(BD0),
    .I2(BD2),
    .I3(BD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q ),
    .Z(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1544_ (.A1(_1346_),
    .A2(_0203_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame2_bit23.Q ),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1545_ (.I0(N1END[2]),
    .I1(N2END[6]),
    .I2(E1END[2]),
    .I3(E2END[6]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q ),
    .Z(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1546_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit22.Q ),
    .A2(_0205_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1547_ (.I0(S1END[2]),
    .I1(S2END[6]),
    .I2(SS4END[2]),
    .I3(W1END[0]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q ),
    .Z(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1548_ (.A1(_1346_),
    .A2(_0207_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1549_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit23.Q ),
    .A2(_0206_),
    .A3(_0208_),
    .B1(_0202_),
    .B2(_0204_),
    .ZN(\Inst_RegFile_switch_matrix.JS2BEG5 ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1550_ (.I0(N2MID[4]),
    .I1(S2MID[4]),
    .S(\Inst_RegFile_ConfigMem.Inst_frame7_bit20.Q ),
    .Z(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1551_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame7_bit20.Q ),
    .A2(\Inst_RegFile_switch_matrix.JS2BEG5 ),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1552_ (.A1(_1267_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame7_bit20.Q ),
    .B(\Inst_RegFile_ConfigMem.Inst_frame7_bit21.Q ),
    .C(_0210_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1553_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame7_bit21.Q ),
    .A2(_0209_),
    .B(_0211_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1554_ (.I0(N2MID[4]),
    .I1(W2MID[4]),
    .I2(S2MID[4]),
    .I3(\Inst_RegFile_switch_matrix.JS2BEG5 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit21.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit20.Q ),
    .Z(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1555_ (.I0(N2MID[5]),
    .I1(E2MID[5]),
    .I2(S2MID[5]),
    .I3(W2MID[5]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit21.Q ),
    .Z(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1556_ (.I(_0214_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1557_ (.A1(_1345_),
    .A2(_0215_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1558_ (.A1(_1345_),
    .A2(_0213_),
    .B(_0216_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame8_bit15.Q ),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1559_ (.A1(_0200_),
    .A2(_0217_),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1560_ (.A1(_0200_),
    .A2(_0217_),
    .Z(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1561_ (.A1(_1296_),
    .A2(A_ADR0),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1562_ (.A1(\Inst_RegFile_32x4.mem[24][0] ),
    .A2(A_ADR0),
    .B(_0220_),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1563_ (.A1(_0180_),
    .A2(_0221_),
    .B(_0218_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1564_ (.I0(W6END[0]),
    .I1(AD0),
    .I2(AD1),
    .I3(AD2),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q ),
    .Z(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1565_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit14.Q ),
    .A2(_0223_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1566_ (.I0(BD0),
    .I1(BD2),
    .I2(BD1),
    .I3(BD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q ),
    .Z(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1567_ (.A1(_1351_),
    .A2(_0225_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame1_bit15.Q ),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1568_ (.I0(N1END[2]),
    .I1(N2END[4]),
    .I2(NN4END[3]),
    .I3(E2END[4]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q ),
    .Z(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1569_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit14.Q ),
    .A2(_0227_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1570_ (.I0(E6END[0]),
    .I1(S2END[4]),
    .I2(S4END[0]),
    .I3(W2END[4]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q ),
    .Z(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1571_ (.A1(_1351_),
    .A2(_0229_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1572_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit15.Q ),
    .A2(_0228_),
    .A3(_0230_),
    .B1(_0224_),
    .B2(_0226_),
    .ZN(\Inst_RegFile_switch_matrix.JW2BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1573_ (.A1(_1276_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame0_bit22.Q ),
    .B(\Inst_RegFile_ConfigMem.Inst_frame0_bit23.Q ),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1574_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit22.Q ),
    .A2(\Inst_RegFile_switch_matrix.JW2BEG3 ),
    .B(_0231_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1575_ (.I0(EE4END[3]),
    .I1(S4END[0]),
    .S(\Inst_RegFile_ConfigMem.Inst_frame0_bit22.Q ),
    .Z(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1576_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit23.Q ),
    .A2(_0233_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q ),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1577_ (.I0(NN4END[2]),
    .I1(E2END[1]),
    .S(\Inst_RegFile_ConfigMem.Inst_frame5_bit22.Q ),
    .Z(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1578_ (.A1(W2END[1]),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame5_bit22.Q ),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1579_ (.A1(_1279_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame5_bit22.Q ),
    .B(\Inst_RegFile_ConfigMem.Inst_frame5_bit23.Q ),
    .C(_0236_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1580_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame5_bit23.Q ),
    .A2(_0235_),
    .B(_0237_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1581_ (.A1(_0232_),
    .A2(_0234_),
    .B1(_0238_),
    .B2(\Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q ),
    .C(\Inst_RegFile_ConfigMem.Inst_frame8_bit17.Q ),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1582_ (.I0(WW4END[2]),
    .I1(AD0),
    .I2(AD1),
    .I3(AD2),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q ),
    .Z(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1583_ (.A1(_1348_),
    .A2(_0240_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1584_ (.I0(AD3),
    .I1(BD0),
    .I2(BD2),
    .I3(BD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q ),
    .Z(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1585_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q ),
    .A2(_0242_),
    .B(_1349_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1586_ (.I0(N1END[2]),
    .I1(N2END[6]),
    .I2(E1END[2]),
    .I3(E2END[6]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q ),
    .Z(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1587_ (.I0(S1END[0]),
    .I1(S2END[6]),
    .I2(S1END[2]),
    .I3(W1END[2]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q ),
    .Z(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1588_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q ),
    .A2(_0245_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1589_ (.A1(_1348_),
    .A2(_0244_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame1_bit23.Q ),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1590_ (.A1(_0241_),
    .A2(_0243_),
    .B1(_0246_),
    .B2(_0247_),
    .ZN(\Inst_RegFile_switch_matrix.JW2BEG5 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1591_ (.I0(E2MID[0]),
    .I1(W2MID[0]),
    .I2(S2MID[0]),
    .I3(\Inst_RegFile_switch_matrix.JW2BEG5 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit23.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit22.Q ),
    .Z(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1592_ (.I0(N2MID[1]),
    .I1(E2MID[1]),
    .I2(S2MID[1]),
    .I3(W2MID[1]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit22.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit23.Q ),
    .Z(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1593_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q ),
    .A2(_0249_),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1594_ (.A1(_1350_),
    .A2(_0248_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame8_bit17.Q ),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1595_ (.A1(_0250_),
    .A2(_0251_),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1596_ (.A1(_0239_),
    .A2(_0252_),
    .Z(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1597_ (.A1(_0239_),
    .A2(_0252_),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1598_ (.A1(\Inst_RegFile_32x4.mem[28][0] ),
    .A2(_0147_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1599_ (.A1(_1298_),
    .A2(_0147_),
    .B(_0255_),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1600_ (.A1(\Inst_RegFile_32x4.mem[30][0] ),
    .A2(_0147_),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1601_ (.A1(_1299_),
    .A2(_0147_),
    .B(_0257_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1602_ (.I0(_0256_),
    .I1(_0258_),
    .S(_0181_),
    .Z(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1603_ (.A1(_0183_),
    .A2(_0222_),
    .B1(_0259_),
    .B2(_0218_),
    .C(_0254_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1604_ (.I0(W1END[2]),
    .I1(AD0),
    .I2(AD1),
    .I3(AD2),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q ),
    .Z(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1605_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit22.Q ),
    .A2(_0261_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1606_ (.I0(AD3),
    .I1(BD0),
    .I2(BD2),
    .I3(BD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q ),
    .Z(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1607_ (.A1(_1341_),
    .A2(_0263_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame4_bit23.Q ),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1608_ (.I0(E2END[6]),
    .I1(S1END[2]),
    .I2(S2END[6]),
    .I3(W1END[0]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q ),
    .Z(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1609_ (.A1(_1341_),
    .A2(_0265_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1610_ (.I0(N1END[2]),
    .I1(NN4END[2]),
    .I2(N2END[6]),
    .I3(E1END[2]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q ),
    .Z(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1611_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit22.Q ),
    .A2(_0267_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1612_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit23.Q ),
    .A2(_0266_),
    .A3(_0268_),
    .B1(_0262_),
    .B2(_0264_),
    .ZN(\Inst_RegFile_switch_matrix.JN2BEG5 ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1613_ (.A1(N2END[0]),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame5_bit14.Q ),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1614_ (.A1(_1255_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame5_bit14.Q ),
    .B(\Inst_RegFile_ConfigMem.Inst_frame5_bit15.Q ),
    .C(_0269_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1615_ (.I0(S2END[0]),
    .I1(W2END[0]),
    .S(\Inst_RegFile_ConfigMem.Inst_frame5_bit14.Q ),
    .Z(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1616_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame5_bit15.Q ),
    .A2(_0271_),
    .B(_0270_),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1617_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q ),
    .A2(_0272_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1618_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q ),
    .A2(\Inst_RegFile_switch_matrix.JN2BEG5 ),
    .B(_0273_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame8_bit19.Q ),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1619_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q ),
    .A2(\Inst_RegFile_switch_matrix.JW2BEG5 ),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1620_ (.A1(_1352_),
    .A2(\Inst_RegFile_switch_matrix.JS2BEG5 ),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1621_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit19.Q ),
    .A2(_0275_),
    .A3(_0276_),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1622_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit20.Q ),
    .A2(_0277_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1623_ (.I0(W1END[3]),
    .I1(AD0),
    .I2(AD1),
    .I3(AD2),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q ),
    .Z(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1624_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit26.Q ),
    .A2(_0279_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1625_ (.I0(AD3),
    .I1(BD0),
    .I2(BD1),
    .I3(BD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q ),
    .Z(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1626_ (.A1(_1256_),
    .A2(_0281_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame3_bit27.Q ),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1627_ (.I0(N1END[3]),
    .I1(N2END[7]),
    .I2(E1END[3]),
    .I3(E2END[7]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q ),
    .Z(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1628_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit26.Q ),
    .A2(_0283_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1629_ (.I0(EE4END[1]),
    .I1(S1END[1]),
    .I2(S1END[3]),
    .I3(S2END[7]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q ),
    .Z(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1630_ (.A1(_1256_),
    .A2(_0285_),
    .B(_1257_),
    .ZN(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1631_ (.A1(_0280_),
    .A2(_0282_),
    .B1(_0284_),
    .B2(_0286_),
    .ZN(\Inst_RegFile_switch_matrix.E2BEG6 ));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1632_ (.A1(_0280_),
    .A2(_0282_),
    .B1(_0284_),
    .B2(_0286_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame7_bit26.Q ),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1633_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame7_bit26.Q ),
    .A2(W2MID[2]),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1634_ (.A1(_1258_),
    .A2(_0288_),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1635_ (.A1(N2MID[2]),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame7_bit26.Q ),
    .ZN(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1636_ (.A1(_1254_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame7_bit26.Q ),
    .B(\Inst_RegFile_ConfigMem.Inst_frame7_bit27.Q ),
    .C(_0290_),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1637_ (.A1(_0287_),
    .A2(_0289_),
    .B(_0291_),
    .ZN(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1638_ (.I0(N2MID[5]),
    .I1(E2MID[5]),
    .I2(S2MID[5]),
    .I3(W2MID[5]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit29.Q ),
    .Z(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1639_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q ),
    .A2(_0293_),
    .Z(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1640_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q ),
    .A2(_0292_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame8_bit19.Q ),
    .ZN(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1641_ (.A1(N2END[1]),
    .A2(_1352_),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1642_ (.A1(S2END[1]),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q ),
    .B(\Inst_RegFile_ConfigMem.Inst_frame8_bit19.Q ),
    .ZN(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1643_ (.A1(_0296_),
    .A2(_0297_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame8_bit20.Q ),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1644_ (.A1(_0294_),
    .A2(_0295_),
    .B(_0298_),
    .ZN(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1645_ (.A1(_0274_),
    .A2(_0278_),
    .B(_0299_),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1646_ (.A1(_1293_),
    .A2(A_ADR0),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1647_ (.A1(\Inst_RegFile_32x4.mem[19][0] ),
    .A2(A_ADR0),
    .B1(_0162_),
    .B2(_0179_),
    .C(_0301_),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1648_ (.A1(_1292_),
    .A2(A_ADR0),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1649_ (.A1(\Inst_RegFile_32x4.mem[16][0] ),
    .A2(A_ADR0),
    .B(_0303_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1650_ (.A1(_0180_),
    .A2(_0304_),
    .B(_0302_),
    .C(_0218_),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1651_ (.A1(_1294_),
    .A2(A_ADR0),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1652_ (.A1(\Inst_RegFile_32x4.mem[20][0] ),
    .A2(A_ADR0),
    .B(_0306_),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1653_ (.A1(_1295_),
    .A2(A_ADR0),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1654_ (.A1(\Inst_RegFile_32x4.mem[23][0] ),
    .A2(A_ADR0),
    .B1(_0162_),
    .B2(_0179_),
    .C(_0308_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1655_ (.A1(_0180_),
    .A2(_0307_),
    .B(_0309_),
    .C(_0219_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1656_ (.A1(_0253_),
    .A2(_0305_),
    .A3(_0310_),
    .B(_0300_),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1657_ (.A1(\Inst_RegFile_32x4.mem[3][0] ),
    .A2(A_ADR0),
    .ZN(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1658_ (.A1(_1264_),
    .A2(A_ADR0),
    .B(_0181_),
    .C(_0312_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1659_ (.A1(_1253_),
    .A2(A_ADR0),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1660_ (.A1(\Inst_RegFile_32x4.mem[0][0] ),
    .A2(A_ADR0),
    .B(_0314_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1661_ (.A1(_0180_),
    .A2(_0315_),
    .B(_0218_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1662_ (.I0(\Inst_RegFile_32x4.mem[4][0] ),
    .I1(\Inst_RegFile_32x4.mem[5][0] ),
    .S(A_ADR0),
    .Z(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1663_ (.A1(\Inst_RegFile_32x4.mem[7][0] ),
    .A2(A_ADR0),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1664_ (.A1(_1272_),
    .A2(A_ADR0),
    .B(_0318_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1665_ (.I0(_0317_),
    .I1(_0319_),
    .S(_0181_),
    .Z(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1666_ (.A1(_0313_),
    .A2(_0316_),
    .B1(_0320_),
    .B2(_0218_),
    .C(_0253_),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1667_ (.A1(\Inst_RegFile_32x4.mem[10][0] ),
    .A2(_0147_),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1668_ (.A1(_1284_),
    .A2(_0147_),
    .B(_0181_),
    .C(_0322_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1669_ (.A1(_1283_),
    .A2(A_ADR0),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1670_ (.A1(\Inst_RegFile_32x4.mem[8][0] ),
    .A2(A_ADR0),
    .B(_0324_),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1671_ (.A1(_0180_),
    .A2(_0325_),
    .B(_0218_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1672_ (.A1(\Inst_RegFile_32x4.mem[12][0] ),
    .A2(_0147_),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1673_ (.A1(_1285_),
    .A2(_0147_),
    .B(_0327_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1674_ (.A1(\Inst_RegFile_32x4.mem[14][0] ),
    .A2(_0147_),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1675_ (.A1(_1286_),
    .A2(_0147_),
    .B(_0329_),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1676_ (.I0(_0328_),
    .I1(_0330_),
    .S(_0181_),
    .Z(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1677_ (.A1(_0323_),
    .A2(_0326_),
    .B1(_0331_),
    .B2(_0218_),
    .C(_0254_),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1678_ (.A1(_0300_),
    .A2(_0321_),
    .A3(_0332_),
    .B1(_0311_),
    .B2(_0260_),
    .ZN(\Inst_RegFile_32x4.AD_comb[0] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1679_ (.I0(\Inst_RegFile_32x4.AD_comb[0] ),
    .I1(\Inst_RegFile_32x4.AD_reg[0] ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q ),
    .Z(AD0));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1680_ (.A1(\Inst_RegFile_32x4.mem[8][1] ),
    .A2(A_ADR0),
    .Z(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1681_ (.A1(\Inst_RegFile_32x4.mem[9][1] ),
    .A2(_0147_),
    .B(_0333_),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1682_ (.A1(\Inst_RegFile_32x4.mem[10][1] ),
    .A2(_0147_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1683_ (.A1(\Inst_RegFile_32x4.mem[11][1] ),
    .A2(A_ADR0),
    .B1(_0162_),
    .B2(_0179_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1684_ (.A1(_0180_),
    .A2(_0334_),
    .B1(_0335_),
    .B2(_0336_),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1685_ (.A1(\Inst_RegFile_32x4.mem[14][1] ),
    .A2(_0147_),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1686_ (.A1(\Inst_RegFile_32x4.mem[15][1] ),
    .A2(A_ADR0),
    .B1(_0162_),
    .B2(_0179_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1687_ (.A1(_1303_),
    .A2(A_ADR0),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1688_ (.A1(\Inst_RegFile_32x4.mem[12][1] ),
    .A2(A_ADR0),
    .B(_0340_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1689_ (.A1(_0338_),
    .A2(_0339_),
    .B1(_0341_),
    .B2(_0180_),
    .C(_0219_),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1690_ (.A1(_0219_),
    .A2(_0337_),
    .B(_0342_),
    .C(_0254_),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1691_ (.A1(\Inst_RegFile_32x4.mem[3][1] ),
    .A2(A_ADR0),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1692_ (.A1(_1300_),
    .A2(A_ADR0),
    .B(_0344_),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1693_ (.I0(\Inst_RegFile_32x4.mem[0][1] ),
    .I1(\Inst_RegFile_32x4.mem[1][1] ),
    .S(A_ADR0),
    .Z(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1694_ (.I0(_0345_),
    .I1(_0346_),
    .S(_0180_),
    .Z(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1695_ (.A1(\Inst_RegFile_32x4.mem[6][1] ),
    .A2(_0147_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1696_ (.A1(\Inst_RegFile_32x4.mem[7][1] ),
    .A2(A_ADR0),
    .B1(_0162_),
    .B2(_0179_),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1697_ (.A1(_1301_),
    .A2(A_ADR0),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1698_ (.A1(\Inst_RegFile_32x4.mem[4][1] ),
    .A2(A_ADR0),
    .B(_0350_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1699_ (.A1(_0348_),
    .A2(_0349_),
    .B1(_0351_),
    .B2(_0180_),
    .C(_0219_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1700_ (.A1(_0219_),
    .A2(_0347_),
    .B(_0352_),
    .C(_0253_),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1701_ (.A1(\Inst_RegFile_32x4.mem[27][1] ),
    .A2(A_ADR0),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1702_ (.A1(_1308_),
    .A2(A_ADR0),
    .B(_0181_),
    .C(_0354_),
    .ZN(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1703_ (.A1(_1307_),
    .A2(A_ADR0),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1704_ (.A1(\Inst_RegFile_32x4.mem[25][1] ),
    .A2(A_ADR0),
    .B(_0356_),
    .ZN(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1705_ (.A1(_0180_),
    .A2(_0357_),
    .B(_0218_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1706_ (.A1(\Inst_RegFile_32x4.mem[29][1] ),
    .A2(A_ADR0),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1707_ (.A1(_1309_),
    .A2(A_ADR0),
    .B(_0359_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1708_ (.A1(\Inst_RegFile_32x4.mem[30][1] ),
    .A2(_0147_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1709_ (.A1(_1310_),
    .A2(_0147_),
    .B(_0361_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1710_ (.I0(_0360_),
    .I1(_0362_),
    .S(_0181_),
    .Z(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1711_ (.A1(_0355_),
    .A2(_0358_),
    .B1(_0363_),
    .B2(_0218_),
    .C(_0254_),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1712_ (.A1(_1305_),
    .A2(A_ADR0),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1713_ (.A1(\Inst_RegFile_32x4.mem[19][1] ),
    .A2(A_ADR0),
    .B1(_0162_),
    .B2(_0179_),
    .C(_0365_),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1714_ (.A1(_1304_),
    .A2(A_ADR0),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1715_ (.A1(\Inst_RegFile_32x4.mem[17][1] ),
    .A2(A_ADR0),
    .B(_0367_),
    .ZN(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1716_ (.A1(_0180_),
    .A2(_0368_),
    .B(_0366_),
    .C(_0218_),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1717_ (.A1(_1306_),
    .A2(A_ADR0),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1718_ (.A1(\Inst_RegFile_32x4.mem[20][1] ),
    .A2(A_ADR0),
    .B(_0370_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1719_ (.A1(\Inst_RegFile_32x4.mem[23][1] ),
    .A2(A_ADR0),
    .Z(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1720_ (.A1(\Inst_RegFile_32x4.mem[22][1] ),
    .A2(_0147_),
    .B1(_0162_),
    .B2(_0179_),
    .C(_0372_),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1721_ (.A1(_0180_),
    .A2(_0371_),
    .B(_0373_),
    .C(_0219_),
    .ZN(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1722_ (.A1(_0253_),
    .A2(_0369_),
    .A3(_0374_),
    .B(_0300_),
    .ZN(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1723_ (.A1(_0300_),
    .A2(_0343_),
    .A3(_0353_),
    .B1(_0364_),
    .B2(_0375_),
    .ZN(\Inst_RegFile_32x4.AD_comb[1] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1724_ (.I0(\Inst_RegFile_32x4.AD_comb[1] ),
    .I1(\Inst_RegFile_32x4.AD_reg[1] ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q ),
    .Z(AD1));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1725_ (.A1(\Inst_RegFile_32x4.mem[10][2] ),
    .A2(_0147_),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1726_ (.A1(_1315_),
    .A2(_0147_),
    .B(_0376_),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1727_ (.A1(\Inst_RegFile_32x4.mem[9][2] ),
    .A2(A_ADR0),
    .ZN(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1728_ (.A1(\Inst_RegFile_32x4.mem[8][2] ),
    .A2(_0147_),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1729_ (.A1(_0162_),
    .A2(_0179_),
    .A3(_0378_),
    .A4(_0379_),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1730_ (.A1(_0180_),
    .A2(_0377_),
    .B(_0380_),
    .C(_0219_),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1731_ (.A1(\Inst_RegFile_32x4.mem[14][2] ),
    .A2(_0147_),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1732_ (.A1(_1317_),
    .A2(_0147_),
    .B(_0382_),
    .ZN(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1733_ (.A1(\Inst_RegFile_32x4.mem[13][2] ),
    .A2(A_ADR0),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1734_ (.A1(\Inst_RegFile_32x4.mem[12][2] ),
    .A2(_0147_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1735_ (.A1(_0162_),
    .A2(_0179_),
    .A3(_0384_),
    .A4(_0385_),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1736_ (.A1(_0180_),
    .A2(_0383_),
    .B(_0386_),
    .C(_0218_),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1737_ (.A1(_0253_),
    .A2(_0381_),
    .A3(_0387_),
    .Z(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1738_ (.A1(\Inst_RegFile_32x4.mem[3][2] ),
    .A2(A_ADR0),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1739_ (.A1(_1312_),
    .A2(A_ADR0),
    .B(_0181_),
    .C(_0389_),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1740_ (.A1(_1311_),
    .A2(A_ADR0),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1741_ (.A1(\Inst_RegFile_32x4.mem[0][2] ),
    .A2(A_ADR0),
    .B(_0391_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1742_ (.A1(_0180_),
    .A2(_0392_),
    .B(_0218_),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1743_ (.I0(\Inst_RegFile_32x4.mem[4][2] ),
    .I1(\Inst_RegFile_32x4.mem[5][2] ),
    .S(A_ADR0),
    .Z(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1744_ (.A1(\Inst_RegFile_32x4.mem[7][2] ),
    .A2(A_ADR0),
    .ZN(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1745_ (.A1(_1313_),
    .A2(A_ADR0),
    .B(_0395_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1746_ (.I0(_0394_),
    .I1(_0396_),
    .S(_0181_),
    .Z(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1747_ (.A1(_0390_),
    .A2(_0393_),
    .B1(_0397_),
    .B2(_0218_),
    .C(_0253_),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1748_ (.A1(\Inst_RegFile_32x4.mem[26][2] ),
    .A2(_0147_),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1749_ (.A1(_1323_),
    .A2(_0147_),
    .B(_0399_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1750_ (.A1(\Inst_RegFile_32x4.mem[25][2] ),
    .A2(A_ADR0),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1751_ (.A1(\Inst_RegFile_32x4.mem[24][2] ),
    .A2(_0147_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1752_ (.A1(_0162_),
    .A2(_0179_),
    .A3(_0401_),
    .A4(_0402_),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1753_ (.A1(_0180_),
    .A2(_0400_),
    .B(_0403_),
    .C(_0219_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1754_ (.A1(\Inst_RegFile_32x4.mem[29][2] ),
    .A2(A_ADR0),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1755_ (.A1(\Inst_RegFile_32x4.mem[28][2] ),
    .A2(_0147_),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1756_ (.A1(_0162_),
    .A2(_0179_),
    .A3(_0405_),
    .A4(_0406_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1757_ (.A1(\Inst_RegFile_32x4.mem[30][2] ),
    .A2(_0147_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1758_ (.A1(_1325_),
    .A2(_0147_),
    .B(_0408_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1759_ (.A1(_0180_),
    .A2(_0409_),
    .B(_0407_),
    .C(_0218_),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1760_ (.A1(_0253_),
    .A2(_0404_),
    .A3(_0410_),
    .Z(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1761_ (.A1(_1319_),
    .A2(A_ADR0),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1762_ (.A1(\Inst_RegFile_32x4.mem[19][2] ),
    .A2(A_ADR0),
    .B1(_0162_),
    .B2(_0179_),
    .C(_0412_),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1763_ (.A1(_1318_),
    .A2(A_ADR0),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1764_ (.A1(\Inst_RegFile_32x4.mem[16][2] ),
    .A2(A_ADR0),
    .B(_0414_),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1765_ (.A1(_0180_),
    .A2(_0415_),
    .B(_0413_),
    .C(_0218_),
    .ZN(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1766_ (.A1(_1320_),
    .A2(A_ADR0),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1767_ (.A1(\Inst_RegFile_32x4.mem[20][2] ),
    .A2(A_ADR0),
    .B(_0417_),
    .ZN(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1768_ (.A1(_1321_),
    .A2(A_ADR0),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1769_ (.A1(\Inst_RegFile_32x4.mem[23][2] ),
    .A2(A_ADR0),
    .B1(_0162_),
    .B2(_0179_),
    .C(_0419_),
    .ZN(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1770_ (.A1(_0180_),
    .A2(_0418_),
    .B(_0420_),
    .C(_0219_),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1771_ (.A1(_0253_),
    .A2(_0416_),
    .A3(_0421_),
    .B(_0300_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1772_ (.A1(_0300_),
    .A2(_0388_),
    .A3(_0398_),
    .B1(_0411_),
    .B2(_0422_),
    .ZN(\Inst_RegFile_32x4.AD_comb[2] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1773_ (.I0(\Inst_RegFile_32x4.AD_comb[2] ),
    .I1(\Inst_RegFile_32x4.AD_reg[2] ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q ),
    .Z(AD2));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1774_ (.A1(\Inst_RegFile_32x4.mem[26][3] ),
    .A2(_0147_),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1775_ (.A1(_1338_),
    .A2(_0147_),
    .B(_0181_),
    .C(_0423_),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1776_ (.A1(_1337_),
    .A2(A_ADR0),
    .ZN(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1777_ (.A1(\Inst_RegFile_32x4.mem[24][3] ),
    .A2(A_ADR0),
    .B(_0425_),
    .ZN(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1778_ (.A1(_0180_),
    .A2(_0426_),
    .B(_0218_),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1779_ (.A1(\Inst_RegFile_32x4.mem[28][3] ),
    .A2(_0147_),
    .ZN(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1780_ (.A1(_1339_),
    .A2(_0147_),
    .B(_0428_),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1781_ (.A1(\Inst_RegFile_32x4.mem[30][3] ),
    .A2(_0147_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1782_ (.A1(_1340_),
    .A2(_0147_),
    .B(_0430_),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1783_ (.I0(_0429_),
    .I1(_0431_),
    .S(_0181_),
    .Z(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1784_ (.A1(_0424_),
    .A2(_0427_),
    .B1(_0432_),
    .B2(_0218_),
    .C(_0254_),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1785_ (.A1(_1334_),
    .A2(A_ADR0),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1786_ (.A1(\Inst_RegFile_32x4.mem[19][3] ),
    .A2(A_ADR0),
    .B1(_0162_),
    .B2(_0179_),
    .C(_0434_),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1787_ (.A1(_1333_),
    .A2(A_ADR0),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1788_ (.A1(\Inst_RegFile_32x4.mem[16][3] ),
    .A2(A_ADR0),
    .B(_0436_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1789_ (.A1(_0180_),
    .A2(_0437_),
    .B(_0435_),
    .C(_0218_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1790_ (.A1(_1335_),
    .A2(A_ADR0),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1791_ (.A1(\Inst_RegFile_32x4.mem[20][3] ),
    .A2(A_ADR0),
    .B(_0439_),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1792_ (.A1(_1336_),
    .A2(A_ADR0),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1793_ (.A1(\Inst_RegFile_32x4.mem[23][3] ),
    .A2(A_ADR0),
    .B1(_0162_),
    .B2(_0179_),
    .C(_0441_),
    .ZN(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1794_ (.A1(_0180_),
    .A2(_0440_),
    .B(_0442_),
    .C(_0219_),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1795_ (.A1(_0253_),
    .A2(_0438_),
    .A3(_0443_),
    .B(_0300_),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1796_ (.A1(_1330_),
    .A2(A_ADR0),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1797_ (.A1(\Inst_RegFile_32x4.mem[10][3] ),
    .A2(A_ADR0),
    .B(_0445_),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1798_ (.A1(\Inst_RegFile_32x4.mem[8][3] ),
    .A2(_0147_),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1799_ (.A1(_1329_),
    .A2(_0147_),
    .B(_0180_),
    .C(_0447_),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1800_ (.A1(_0181_),
    .A2(_0446_),
    .B(_0218_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1801_ (.A1(\Inst_RegFile_32x4.mem[14][3] ),
    .A2(_0147_),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1802_ (.A1(\Inst_RegFile_32x4.mem[15][3] ),
    .A2(A_ADR0),
    .B1(_0162_),
    .B2(_0179_),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1803_ (.A1(_1331_),
    .A2(A_ADR0),
    .ZN(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1804_ (.A1(\Inst_RegFile_32x4.mem[12][3] ),
    .A2(A_ADR0),
    .B(_0452_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1805_ (.A1(_0450_),
    .A2(_0451_),
    .B1(_0453_),
    .B2(_0180_),
    .C(_0219_),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1806_ (.A1(_0448_),
    .A2(_0449_),
    .B(_0454_),
    .C(_0254_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1807_ (.A1(\Inst_RegFile_32x4.mem[0][3] ),
    .A2(A_ADR0),
    .Z(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1808_ (.A1(\Inst_RegFile_32x4.mem[1][3] ),
    .A2(_0147_),
    .B(_0456_),
    .ZN(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1809_ (.A1(\Inst_RegFile_32x4.mem[2][3] ),
    .A2(_0147_),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1810_ (.A1(\Inst_RegFile_32x4.mem[3][3] ),
    .A2(A_ADR0),
    .B1(_0162_),
    .B2(_0179_),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1811_ (.A1(_0180_),
    .A2(_0457_),
    .B1(_0458_),
    .B2(_0459_),
    .C(_0218_),
    .ZN(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1812_ (.A1(\Inst_RegFile_32x4.mem[6][3] ),
    .A2(_0147_),
    .ZN(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1813_ (.A1(\Inst_RegFile_32x4.mem[7][3] ),
    .A2(A_ADR0),
    .B1(_0162_),
    .B2(_0179_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1814_ (.A1(_1327_),
    .A2(A_ADR0),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1815_ (.A1(\Inst_RegFile_32x4.mem[4][3] ),
    .A2(A_ADR0),
    .B(_0463_),
    .ZN(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1816_ (.A1(_0461_),
    .A2(_0462_),
    .B1(_0464_),
    .B2(_0180_),
    .C(_0219_),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1817_ (.A1(_0253_),
    .A2(_0460_),
    .A3(_0465_),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1818_ (.A1(_0300_),
    .A2(_0455_),
    .A3(_0466_),
    .B1(_0433_),
    .B2(_0444_),
    .ZN(\Inst_RegFile_32x4.AD_comb[3] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1819_ (.I0(\Inst_RegFile_32x4.AD_comb[3] ),
    .I1(\Inst_RegFile_32x4.AD_reg[3] ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q ),
    .Z(AD3));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1820_ (.A1(_0287_),
    .A2(_0289_),
    .B(_0291_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame8_bit23.Q ),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1821_ (.I0(N2MID[3]),
    .I1(E2MID[3]),
    .I2(S2MID[3]),
    .I3(W2MID[3]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit26.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit27.Q ),
    .Z(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1822_ (.A1(_1260_),
    .A2(_0468_),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1823_ (.I0(W1END[1]),
    .I1(AD0),
    .I2(AD1),
    .I3(AD2),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q ),
    .Z(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1824_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit18.Q ),
    .A2(_0470_),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1825_ (.I0(AD3),
    .I1(BD2),
    .I2(BD1),
    .I3(BD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q ),
    .Z(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1826_ (.A1(_1262_),
    .A2(_0472_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame3_bit19.Q ),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1827_ (.I0(N1END[1]),
    .I1(N2END[5]),
    .I2(E1END[1]),
    .I3(E2END[5]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q ),
    .Z(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1828_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit18.Q ),
    .A2(_0474_),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1829_ (.I0(EE4END[3]),
    .I1(S1END[1]),
    .I2(S1END[3]),
    .I3(S2END[5]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q ),
    .Z(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1830_ (.A1(_1262_),
    .A2(_0476_),
    .B(_1263_),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1831_ (.A1(_0471_),
    .A2(_0473_),
    .B1(_0475_),
    .B2(_0477_),
    .ZN(\Inst_RegFile_switch_matrix.E2BEG4 ));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1832_ (.A1(_0471_),
    .A2(_0473_),
    .B1(_0475_),
    .B2(_0477_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q ),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1833_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q ),
    .A2(W2END[2]),
    .B(\Inst_RegFile_ConfigMem.Inst_frame0_bit27.Q ),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1834_ (.I(_0479_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1835_ (.A1(N4END[2]),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q ),
    .ZN(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1836_ (.A1(_1261_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q ),
    .B(\Inst_RegFile_ConfigMem.Inst_frame0_bit27.Q ),
    .C(_0481_),
    .ZN(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1837_ (.A1(_0478_),
    .A2(_0480_),
    .B(_0482_),
    .C(_1260_),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1838_ (.I0(N2END[3]),
    .I1(E2END[3]),
    .I2(SS4END[0]),
    .I3(W2END[3]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit26.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit27.Q ),
    .Z(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1839_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit23.Q ),
    .A2(_0484_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame8_bit24.Q ),
    .ZN(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1840_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit24.Q ),
    .A2(_0467_),
    .A3(_0469_),
    .B1(_0483_),
    .B2(_0485_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1841_ (.A1(\Inst_RegFile_32x4.mem[19][0] ),
    .A2(B_ADR0),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1842_ (.A1(_1293_),
    .A2(B_ADR0),
    .B(_0486_),
    .C(_0487_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1843_ (.I0(W1END[3]),
    .I1(AD0),
    .I2(AD1),
    .I3(AD2),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q ),
    .Z(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1844_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit26.Q ),
    .A2(_0489_),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1845_ (.I0(AD3),
    .I1(BD0),
    .I2(BD1),
    .I3(BD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q ),
    .Z(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1846_ (.A1(_1266_),
    .A2(_0491_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame2_bit27.Q ),
    .ZN(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1847_ (.I0(N1END[3]),
    .I1(N2END[7]),
    .I2(E1END[3]),
    .I3(E2END[7]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q ),
    .Z(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1848_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit26.Q ),
    .A2(_0493_),
    .ZN(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1849_ (.I0(S1END[3]),
    .I1(S2END[7]),
    .I2(SS4END[1]),
    .I3(W1END[1]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q ),
    .Z(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1850_ (.A1(_1266_),
    .A2(_0495_),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1851_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit27.Q ),
    .A2(_0494_),
    .A3(_0496_),
    .B1(_0490_),
    .B2(_0492_),
    .ZN(\Inst_RegFile_switch_matrix.JS2BEG6 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1852_ (.I0(E2MID[4]),
    .I1(S2MID[4]),
    .I2(W2MID[4]),
    .I3(\Inst_RegFile_switch_matrix.JS2BEG6 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit29.Q ),
    .Z(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1853_ (.A1(_1265_),
    .A2(_0497_),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1854_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit25.Q ),
    .A2(_0293_),
    .Z(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1855_ (.A1(_1265_),
    .A2(_0497_),
    .B(_0499_),
    .ZN(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1856_ (.I0(W1END[3]),
    .I1(AD0),
    .I2(AD1),
    .I3(AD2),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q ),
    .Z(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1857_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit18.Q ),
    .A2(_0501_),
    .ZN(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1858_ (.I0(AD3),
    .I1(BD2),
    .I2(BD1),
    .I3(BD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q ),
    .Z(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1859_ (.A1(_1270_),
    .A2(_0503_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame2_bit19.Q ),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1860_ (.I0(N1END[1]),
    .I1(N2END[5]),
    .I2(E1END[1]),
    .I3(E2END[5]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q ),
    .Z(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1861_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit18.Q ),
    .A2(_0505_),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1862_ (.I0(S1END[1]),
    .I1(S2END[5]),
    .I2(SS4END[3]),
    .I3(W1END[1]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q ),
    .Z(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1863_ (.A1(_1270_),
    .A2(_0507_),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1864_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit19.Q ),
    .A2(_0506_),
    .A3(_0508_),
    .B1(_0502_),
    .B2(_0504_),
    .ZN(\Inst_RegFile_switch_matrix.JS2BEG4 ));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1865_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit28.Q ),
    .A2(_1268_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame0_bit29.Q ),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1866_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit28.Q ),
    .A2(\Inst_RegFile_switch_matrix.JS2BEG4 ),
    .B(_0509_),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1867_ (.I0(E6END[1]),
    .I1(S4END[1]),
    .S(\Inst_RegFile_ConfigMem.Inst_frame0_bit28.Q ),
    .Z(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1868_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit29.Q ),
    .A2(_0511_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame8_bit25.Q ),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1869_ (.A1(_0510_),
    .A2(_0512_),
    .Z(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1870_ (.I0(NN4END[1]),
    .I1(E2END[5]),
    .I2(S2END[5]),
    .I3(W2END[5]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit29.Q ),
    .Z(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1871_ (.A1(_1265_),
    .A2(_0514_),
    .B(_1271_),
    .ZN(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1872_ (.A1(_0510_),
    .A2(_0512_),
    .B(_0515_),
    .ZN(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1873_ (.A1(_1271_),
    .A2(_0500_),
    .B1(_0513_),
    .B2(_0515_),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1874_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit26.Q ),
    .A2(_0498_),
    .A3(_0499_),
    .B(_0516_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1875_ (.A1(\Inst_RegFile_32x4.mem[16][0] ),
    .A2(B_ADR0),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1876_ (.A1(_1292_),
    .A2(B_ADR0),
    .B(_0519_),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1877_ (.A1(_0486_),
    .A2(_0520_),
    .B(_0518_),
    .C(_0488_),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1878_ (.I0(WW4END[3]),
    .I1(AD0),
    .I2(AD1),
    .I3(AD2),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q ),
    .Z(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1879_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit18.Q ),
    .A2(_0522_),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1880_ (.I0(AD3),
    .I1(BD2),
    .I2(BD1),
    .I3(BD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q ),
    .Z(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1881_ (.A1(_1281_),
    .A2(_0524_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame1_bit19.Q ),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1882_ (.I0(N1END[1]),
    .I1(N2END[5]),
    .I2(E1END[1]),
    .I3(E2END[5]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q ),
    .Z(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1883_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit18.Q ),
    .A2(_0526_),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1884_ (.I0(S1END[1]),
    .I1(S2END[5]),
    .I2(S1END[3]),
    .I3(W1END[1]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q ),
    .Z(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1885_ (.A1(_1281_),
    .A2(_0528_),
    .ZN(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1886_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit19.Q ),
    .A2(_0527_),
    .A3(_0529_),
    .B1(_0523_),
    .B2(_0525_),
    .ZN(\Inst_RegFile_switch_matrix.JW2BEG4 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1887_ (.I0(NN4END[0]),
    .I1(E6END[0]),
    .I2(W2END[0]),
    .I3(\Inst_RegFile_switch_matrix.JW2BEG4 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame0_bit30.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame0_bit31.Q ),
    .Z(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1888_ (.I0(N2END[1]),
    .I1(S2END[1]),
    .I2(EE4END[3]),
    .I3(W2END[1]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit31.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit30.Q ),
    .Z(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1889_ (.I0(_0530_),
    .I1(_0531_),
    .S(_1273_),
    .Z(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1890_ (.A1(_1282_),
    .A2(_0532_),
    .Z(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1891_ (.I0(AD3),
    .I1(BD0),
    .I2(BD1),
    .I3(BD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q ),
    .Z(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1892_ (.I0(WW4END[1]),
    .I1(AD0),
    .I2(AD1),
    .I3(AD2),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q ),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1893_ (.A1(_1275_),
    .A2(_0535_),
    .ZN(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1894_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q ),
    .A2(_0534_),
    .B(_1277_),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1895_ (.I0(N1END[3]),
    .I1(N2END[7]),
    .I2(E1END[3]),
    .I3(E2END[7]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q ),
    .Z(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1896_ (.I0(S1END[1]),
    .I1(S2END[7]),
    .I2(S1END[3]),
    .I3(W1END[3]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q ),
    .Z(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1897_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q ),
    .A2(_0539_),
    .ZN(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1898_ (.A1(_1275_),
    .A2(_0538_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame1_bit27.Q ),
    .ZN(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1899_ (.A1(_0536_),
    .A2(_0537_),
    .B1(_0540_),
    .B2(_0541_),
    .ZN(\Inst_RegFile_switch_matrix.JW2BEG6 ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1900_ (.I0(W2MID[0]),
    .I1(\Inst_RegFile_switch_matrix.JW2BEG6 ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame7_bit30.Q ),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1901_ (.A1(N2MID[0]),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame7_bit30.Q ),
    .ZN(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1902_ (.A1(_1274_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame7_bit30.Q ),
    .B(\Inst_RegFile_ConfigMem.Inst_frame7_bit31.Q ),
    .C(_0543_),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1903_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame7_bit31.Q ),
    .A2(_0542_),
    .B(_0544_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame8_bit27.Q ),
    .ZN(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1904_ (.I0(N2MID[1]),
    .I1(E2MID[1]),
    .I2(S2MID[1]),
    .I3(W2MID[1]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit30.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit31.Q ),
    .Z(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1905_ (.A1(_1273_),
    .A2(_0546_),
    .ZN(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1906_ (.A1(_0545_),
    .A2(_0547_),
    .ZN(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1907_ (.I0(_0532_),
    .I1(_0548_),
    .S(_1282_),
    .Z(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1908_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit28.Q ),
    .A2(_0548_),
    .B(_0533_),
    .ZN(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1909_ (.A1(\Inst_RegFile_32x4.mem[23][0] ),
    .A2(B_ADR0),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1910_ (.A1(_1295_),
    .A2(B_ADR0),
    .B(_0486_),
    .C(_0551_),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1911_ (.A1(\Inst_RegFile_32x4.mem[20][0] ),
    .A2(B_ADR0),
    .ZN(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1912_ (.A1(_1294_),
    .A2(B_ADR0),
    .B(_0553_),
    .ZN(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1913_ (.A1(_0486_),
    .A2(_0554_),
    .B(_0552_),
    .C(_0517_),
    .ZN(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1914_ (.A1(_0521_),
    .A2(_0550_),
    .A3(_0555_),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1915_ (.I0(W1END[3]),
    .I1(AD0),
    .I2(AD1),
    .I3(AD2),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q ),
    .Z(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1916_ (.I0(AD3),
    .I1(BD0),
    .I2(BD1),
    .I3(BD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q ),
    .Z(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1917_ (.I0(_0557_),
    .I1(_0558_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit26.Q ),
    .Z(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1918_ (.I0(N1END[3]),
    .I1(N2END[7]),
    .I2(NN4END[1]),
    .I3(E1END[3]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q ),
    .Z(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1919_ (.I0(E2END[7]),
    .I1(S1END[3]),
    .I2(S2END[7]),
    .I3(W1END[1]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q ),
    .Z(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1920_ (.I0(_0560_),
    .I1(_0561_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit26.Q ),
    .Z(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1921_ (.I0(_0562_),
    .I1(_0559_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit27.Q ),
    .Z(\Inst_RegFile_switch_matrix.JN2BEG6 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1922_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q ),
    .A2(\Inst_RegFile_switch_matrix.JW2BEG6 ),
    .ZN(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1923_ (.A1(_1287_),
    .A2(\Inst_RegFile_switch_matrix.JS2BEG6 ),
    .ZN(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1924_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit30.Q ),
    .A2(_0563_),
    .A3(_0564_),
    .Z(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1925_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q ),
    .A2(_0238_),
    .ZN(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1926_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q ),
    .A2(\Inst_RegFile_switch_matrix.JN2BEG6 ),
    .Z(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1927_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit30.Q ),
    .A2(_0566_),
    .A3(_0567_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame8_bit31.Q ),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1928_ (.A1(_0565_),
    .A2(_0568_),
    .ZN(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1929_ (.I0(E2MID[2]),
    .I1(W2MID[2]),
    .I2(S2MID[2]),
    .I3(\Inst_RegFile_switch_matrix.E2BEG3 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit3.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit2.Q ),
    .Z(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1930_ (.A1(_1287_),
    .A2(_0570_),
    .ZN(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1931_ (.I0(N2MID[5]),
    .I1(E2MID[5]),
    .I2(S2MID[5]),
    .I3(W2MID[5]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit4.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit5.Q ),
    .Z(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1932_ (.I(_0572_),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1933_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q ),
    .A2(_0572_),
    .ZN(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1934_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit30.Q ),
    .A2(_0571_),
    .A3(_0574_),
    .Z(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1935_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit30.Q ),
    .A2(_0571_),
    .A3(_0574_),
    .ZN(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1936_ (.A1(S2END[2]),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q ),
    .Z(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1937_ (.A1(N2END[2]),
    .A2(_1287_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame8_bit30.Q ),
    .C(_0577_),
    .ZN(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1938_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit31.Q ),
    .A2(_0578_),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1939_ (.A1(_0576_),
    .A2(_0579_),
    .B(_0569_),
    .ZN(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1940_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit31.Q ),
    .A2(_0575_),
    .A3(_0578_),
    .B1(_0565_),
    .B2(_0568_),
    .ZN(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1941_ (.A1(_1296_),
    .A2(B_ADR0),
    .ZN(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1942_ (.A1(\Inst_RegFile_32x4.mem[24][0] ),
    .A2(B_ADR0),
    .B(_0582_),
    .ZN(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1943_ (.A1(_1297_),
    .A2(B_ADR0),
    .ZN(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1944_ (.A1(\Inst_RegFile_32x4.mem[26][0] ),
    .A2(B_ADR0),
    .B(_0584_),
    .ZN(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1945_ (.I0(_0583_),
    .I1(_0585_),
    .S(_0486_),
    .Z(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1946_ (.A1(_1299_),
    .A2(B_ADR0),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1947_ (.A1(\Inst_RegFile_32x4.mem[30][0] ),
    .A2(B_ADR0),
    .B(_0587_),
    .ZN(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1948_ (.A1(_1298_),
    .A2(B_ADR0),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1949_ (.A1(\Inst_RegFile_32x4.mem[28][0] ),
    .A2(B_ADR0),
    .B(_0589_),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1950_ (.I0(_0590_),
    .I1(_0588_),
    .S(_0486_),
    .Z(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1951_ (.I0(_0586_),
    .I1(_0591_),
    .S(_0517_),
    .Z(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1952_ (.A1(_0549_),
    .A2(_0592_),
    .B(_0580_),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1953_ (.A1(\Inst_RegFile_32x4.mem[0][0] ),
    .A2(B_ADR0),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1954_ (.A1(_1253_),
    .A2(B_ADR0),
    .B(_0594_),
    .ZN(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1955_ (.A1(\Inst_RegFile_32x4.mem[3][0] ),
    .A2(B_ADR0),
    .ZN(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1956_ (.A1(_1264_),
    .A2(B_ADR0),
    .B(_0486_),
    .C(_0596_),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1957_ (.A1(_0486_),
    .A2(_0595_),
    .B(_0597_),
    .C(_0518_),
    .ZN(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1958_ (.A1(\Inst_RegFile_32x4.mem[7][0] ),
    .A2(B_ADR0),
    .ZN(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1959_ (.A1(_1272_),
    .A2(B_ADR0),
    .B(_0486_),
    .C(_0599_),
    .ZN(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1960_ (.I0(\Inst_RegFile_32x4.mem[4][0] ),
    .I1(\Inst_RegFile_32x4.mem[5][0] ),
    .S(B_ADR0),
    .Z(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1961_ (.A1(_0486_),
    .A2(_0601_),
    .B(_0600_),
    .C(_0517_),
    .ZN(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1962_ (.A1(_0550_),
    .A2(_0598_),
    .A3(_0602_),
    .ZN(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1963_ (.A1(_1283_),
    .A2(B_ADR0),
    .ZN(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1964_ (.A1(\Inst_RegFile_32x4.mem[8][0] ),
    .A2(B_ADR0),
    .B(_0604_),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1965_ (.A1(_1284_),
    .A2(B_ADR0),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1966_ (.A1(\Inst_RegFile_32x4.mem[10][0] ),
    .A2(B_ADR0),
    .B(_0606_),
    .ZN(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1967_ (.I0(_0605_),
    .I1(_0607_),
    .S(_0486_),
    .Z(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1968_ (.A1(_1286_),
    .A2(B_ADR0),
    .ZN(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1969_ (.A1(\Inst_RegFile_32x4.mem[14][0] ),
    .A2(B_ADR0),
    .B(_0609_),
    .ZN(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1970_ (.A1(_1285_),
    .A2(B_ADR0),
    .ZN(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1971_ (.A1(\Inst_RegFile_32x4.mem[12][0] ),
    .A2(B_ADR0),
    .B(_0611_),
    .ZN(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1972_ (.I0(_0612_),
    .I1(_0610_),
    .S(_0486_),
    .Z(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1973_ (.I0(_0608_),
    .I1(_0613_),
    .S(_0517_),
    .Z(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1974_ (.A1(_0549_),
    .A2(_0614_),
    .B(_0581_),
    .ZN(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1975_ (.A1(_0556_),
    .A2(_0593_),
    .B1(_0603_),
    .B2(_0615_),
    .ZN(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1976_ (.I(_0616_),
    .ZN(\Inst_RegFile_32x4.BD_comb[0] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1977_ (.A1(\Inst_RegFile_32x4.BD_reg[0] ),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q ),
    .ZN(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1978_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q ),
    .A2(_0616_),
    .B(_0617_),
    .ZN(BD0));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1979_ (.A1(_1304_),
    .A2(B_ADR0),
    .ZN(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1980_ (.A1(\Inst_RegFile_32x4.mem[17][1] ),
    .A2(B_ADR0),
    .B(_0486_),
    .C(_0618_),
    .ZN(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1981_ (.A1(\Inst_RegFile_32x4.mem[19][1] ),
    .A2(B_ADR0),
    .ZN(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1982_ (.A1(_1305_),
    .A2(B_ADR0),
    .B(_0486_),
    .C(_0620_),
    .ZN(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1983_ (.A1(_0517_),
    .A2(_0619_),
    .ZN(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1984_ (.I0(\Inst_RegFile_32x4.mem[22][1] ),
    .I1(\Inst_RegFile_32x4.mem[23][1] ),
    .S(B_ADR0),
    .Z(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1985_ (.A1(\Inst_RegFile_32x4.mem[20][1] ),
    .A2(B_ADR0),
    .ZN(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1986_ (.A1(_1306_),
    .A2(B_ADR0),
    .B(_0624_),
    .ZN(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1987_ (.I0(_0625_),
    .I1(_0623_),
    .S(_0486_),
    .Z(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1988_ (.A1(_0621_),
    .A2(_0622_),
    .B1(_0626_),
    .B2(_0517_),
    .C(_0549_),
    .ZN(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1989_ (.A1(_1307_),
    .A2(B_ADR0),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1990_ (.A1(\Inst_RegFile_32x4.mem[25][1] ),
    .A2(B_ADR0),
    .B(_0486_),
    .C(_0628_),
    .ZN(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1991_ (.A1(\Inst_RegFile_32x4.mem[27][1] ),
    .A2(B_ADR0),
    .ZN(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1992_ (.A1(_1308_),
    .A2(B_ADR0),
    .B(_0486_),
    .C(_0630_),
    .ZN(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1993_ (.A1(_0517_),
    .A2(_0629_),
    .ZN(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1994_ (.A1(_1310_),
    .A2(B_ADR0),
    .ZN(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1995_ (.A1(\Inst_RegFile_32x4.mem[30][1] ),
    .A2(B_ADR0),
    .B(_0633_),
    .ZN(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1996_ (.A1(_1309_),
    .A2(B_ADR0),
    .ZN(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1997_ (.A1(\Inst_RegFile_32x4.mem[29][1] ),
    .A2(B_ADR0),
    .B(_0486_),
    .C(_0635_),
    .ZN(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1998_ (.A1(_0486_),
    .A2(_0634_),
    .B(_0636_),
    .ZN(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1999_ (.A1(_0631_),
    .A2(_0632_),
    .B1(_0637_),
    .B2(_0517_),
    .C(_0550_),
    .ZN(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2000_ (.I0(\Inst_RegFile_32x4.mem[0][1] ),
    .I1(\Inst_RegFile_32x4.mem[1][1] ),
    .S(B_ADR0),
    .Z(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2001_ (.A1(\Inst_RegFile_32x4.mem[3][1] ),
    .A2(B_ADR0),
    .ZN(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2002_ (.A1(_1300_),
    .A2(B_ADR0),
    .B(_0486_),
    .C(_0640_),
    .ZN(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2003_ (.A1(_0486_),
    .A2(_0639_),
    .B(_0641_),
    .C(_0518_),
    .ZN(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2004_ (.A1(\Inst_RegFile_32x4.mem[7][1] ),
    .A2(B_ADR0),
    .ZN(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2005_ (.A1(_1302_),
    .A2(B_ADR0),
    .B(_0486_),
    .C(_0643_),
    .ZN(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2006_ (.A1(\Inst_RegFile_32x4.mem[4][1] ),
    .A2(B_ADR0),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2007_ (.A1(_1301_),
    .A2(B_ADR0),
    .B(_0645_),
    .ZN(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2008_ (.A1(_0486_),
    .A2(_0646_),
    .B(_0644_),
    .C(_0517_),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2009_ (.A1(_0550_),
    .A2(_0642_),
    .A3(_0647_),
    .Z(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2010_ (.I0(\Inst_RegFile_32x4.mem[10][1] ),
    .I1(\Inst_RegFile_32x4.mem[11][1] ),
    .S(B_ADR0),
    .Z(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2011_ (.I0(\Inst_RegFile_32x4.mem[8][1] ),
    .I1(\Inst_RegFile_32x4.mem[9][1] ),
    .S(B_ADR0),
    .Z(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2012_ (.I0(_0650_),
    .I1(_0649_),
    .S(_0486_),
    .Z(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2013_ (.I0(\Inst_RegFile_32x4.mem[14][1] ),
    .I1(\Inst_RegFile_32x4.mem[15][1] ),
    .S(B_ADR0),
    .Z(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2014_ (.A1(\Inst_RegFile_32x4.mem[12][1] ),
    .A2(B_ADR0),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2015_ (.A1(_1303_),
    .A2(B_ADR0),
    .B(_0653_),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2016_ (.I0(_0654_),
    .I1(_0652_),
    .S(_0486_),
    .Z(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2017_ (.I0(_0651_),
    .I1(_0655_),
    .S(_0517_),
    .Z(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2018_ (.A1(_0550_),
    .A2(_0656_),
    .B(_0580_),
    .ZN(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2019_ (.A1(_0580_),
    .A2(_0627_),
    .A3(_0638_),
    .B1(_0648_),
    .B2(_0657_),
    .ZN(\Inst_RegFile_32x4.BD_comb[1] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2020_ (.I0(\Inst_RegFile_32x4.BD_comb[1] ),
    .I1(\Inst_RegFile_32x4.BD_reg[1] ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q ),
    .Z(BD1));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2021_ (.A1(\Inst_RegFile_32x4.mem[16][3] ),
    .A2(B_ADR0),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2022_ (.A1(_1333_),
    .A2(B_ADR0),
    .B(_0658_),
    .ZN(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2023_ (.A1(\Inst_RegFile_32x4.mem[19][3] ),
    .A2(B_ADR0),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2024_ (.A1(_1334_),
    .A2(B_ADR0),
    .B(_0486_),
    .C(_0660_),
    .ZN(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2025_ (.A1(_0486_),
    .A2(_0659_),
    .B(_0661_),
    .C(_0518_),
    .ZN(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2026_ (.A1(\Inst_RegFile_32x4.mem[23][3] ),
    .A2(B_ADR0),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2027_ (.A1(_1336_),
    .A2(B_ADR0),
    .B(_0486_),
    .C(_0663_),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2028_ (.A1(\Inst_RegFile_32x4.mem[20][3] ),
    .A2(B_ADR0),
    .ZN(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2029_ (.A1(_1335_),
    .A2(B_ADR0),
    .B(_0665_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2030_ (.A1(_0486_),
    .A2(_0666_),
    .B(_0664_),
    .C(_0517_),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2031_ (.A1(_0550_),
    .A2(_0662_),
    .A3(_0667_),
    .ZN(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2032_ (.A1(_1337_),
    .A2(B_ADR0),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2033_ (.A1(\Inst_RegFile_32x4.mem[24][3] ),
    .A2(B_ADR0),
    .B(_0669_),
    .ZN(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2034_ (.A1(_1338_),
    .A2(B_ADR0),
    .ZN(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2035_ (.A1(\Inst_RegFile_32x4.mem[26][3] ),
    .A2(B_ADR0),
    .B(_0671_),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2036_ (.I0(_0670_),
    .I1(_0672_),
    .S(_0486_),
    .Z(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2037_ (.A1(_1340_),
    .A2(B_ADR0),
    .ZN(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2038_ (.A1(\Inst_RegFile_32x4.mem[30][3] ),
    .A2(B_ADR0),
    .B(_0674_),
    .ZN(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2039_ (.A1(_1339_),
    .A2(B_ADR0),
    .ZN(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2040_ (.A1(\Inst_RegFile_32x4.mem[28][3] ),
    .A2(B_ADR0),
    .B(_0676_),
    .ZN(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2041_ (.I0(_0677_),
    .I1(_0675_),
    .S(_0486_),
    .Z(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2042_ (.I0(_0673_),
    .I1(_0678_),
    .S(_0517_),
    .Z(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2043_ (.A1(_0549_),
    .A2(_0679_),
    .B(_0580_),
    .ZN(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2044_ (.I0(\Inst_RegFile_32x4.mem[0][3] ),
    .I1(\Inst_RegFile_32x4.mem[1][3] ),
    .S(B_ADR0),
    .Z(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2045_ (.A1(\Inst_RegFile_32x4.mem[3][3] ),
    .A2(B_ADR0),
    .ZN(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2046_ (.A1(_1326_),
    .A2(B_ADR0),
    .B(_0486_),
    .C(_0682_),
    .ZN(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2047_ (.A1(_0486_),
    .A2(_0681_),
    .B(_0683_),
    .C(_0518_),
    .ZN(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2048_ (.A1(\Inst_RegFile_32x4.mem[7][3] ),
    .A2(B_ADR0),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2049_ (.A1(_1328_),
    .A2(B_ADR0),
    .B(_0486_),
    .C(_0685_),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2050_ (.A1(\Inst_RegFile_32x4.mem[4][3] ),
    .A2(B_ADR0),
    .ZN(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2051_ (.A1(_1327_),
    .A2(B_ADR0),
    .B(_0687_),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2052_ (.A1(_0486_),
    .A2(_0688_),
    .B(_0686_),
    .C(_0517_),
    .ZN(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2053_ (.A1(_0550_),
    .A2(_0684_),
    .A3(_0689_),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2054_ (.A1(_1329_),
    .A2(B_ADR0),
    .ZN(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2055_ (.A1(\Inst_RegFile_32x4.mem[8][3] ),
    .A2(B_ADR0),
    .B(_0691_),
    .ZN(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2056_ (.A1(_1330_),
    .A2(B_ADR0),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2057_ (.A1(\Inst_RegFile_32x4.mem[10][3] ),
    .A2(B_ADR0),
    .B(_0693_),
    .ZN(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2058_ (.I0(_0692_),
    .I1(_0694_),
    .S(_0486_),
    .Z(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2059_ (.A1(_1332_),
    .A2(B_ADR0),
    .ZN(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2060_ (.A1(\Inst_RegFile_32x4.mem[14][3] ),
    .A2(B_ADR0),
    .B(_0696_),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2061_ (.A1(_1331_),
    .A2(B_ADR0),
    .ZN(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2062_ (.A1(\Inst_RegFile_32x4.mem[12][3] ),
    .A2(B_ADR0),
    .B(_0698_),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2063_ (.I0(_0699_),
    .I1(_0697_),
    .S(_0486_),
    .Z(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2064_ (.I0(_0695_),
    .I1(_0700_),
    .S(_0517_),
    .Z(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2065_ (.A1(_0549_),
    .A2(_0701_),
    .B(_0581_),
    .ZN(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2066_ (.A1(_0668_),
    .A2(_0680_),
    .B1(_0690_),
    .B2(_0702_),
    .ZN(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2067_ (.I(_0703_),
    .ZN(\Inst_RegFile_32x4.BD_comb[3] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2068_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q ),
    .A2(\Inst_RegFile_32x4.BD_reg[3] ),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2069_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q ),
    .A2(_0703_),
    .B(_0704_),
    .ZN(BD3));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2070_ (.A1(\Inst_RegFile_32x4.mem[0][2] ),
    .A2(B_ADR0),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2071_ (.A1(_1311_),
    .A2(B_ADR0),
    .B(_0705_),
    .ZN(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2072_ (.A1(\Inst_RegFile_32x4.mem[3][2] ),
    .A2(B_ADR0),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2073_ (.A1(_1312_),
    .A2(B_ADR0),
    .B(_0486_),
    .C(_0707_),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2074_ (.A1(_0486_),
    .A2(_0706_),
    .B(_0708_),
    .C(_0518_),
    .ZN(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2075_ (.A1(\Inst_RegFile_32x4.mem[7][2] ),
    .A2(B_ADR0),
    .ZN(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2076_ (.A1(_1313_),
    .A2(B_ADR0),
    .B(_0486_),
    .C(_0710_),
    .ZN(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2077_ (.I0(\Inst_RegFile_32x4.mem[4][2] ),
    .I1(\Inst_RegFile_32x4.mem[5][2] ),
    .S(B_ADR0),
    .Z(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2078_ (.A1(_0486_),
    .A2(_0712_),
    .B(_0711_),
    .C(_0517_),
    .ZN(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2079_ (.A1(_0550_),
    .A2(_0709_),
    .A3(_0713_),
    .ZN(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2080_ (.A1(_1314_),
    .A2(B_ADR0),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2081_ (.A1(\Inst_RegFile_32x4.mem[8][2] ),
    .A2(B_ADR0),
    .B(_0715_),
    .ZN(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2082_ (.A1(_1315_),
    .A2(B_ADR0),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2083_ (.A1(\Inst_RegFile_32x4.mem[10][2] ),
    .A2(B_ADR0),
    .B(_0717_),
    .ZN(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2084_ (.I0(_0716_),
    .I1(_0718_),
    .S(_0486_),
    .Z(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2085_ (.A1(_1317_),
    .A2(B_ADR0),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2086_ (.A1(\Inst_RegFile_32x4.mem[14][2] ),
    .A2(B_ADR0),
    .B(_0720_),
    .ZN(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2087_ (.A1(_1316_),
    .A2(B_ADR0),
    .ZN(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2088_ (.A1(\Inst_RegFile_32x4.mem[12][2] ),
    .A2(B_ADR0),
    .B(_0722_),
    .ZN(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2089_ (.I0(_0723_),
    .I1(_0721_),
    .S(_0486_),
    .Z(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2090_ (.I0(_0719_),
    .I1(_0724_),
    .S(_0517_),
    .Z(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2091_ (.A1(_0549_),
    .A2(_0725_),
    .B(_0581_),
    .ZN(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2092_ (.A1(\Inst_RegFile_32x4.mem[16][2] ),
    .A2(B_ADR0),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2093_ (.A1(_1318_),
    .A2(B_ADR0),
    .B(_0727_),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2094_ (.A1(\Inst_RegFile_32x4.mem[19][2] ),
    .A2(B_ADR0),
    .ZN(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2095_ (.A1(_1319_),
    .A2(B_ADR0),
    .B(_0486_),
    .C(_0729_),
    .ZN(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2096_ (.A1(_0486_),
    .A2(_0728_),
    .B(_0730_),
    .C(_0518_),
    .ZN(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2097_ (.A1(\Inst_RegFile_32x4.mem[23][2] ),
    .A2(B_ADR0),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2098_ (.A1(_1321_),
    .A2(B_ADR0),
    .B(_0486_),
    .C(_0732_),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2099_ (.A1(\Inst_RegFile_32x4.mem[20][2] ),
    .A2(B_ADR0),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2100_ (.A1(_1320_),
    .A2(B_ADR0),
    .B(_0734_),
    .ZN(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2101_ (.A1(_0486_),
    .A2(_0735_),
    .B(_0733_),
    .C(_0517_),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2102_ (.A1(_0550_),
    .A2(_0731_),
    .A3(_0736_),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2103_ (.A1(_1322_),
    .A2(B_ADR0),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2104_ (.A1(\Inst_RegFile_32x4.mem[24][2] ),
    .A2(B_ADR0),
    .B(_0738_),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2105_ (.A1(_1323_),
    .A2(B_ADR0),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2106_ (.A1(\Inst_RegFile_32x4.mem[26][2] ),
    .A2(B_ADR0),
    .B(_0740_),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2107_ (.I0(_0739_),
    .I1(_0741_),
    .S(_0486_),
    .Z(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2108_ (.A1(_1325_),
    .A2(B_ADR0),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2109_ (.A1(\Inst_RegFile_32x4.mem[30][2] ),
    .A2(B_ADR0),
    .B(_0743_),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2110_ (.A1(_1324_),
    .A2(B_ADR0),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2111_ (.A1(\Inst_RegFile_32x4.mem[28][2] ),
    .A2(B_ADR0),
    .B(_0745_),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2112_ (.I0(_0746_),
    .I1(_0744_),
    .S(_0486_),
    .Z(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2113_ (.I0(_0742_),
    .I1(_0747_),
    .S(_0517_),
    .Z(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2114_ (.A1(_0549_),
    .A2(_0748_),
    .B(_0580_),
    .ZN(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2115_ (.A1(_0714_),
    .A2(_0726_),
    .B1(_0737_),
    .B2(_0749_),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2116_ (.I(_0750_),
    .ZN(\Inst_RegFile_32x4.BD_comb[2] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2117_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q ),
    .A2(\Inst_RegFile_32x4.BD_reg[2] ),
    .ZN(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2118_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q ),
    .A2(_0750_),
    .B(_0751_),
    .ZN(BD2));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2119_ (.I0(W1END[3]),
    .I1(AD0),
    .I2(AD1),
    .I3(AD2),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q ),
    .Z(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2120_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q ),
    .A2(_0752_),
    .ZN(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2121_ (.I0(AD3),
    .I1(BD2),
    .I2(BD1),
    .I3(BD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q ),
    .Z(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2122_ (.A1(_1252_),
    .A2(_0754_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame4_bit19.Q ),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2123_ (.I0(N1END[1]),
    .I1(N2END[5]),
    .I2(NN4END[3]),
    .I3(E1END[1]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q ),
    .Z(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2124_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q ),
    .A2(_0756_),
    .ZN(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2125_ (.I0(E2END[5]),
    .I1(S1END[1]),
    .I2(S2END[5]),
    .I3(W1END[1]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q ),
    .Z(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2126_ (.A1(_1252_),
    .A2(_0758_),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2127_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit19.Q ),
    .A2(_0757_),
    .A3(_0759_),
    .B1(_0753_),
    .B2(_0755_),
    .ZN(\Inst_RegFile_switch_matrix.JN2BEG4 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2128_ (.I(\Inst_RegFile_switch_matrix.JN2BEG4 ),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2129_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit24.Q ),
    .A2(_0760_),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2130_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit24.Q ),
    .A2(S4END[3]),
    .B(\Inst_RegFile_ConfigMem.Inst_frame0_bit25.Q ),
    .C(_0761_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2131_ (.A1(_1251_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame0_bit24.Q ),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2132_ (.A1(N4END[3]),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame0_bit24.Q ),
    .B(_0763_),
    .ZN(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2133_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit25.Q ),
    .A2(_0764_),
    .B(_0762_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame8_bit21.Q ),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2134_ (.I0(N2END[7]),
    .I1(E2END[7]),
    .I2(S2END[7]),
    .I3(WW4END[0]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit25.Q ),
    .Z(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2135_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit21.Q ),
    .A2(_0766_),
    .B(_0765_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame8_bit22.Q ),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2136_ (.I0(S2MID[6]),
    .I1(\Inst_RegFile_switch_matrix.JN2BEG6 ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame7_bit24.Q ),
    .Z(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2137_ (.A1(N2MID[6]),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame7_bit24.Q ),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2138_ (.A1(_1247_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame7_bit24.Q ),
    .B(\Inst_RegFile_ConfigMem.Inst_frame7_bit25.Q ),
    .C(_0769_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2139_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame7_bit25.Q ),
    .A2(_0768_),
    .B(_0770_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame8_bit21.Q ),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2140_ (.I0(N2MID[7]),
    .I1(E2MID[7]),
    .I2(S2MID[7]),
    .I3(W2MID[7]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit24.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit25.Q ),
    .Z(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2141_ (.A1(_1249_),
    .A2(_0772_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2142_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit22.Q ),
    .A2(_0771_),
    .A3(_0773_),
    .B(_0767_),
    .ZN(B_ADR0));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2143_ (.I0(W6END[0]),
    .I1(AD0),
    .I2(AD1),
    .I3(AD2),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q ),
    .Z(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2144_ (.I0(BD0),
    .I1(BD2),
    .I2(BD1),
    .I3(BD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q ),
    .Z(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2145_ (.I0(_0774_),
    .I1(_0775_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit14.Q ),
    .Z(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2146_ (.I0(N2END[4]),
    .I1(N4END[0]),
    .I2(E1END[2]),
    .I3(E2END[4]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q ),
    .Z(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2147_ (.I0(E6END[0]),
    .I1(S2END[4]),
    .I2(W2END[4]),
    .I3(WW4END[3]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q ),
    .Z(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2148_ (.I0(_0777_),
    .I1(_0778_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit14.Q ),
    .Z(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2149_ (.I0(_0779_),
    .I1(_0776_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit15.Q ),
    .Z(\Inst_RegFile_switch_matrix.JN2BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2150_ (.I0(N4END[3]),
    .I1(E2END[3]),
    .I2(W2END[3]),
    .I3(\Inst_RegFile_switch_matrix.JN2BEG3 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame0_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame0_bit17.Q ),
    .Z(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2151_ (.I(_0780_),
    .ZN(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2152_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit10.Q ),
    .A2(_0781_),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2153_ (.I0(N2END[7]),
    .I1(S2END[7]),
    .I2(EE4END[2]),
    .I3(W2END[7]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit17.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit16.Q ),
    .Z(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2154_ (.I(_0783_),
    .ZN(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2155_ (.I0(N2MID[6]),
    .I1(E2MID[6]),
    .I2(W2MID[6]),
    .I3(\Inst_RegFile_switch_matrix.JN2BEG5 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit17.Q ),
    .Z(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2156_ (.A1(W2MID[7]),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame6_bit16.Q ),
    .ZN(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2157_ (.A1(_1248_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame6_bit16.Q ),
    .B(\Inst_RegFile_ConfigMem.Inst_frame6_bit17.Q ),
    .C(_0786_),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2158_ (.I0(N2MID[7]),
    .I1(E2MID[7]),
    .S(\Inst_RegFile_ConfigMem.Inst_frame6_bit16.Q ),
    .Z(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2159_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame6_bit17.Q ),
    .A2(_0788_),
    .B(_0787_),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2160_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit10.Q ),
    .A2(_0789_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame8_bit11.Q ),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2161_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit10.Q ),
    .A2(_0785_),
    .B(_0790_),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2162_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit10.Q ),
    .A2(_0783_),
    .B(_0782_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame8_bit11.Q ),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2163_ (.A1(_0791_),
    .A2(_0792_),
    .ZN(A_ADR0));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2164_ (.I0(W6END[1]),
    .I1(AD0),
    .I2(AD1),
    .I3(AD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q ),
    .Z(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2165_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit10.Q ),
    .A2(_0793_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2166_ (.I0(BD0),
    .I1(BD2),
    .I2(BD1),
    .I3(BD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q ),
    .Z(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2167_ (.A1(_1354_),
    .A2(_0795_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame1_bit11.Q ),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2168_ (.I0(N1END[1]),
    .I1(N2END[3]),
    .I2(NN4END[2]),
    .I3(E2END[3]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q ),
    .Z(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2169_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit10.Q ),
    .A2(_0797_),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2170_ (.I0(E6END[1]),
    .I1(S2END[3]),
    .I2(S4END[3]),
    .I3(W2END[3]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q ),
    .Z(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2171_ (.A1(_1354_),
    .A2(_0799_),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2172_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit11.Q ),
    .A2(_0798_),
    .A3(_0800_),
    .B1(_0794_),
    .B2(_0796_),
    .ZN(\Inst_RegFile_switch_matrix.JW2BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2173_ (.I0(BD0),
    .I1(BD2),
    .I2(BD1),
    .I3(BD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q ),
    .Z(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2174_ (.I0(W6END[1]),
    .I1(AD0),
    .I2(AD1),
    .I3(AD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q ),
    .Z(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2175_ (.I0(_0802_),
    .I1(_0801_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit10.Q ),
    .Z(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2176_ (.I0(E6END[1]),
    .I1(S2END[3]),
    .I2(S4END[3]),
    .I3(W2END[3]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q ),
    .Z(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2177_ (.I0(N2END[3]),
    .I1(E2END[3]),
    .I2(E1END[1]),
    .I3(EE4END[2]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q ),
    .Z(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2178_ (.I0(_0805_),
    .I1(_0804_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit10.Q ),
    .Z(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2179_ (.I0(_0806_),
    .I1(_0803_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit11.Q ),
    .Z(\Inst_RegFile_switch_matrix.JS2BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2180_ (.I0(W6END[1]),
    .I1(AD0),
    .I2(AD1),
    .I3(AD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q ),
    .Z(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2181_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit10.Q ),
    .A2(_0807_),
    .ZN(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2182_ (.I0(BD0),
    .I1(BD2),
    .I2(BD1),
    .I3(BD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q ),
    .Z(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2183_ (.A1(_1355_),
    .A2(_0809_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame3_bit11.Q ),
    .ZN(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2184_ (.I0(N1END[1]),
    .I1(N2END[3]),
    .I2(N4END[3]),
    .I3(E2END[3]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q ),
    .Z(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2185_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit10.Q ),
    .A2(_0811_),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2186_ (.I0(E6END[1]),
    .I1(S2END[3]),
    .I2(SS4END[2]),
    .I3(W2END[3]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q ),
    .Z(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2187_ (.A1(_1355_),
    .A2(_0813_),
    .ZN(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2188_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit11.Q ),
    .A2(_0812_),
    .A3(_0814_),
    .B1(_0808_),
    .B2(_0810_),
    .ZN(\Inst_RegFile_switch_matrix.E2BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2189_ (.I0(W6END[1]),
    .I1(AD0),
    .I2(AD1),
    .I3(AD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q ),
    .Z(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2190_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit10.Q ),
    .A2(_0815_),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2191_ (.I0(BD0),
    .I1(BD2),
    .I2(BD1),
    .I3(BD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q ),
    .Z(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2192_ (.A1(_0128_),
    .A2(_0817_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame4_bit11.Q ),
    .ZN(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2193_ (.I0(N2END[3]),
    .I1(E1END[1]),
    .I2(N4END[3]),
    .I3(E2END[3]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q ),
    .Z(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2194_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame4_bit10.Q ),
    .A2(_0819_),
    .ZN(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2195_ (.I0(E6END[1]),
    .I1(S2END[3]),
    .I2(W2END[3]),
    .I3(WW4END[2]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q ),
    .Z(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2196_ (.A1(_0128_),
    .A2(_0821_),
    .B(_0129_),
    .ZN(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2197_ (.A1(_0816_),
    .A2(_0818_),
    .B1(_0820_),
    .B2(_0822_),
    .ZN(\Inst_RegFile_switch_matrix.JN2BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2198_ (.I0(W6END[0]),
    .I1(AD0),
    .I2(AD2),
    .I3(AD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q ),
    .Z(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2199_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q ),
    .A2(_0823_),
    .ZN(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2200_ (.I0(BD0),
    .I1(BD2),
    .I2(BD1),
    .I3(BD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q ),
    .Z(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2201_ (.A1(_0130_),
    .A2(_0825_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame1_bit7.Q ),
    .ZN(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2202_ (.I0(S2END[2]),
    .I1(S4END[2]),
    .I2(SS4END[1]),
    .I3(W2END[2]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q ),
    .Z(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2203_ (.A1(_0130_),
    .A2(_0827_),
    .ZN(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2204_ (.I0(N1END[0]),
    .I1(E2END[2]),
    .I2(N2END[2]),
    .I3(E6END[0]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q ),
    .Z(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2205_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q ),
    .A2(_0829_),
    .ZN(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2206_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit7.Q ),
    .A2(_0828_),
    .A3(_0830_),
    .B1(_0824_),
    .B2(_0826_),
    .ZN(\Inst_RegFile_switch_matrix.JW2BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2207_ (.I0(W6END[0]),
    .I1(AD0),
    .I2(AD2),
    .I3(AD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q ),
    .Z(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2208_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q ),
    .A2(_0831_),
    .ZN(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2209_ (.I0(BD0),
    .I1(BD2),
    .I2(BD1),
    .I3(BD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q ),
    .Z(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2210_ (.A1(_0131_),
    .A2(_0833_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame2_bit7.Q ),
    .ZN(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2211_ (.I0(N2END[2]),
    .I1(E2END[2]),
    .I2(E1END[0]),
    .I3(E6END[0]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q ),
    .Z(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2212_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q ),
    .A2(_0835_),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2213_ (.I0(S2END[2]),
    .I1(S4END[2]),
    .I2(W2END[2]),
    .I3(WW4END[1]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q ),
    .Z(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2214_ (.A1(_0131_),
    .A2(_0837_),
    .ZN(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2215_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit7.Q ),
    .A2(_0836_),
    .A3(_0838_),
    .B1(_0832_),
    .B2(_0834_),
    .ZN(\Inst_RegFile_switch_matrix.JS2BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2216_ (.I0(W6END[0]),
    .I1(AD0),
    .I2(AD2),
    .I3(AD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q ),
    .Z(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2217_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit6.Q ),
    .A2(_0839_),
    .ZN(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2218_ (.I0(BD0),
    .I1(BD2),
    .I2(BD1),
    .I3(BD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q ),
    .Z(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2219_ (.A1(_0132_),
    .A2(_0841_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame3_bit7.Q ),
    .ZN(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2220_ (.I0(E2END[2]),
    .I1(S2END[2]),
    .I2(E6END[0]),
    .I3(W2END[2]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q ),
    .Z(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2221_ (.A1(_0132_),
    .A2(_0843_),
    .ZN(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2222_ (.I0(N1END[0]),
    .I1(N2END[2]),
    .I2(N4END[2]),
    .I3(NN4END[1]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q ),
    .Z(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2223_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit6.Q ),
    .A2(_0845_),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2224_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit7.Q ),
    .A2(_0844_),
    .A3(_0846_),
    .B1(_0840_),
    .B2(_0842_),
    .ZN(\Inst_RegFile_switch_matrix.E2BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2225_ (.I0(W6END[0]),
    .I1(AD0),
    .I2(AD2),
    .I3(AD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q ),
    .Z(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2226_ (.I0(BD0),
    .I1(BD2),
    .I2(BD1),
    .I3(BD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q ),
    .Z(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2227_ (.I0(_0847_),
    .I1(_0848_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit6.Q ),
    .Z(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2228_ (.I0(N2END[2]),
    .I1(E1END[0]),
    .I2(N4END[2]),
    .I3(E2END[2]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q ),
    .Z(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2229_ (.I0(EE4END[1]),
    .I1(E6END[0]),
    .I2(S2END[2]),
    .I3(W2END[2]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q ),
    .Z(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2230_ (.I0(_0850_),
    .I1(_0851_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit6.Q ),
    .Z(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2231_ (.I0(_0852_),
    .I1(_0849_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit7.Q ),
    .Z(\Inst_RegFile_switch_matrix.JN2BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2232_ (.I0(WW4END[0]),
    .I1(AD0),
    .I2(AD1),
    .I3(AD2),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q ),
    .Z(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2233_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit30.Q ),
    .A2(_0853_),
    .ZN(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2234_ (.I0(AD3),
    .I1(BD0),
    .I2(BD1),
    .I3(BD2),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q ),
    .Z(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2235_ (.A1(_0133_),
    .A2(_0855_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame1_bit31.Q ),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2236_ (.I0(S1END[0]),
    .I1(S2END[0]),
    .I2(S1END[2]),
    .I3(W1END[0]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q ),
    .Z(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2237_ (.A1(_0133_),
    .A2(_0857_),
    .ZN(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2238_ (.I0(N1END[0]),
    .I1(E1END[0]),
    .I2(N2END[0]),
    .I3(E2END[0]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q ),
    .Z(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2239_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit30.Q ),
    .A2(_0859_),
    .ZN(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2240_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame1_bit31.Q ),
    .A2(_0858_),
    .A3(_0860_),
    .B1(_0854_),
    .B2(_0856_),
    .ZN(\Inst_RegFile_switch_matrix.JW2BEG7 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2241_ (.I0(W6END[1]),
    .I1(AD2),
    .I2(AD1),
    .I3(AD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q ),
    .Z(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2242_ (.I0(BD0),
    .I1(BD2),
    .I2(BD1),
    .I3(BD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q ),
    .Z(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2243_ (.I0(_0861_),
    .I1(_0862_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame1_bit2.Q ),
    .Z(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2244_ (.I0(N1END[3]),
    .I1(N2END[1]),
    .I2(E2END[1]),
    .I3(E6END[1]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q ),
    .Z(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2245_ (.I0(S2END[1]),
    .I1(S4END[1]),
    .I2(SS4END[0]),
    .I3(W2END[1]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q ),
    .Z(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2246_ (.I0(_0864_),
    .I1(_0865_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame1_bit2.Q ),
    .Z(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2247_ (.I0(_0866_),
    .I1(_0863_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame1_bit3.Q ),
    .Z(\Inst_RegFile_switch_matrix.JW2BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2248_ (.I0(AD3),
    .I1(BD0),
    .I2(BD1),
    .I3(BD2),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q ),
    .Z(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2249_ (.I0(W1END[2]),
    .I1(AD0),
    .I2(AD1),
    .I3(AD2),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q ),
    .Z(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2250_ (.I0(_0868_),
    .I1(_0867_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit30.Q ),
    .Z(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2251_ (.I0(S1END[0]),
    .I1(S2END[0]),
    .I2(SS4END[0]),
    .I3(W1END[0]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q ),
    .Z(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2252_ (.I0(N1END[0]),
    .I1(E1END[0]),
    .I2(N2END[0]),
    .I3(E2END[0]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q ),
    .Z(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2253_ (.I0(_0871_),
    .I1(_0870_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit30.Q ),
    .Z(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2254_ (.I0(_0872_),
    .I1(_0869_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame2_bit31.Q ),
    .Z(\Inst_RegFile_switch_matrix.JS2BEG7 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2255_ (.I0(BD0),
    .I1(BD2),
    .I2(BD1),
    .I3(BD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q ),
    .Z(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2256_ (.A1(_0134_),
    .A2(_0873_),
    .ZN(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2257_ (.I0(W6END[1]),
    .I1(AD2),
    .I2(AD1),
    .I3(AD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q ),
    .Z(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2258_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit2.Q ),
    .A2(_0875_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame2_bit3.Q ),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2259_ (.I0(S2END[1]),
    .I1(W2END[1]),
    .I2(S4END[1]),
    .I3(WW4END[0]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q ),
    .Z(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2260_ (.A1(_0134_),
    .A2(_0877_),
    .ZN(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2261_ (.I0(N2END[1]),
    .I1(E2END[1]),
    .I2(E1END[3]),
    .I3(E6END[1]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q ),
    .Z(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2262_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit2.Q ),
    .A2(_0879_),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2263_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame2_bit3.Q ),
    .A2(_0878_),
    .A3(_0880_),
    .B1(_0874_),
    .B2(_0876_),
    .ZN(\Inst_RegFile_switch_matrix.JS2BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2264_ (.I0(AD3),
    .I1(BD0),
    .I2(BD1),
    .I3(BD2),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q ),
    .Z(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2265_ (.I(_0881_),
    .ZN(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2266_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit30.Q ),
    .A2(_0882_),
    .ZN(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2267_ (.I0(W1END[0]),
    .I1(AD0),
    .I2(AD1),
    .I3(AD2),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q ),
    .Z(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2268_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit30.Q ),
    .A2(_0884_),
    .B(_0883_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame3_bit31.Q ),
    .ZN(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2269_ (.I0(EE4END[0]),
    .I1(S1END[2]),
    .I2(S1END[0]),
    .I3(S2END[0]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q ),
    .Z(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2270_ (.I(_0886_),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2271_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit30.Q ),
    .A2(_0887_),
    .ZN(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2272_ (.I0(N1END[0]),
    .I1(E1END[0]),
    .I2(N2END[0]),
    .I3(E2END[0]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q ),
    .Z(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2273_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit30.Q ),
    .A2(_0889_),
    .B(_0888_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2274_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit31.Q ),
    .A2(_0890_),
    .B(_0885_),
    .ZN(\Inst_RegFile_switch_matrix.E2BEG7 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2275_ (.I0(BD0),
    .I1(BD2),
    .I2(BD1),
    .I3(BD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q ),
    .Z(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2276_ (.A1(_0135_),
    .A2(_0891_),
    .ZN(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2277_ (.I0(W6END[1]),
    .I1(AD2),
    .I2(AD1),
    .I3(AD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q ),
    .Z(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2278_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit2.Q ),
    .A2(_0893_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame3_bit3.Q ),
    .ZN(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2279_ (.I0(N1END[3]),
    .I1(N2END[1]),
    .I2(N4END[1]),
    .I3(NN4END[0]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q ),
    .Z(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2280_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit2.Q ),
    .A2(_0895_),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2281_ (.I0(E2END[1]),
    .I1(S2END[1]),
    .I2(E6END[1]),
    .I3(W2END[1]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q ),
    .Z(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2282_ (.A1(_0135_),
    .A2(_0897_),
    .ZN(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2283_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame3_bit3.Q ),
    .A2(_0896_),
    .A3(_0898_),
    .B1(_0892_),
    .B2(_0894_),
    .ZN(\Inst_RegFile_switch_matrix.E2BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2284_ (.I0(W1END[2]),
    .I1(AD0),
    .I2(AD1),
    .I3(AD2),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q ),
    .Z(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2285_ (.I0(AD3),
    .I1(BD0),
    .I2(BD1),
    .I3(BD2),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q ),
    .Z(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2286_ (.I0(_0899_),
    .I1(_0900_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit30.Q ),
    .Z(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2287_ (.I0(E2END[0]),
    .I1(S2END[0]),
    .I2(S1END[0]),
    .I3(W1END[0]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q ),
    .Z(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2288_ (.I0(N1END[0]),
    .I1(N2END[0]),
    .I2(NN4END[0]),
    .I3(E1END[0]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q ),
    .Z(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2289_ (.I0(_0903_),
    .I1(_0902_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit30.Q ),
    .Z(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2290_ (.I0(_0904_),
    .I1(_0901_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit31.Q ),
    .Z(\Inst_RegFile_switch_matrix.JN2BEG7 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2291_ (.I0(W6END[1]),
    .I1(AD2),
    .I2(AD1),
    .I3(AD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q ),
    .Z(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2292_ (.I0(BD0),
    .I1(BD2),
    .I2(BD1),
    .I3(BD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q ),
    .Z(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2293_ (.I0(_0905_),
    .I1(_0906_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit2.Q ),
    .Z(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2294_ (.I0(EE4END[0]),
    .I1(E6END[1]),
    .I2(S2END[1]),
    .I3(W2END[1]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q ),
    .Z(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2295_ (.I0(N2END[1]),
    .I1(N4END[1]),
    .I2(E1END[3]),
    .I3(E2END[1]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q ),
    .Z(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2296_ (.I0(_0909_),
    .I1(_0908_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit2.Q ),
    .Z(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2297_ (.I0(_0910_),
    .I1(_0907_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame4_bit3.Q ),
    .Z(\Inst_RegFile_switch_matrix.JN2BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2298_ (.I0(NN4END[2]),
    .I1(E1END[2]),
    .I2(SS4END[2]),
    .I3(W1END[2]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q ),
    .Z(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2299_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit18.Q ),
    .A2(_0911_),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2300_ (.I0(AD0),
    .I1(AD2),
    .I2(AD1),
    .I3(AD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q ),
    .Z(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2301_ (.A1(_0136_),
    .A2(_0913_),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2302_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q ),
    .A2(_0497_),
    .ZN(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2303_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q ),
    .A2(_0212_),
    .B(_0915_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q ),
    .ZN(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2304_ (.I0(N2MID[4]),
    .I1(E2MID[4]),
    .S(\Inst_RegFile_ConfigMem.Inst_frame7_bit4.Q ),
    .Z(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2305_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame7_bit4.Q ),
    .A2(\Inst_RegFile_switch_matrix.JS2BEG3 ),
    .ZN(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2306_ (.A1(_1267_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame7_bit4.Q ),
    .B(\Inst_RegFile_ConfigMem.Inst_frame7_bit5.Q ),
    .C(_0918_),
    .ZN(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2307_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame7_bit5.Q ),
    .A2(_0917_),
    .B(_0919_),
    .ZN(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2308_ (.I(_0920_),
    .ZN(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2309_ (.I0(N2MID[4]),
    .I1(S2MID[4]),
    .I2(E2MID[4]),
    .I3(\Inst_RegFile_switch_matrix.JS2BEG4 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit13.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit12.Q ),
    .Z(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2310_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q ),
    .A2(_0922_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q ),
    .ZN(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2311_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q ),
    .A2(_0920_),
    .B(_0923_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2312_ (.A1(_0916_),
    .A2(_0924_),
    .B(_0136_),
    .ZN(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2313_ (.I0(BD0),
    .I1(BD2),
    .I2(BD1),
    .I3(BD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q ),
    .Z(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2314_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit18.Q ),
    .A2(_0926_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame9_bit19.Q ),
    .ZN(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2315_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit19.Q ),
    .A2(_0912_),
    .A3(_0914_),
    .B1(_0925_),
    .B2(_0927_),
    .ZN(\Inst_RegFile_switch_matrix.W6BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2316_ (.I0(NN4END[1]),
    .I1(E1END[3]),
    .I2(SS4END[1]),
    .I3(W1END[3]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q ),
    .Z(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2317_ (.I0(AD0),
    .I1(AD2),
    .I2(AD1),
    .I3(AD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q ),
    .Z(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2318_ (.I0(N2MID[3]),
    .I1(E2MID[3]),
    .I2(S2MID[3]),
    .I3(W2MID[3]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit10.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit11.Q ),
    .Z(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2319_ (.I(_0930_),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2320_ (.I0(N2MID[3]),
    .I1(E2MID[3]),
    .S(\Inst_RegFile_ConfigMem.Inst_frame6_bit2.Q ),
    .Z(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2321_ (.A1(W2MID[3]),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame6_bit2.Q ),
    .ZN(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2322_ (.A1(_1259_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame6_bit2.Q ),
    .B(\Inst_RegFile_ConfigMem.Inst_frame6_bit3.Q ),
    .C(_0933_),
    .ZN(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2323_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame6_bit3.Q ),
    .A2(_0932_),
    .B(_0934_),
    .ZN(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2324_ (.I(_0935_),
    .ZN(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2325_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q ),
    .A2(_0935_),
    .ZN(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2326_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q ),
    .A2(_0930_),
    .B(_0937_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q ),
    .ZN(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2327_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q ),
    .A2(_0160_),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2328_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q ),
    .A2(_0468_),
    .B(_0939_),
    .ZN(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2329_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q ),
    .A2(_0940_),
    .B(_0938_),
    .ZN(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2330_ (.I0(BD0),
    .I1(BD2),
    .I2(BD1),
    .I3(BD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q ),
    .Z(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2331_ (.I0(_0928_),
    .I1(_0929_),
    .I2(_0942_),
    .I3(_0941_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit14.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit15.Q ),
    .Z(\Inst_RegFile_switch_matrix.W6BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2332_ (.I0(N2END[4]),
    .I1(S2END[4]),
    .I2(EE4END[0]),
    .I3(W2END[4]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit5.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit4.Q ),
    .Z(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2333_ (.I0(BD0),
    .I1(_0213_),
    .I2(_0497_),
    .I3(_0943_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit9.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit10.Q ),
    .Z(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2334_ (.I0(N1END[1]),
    .I1(S1END[1]),
    .I2(W1END[1]),
    .I3(AD0),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit9.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit10.Q ),
    .Z(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2335_ (.I0(_0945_),
    .I1(_0944_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit11.Q ),
    .Z(\Inst_RegFile_switch_matrix.WW4BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2336_ (.I0(N2END[4]),
    .I1(E2END[4]),
    .I2(SS4END[2]),
    .I3(W2END[4]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit13.Q ),
    .Z(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2337_ (.I0(_0468_),
    .I1(_0946_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q ),
    .Z(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2338_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q ),
    .A2(BD3),
    .ZN(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2339_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q ),
    .A2(_0160_),
    .B(_0948_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame9_bit7.Q ),
    .ZN(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2340_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit7.Q ),
    .A2(_0947_),
    .B(_0949_),
    .ZN(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2341_ (.I0(N1END[0]),
    .I1(S1END[0]),
    .I2(W1END[0]),
    .I3(AD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit7.Q ),
    .Z(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2342_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit8.Q ),
    .A2(_0951_),
    .ZN(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2343_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit8.Q ),
    .A2(_0950_),
    .B(_0952_),
    .ZN(\Inst_RegFile_switch_matrix.WW4BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2344_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit3.Q ),
    .A2(_0920_),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2345_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit3.Q ),
    .A2(BD2),
    .B(_0953_),
    .ZN(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2346_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit3.Q ),
    .A2(_0198_),
    .ZN(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2347_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit3.Q ),
    .A2(_0922_),
    .B(_0955_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame9_bit4.Q ),
    .ZN(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2348_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit4.Q ),
    .A2(_0954_),
    .B(_0956_),
    .ZN(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2349_ (.I0(N1END[3]),
    .I1(S1END[3]),
    .I2(W1END[3]),
    .I3(AD2),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit3.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit4.Q ),
    .Z(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2350_ (.I0(_0958_),
    .I1(_0957_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit5.Q ),
    .Z(\Inst_RegFile_switch_matrix.WW4BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2351_ (.I0(BD1),
    .I1(_0930_),
    .I2(_0936_),
    .I3(_0514_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit1.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit0.Q ),
    .Z(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2352_ (.I0(N1END[2]),
    .I1(S1END[2]),
    .I2(W1END[2]),
    .I3(AD1),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit0.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit1.Q ),
    .Z(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2353_ (.I0(_0960_),
    .I1(_0959_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame9_bit2.Q ),
    .Z(\Inst_RegFile_switch_matrix.WW4BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2354_ (.I0(N2END[0]),
    .I1(S2END[0]),
    .I2(E2END[0]),
    .I3(WW4END[3]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit7.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit6.Q ),
    .Z(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2355_ (.I0(BD0),
    .I1(_0213_),
    .I2(_0497_),
    .I3(_0961_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit21.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit22.Q ),
    .Z(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2356_ (.I0(N1END[1]),
    .I1(E1END[1]),
    .I2(W1END[1]),
    .I3(AD0),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit21.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit22.Q ),
    .Z(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2357_ (.I0(_0963_),
    .I1(_0962_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame10_bit23.Q ),
    .Z(\Inst_RegFile_switch_matrix.SS4BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2358_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q ),
    .A2(_0272_),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2359_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q ),
    .A2(_0468_),
    .B(_0964_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame10_bit19.Q ),
    .ZN(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2360_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q ),
    .A2(_0160_),
    .ZN(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2361_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q ),
    .A2(BD3),
    .B(_0966_),
    .ZN(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2362_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit19.Q ),
    .A2(_0967_),
    .B(_0965_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame10_bit20.Q ),
    .ZN(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2363_ (.I0(N1END[0]),
    .I1(E1END[0]),
    .I2(W1END[0]),
    .I3(AD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit19.Q ),
    .Z(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2364_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit20.Q ),
    .A2(_0969_),
    .B(_0968_),
    .ZN(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2365_ (.I(_0970_),
    .ZN(\Inst_RegFile_switch_matrix.SS4BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2366_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q ),
    .A2(_0920_),
    .ZN(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2367_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q ),
    .A2(BD2),
    .B(_0971_),
    .ZN(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2368_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q ),
    .A2(_0238_),
    .ZN(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2369_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q ),
    .A2(_0922_),
    .B(_0973_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame10_bit16.Q ),
    .ZN(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2370_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit16.Q ),
    .A2(_0972_),
    .B(_0974_),
    .ZN(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2371_ (.I0(N1END[3]),
    .I1(E1END[3]),
    .I2(W1END[3]),
    .I3(AD2),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit16.Q ),
    .Z(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2372_ (.I0(_0976_),
    .I1(_0975_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame10_bit17.Q ),
    .Z(\Inst_RegFile_switch_matrix.SS4BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2373_ (.I0(BD1),
    .I1(_0930_),
    .I2(_0936_),
    .I3(_0531_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit13.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit12.Q ),
    .Z(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2374_ (.I0(N1END[2]),
    .I1(E1END[2]),
    .I2(W1END[2]),
    .I3(AD1),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit13.Q ),
    .Z(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2375_ (.I0(_0978_),
    .I1(_0977_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame10_bit14.Q ),
    .Z(\Inst_RegFile_switch_matrix.SS4BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2376_ (.I0(NN4END[3]),
    .I1(SS4END[3]),
    .I2(E1END[2]),
    .I3(W1END[2]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q ),
    .Z(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2377_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit26.Q ),
    .A2(_0979_),
    .ZN(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2378_ (.I0(AD0),
    .I1(AD2),
    .I2(AD1),
    .I3(AD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q ),
    .Z(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2379_ (.A1(_0137_),
    .A2(_0981_),
    .ZN(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2380_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q ),
    .A2(_0497_),
    .ZN(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2381_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q ),
    .A2(_0212_),
    .B(_0983_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q ),
    .ZN(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2382_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q ),
    .A2(_0922_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q ),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2383_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q ),
    .A2(_0920_),
    .B(_0985_),
    .ZN(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2384_ (.A1(_0984_),
    .A2(_0986_),
    .B(_0137_),
    .ZN(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2385_ (.I0(BD0),
    .I1(BD2),
    .I2(BD1),
    .I3(BD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q ),
    .Z(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2386_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit26.Q ),
    .A2(_0988_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame11_bit27.Q ),
    .ZN(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2387_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit27.Q ),
    .A2(_0980_),
    .A3(_0982_),
    .B1(_0987_),
    .B2(_0989_),
    .ZN(\Inst_RegFile_switch_matrix.E6BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2388_ (.I0(NN4END[0]),
    .I1(SS4END[0]),
    .I2(E1END[3]),
    .I3(W1END[3]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q ),
    .Z(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2389_ (.I0(AD0),
    .I1(AD2),
    .I2(AD1),
    .I3(AD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q ),
    .Z(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2390_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q ),
    .A2(_0935_),
    .ZN(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2391_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q ),
    .A2(_0930_),
    .B(_0992_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q ),
    .ZN(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2392_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q ),
    .A2(_0160_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q ),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2393_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q ),
    .A2(_0468_),
    .B(_0994_),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2394_ (.A1(_0993_),
    .A2(_0995_),
    .ZN(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2395_ (.I0(BD0),
    .I1(BD2),
    .I2(BD1),
    .I3(BD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q ),
    .Z(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2396_ (.I0(_0990_),
    .I1(_0991_),
    .I2(_0997_),
    .I3(_0996_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit22.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit23.Q ),
    .Z(\Inst_RegFile_switch_matrix.E6BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2397_ (.I0(N2END[6]),
    .I1(E2END[6]),
    .I2(SS4END[3]),
    .I3(W2END[6]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit0.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit1.Q ),
    .Z(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2398_ (.I0(BD0),
    .I1(_0213_),
    .I2(_0497_),
    .I3(_0998_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit17.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit18.Q ),
    .Z(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2399_ (.I0(N1END[1]),
    .I1(E1END[1]),
    .I2(S1END[1]),
    .I3(AD0),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit17.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit18.Q ),
    .Z(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2400_ (.I0(_1000_),
    .I1(_0999_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame11_bit19.Q ),
    .Z(\Inst_RegFile_switch_matrix.EE4BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2401_ (.I0(NN4END[3]),
    .I1(E2END[6]),
    .I2(S2END[6]),
    .I3(W2END[6]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit9.Q ),
    .Z(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2402_ (.I0(_0468_),
    .I1(_1001_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q ),
    .Z(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2403_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q ),
    .A2(BD3),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2404_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q ),
    .A2(_0160_),
    .B(_1003_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q ),
    .ZN(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2405_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q ),
    .A2(_1002_),
    .B(_1004_),
    .ZN(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2406_ (.I0(N1END[0]),
    .I1(E1END[0]),
    .I2(S1END[0]),
    .I3(AD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q ),
    .Z(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2407_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit16.Q ),
    .A2(_1006_),
    .ZN(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2408_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit16.Q ),
    .A2(_1005_),
    .B(_1007_),
    .ZN(\Inst_RegFile_switch_matrix.EE4BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2409_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q ),
    .A2(_0920_),
    .ZN(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2410_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q ),
    .A2(BD2),
    .B(_1008_),
    .ZN(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2411_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q ),
    .A2(_0784_),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2412_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q ),
    .A2(_0922_),
    .B(_1010_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame11_bit12.Q ),
    .ZN(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2413_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit12.Q ),
    .A2(_1009_),
    .B(_1011_),
    .ZN(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2414_ (.I0(N1END[3]),
    .I1(E1END[3]),
    .I2(S1END[3]),
    .I3(AD2),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit12.Q ),
    .Z(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2415_ (.I0(_1013_),
    .I1(_1012_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame11_bit13.Q ),
    .Z(\Inst_RegFile_switch_matrix.EE4BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2416_ (.I0(BD1),
    .I1(_0930_),
    .I2(_0936_),
    .I3(_0766_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit9.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit8.Q ),
    .Z(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2417_ (.I0(N1END[2]),
    .I1(E1END[2]),
    .I2(S1END[2]),
    .I3(AD1),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit9.Q ),
    .Z(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2418_ (.I0(_1015_),
    .I1(_1014_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame11_bit10.Q ),
    .Z(\Inst_RegFile_switch_matrix.EE4BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2419_ (.I0(NN4END[0]),
    .I1(S2END[2]),
    .I2(E2END[2]),
    .I3(W2END[2]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit3.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit2.Q ),
    .Z(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2420_ (.I0(BD0),
    .I1(_0213_),
    .I2(_0497_),
    .I3(_1016_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit29.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit30.Q ),
    .Z(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2421_ (.I0(N1END[1]),
    .I1(E1END[1]),
    .I2(W1END[1]),
    .I3(AD0),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit29.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit30.Q ),
    .Z(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2422_ (.I0(_1018_),
    .I1(_1017_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit31.Q ),
    .Z(\Inst_RegFile_switch_matrix.NN4BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2423_ (.I0(N2END[2]),
    .I1(S2END[2]),
    .I2(E2END[2]),
    .I3(WW4END[2]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame5_bit11.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame5_bit10.Q ),
    .Z(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2424_ (.I0(_0468_),
    .I1(_1019_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q ),
    .Z(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2425_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q ),
    .A2(BD3),
    .ZN(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2426_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q ),
    .A2(_0160_),
    .B(_1021_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame12_bit27.Q ),
    .ZN(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2427_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit27.Q ),
    .A2(_1020_),
    .B(_1022_),
    .ZN(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2428_ (.I0(N1END[0]),
    .I1(E1END[0]),
    .I2(W1END[0]),
    .I3(AD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit27.Q ),
    .Z(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2429_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit28.Q ),
    .A2(_1024_),
    .ZN(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2430_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit28.Q ),
    .A2(_1023_),
    .B(_1025_),
    .ZN(\Inst_RegFile_switch_matrix.NN4BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2431_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q ),
    .A2(_0920_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame12_bit24.Q ),
    .ZN(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2432_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q ),
    .A2(BD2),
    .B(_1026_),
    .ZN(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2433_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q ),
    .A2(_0178_),
    .ZN(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2434_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q ),
    .A2(_0922_),
    .B(_1028_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame12_bit24.Q ),
    .ZN(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2435_ (.A1(_1027_),
    .A2(_1029_),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2436_ (.I0(N1END[3]),
    .I1(E1END[3]),
    .I2(W1END[3]),
    .I3(AD2),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit24.Q ),
    .Z(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2437_ (.I0(_1031_),
    .I1(_1030_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit25.Q ),
    .Z(\Inst_RegFile_switch_matrix.NN4BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2438_ (.I0(_0930_),
    .I1(_0484_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q ),
    .Z(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2439_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q ),
    .A2(BD1),
    .ZN(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2440_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q ),
    .A2(_0935_),
    .B(_1033_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame12_bit21.Q ),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2441_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit21.Q ),
    .A2(_1032_),
    .B(_1034_),
    .ZN(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2442_ (.I0(N1END[2]),
    .I1(E1END[2]),
    .I2(W1END[2]),
    .I3(AD1),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit21.Q ),
    .Z(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2443_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit22.Q ),
    .A2(_1036_),
    .ZN(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2444_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit22.Q ),
    .A2(_1035_),
    .B(_1037_),
    .ZN(\Inst_RegFile_switch_matrix.NN4BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2445_ (.I0(NN4END[3]),
    .I1(S4END[3]),
    .S(\Inst_RegFile_ConfigMem.Inst_frame0_bit0.Q ),
    .Z(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2446_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit0.Q ),
    .A2(\Inst_RegFile_switch_matrix.JN2BEG1 ),
    .ZN(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2447_ (.A1(_1250_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame0_bit0.Q ),
    .B(\Inst_RegFile_ConfigMem.Inst_frame0_bit1.Q ),
    .C(_1039_),
    .ZN(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2448_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit1.Q ),
    .A2(_1038_),
    .B(_1040_),
    .ZN(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2449_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit30.Q ),
    .A2(_1041_),
    .ZN(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2450_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit30.Q ),
    .A2(\Inst_RegFile_switch_matrix.JS2BEG2 ),
    .B(_1042_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame10_bit31.Q ),
    .ZN(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2451_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit30.Q ),
    .A2(_0573_),
    .ZN(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2452_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit30.Q ),
    .A2(AD0),
    .B(_1044_),
    .ZN(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2453_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit31.Q ),
    .A2(_1045_),
    .B(_1043_),
    .ZN(\Inst_RegFile_switch_matrix.W1BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2454_ (.I0(BD3),
    .I1(_0468_),
    .I2(\Inst_RegFile_switch_matrix.JS2BEG1 ),
    .I3(_0530_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit28.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit29.Q ),
    .Z(\Inst_RegFile_switch_matrix.W1BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2455_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit26.Q ),
    .A2(_0789_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame10_bit27.Q ),
    .ZN(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2456_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit26.Q ),
    .A2(BD2),
    .B(_1046_),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2457_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit26.Q ),
    .A2(_0195_),
    .ZN(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2458_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit26.Q ),
    .A2(\Inst_RegFile_switch_matrix.JS2BEG0 ),
    .B(_1048_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame10_bit27.Q ),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2459_ (.A1(_1047_),
    .A2(_1049_),
    .ZN(\Inst_RegFile_switch_matrix.W1BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2460_ (.I0(N4END[2]),
    .I1(E2END[2]),
    .S(\Inst_RegFile_ConfigMem.Inst_frame0_bit10.Q ),
    .Z(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2461_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit10.Q ),
    .A2(\Inst_RegFile_switch_matrix.E2BEG2 ),
    .Z(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2462_ (.A1(_1342_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame0_bit10.Q ),
    .B(\Inst_RegFile_ConfigMem.Inst_frame0_bit11.Q ),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2463_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit11.Q ),
    .A2(_1050_),
    .B1(_1051_),
    .B2(_1052_),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2464_ (.A1(_1278_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame6_bit14.Q ),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2465_ (.A1(W2MID[1]),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame6_bit14.Q ),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2466_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame6_bit15.Q ),
    .A2(_1055_),
    .ZN(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2467_ (.I0(N2MID[1]),
    .I1(E2MID[1]),
    .S(\Inst_RegFile_ConfigMem.Inst_frame6_bit14.Q ),
    .Z(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2468_ (.A1(_1054_),
    .A2(_1056_),
    .B1(_1057_),
    .B2(\Inst_RegFile_ConfigMem.Inst_frame6_bit15.Q ),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2469_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit24.Q ),
    .A2(_1058_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame10_bit25.Q ),
    .ZN(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2470_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit24.Q ),
    .A2(BD1),
    .B(_1059_),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2471_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit24.Q ),
    .A2(_1053_),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2472_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit24.Q ),
    .A2(\Inst_RegFile_switch_matrix.JS2BEG3 ),
    .B(_1061_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame10_bit25.Q ),
    .ZN(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2473_ (.A1(_1060_),
    .A2(_1062_),
    .ZN(\Inst_RegFile_switch_matrix.W1BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2474_ (.I0(S2END[1]),
    .I1(W6END[0]),
    .I2(S4END[0]),
    .I3(AD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit11.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit10.Q ),
    .Z(\Inst_RegFile_switch_matrix.S4BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2475_ (.I0(S2END[0]),
    .I1(W6END[1]),
    .I2(S4END[3]),
    .I3(AD2),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit9.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit8.Q ),
    .Z(\Inst_RegFile_switch_matrix.S4BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2476_ (.I0(E6END[0]),
    .I1(S2END[3]),
    .I2(S4END[2]),
    .I3(AD1),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit6.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit7.Q ),
    .Z(\Inst_RegFile_switch_matrix.S4BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2477_ (.I0(E6END[1]),
    .I1(S4END[1]),
    .I2(S2END[2]),
    .I3(AD0),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit5.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit4.Q ),
    .Z(\Inst_RegFile_switch_matrix.S4BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2478_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit2.Q ),
    .A2(_0573_),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2479_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit2.Q ),
    .A2(BD3),
    .B(_1063_),
    .C(_0139_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2480_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit2.Q ),
    .A2(_1041_),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2481_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame10_bit2.Q ),
    .A2(\Inst_RegFile_switch_matrix.E2BEG2 ),
    .B(_1065_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame10_bit3.Q ),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2482_ (.A1(_1064_),
    .A2(_1066_),
    .ZN(\Inst_RegFile_switch_matrix.S1BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2483_ (.I0(BD2),
    .I1(_0468_),
    .I2(\Inst_RegFile_switch_matrix.E2BEG1 ),
    .I3(_0530_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame10_bit0.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame10_bit1.Q ),
    .Z(\Inst_RegFile_switch_matrix.S1BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2484_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit30.Q ),
    .A2(_0195_),
    .ZN(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2485_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit30.Q ),
    .A2(\Inst_RegFile_switch_matrix.E2BEG0 ),
    .B(_1067_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame11_bit31.Q ),
    .ZN(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2486_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit30.Q ),
    .A2(_0789_),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2487_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit30.Q ),
    .A2(BD1),
    .B(_1069_),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2488_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit31.Q ),
    .A2(_1070_),
    .B(_1068_),
    .ZN(\Inst_RegFile_switch_matrix.S1BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2489_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit28.Q ),
    .A2(_1058_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame11_bit29.Q ),
    .ZN(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2490_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit28.Q ),
    .A2(BD0),
    .B(_1071_),
    .ZN(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2491_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit28.Q ),
    .A2(_1053_),
    .ZN(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2492_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit28.Q ),
    .A2(\Inst_RegFile_switch_matrix.E2BEG3 ),
    .B(_1073_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame11_bit29.Q ),
    .ZN(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2493_ (.A1(_1072_),
    .A2(_1074_),
    .ZN(\Inst_RegFile_switch_matrix.S1BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2494_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit6.Q ),
    .A2(_1041_),
    .ZN(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2495_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit6.Q ),
    .A2(\Inst_RegFile_switch_matrix.JN2BEG2 ),
    .B(_1075_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame11_bit7.Q ),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2496_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit6.Q ),
    .A2(_0573_),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2497_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit6.Q ),
    .A2(BD2),
    .B(_1077_),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2498_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit7.Q ),
    .A2(_1078_),
    .B(_1076_),
    .ZN(\Inst_RegFile_switch_matrix.E1BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2499_ (.I0(BD1),
    .I1(_0468_),
    .I2(\Inst_RegFile_switch_matrix.JN2BEG1 ),
    .I3(_0530_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame11_bit4.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame11_bit5.Q ),
    .Z(\Inst_RegFile_switch_matrix.E1BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2500_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit2.Q ),
    .A2(_0789_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame11_bit3.Q ),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2501_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit2.Q ),
    .A2(BD0),
    .B(_1079_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2502_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit2.Q ),
    .A2(_0195_),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2503_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit2.Q ),
    .A2(\Inst_RegFile_switch_matrix.JN2BEG0 ),
    .B(_1081_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame11_bit3.Q ),
    .ZN(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2504_ (.A1(_1080_),
    .A2(_1082_),
    .ZN(\Inst_RegFile_switch_matrix.E1BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2505_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit0.Q ),
    .A2(_1058_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame11_bit1.Q ),
    .ZN(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2506_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit0.Q ),
    .A2(AD3),
    .B(_1083_),
    .ZN(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2507_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit0.Q ),
    .A2(_1053_),
    .ZN(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2508_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame11_bit0.Q ),
    .A2(\Inst_RegFile_switch_matrix.JN2BEG3 ),
    .B(_1085_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame11_bit1.Q ),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2509_ (.A1(_1084_),
    .A2(_1086_),
    .ZN(\Inst_RegFile_switch_matrix.E1BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2510_ (.I0(N2END[1]),
    .I1(N4END[0]),
    .I2(W6END[0]),
    .I3(BD3),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit18.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit19.Q ),
    .Z(\Inst_RegFile_switch_matrix.N4BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2511_ (.I0(N2END[0]),
    .I1(W6END[1]),
    .I2(N4END[3]),
    .I3(BD2),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit17.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit16.Q ),
    .Z(\Inst_RegFile_switch_matrix.N4BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2512_ (.I0(N2END[3]),
    .I1(N4END[2]),
    .I2(E6END[0]),
    .I3(BD1),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit14.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit15.Q ),
    .Z(\Inst_RegFile_switch_matrix.N4BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2513_ (.I0(N2END[2]),
    .I1(N4END[1]),
    .I2(E6END[1]),
    .I3(BD0),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit13.Q ),
    .Z(\Inst_RegFile_switch_matrix.N4BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2514_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit10.Q ),
    .A2(_1041_),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2515_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit10.Q ),
    .A2(\Inst_RegFile_switch_matrix.JW2BEG2 ),
    .B(_1087_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame12_bit11.Q ),
    .ZN(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2516_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit10.Q ),
    .A2(_0573_),
    .ZN(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2517_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit10.Q ),
    .A2(BD1),
    .B(_1089_),
    .ZN(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2518_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit11.Q ),
    .A2(_1090_),
    .B(_1088_),
    .ZN(\Inst_RegFile_switch_matrix.N1BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2519_ (.I0(BD0),
    .I1(_0468_),
    .I2(\Inst_RegFile_switch_matrix.JW2BEG1 ),
    .I3(_0530_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame12_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame12_bit9.Q ),
    .Z(\Inst_RegFile_switch_matrix.N1BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2520_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit6.Q ),
    .A2(\Inst_RegFile_switch_matrix.JW2BEG0 ),
    .ZN(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2521_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit6.Q ),
    .A2(_0195_),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2522_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit7.Q ),
    .A2(_1092_),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2523_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit6.Q ),
    .A2(_0789_),
    .ZN(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2524_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit6.Q ),
    .A2(AD3),
    .B(_1094_),
    .ZN(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2525_ (.A1(_1091_),
    .A2(_1093_),
    .B1(_1095_),
    .B2(\Inst_RegFile_ConfigMem.Inst_frame12_bit7.Q ),
    .ZN(\Inst_RegFile_switch_matrix.N1BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2526_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit4.Q ),
    .A2(_1058_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame12_bit5.Q ),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2527_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit4.Q ),
    .A2(AD2),
    .B(_1096_),
    .ZN(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2528_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit4.Q ),
    .A2(_1053_),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2529_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame12_bit4.Q ),
    .A2(\Inst_RegFile_switch_matrix.JW2BEG3 ),
    .B(_1098_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame12_bit5.Q ),
    .ZN(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2530_ (.A1(_1097_),
    .A2(_1099_),
    .ZN(\Inst_RegFile_switch_matrix.N1BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2531_ (.I0(_0961_),
    .I1(\Inst_RegFile_switch_matrix.JN2BEG7 ),
    .I2(\Inst_RegFile_switch_matrix.JS2BEG7 ),
    .I3(\Inst_RegFile_switch_matrix.JW2BEG7 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame8_bit4.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame8_bit5.Q ),
    .Z(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2532_ (.I(_1100_),
    .ZN(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2533_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit4.Q ),
    .A2(_0215_),
    .ZN(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2534_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit4.Q ),
    .A2(_0156_),
    .B(_1102_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame8_bit5.Q ),
    .ZN(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2535_ (.A1(N2END[0]),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame8_bit4.Q ),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2536_ (.A1(_1353_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame8_bit4.Q ),
    .B(\Inst_RegFile_ConfigMem.Inst_frame8_bit5.Q ),
    .C(_1104_),
    .ZN(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2537_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit6.Q ),
    .A2(_1105_),
    .ZN(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2538_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit6.Q ),
    .A2(_1101_),
    .B1(_1103_),
    .B2(_1106_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2539_ (.A1(_1290_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame0_bit14.Q ),
    .B(\Inst_RegFile_ConfigMem.Inst_frame0_bit15.Q ),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2540_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit14.Q ),
    .A2(\Inst_RegFile_switch_matrix.JW2BEG2 ),
    .B(_1108_),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2541_ (.I0(N4END[0]),
    .I1(SS4END[0]),
    .S(\Inst_RegFile_ConfigMem.Inst_frame0_bit14.Q ),
    .Z(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2542_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit15.Q ),
    .A2(_1110_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame8_bit2.Q ),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2543_ (.A1(_1109_),
    .A2(_1111_),
    .Z(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2544_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit2.Q ),
    .A2(_0272_),
    .Z(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2545_ (.I0(N2MID[0]),
    .I1(W2MID[0]),
    .I2(S2MID[0]),
    .I3(\Inst_RegFile_switch_matrix.JW2BEG4 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit15.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit14.Q ),
    .Z(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2546_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit3.Q ),
    .A2(_1113_),
    .Z(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2547_ (.A1(_1109_),
    .A2(_1111_),
    .B(_1113_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame8_bit3.Q ),
    .ZN(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2548_ (.A1(_0144_),
    .A2(_1114_),
    .Z(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2549_ (.A1(_0144_),
    .A2(_1058_),
    .ZN(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2550_ (.A1(_0144_),
    .A2(_1114_),
    .B(_1118_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame8_bit3.Q ),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2551_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit3.Q ),
    .A2(_1117_),
    .A3(_1118_),
    .B(_1116_),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2552_ (.A1(_1112_),
    .A2(_1115_),
    .B(_1119_),
    .ZN(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2553_ (.A1(_1107_),
    .A2(_1121_),
    .Z(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2554_ (.I0(N2MID[5]),
    .I1(E2MID[5]),
    .I2(S2MID[5]),
    .I3(W2MID[5]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit12.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit13.Q ),
    .Z(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2555_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit0.Q ),
    .A2(_1123_),
    .Z(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2556_ (.A1(_0142_),
    .A2(_0922_),
    .B(_1124_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q ),
    .ZN(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2557_ (.A1(_0143_),
    .A2(\Inst_RegFile_switch_matrix.JS2BEG2 ),
    .ZN(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2558_ (.A1(S4END[1]),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame0_bit12.Q ),
    .B(\Inst_RegFile_ConfigMem.Inst_frame0_bit13.Q ),
    .ZN(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2559_ (.A1(_1255_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame0_bit12.Q ),
    .ZN(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2560_ (.A1(NN4END[1]),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame0_bit12.Q ),
    .B(_1128_),
    .ZN(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2561_ (.A1(_1126_),
    .A2(_1127_),
    .B1(_1129_),
    .B2(\Inst_RegFile_ConfigMem.Inst_frame0_bit13.Q ),
    .C(\Inst_RegFile_ConfigMem.Inst_frame8_bit0.Q ),
    .ZN(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2562_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit0.Q ),
    .A2(_0946_),
    .B(_1130_),
    .ZN(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2563_ (.A1(_0142_),
    .A2(_0922_),
    .B(_1124_),
    .ZN(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2564_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q ),
    .A2(_1131_),
    .B(_1125_),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2565_ (.I0(_1132_),
    .I1(_1131_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q ),
    .Z(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2566_ (.A1(_1122_),
    .A2(_1134_),
    .ZN(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2567_ (.I0(N2MID[2]),
    .I1(W2MID[2]),
    .I2(E2MID[2]),
    .I3(\Inst_RegFile_switch_matrix.E2BEG4 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit11.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit10.Q ),
    .Z(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2568_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit30.Q ),
    .A2(_1136_),
    .ZN(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2569_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit30.Q ),
    .A2(_0931_),
    .B(_1137_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q ),
    .ZN(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2570_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit30.Q ),
    .A2(_1019_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q ),
    .ZN(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2571_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit30.Q ),
    .A2(_1053_),
    .B(_1139_),
    .ZN(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2572_ (.A1(_1138_),
    .A2(_1140_),
    .Z(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2573_ (.A1(_1138_),
    .A2(_1140_),
    .ZN(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2574_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q ),
    .A2(\Inst_RegFile_switch_matrix.JW2BEG0 ),
    .ZN(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2575_ (.A1(_0145_),
    .A2(\Inst_RegFile_switch_matrix.JS2BEG0 ),
    .B(_0146_),
    .ZN(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2576_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q ),
    .A2(\Inst_RegFile_switch_matrix.JN2BEG0 ),
    .ZN(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2577_ (.A1(_0145_),
    .A2(_0531_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame8_bit8.Q ),
    .ZN(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2578_ (.A1(_1143_),
    .A2(_1144_),
    .B1(_1145_),
    .B2(_1146_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2579_ (.I0(N2END[3]),
    .I1(S2END[3]),
    .I2(_1136_),
    .I3(_1123_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame8_bit8.Q ),
    .Z(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2580_ (.I0(_1148_),
    .I1(_1147_),
    .S(\Inst_RegFile_ConfigMem.Inst_frame8_bit9.Q ),
    .Z(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2581_ (.A1(_0816_),
    .A2(_0818_),
    .B1(_0820_),
    .B2(_0822_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame0_bit8.Q ),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2582_ (.A1(WW4END[2]),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame0_bit8.Q ),
    .B(\Inst_RegFile_ConfigMem.Inst_frame0_bit9.Q ),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2583_ (.I(_1151_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2584_ (.A1(E2END[3]),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame0_bit8.Q ),
    .ZN(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2585_ (.A1(_1269_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame0_bit8.Q ),
    .B(\Inst_RegFile_ConfigMem.Inst_frame0_bit9.Q ),
    .C(_1153_),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2586_ (.A1(_1150_),
    .A2(_1152_),
    .B(_1154_),
    .C(_0141_),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2587_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q ),
    .A2(_1001_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame9_bit29.Q ),
    .ZN(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2588_ (.A1(_1155_),
    .A2(_1156_),
    .ZN(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2589_ (.A1(_0140_),
    .A2(\Inst_RegFile_switch_matrix.JN2BEG4 ),
    .ZN(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2590_ (.A1(W2MID[6]),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame7_bit8.Q ),
    .B(\Inst_RegFile_ConfigMem.Inst_frame7_bit9.Q ),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2591_ (.I0(W2MID[6]),
    .I1(\Inst_RegFile_switch_matrix.JN2BEG4 ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame7_bit8.Q ),
    .Z(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2592_ (.A1(S2MID[6]),
    .A2(_0140_),
    .ZN(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2593_ (.A1(_1247_),
    .A2(_0140_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame7_bit9.Q ),
    .C(_1161_),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2594_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q ),
    .A2(_1162_),
    .ZN(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2595_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame7_bit9.Q ),
    .A2(_1160_),
    .B(_1162_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q ),
    .ZN(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2596_ (.A1(_1158_),
    .A2(_1159_),
    .B(_1163_),
    .ZN(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2597_ (.I0(N2MID[7]),
    .I1(E2MID[7]),
    .I2(S2MID[7]),
    .I3(W2MID[7]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit8.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit9.Q ),
    .Z(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2598_ (.A1(_0141_),
    .A2(_1166_),
    .ZN(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2599_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit29.Q ),
    .A2(_1167_),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2600_ (.A1(_1165_),
    .A2(_1168_),
    .B(_1157_),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2601_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit29.Q ),
    .A2(_1164_),
    .A3(_1167_),
    .B1(_1155_),
    .B2(_1156_),
    .ZN(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2602_ (.A1(_1149_),
    .A2(_1169_),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2603_ (.A1(_1141_),
    .A2(_1171_),
    .ZN(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2604_ (.A1(_1142_),
    .A2(_1149_),
    .A3(_1169_),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2605_ (.A1(_1135_),
    .A2(_1173_),
    .ZN(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2606_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit20.Q ),
    .A2(_1041_),
    .ZN(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2607_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit20.Q ),
    .A2(_0998_),
    .B(_1175_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame9_bit21.Q ),
    .ZN(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2608_ (.I0(N2MID[6]),
    .I1(S2MID[6]),
    .I2(W2MID[6]),
    .I3(\Inst_RegFile_switch_matrix.JN2BEG3 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame7_bit0.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame7_bit1.Q ),
    .Z(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2609_ (.I0(N2MID[7]),
    .I1(E2MID[7]),
    .I2(S2MID[7]),
    .I3(W2MID[7]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit0.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit1.Q ),
    .Z(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2610_ (.I(_1178_),
    .ZN(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2611_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit20.Q ),
    .A2(_1179_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame9_bit21.Q ),
    .ZN(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2612_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit20.Q ),
    .A2(_1177_),
    .B(_1180_),
    .ZN(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2613_ (.A1(_1176_),
    .A2(_1181_),
    .ZN(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2614_ (.I0(\Inst_RegFile_32x4.mem[24][0] ),
    .I1(_1182_),
    .S(_1174_),
    .Z(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2615_ (.I0(EE4END[2]),
    .I1(W2END[7]),
    .I2(S4END[2]),
    .I3(\Inst_RegFile_switch_matrix.E2BEG1 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame0_bit3.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame0_bit2.Q ),
    .Z(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2616_ (.I0(_0570_),
    .I1(_0936_),
    .I2(_1016_),
    .I3(_1183_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit22.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit23.Q ),
    .Z(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2617_ (.I0(\Inst_RegFile_32x4.mem[24][1] ),
    .I1(_1184_),
    .S(_1174_),
    .Z(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2618_ (.I0(N4END[1]),
    .I1(W6END[1]),
    .I2(E6END[1]),
    .I3(\Inst_RegFile_switch_matrix.JS2BEG1 ),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame0_bit5.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame0_bit4.Q ),
    .Z(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2619_ (.I0(_0921_),
    .I1(_0943_),
    .I2(_0572_),
    .I3(_1185_),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame9_bit25.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame9_bit24.Q ),
    .Z(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2620_ (.I0(\Inst_RegFile_32x4.mem[24][2] ),
    .I1(_1186_),
    .S(_1174_),
    .Z(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2621_ (.I0(S4END[0]),
    .I1(\Inst_RegFile_switch_matrix.JW2BEG1 ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame0_bit6.Q ),
    .Z(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2622_ (.A1(N4END[0]),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame0_bit6.Q ),
    .ZN(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2623_ (.A1(_1280_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame0_bit6.Q ),
    .B(\Inst_RegFile_ConfigMem.Inst_frame0_bit7.Q ),
    .C(_1188_),
    .ZN(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2624_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame0_bit7.Q ),
    .A2(_1187_),
    .B(_1189_),
    .C(_0138_),
    .ZN(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2625_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q ),
    .A2(_0961_),
    .B(\Inst_RegFile_ConfigMem.Inst_frame9_bit27.Q ),
    .ZN(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2626_ (.I0(S2MID[0]),
    .I1(\Inst_RegFile_switch_matrix.JW2BEG3 ),
    .S(\Inst_RegFile_ConfigMem.Inst_frame7_bit6.Q ),
    .Z(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2627_ (.A1(N2MID[0]),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame7_bit6.Q ),
    .ZN(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2628_ (.A1(_1274_),
    .A2(\Inst_RegFile_ConfigMem.Inst_frame7_bit6.Q ),
    .B(\Inst_RegFile_ConfigMem.Inst_frame7_bit7.Q ),
    .C(_1193_),
    .ZN(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2629_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame7_bit7.Q ),
    .A2(_1192_),
    .B(_1194_),
    .C(\Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q ),
    .ZN(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _2630_ (.I0(N2MID[1]),
    .I1(E2MID[1]),
    .I2(S2MID[1]),
    .I3(W2MID[1]),
    .S0(\Inst_RegFile_ConfigMem.Inst_frame6_bit6.Q ),
    .S1(\Inst_RegFile_ConfigMem.Inst_frame6_bit7.Q ),
    .Z(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2631_ (.A1(_0138_),
    .A2(_1196_),
    .ZN(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2632_ (.A1(\Inst_RegFile_ConfigMem.Inst_frame9_bit27.Q ),
    .A2(_1195_),
    .A3(_1197_),
    .B1(_1190_),
    .B2(_1191_),
    .ZN(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2633_ (.I0(\Inst_RegFile_32x4.mem[24][3] ),
    .I1(_1198_),
    .S(_1174_),
    .Z(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2634_ (.A1(_1149_),
    .A2(_1170_),
    .ZN(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2635_ (.A1(_1141_),
    .A2(_1199_),
    .ZN(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2636_ (.A1(_1142_),
    .A2(_1149_),
    .A3(_1170_),
    .ZN(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2637_ (.A1(_1135_),
    .A2(_1201_),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2638_ (.I0(\Inst_RegFile_32x4.mem[25][0] ),
    .I1(_1182_),
    .S(_1202_),
    .Z(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2639_ (.I0(\Inst_RegFile_32x4.mem[25][1] ),
    .I1(_1184_),
    .S(_1202_),
    .Z(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2640_ (.I0(\Inst_RegFile_32x4.mem[25][2] ),
    .I1(_1186_),
    .S(_1202_),
    .Z(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2641_ (.I0(\Inst_RegFile_32x4.mem[25][3] ),
    .I1(_1198_),
    .S(_1202_),
    .Z(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2642_ (.A1(_1142_),
    .A2(_1171_),
    .ZN(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2643_ (.A1(_1141_),
    .A2(_1149_),
    .A3(_1169_),
    .ZN(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2644_ (.A1(_1135_),
    .A2(_1204_),
    .ZN(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2645_ (.I0(\Inst_RegFile_32x4.mem[26][0] ),
    .I1(_1182_),
    .S(_1205_),
    .Z(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2646_ (.I0(\Inst_RegFile_32x4.mem[26][1] ),
    .I1(_1184_),
    .S(_1205_),
    .Z(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2647_ (.I0(\Inst_RegFile_32x4.mem[26][2] ),
    .I1(_1186_),
    .S(_1205_),
    .Z(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2648_ (.I0(\Inst_RegFile_32x4.mem[26][3] ),
    .I1(_1198_),
    .S(_1205_),
    .Z(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2649_ (.A1(_1142_),
    .A2(_1199_),
    .ZN(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2650_ (.A1(_1141_),
    .A2(_1149_),
    .A3(_1170_),
    .ZN(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2651_ (.A1(_1135_),
    .A2(_1207_),
    .ZN(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2652_ (.I0(\Inst_RegFile_32x4.mem[27][0] ),
    .I1(_1182_),
    .S(_1208_),
    .Z(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2653_ (.I0(\Inst_RegFile_32x4.mem[27][1] ),
    .I1(_1184_),
    .S(_1208_),
    .Z(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2654_ (.I0(\Inst_RegFile_32x4.mem[27][2] ),
    .I1(_1186_),
    .S(_1208_),
    .Z(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2655_ (.I0(\Inst_RegFile_32x4.mem[27][3] ),
    .I1(_1198_),
    .S(_1208_),
    .Z(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2656_ (.A1(_1122_),
    .A2(_1133_),
    .ZN(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2657_ (.A1(_1173_),
    .A2(_1209_),
    .ZN(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2658_ (.I0(\Inst_RegFile_32x4.mem[28][0] ),
    .I1(_1182_),
    .S(_1210_),
    .Z(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2659_ (.I0(\Inst_RegFile_32x4.mem[28][1] ),
    .I1(_1184_),
    .S(_1210_),
    .Z(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2660_ (.I0(\Inst_RegFile_32x4.mem[28][2] ),
    .I1(_1186_),
    .S(_1210_),
    .Z(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2661_ (.I0(\Inst_RegFile_32x4.mem[28][3] ),
    .I1(_1198_),
    .S(_1210_),
    .Z(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2662_ (.A1(_1107_),
    .A2(_1121_),
    .Z(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2663_ (.A1(_1133_),
    .A2(_1211_),
    .ZN(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2664_ (.A1(_1203_),
    .A2(_1212_),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2665_ (.I0(_1182_),
    .I1(\Inst_RegFile_32x4.mem[2][0] ),
    .S(_1213_),
    .Z(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2666_ (.I0(_1184_),
    .I1(\Inst_RegFile_32x4.mem[2][1] ),
    .S(_1213_),
    .Z(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2667_ (.I0(_1186_),
    .I1(\Inst_RegFile_32x4.mem[2][2] ),
    .S(_1213_),
    .Z(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2668_ (.I0(_1198_),
    .I1(\Inst_RegFile_32x4.mem[2][3] ),
    .S(_1213_),
    .Z(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2669_ (.A1(_1204_),
    .A2(_1209_),
    .ZN(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2670_ (.I0(\Inst_RegFile_32x4.mem[30][0] ),
    .I1(_1182_),
    .S(_1214_),
    .Z(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2671_ (.I0(\Inst_RegFile_32x4.mem[30][1] ),
    .I1(_1184_),
    .S(_1214_),
    .Z(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2672_ (.I0(\Inst_RegFile_32x4.mem[30][2] ),
    .I1(_1186_),
    .S(_1214_),
    .Z(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2673_ (.I0(\Inst_RegFile_32x4.mem[30][3] ),
    .I1(_1198_),
    .S(_1214_),
    .Z(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2674_ (.A1(_1107_),
    .A2(_1120_),
    .Z(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2675_ (.A1(_1133_),
    .A2(_1215_),
    .ZN(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2676_ (.A1(_1200_),
    .A2(_1216_),
    .ZN(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2677_ (.I0(_1182_),
    .I1(\Inst_RegFile_32x4.mem[9][0] ),
    .S(_1217_),
    .Z(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2678_ (.I0(_1184_),
    .I1(\Inst_RegFile_32x4.mem[9][1] ),
    .S(_1217_),
    .Z(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2679_ (.I0(_1186_),
    .I1(\Inst_RegFile_32x4.mem[9][2] ),
    .S(_1217_),
    .Z(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2680_ (.I0(_1198_),
    .I1(\Inst_RegFile_32x4.mem[9][3] ),
    .S(_1217_),
    .Z(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2681_ (.A1(_1134_),
    .A2(_1215_),
    .ZN(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2682_ (.A1(_1200_),
    .A2(_1218_),
    .ZN(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2683_ (.I0(_1182_),
    .I1(\Inst_RegFile_32x4.mem[13][0] ),
    .S(_1219_),
    .Z(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2684_ (.I0(_1184_),
    .I1(\Inst_RegFile_32x4.mem[13][1] ),
    .S(_1219_),
    .Z(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2685_ (.I0(_1186_),
    .I1(\Inst_RegFile_32x4.mem[13][2] ),
    .S(_1219_),
    .Z(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2686_ (.I0(_1198_),
    .I1(\Inst_RegFile_32x4.mem[13][3] ),
    .S(_1219_),
    .Z(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2687_ (.A1(_1107_),
    .A2(_1120_),
    .Z(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2688_ (.A1(_1134_),
    .A2(_1220_),
    .ZN(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2689_ (.A1(_1201_),
    .A2(_1221_),
    .ZN(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2690_ (.I0(\Inst_RegFile_32x4.mem[17][0] ),
    .I1(_1182_),
    .S(_1222_),
    .Z(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2691_ (.I0(\Inst_RegFile_32x4.mem[17][1] ),
    .I1(_1184_),
    .S(_1222_),
    .Z(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2692_ (.I0(\Inst_RegFile_32x4.mem[17][2] ),
    .I1(_1186_),
    .S(_1222_),
    .Z(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2693_ (.I0(\Inst_RegFile_32x4.mem[17][3] ),
    .I1(_1198_),
    .S(_1222_),
    .Z(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2694_ (.A1(_1133_),
    .A2(_1220_),
    .ZN(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2695_ (.A1(_1204_),
    .A2(_1223_),
    .ZN(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2696_ (.I0(\Inst_RegFile_32x4.mem[22][0] ),
    .I1(_1182_),
    .S(_1224_),
    .Z(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2697_ (.I0(\Inst_RegFile_32x4.mem[22][1] ),
    .I1(_1184_),
    .S(_1224_),
    .Z(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2698_ (.I0(\Inst_RegFile_32x4.mem[22][2] ),
    .I1(_1186_),
    .S(_1224_),
    .Z(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2699_ (.I0(\Inst_RegFile_32x4.mem[22][3] ),
    .I1(_1198_),
    .S(_1224_),
    .Z(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2700_ (.A1(_1207_),
    .A2(_1223_),
    .ZN(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2701_ (.I0(\Inst_RegFile_32x4.mem[23][0] ),
    .I1(_1182_),
    .S(_1225_),
    .Z(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2702_ (.I0(\Inst_RegFile_32x4.mem[23][1] ),
    .I1(_1184_),
    .S(_1225_),
    .Z(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2703_ (.I0(\Inst_RegFile_32x4.mem[23][2] ),
    .I1(_1186_),
    .S(_1225_),
    .Z(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2704_ (.I0(\Inst_RegFile_32x4.mem[23][3] ),
    .I1(_1198_),
    .S(_1225_),
    .Z(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2705_ (.A1(_1203_),
    .A2(_1218_),
    .ZN(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2706_ (.I0(_1182_),
    .I1(\Inst_RegFile_32x4.mem[14][0] ),
    .S(_1226_),
    .Z(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2707_ (.I0(_1184_),
    .I1(\Inst_RegFile_32x4.mem[14][1] ),
    .S(_1226_),
    .Z(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2708_ (.I0(_1186_),
    .I1(\Inst_RegFile_32x4.mem[14][2] ),
    .S(_1226_),
    .Z(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2709_ (.I0(_1198_),
    .I1(\Inst_RegFile_32x4.mem[14][3] ),
    .S(_1226_),
    .Z(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2710_ (.A1(_1206_),
    .A2(_1218_),
    .ZN(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2711_ (.I0(_1182_),
    .I1(\Inst_RegFile_32x4.mem[15][0] ),
    .S(_1227_),
    .Z(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2712_ (.I0(_1184_),
    .I1(\Inst_RegFile_32x4.mem[15][1] ),
    .S(_1227_),
    .Z(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2713_ (.I0(_1186_),
    .I1(\Inst_RegFile_32x4.mem[15][2] ),
    .S(_1227_),
    .Z(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2714_ (.I0(_1198_),
    .I1(\Inst_RegFile_32x4.mem[15][3] ),
    .S(_1227_),
    .Z(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2715_ (.A1(_1173_),
    .A2(_1221_),
    .ZN(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2716_ (.I0(\Inst_RegFile_32x4.mem[16][0] ),
    .I1(_1182_),
    .S(_1228_),
    .Z(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2717_ (.I0(\Inst_RegFile_32x4.mem[16][1] ),
    .I1(_1184_),
    .S(_1228_),
    .Z(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2718_ (.I0(\Inst_RegFile_32x4.mem[16][2] ),
    .I1(_1186_),
    .S(_1228_),
    .Z(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2719_ (.I0(\Inst_RegFile_32x4.mem[16][3] ),
    .I1(_1198_),
    .S(_1228_),
    .Z(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2720_ (.A1(_1204_),
    .A2(_1221_),
    .ZN(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2721_ (.I0(\Inst_RegFile_32x4.mem[18][0] ),
    .I1(_1182_),
    .S(_1229_),
    .Z(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2722_ (.I0(\Inst_RegFile_32x4.mem[18][1] ),
    .I1(_1184_),
    .S(_1229_),
    .Z(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2723_ (.I0(\Inst_RegFile_32x4.mem[18][2] ),
    .I1(_1186_),
    .S(_1229_),
    .Z(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2724_ (.I0(\Inst_RegFile_32x4.mem[18][3] ),
    .I1(_1198_),
    .S(_1229_),
    .Z(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2725_ (.A1(_1200_),
    .A2(_1212_),
    .ZN(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2726_ (.I0(_1182_),
    .I1(\Inst_RegFile_32x4.mem[1][0] ),
    .S(_1230_),
    .Z(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2727_ (.I0(_1184_),
    .I1(\Inst_RegFile_32x4.mem[1][1] ),
    .S(_1230_),
    .Z(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2728_ (.I0(_1186_),
    .I1(\Inst_RegFile_32x4.mem[1][2] ),
    .S(_1230_),
    .Z(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2729_ (.I0(_1198_),
    .I1(\Inst_RegFile_32x4.mem[1][3] ),
    .S(_1230_),
    .Z(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2730_ (.A1(_1173_),
    .A2(_1223_),
    .ZN(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2731_ (.I0(\Inst_RegFile_32x4.mem[20][0] ),
    .I1(_1182_),
    .S(_1231_),
    .Z(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2732_ (.I0(\Inst_RegFile_32x4.mem[20][1] ),
    .I1(_1184_),
    .S(_1231_),
    .Z(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2733_ (.I0(\Inst_RegFile_32x4.mem[20][2] ),
    .I1(_1186_),
    .S(_1231_),
    .Z(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2734_ (.I0(\Inst_RegFile_32x4.mem[20][3] ),
    .I1(_1198_),
    .S(_1231_),
    .Z(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2735_ (.A1(_1201_),
    .A2(_1223_),
    .ZN(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2736_ (.I0(\Inst_RegFile_32x4.mem[21][0] ),
    .I1(_1182_),
    .S(_1232_),
    .Z(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2737_ (.I0(\Inst_RegFile_32x4.mem[21][1] ),
    .I1(_1184_),
    .S(_1232_),
    .Z(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2738_ (.I0(\Inst_RegFile_32x4.mem[21][2] ),
    .I1(_1186_),
    .S(_1232_),
    .Z(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2739_ (.I0(\Inst_RegFile_32x4.mem[21][3] ),
    .I1(_1198_),
    .S(_1232_),
    .Z(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2740_ (.A1(_1207_),
    .A2(_1221_),
    .ZN(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2741_ (.I0(\Inst_RegFile_32x4.mem[19][0] ),
    .I1(_1182_),
    .S(_1233_),
    .Z(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2742_ (.I0(\Inst_RegFile_32x4.mem[19][1] ),
    .I1(_1184_),
    .S(_1233_),
    .Z(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2743_ (.I0(\Inst_RegFile_32x4.mem[19][2] ),
    .I1(_1186_),
    .S(_1233_),
    .Z(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2744_ (.I0(\Inst_RegFile_32x4.mem[19][3] ),
    .I1(_1198_),
    .S(_1233_),
    .Z(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2745_ (.A1(_1201_),
    .A2(_1209_),
    .ZN(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2746_ (.I0(\Inst_RegFile_32x4.mem[29][0] ),
    .I1(_1182_),
    .S(_1234_),
    .Z(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2747_ (.I0(\Inst_RegFile_32x4.mem[29][1] ),
    .I1(_1184_),
    .S(_1234_),
    .Z(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2748_ (.I0(\Inst_RegFile_32x4.mem[29][2] ),
    .I1(_1186_),
    .S(_1234_),
    .Z(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2749_ (.I0(\Inst_RegFile_32x4.mem[29][3] ),
    .I1(_1198_),
    .S(_1234_),
    .Z(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2750_ (.A1(_1207_),
    .A2(_1209_),
    .ZN(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2751_ (.I0(\Inst_RegFile_32x4.mem[31][0] ),
    .I1(_1182_),
    .S(_1235_),
    .Z(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2752_ (.I0(\Inst_RegFile_32x4.mem[31][1] ),
    .I1(_1184_),
    .S(_1235_),
    .Z(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2753_ (.I0(\Inst_RegFile_32x4.mem[31][2] ),
    .I1(_1186_),
    .S(_1235_),
    .Z(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2754_ (.I0(\Inst_RegFile_32x4.mem[31][3] ),
    .I1(_1198_),
    .S(_1235_),
    .Z(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2755_ (.A1(_1206_),
    .A2(_1212_),
    .ZN(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2756_ (.I0(_1182_),
    .I1(\Inst_RegFile_32x4.mem[3][0] ),
    .S(_1236_),
    .Z(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2757_ (.I0(_1184_),
    .I1(\Inst_RegFile_32x4.mem[3][1] ),
    .S(_1236_),
    .Z(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2758_ (.I0(_1186_),
    .I1(\Inst_RegFile_32x4.mem[3][2] ),
    .S(_1236_),
    .Z(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2759_ (.I0(_1198_),
    .I1(\Inst_RegFile_32x4.mem[3][3] ),
    .S(_1236_),
    .Z(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2760_ (.A1(_1134_),
    .A2(_1211_),
    .ZN(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2761_ (.A1(_1172_),
    .A2(_1237_),
    .ZN(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2762_ (.I0(_1182_),
    .I1(\Inst_RegFile_32x4.mem[4][0] ),
    .S(_1238_),
    .Z(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2763_ (.I0(_1184_),
    .I1(\Inst_RegFile_32x4.mem[4][1] ),
    .S(_1238_),
    .Z(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2764_ (.I0(_1186_),
    .I1(\Inst_RegFile_32x4.mem[4][2] ),
    .S(_1238_),
    .Z(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2765_ (.I0(_1198_),
    .I1(\Inst_RegFile_32x4.mem[4][3] ),
    .S(_1238_),
    .Z(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2766_ (.A1(_1200_),
    .A2(_1237_),
    .ZN(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2767_ (.I0(_1182_),
    .I1(\Inst_RegFile_32x4.mem[5][0] ),
    .S(_1239_),
    .Z(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2768_ (.I0(_1184_),
    .I1(\Inst_RegFile_32x4.mem[5][1] ),
    .S(_1239_),
    .Z(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2769_ (.I0(_1186_),
    .I1(\Inst_RegFile_32x4.mem[5][2] ),
    .S(_1239_),
    .Z(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2770_ (.I0(_1198_),
    .I1(\Inst_RegFile_32x4.mem[5][3] ),
    .S(_1239_),
    .Z(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2771_ (.A1(_1203_),
    .A2(_1237_),
    .ZN(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2772_ (.I0(_1182_),
    .I1(\Inst_RegFile_32x4.mem[6][0] ),
    .S(_1240_),
    .Z(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2773_ (.I0(_1184_),
    .I1(\Inst_RegFile_32x4.mem[6][1] ),
    .S(_1240_),
    .Z(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2774_ (.I0(_1186_),
    .I1(\Inst_RegFile_32x4.mem[6][2] ),
    .S(_1240_),
    .Z(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2775_ (.I0(_1198_),
    .I1(\Inst_RegFile_32x4.mem[6][3] ),
    .S(_1240_),
    .Z(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2776_ (.A1(_1206_),
    .A2(_1237_),
    .ZN(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2777_ (.I0(_1182_),
    .I1(\Inst_RegFile_32x4.mem[7][0] ),
    .S(_1241_),
    .Z(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2778_ (.I0(_1184_),
    .I1(\Inst_RegFile_32x4.mem[7][1] ),
    .S(_1241_),
    .Z(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2779_ (.I0(_1186_),
    .I1(\Inst_RegFile_32x4.mem[7][2] ),
    .S(_1241_),
    .Z(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2780_ (.I0(_1198_),
    .I1(\Inst_RegFile_32x4.mem[7][3] ),
    .S(_1241_),
    .Z(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2781_ (.A1(_1172_),
    .A2(_1216_),
    .ZN(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2782_ (.I0(_1182_),
    .I1(\Inst_RegFile_32x4.mem[8][0] ),
    .S(_1242_),
    .Z(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2783_ (.I0(_1184_),
    .I1(\Inst_RegFile_32x4.mem[8][1] ),
    .S(_1242_),
    .Z(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2784_ (.I0(_1186_),
    .I1(\Inst_RegFile_32x4.mem[8][2] ),
    .S(_1242_),
    .Z(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2785_ (.I0(_1198_),
    .I1(\Inst_RegFile_32x4.mem[8][3] ),
    .S(_1242_),
    .Z(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2786_ (.A1(_1172_),
    .A2(_1212_),
    .ZN(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2787_ (.I0(_1182_),
    .I1(\Inst_RegFile_32x4.mem[0][0] ),
    .S(_1243_),
    .Z(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2788_ (.I0(_1184_),
    .I1(\Inst_RegFile_32x4.mem[0][1] ),
    .S(_1243_),
    .Z(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2789_ (.I0(_1186_),
    .I1(\Inst_RegFile_32x4.mem[0][2] ),
    .S(_1243_),
    .Z(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2790_ (.I0(_1198_),
    .I1(\Inst_RegFile_32x4.mem[0][3] ),
    .S(_1243_),
    .Z(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2791_ (.A1(_1203_),
    .A2(_1216_),
    .ZN(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2792_ (.I0(_1182_),
    .I1(\Inst_RegFile_32x4.mem[10][0] ),
    .S(_1244_),
    .Z(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2793_ (.I0(_1184_),
    .I1(\Inst_RegFile_32x4.mem[10][1] ),
    .S(_1244_),
    .Z(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2794_ (.I0(_1186_),
    .I1(\Inst_RegFile_32x4.mem[10][2] ),
    .S(_1244_),
    .Z(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2795_ (.I0(_1198_),
    .I1(\Inst_RegFile_32x4.mem[10][3] ),
    .S(_1244_),
    .Z(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2796_ (.A1(_1206_),
    .A2(_1216_),
    .ZN(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2797_ (.I0(_1182_),
    .I1(\Inst_RegFile_32x4.mem[11][0] ),
    .S(_1245_),
    .Z(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2798_ (.I0(_1184_),
    .I1(\Inst_RegFile_32x4.mem[11][1] ),
    .S(_1245_),
    .Z(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2799_ (.I0(_1186_),
    .I1(\Inst_RegFile_32x4.mem[11][2] ),
    .S(_1245_),
    .Z(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2800_ (.I0(_1198_),
    .I1(\Inst_RegFile_32x4.mem[11][3] ),
    .S(_1245_),
    .Z(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2801_ (.A1(_1172_),
    .A2(_1218_),
    .ZN(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2802_ (.I0(_1182_),
    .I1(\Inst_RegFile_32x4.mem[12][0] ),
    .S(_1246_),
    .Z(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2803_ (.I0(_1184_),
    .I1(\Inst_RegFile_32x4.mem[12][1] ),
    .S(_1246_),
    .Z(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2804_ (.I0(_1186_),
    .I1(\Inst_RegFile_32x4.mem[12][2] ),
    .S(_1246_),
    .Z(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2805_ (.I0(_1198_),
    .I1(\Inst_RegFile_32x4.mem[12][3] ),
    .S(_1246_),
    .Z(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2806_ (.D(_0000_),
    .CLK(clknet_4_9_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[24][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2807_ (.D(_0001_),
    .CLK(clknet_4_8_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[24][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2808_ (.D(_0002_),
    .CLK(clknet_4_8_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[24][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2809_ (.D(_0003_),
    .CLK(clknet_4_3_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[24][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2810_ (.D(_0004_),
    .CLK(clknet_4_3_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[25][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2811_ (.D(_0005_),
    .CLK(clknet_4_8_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[25][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2812_ (.D(_0006_),
    .CLK(clknet_4_8_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[25][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2813_ (.D(_0007_),
    .CLK(clknet_4_3_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[25][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2814_ (.D(_0008_),
    .CLK(clknet_4_9_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[26][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2815_ (.D(_0009_),
    .CLK(clknet_4_9_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[26][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2816_ (.D(_0010_),
    .CLK(clknet_4_8_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[26][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2817_ (.D(_0011_),
    .CLK(clknet_4_6_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[26][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2818_ (.D(_0012_),
    .CLK(clknet_4_6_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[27][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2819_ (.D(_0013_),
    .CLK(clknet_4_9_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[27][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2820_ (.D(_0014_),
    .CLK(clknet_4_8_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[27][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2821_ (.D(_0015_),
    .CLK(clknet_4_9_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[27][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2822_ (.D(_0016_),
    .CLK(clknet_4_13_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[28][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2823_ (.D(_0017_),
    .CLK(clknet_4_13_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[28][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2824_ (.D(_0018_),
    .CLK(clknet_4_8_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[28][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2825_ (.D(_0019_),
    .CLK(clknet_4_13_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[28][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2826_ (.D(_0020_),
    .CLK(clknet_4_0_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2827_ (.D(_0021_),
    .CLK(clknet_4_0_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2828_ (.D(_0022_),
    .CLK(clknet_4_2_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2829_ (.D(_0023_),
    .CLK(clknet_4_2_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2830_ (.D(_0024_),
    .CLK(clknet_4_12_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[30][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2831_ (.D(_0025_),
    .CLK(clknet_4_9_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[30][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2832_ (.D(_0026_),
    .CLK(clknet_4_3_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[30][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2833_ (.D(_0027_),
    .CLK(clknet_4_9_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[30][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2834_ (.D(_0028_),
    .CLK(clknet_4_7_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2835_ (.D(_0029_),
    .CLK(clknet_4_7_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2836_ (.D(_0030_),
    .CLK(clknet_4_5_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2837_ (.D(_0031_),
    .CLK(clknet_4_7_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2838_ (.D(_0032_),
    .CLK(clknet_4_5_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2839_ (.D(_0033_),
    .CLK(clknet_4_5_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2840_ (.D(_0034_),
    .CLK(clknet_4_4_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2841_ (.D(_0035_),
    .CLK(clknet_4_5_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2842_ (.D(_0036_),
    .CLK(clknet_4_10_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[17][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2843_ (.D(_0037_),
    .CLK(clknet_4_11_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[17][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2844_ (.D(_0038_),
    .CLK(clknet_4_10_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[17][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2845_ (.D(_0039_),
    .CLK(clknet_4_10_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[17][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2846_ (.D(_0040_),
    .CLK(clknet_4_15_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[22][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2847_ (.D(_0041_),
    .CLK(clknet_4_13_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[22][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2848_ (.D(_0042_),
    .CLK(clknet_4_14_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[22][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2849_ (.D(_0043_),
    .CLK(clknet_4_15_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[22][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2850_ (.D(_0044_),
    .CLK(clknet_4_15_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[23][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2851_ (.D(_0045_),
    .CLK(clknet_4_11_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[23][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2852_ (.D(_0046_),
    .CLK(clknet_4_14_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[23][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2853_ (.D(_0047_),
    .CLK(clknet_4_15_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[23][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2854_ (.D(_0048_),
    .CLK(clknet_4_5_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2855_ (.D(_0049_),
    .CLK(clknet_4_4_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2856_ (.D(_0050_),
    .CLK(clknet_4_4_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2857_ (.D(_0051_),
    .CLK(clknet_4_5_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2858_ (.D(_0052_),
    .CLK(clknet_4_5_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2859_ (.D(_0053_),
    .CLK(clknet_4_4_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2860_ (.D(_0054_),
    .CLK(clknet_4_4_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2861_ (.D(_0055_),
    .CLK(clknet_4_5_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2862_ (.D(_0056_),
    .CLK(clknet_4_10_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[16][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2863_ (.D(_0057_),
    .CLK(clknet_4_11_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[16][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2864_ (.D(_0058_),
    .CLK(clknet_4_10_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[16][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2865_ (.D(_0059_),
    .CLK(clknet_4_10_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[16][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2866_ (.D(_0060_),
    .CLK(clknet_4_14_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[18][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2867_ (.D(_0061_),
    .CLK(clknet_4_11_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[18][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2868_ (.D(_0062_),
    .CLK(clknet_4_10_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[18][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2869_ (.D(_0063_),
    .CLK(clknet_4_14_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[18][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2870_ (.D(_0064_),
    .CLK(clknet_4_2_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2871_ (.D(_0065_),
    .CLK(clknet_4_0_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2872_ (.D(_0066_),
    .CLK(clknet_4_2_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2873_ (.D(_0067_),
    .CLK(clknet_4_2_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2874_ (.D(_0068_),
    .CLK(clknet_4_13_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[20][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2875_ (.D(_0069_),
    .CLK(clknet_4_12_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[20][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2876_ (.D(_0070_),
    .CLK(clknet_4_12_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[20][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2877_ (.D(_0071_),
    .CLK(clknet_4_12_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[20][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2878_ (.D(_0072_),
    .CLK(clknet_4_15_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[21][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2879_ (.D(_0073_),
    .CLK(clknet_4_12_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[21][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2880_ (.D(_0074_),
    .CLK(clknet_4_11_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[21][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2881_ (.D(_0075_),
    .CLK(clknet_4_14_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[21][3] ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2882_ (.D(FrameData[2]),
    .E(FrameStrobe[12]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2883_ (.D(FrameData[3]),
    .E(FrameStrobe[12]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2884_ (.D(FrameData[4]),
    .E(FrameStrobe[12]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2885_ (.D(FrameData[5]),
    .E(FrameStrobe[12]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2886_ (.D(FrameData[6]),
    .E(FrameStrobe[12]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2887_ (.D(FrameData[7]),
    .E(FrameStrobe[12]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2888_ (.D(FrameData[8]),
    .E(FrameStrobe[12]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2889_ (.D(FrameData[9]),
    .E(FrameStrobe[12]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2890_ (.D(FrameData[10]),
    .E(FrameStrobe[12]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2891_ (.D(FrameData[11]),
    .E(FrameStrobe[12]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2892_ (.D(FrameData[12]),
    .E(FrameStrobe[12]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2893_ (.D(FrameData[13]),
    .E(FrameStrobe[12]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2894_ (.D(FrameData[14]),
    .E(FrameStrobe[12]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2895_ (.D(FrameData[15]),
    .E(FrameStrobe[12]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2896_ (.D(FrameData[16]),
    .E(FrameStrobe[12]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2897_ (.D(FrameData[17]),
    .E(FrameStrobe[12]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2898_ (.D(FrameData[18]),
    .E(FrameStrobe[12]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2899_ (.D(FrameData[19]),
    .E(FrameStrobe[12]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2900_ (.D(FrameData[20]),
    .E(FrameStrobe[12]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2901_ (.D(FrameData[21]),
    .E(FrameStrobe[12]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2902_ (.D(FrameData[22]),
    .E(FrameStrobe[12]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2903_ (.D(FrameData[23]),
    .E(FrameStrobe[12]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2904_ (.D(FrameData[24]),
    .E(FrameStrobe[12]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2905_ (.D(FrameData[25]),
    .E(FrameStrobe[12]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2906_ (.D(FrameData[26]),
    .E(FrameStrobe[12]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2907_ (.D(FrameData[27]),
    .E(FrameStrobe[12]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2908_ (.D(FrameData[28]),
    .E(FrameStrobe[12]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2909_ (.D(FrameData[29]),
    .E(FrameStrobe[12]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2910_ (.D(FrameData[30]),
    .E(FrameStrobe[12]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2911_ (.D(FrameData[31]),
    .E(FrameStrobe[12]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame12_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2912_ (.D(FrameData[0]),
    .E(FrameStrobe[11]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2913_ (.D(FrameData[1]),
    .E(FrameStrobe[11]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2914_ (.D(FrameData[2]),
    .E(FrameStrobe[11]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2915_ (.D(FrameData[3]),
    .E(FrameStrobe[11]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2916_ (.D(FrameData[4]),
    .E(FrameStrobe[11]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2917_ (.D(FrameData[5]),
    .E(FrameStrobe[11]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2918_ (.D(FrameData[6]),
    .E(FrameStrobe[11]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2919_ (.D(FrameData[7]),
    .E(FrameStrobe[11]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2920_ (.D(FrameData[8]),
    .E(FrameStrobe[11]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2921_ (.D(FrameData[9]),
    .E(FrameStrobe[11]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2922_ (.D(FrameData[10]),
    .E(FrameStrobe[11]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2923_ (.D(FrameData[11]),
    .E(FrameStrobe[11]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2924_ (.D(FrameData[12]),
    .E(FrameStrobe[11]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2925_ (.D(FrameData[13]),
    .E(FrameStrobe[11]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2926_ (.D(FrameData[14]),
    .E(FrameStrobe[11]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2927_ (.D(FrameData[15]),
    .E(FrameStrobe[11]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2928_ (.D(FrameData[16]),
    .E(FrameStrobe[11]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2929_ (.D(FrameData[17]),
    .E(FrameStrobe[11]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2930_ (.D(FrameData[18]),
    .E(FrameStrobe[11]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2931_ (.D(FrameData[19]),
    .E(FrameStrobe[11]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2932_ (.D(FrameData[20]),
    .E(FrameStrobe[11]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2933_ (.D(FrameData[21]),
    .E(FrameStrobe[11]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2934_ (.D(FrameData[22]),
    .E(FrameStrobe[11]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2935_ (.D(FrameData[23]),
    .E(FrameStrobe[11]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2936_ (.D(FrameData[24]),
    .E(FrameStrobe[11]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2937_ (.D(FrameData[25]),
    .E(FrameStrobe[11]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2938_ (.D(FrameData[26]),
    .E(FrameStrobe[11]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2939_ (.D(FrameData[27]),
    .E(FrameStrobe[11]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2940_ (.D(FrameData[28]),
    .E(FrameStrobe[11]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2941_ (.D(FrameData[29]),
    .E(FrameStrobe[11]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2942_ (.D(FrameData[30]),
    .E(FrameStrobe[11]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2943_ (.D(FrameData[31]),
    .E(FrameStrobe[11]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame11_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2944_ (.D(FrameData[0]),
    .E(FrameStrobe[10]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2945_ (.D(FrameData[1]),
    .E(FrameStrobe[10]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2946_ (.D(FrameData[2]),
    .E(FrameStrobe[10]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2947_ (.D(FrameData[3]),
    .E(FrameStrobe[10]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2948_ (.D(FrameData[4]),
    .E(FrameStrobe[10]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2949_ (.D(FrameData[5]),
    .E(FrameStrobe[10]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2950_ (.D(FrameData[6]),
    .E(FrameStrobe[10]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2951_ (.D(FrameData[7]),
    .E(FrameStrobe[10]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2952_ (.D(FrameData[8]),
    .E(FrameStrobe[10]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2953_ (.D(FrameData[9]),
    .E(FrameStrobe[10]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2954_ (.D(FrameData[10]),
    .E(FrameStrobe[10]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2955_ (.D(FrameData[11]),
    .E(FrameStrobe[10]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2956_ (.D(FrameData[12]),
    .E(FrameStrobe[10]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2957_ (.D(FrameData[13]),
    .E(FrameStrobe[10]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2958_ (.D(FrameData[14]),
    .E(FrameStrobe[10]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2959_ (.D(FrameData[15]),
    .E(FrameStrobe[10]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2960_ (.D(FrameData[16]),
    .E(FrameStrobe[10]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2961_ (.D(FrameData[17]),
    .E(FrameStrobe[10]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2962_ (.D(FrameData[18]),
    .E(FrameStrobe[10]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2963_ (.D(FrameData[19]),
    .E(FrameStrobe[10]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2964_ (.D(FrameData[20]),
    .E(FrameStrobe[10]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2965_ (.D(FrameData[21]),
    .E(FrameStrobe[10]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2966_ (.D(FrameData[22]),
    .E(FrameStrobe[10]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2967_ (.D(FrameData[23]),
    .E(FrameStrobe[10]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2968_ (.D(FrameData[24]),
    .E(FrameStrobe[10]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2969_ (.D(FrameData[25]),
    .E(FrameStrobe[10]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2970_ (.D(FrameData[26]),
    .E(FrameStrobe[10]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2971_ (.D(FrameData[27]),
    .E(FrameStrobe[10]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2972_ (.D(FrameData[28]),
    .E(FrameStrobe[10]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2973_ (.D(FrameData[29]),
    .E(FrameStrobe[10]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2974_ (.D(FrameData[30]),
    .E(FrameStrobe[10]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2975_ (.D(FrameData[31]),
    .E(FrameStrobe[10]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame10_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2976_ (.D(FrameData[0]),
    .E(FrameStrobe[9]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2977_ (.D(FrameData[1]),
    .E(FrameStrobe[9]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2978_ (.D(FrameData[2]),
    .E(FrameStrobe[9]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2979_ (.D(FrameData[3]),
    .E(FrameStrobe[9]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2980_ (.D(FrameData[4]),
    .E(FrameStrobe[9]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2981_ (.D(FrameData[5]),
    .E(FrameStrobe[9]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2982_ (.D(FrameData[6]),
    .E(FrameStrobe[9]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2983_ (.D(FrameData[7]),
    .E(FrameStrobe[9]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2984_ (.D(FrameData[8]),
    .E(FrameStrobe[9]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2985_ (.D(FrameData[9]),
    .E(FrameStrobe[9]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2986_ (.D(FrameData[10]),
    .E(FrameStrobe[9]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2987_ (.D(FrameData[11]),
    .E(FrameStrobe[9]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2988_ (.D(FrameData[12]),
    .E(FrameStrobe[9]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2989_ (.D(FrameData[13]),
    .E(FrameStrobe[9]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2990_ (.D(FrameData[14]),
    .E(FrameStrobe[9]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2991_ (.D(FrameData[15]),
    .E(FrameStrobe[9]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2992_ (.D(FrameData[16]),
    .E(FrameStrobe[9]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2993_ (.D(FrameData[17]),
    .E(FrameStrobe[9]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2994_ (.D(FrameData[18]),
    .E(FrameStrobe[9]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2995_ (.D(FrameData[19]),
    .E(FrameStrobe[9]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2996_ (.D(FrameData[20]),
    .E(FrameStrobe[9]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2997_ (.D(FrameData[21]),
    .E(FrameStrobe[9]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2998_ (.D(FrameData[22]),
    .E(FrameStrobe[9]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2999_ (.D(FrameData[23]),
    .E(FrameStrobe[9]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3000_ (.D(FrameData[24]),
    .E(FrameStrobe[9]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3001_ (.D(FrameData[25]),
    .E(FrameStrobe[9]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3002_ (.D(FrameData[26]),
    .E(FrameStrobe[9]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3003_ (.D(FrameData[27]),
    .E(FrameStrobe[9]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3004_ (.D(FrameData[28]),
    .E(FrameStrobe[9]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3005_ (.D(FrameData[29]),
    .E(FrameStrobe[9]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3006_ (.D(FrameData[30]),
    .E(FrameStrobe[9]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3007_ (.D(FrameData[31]),
    .E(FrameStrobe[9]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame9_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3008_ (.D(FrameData[0]),
    .E(FrameStrobe[8]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3009_ (.D(FrameData[1]),
    .E(FrameStrobe[8]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3010_ (.D(FrameData[2]),
    .E(FrameStrobe[8]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3011_ (.D(FrameData[3]),
    .E(FrameStrobe[8]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3012_ (.D(FrameData[4]),
    .E(FrameStrobe[8]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3013_ (.D(FrameData[5]),
    .E(FrameStrobe[8]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3014_ (.D(FrameData[6]),
    .E(FrameStrobe[8]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3015_ (.D(FrameData[7]),
    .E(FrameStrobe[8]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3016_ (.D(FrameData[8]),
    .E(FrameStrobe[8]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3017_ (.D(FrameData[9]),
    .E(FrameStrobe[8]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3018_ (.D(FrameData[10]),
    .E(FrameStrobe[8]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3019_ (.D(FrameData[11]),
    .E(FrameStrobe[8]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3020_ (.D(FrameData[12]),
    .E(FrameStrobe[8]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3021_ (.D(FrameData[13]),
    .E(FrameStrobe[8]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3022_ (.D(FrameData[14]),
    .E(FrameStrobe[8]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3023_ (.D(FrameData[15]),
    .E(FrameStrobe[8]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3024_ (.D(FrameData[16]),
    .E(FrameStrobe[8]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3025_ (.D(FrameData[17]),
    .E(FrameStrobe[8]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3026_ (.D(FrameData[18]),
    .E(FrameStrobe[8]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3027_ (.D(FrameData[19]),
    .E(FrameStrobe[8]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3028_ (.D(FrameData[20]),
    .E(FrameStrobe[8]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3029_ (.D(FrameData[21]),
    .E(FrameStrobe[8]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3030_ (.D(FrameData[22]),
    .E(FrameStrobe[8]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3031_ (.D(FrameData[23]),
    .E(FrameStrobe[8]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3032_ (.D(FrameData[24]),
    .E(FrameStrobe[8]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3033_ (.D(FrameData[25]),
    .E(FrameStrobe[8]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3034_ (.D(FrameData[26]),
    .E(FrameStrobe[8]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3035_ (.D(FrameData[27]),
    .E(FrameStrobe[8]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3036_ (.D(FrameData[28]),
    .E(FrameStrobe[8]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3037_ (.D(FrameData[29]),
    .E(FrameStrobe[8]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3038_ (.D(FrameData[30]),
    .E(FrameStrobe[8]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3039_ (.D(FrameData[31]),
    .E(FrameStrobe[8]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame8_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3040_ (.D(FrameData[0]),
    .E(FrameStrobe[7]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3041_ (.D(FrameData[1]),
    .E(FrameStrobe[7]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3042_ (.D(FrameData[2]),
    .E(FrameStrobe[7]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3043_ (.D(FrameData[3]),
    .E(FrameStrobe[7]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3044_ (.D(FrameData[4]),
    .E(FrameStrobe[7]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3045_ (.D(FrameData[5]),
    .E(FrameStrobe[7]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3046_ (.D(FrameData[6]),
    .E(FrameStrobe[7]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3047_ (.D(FrameData[7]),
    .E(FrameStrobe[7]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3048_ (.D(FrameData[8]),
    .E(FrameStrobe[7]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3049_ (.D(FrameData[9]),
    .E(FrameStrobe[7]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3050_ (.D(FrameData[10]),
    .E(FrameStrobe[7]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3051_ (.D(FrameData[11]),
    .E(FrameStrobe[7]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3052_ (.D(FrameData[12]),
    .E(FrameStrobe[7]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3053_ (.D(FrameData[13]),
    .E(FrameStrobe[7]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3054_ (.D(FrameData[14]),
    .E(FrameStrobe[7]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3055_ (.D(FrameData[15]),
    .E(FrameStrobe[7]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3056_ (.D(FrameData[16]),
    .E(FrameStrobe[7]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3057_ (.D(FrameData[17]),
    .E(FrameStrobe[7]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3058_ (.D(FrameData[18]),
    .E(FrameStrobe[7]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3059_ (.D(FrameData[19]),
    .E(FrameStrobe[7]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3060_ (.D(FrameData[20]),
    .E(FrameStrobe[7]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3061_ (.D(FrameData[21]),
    .E(FrameStrobe[7]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3062_ (.D(FrameData[22]),
    .E(FrameStrobe[7]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3063_ (.D(FrameData[23]),
    .E(FrameStrobe[7]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3064_ (.D(FrameData[24]),
    .E(FrameStrobe[7]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3065_ (.D(FrameData[25]),
    .E(FrameStrobe[7]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3066_ (.D(FrameData[26]),
    .E(FrameStrobe[7]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3067_ (.D(FrameData[27]),
    .E(FrameStrobe[7]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3068_ (.D(FrameData[28]),
    .E(FrameStrobe[7]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3069_ (.D(FrameData[29]),
    .E(FrameStrobe[7]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3070_ (.D(FrameData[30]),
    .E(FrameStrobe[7]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3071_ (.D(FrameData[31]),
    .E(FrameStrobe[7]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame7_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3072_ (.D(FrameData[0]),
    .E(FrameStrobe[6]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3073_ (.D(FrameData[1]),
    .E(FrameStrobe[6]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3074_ (.D(FrameData[2]),
    .E(FrameStrobe[6]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3075_ (.D(FrameData[3]),
    .E(FrameStrobe[6]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3076_ (.D(FrameData[4]),
    .E(FrameStrobe[6]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3077_ (.D(FrameData[5]),
    .E(FrameStrobe[6]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3078_ (.D(FrameData[6]),
    .E(FrameStrobe[6]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3079_ (.D(FrameData[7]),
    .E(FrameStrobe[6]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3080_ (.D(FrameData[8]),
    .E(FrameStrobe[6]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3081_ (.D(FrameData[9]),
    .E(FrameStrobe[6]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3082_ (.D(FrameData[10]),
    .E(FrameStrobe[6]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3083_ (.D(FrameData[11]),
    .E(FrameStrobe[6]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3084_ (.D(FrameData[12]),
    .E(FrameStrobe[6]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3085_ (.D(FrameData[13]),
    .E(FrameStrobe[6]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3086_ (.D(FrameData[14]),
    .E(FrameStrobe[6]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3087_ (.D(FrameData[15]),
    .E(FrameStrobe[6]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3088_ (.D(FrameData[16]),
    .E(FrameStrobe[6]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3089_ (.D(FrameData[17]),
    .E(FrameStrobe[6]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3090_ (.D(FrameData[18]),
    .E(FrameStrobe[6]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3091_ (.D(FrameData[19]),
    .E(FrameStrobe[6]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3092_ (.D(FrameData[20]),
    .E(FrameStrobe[6]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3093_ (.D(FrameData[21]),
    .E(FrameStrobe[6]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3094_ (.D(FrameData[22]),
    .E(FrameStrobe[6]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3095_ (.D(FrameData[23]),
    .E(FrameStrobe[6]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3096_ (.D(FrameData[24]),
    .E(FrameStrobe[6]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3097_ (.D(FrameData[25]),
    .E(FrameStrobe[6]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3098_ (.D(FrameData[26]),
    .E(FrameStrobe[6]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3099_ (.D(FrameData[27]),
    .E(FrameStrobe[6]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3100_ (.D(FrameData[28]),
    .E(FrameStrobe[6]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3101_ (.D(FrameData[29]),
    .E(FrameStrobe[6]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3102_ (.D(FrameData[30]),
    .E(FrameStrobe[6]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3103_ (.D(FrameData[31]),
    .E(FrameStrobe[6]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame6_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3104_ (.D(FrameData[0]),
    .E(FrameStrobe[5]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3105_ (.D(FrameData[1]),
    .E(FrameStrobe[5]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3106_ (.D(FrameData[2]),
    .E(FrameStrobe[5]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3107_ (.D(FrameData[3]),
    .E(FrameStrobe[5]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3108_ (.D(FrameData[4]),
    .E(FrameStrobe[5]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3109_ (.D(FrameData[5]),
    .E(FrameStrobe[5]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3110_ (.D(FrameData[6]),
    .E(FrameStrobe[5]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3111_ (.D(FrameData[7]),
    .E(FrameStrobe[5]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3112_ (.D(FrameData[8]),
    .E(FrameStrobe[5]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3113_ (.D(FrameData[9]),
    .E(FrameStrobe[5]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3114_ (.D(FrameData[10]),
    .E(FrameStrobe[5]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3115_ (.D(FrameData[11]),
    .E(FrameStrobe[5]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3116_ (.D(FrameData[12]),
    .E(FrameStrobe[5]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3117_ (.D(FrameData[13]),
    .E(FrameStrobe[5]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3118_ (.D(FrameData[14]),
    .E(FrameStrobe[5]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3119_ (.D(FrameData[15]),
    .E(FrameStrobe[5]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3120_ (.D(FrameData[16]),
    .E(FrameStrobe[5]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3121_ (.D(FrameData[17]),
    .E(FrameStrobe[5]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3122_ (.D(FrameData[18]),
    .E(FrameStrobe[5]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3123_ (.D(FrameData[19]),
    .E(FrameStrobe[5]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3124_ (.D(FrameData[20]),
    .E(FrameStrobe[5]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3125_ (.D(FrameData[21]),
    .E(FrameStrobe[5]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3126_ (.D(FrameData[22]),
    .E(FrameStrobe[5]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3127_ (.D(FrameData[23]),
    .E(FrameStrobe[5]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3128_ (.D(FrameData[24]),
    .E(FrameStrobe[5]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3129_ (.D(FrameData[25]),
    .E(FrameStrobe[5]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3130_ (.D(FrameData[26]),
    .E(FrameStrobe[5]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3131_ (.D(FrameData[27]),
    .E(FrameStrobe[5]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3132_ (.D(FrameData[28]),
    .E(FrameStrobe[5]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3133_ (.D(FrameData[29]),
    .E(FrameStrobe[5]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3134_ (.D(FrameData[30]),
    .E(FrameStrobe[5]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3135_ (.D(FrameData[31]),
    .E(FrameStrobe[5]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame5_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3136_ (.D(FrameData[0]),
    .E(FrameStrobe[4]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3137_ (.D(FrameData[1]),
    .E(FrameStrobe[4]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3138_ (.D(FrameData[2]),
    .E(FrameStrobe[4]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3139_ (.D(FrameData[3]),
    .E(FrameStrobe[4]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3140_ (.D(FrameData[4]),
    .E(FrameStrobe[4]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3141_ (.D(FrameData[5]),
    .E(FrameStrobe[4]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3142_ (.D(FrameData[6]),
    .E(FrameStrobe[4]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3143_ (.D(FrameData[7]),
    .E(FrameStrobe[4]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3144_ (.D(FrameData[8]),
    .E(FrameStrobe[4]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3145_ (.D(FrameData[9]),
    .E(FrameStrobe[4]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3146_ (.D(FrameData[10]),
    .E(FrameStrobe[4]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3147_ (.D(FrameData[11]),
    .E(FrameStrobe[4]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3148_ (.D(FrameData[12]),
    .E(FrameStrobe[4]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3149_ (.D(FrameData[13]),
    .E(FrameStrobe[4]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3150_ (.D(FrameData[14]),
    .E(FrameStrobe[4]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3151_ (.D(FrameData[15]),
    .E(FrameStrobe[4]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3152_ (.D(FrameData[16]),
    .E(FrameStrobe[4]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3153_ (.D(FrameData[17]),
    .E(FrameStrobe[4]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3154_ (.D(FrameData[18]),
    .E(FrameStrobe[4]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3155_ (.D(FrameData[19]),
    .E(FrameStrobe[4]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3156_ (.D(FrameData[20]),
    .E(FrameStrobe[4]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3157_ (.D(FrameData[21]),
    .E(FrameStrobe[4]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3158_ (.D(FrameData[22]),
    .E(FrameStrobe[4]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3159_ (.D(FrameData[23]),
    .E(FrameStrobe[4]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3160_ (.D(FrameData[24]),
    .E(FrameStrobe[4]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3161_ (.D(FrameData[25]),
    .E(FrameStrobe[4]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3162_ (.D(FrameData[26]),
    .E(FrameStrobe[4]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3163_ (.D(FrameData[27]),
    .E(FrameStrobe[4]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3164_ (.D(FrameData[28]),
    .E(FrameStrobe[4]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3165_ (.D(FrameData[29]),
    .E(FrameStrobe[4]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3166_ (.D(FrameData[30]),
    .E(FrameStrobe[4]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3167_ (.D(FrameData[31]),
    .E(FrameStrobe[4]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame4_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3168_ (.D(FrameData[0]),
    .E(FrameStrobe[3]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3169_ (.D(FrameData[1]),
    .E(FrameStrobe[3]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3170_ (.D(FrameData[2]),
    .E(FrameStrobe[3]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3171_ (.D(FrameData[3]),
    .E(FrameStrobe[3]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3172_ (.D(FrameData[4]),
    .E(FrameStrobe[3]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3173_ (.D(FrameData[5]),
    .E(FrameStrobe[3]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3174_ (.D(FrameData[6]),
    .E(FrameStrobe[3]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3175_ (.D(FrameData[7]),
    .E(FrameStrobe[3]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3176_ (.D(FrameData[8]),
    .E(FrameStrobe[3]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3177_ (.D(FrameData[9]),
    .E(FrameStrobe[3]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3178_ (.D(FrameData[10]),
    .E(FrameStrobe[3]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3179_ (.D(FrameData[11]),
    .E(FrameStrobe[3]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3180_ (.D(FrameData[12]),
    .E(FrameStrobe[3]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3181_ (.D(FrameData[13]),
    .E(FrameStrobe[3]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3182_ (.D(FrameData[14]),
    .E(FrameStrobe[3]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3183_ (.D(FrameData[15]),
    .E(FrameStrobe[3]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3184_ (.D(FrameData[16]),
    .E(FrameStrobe[3]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3185_ (.D(FrameData[17]),
    .E(FrameStrobe[3]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3186_ (.D(FrameData[18]),
    .E(FrameStrobe[3]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3187_ (.D(FrameData[19]),
    .E(FrameStrobe[3]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3188_ (.D(FrameData[20]),
    .E(FrameStrobe[3]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3189_ (.D(FrameData[21]),
    .E(FrameStrobe[3]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3190_ (.D(FrameData[22]),
    .E(FrameStrobe[3]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3191_ (.D(FrameData[23]),
    .E(FrameStrobe[3]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3192_ (.D(FrameData[24]),
    .E(FrameStrobe[3]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3193_ (.D(FrameData[25]),
    .E(FrameStrobe[3]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3194_ (.D(FrameData[26]),
    .E(FrameStrobe[3]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3195_ (.D(FrameData[27]),
    .E(FrameStrobe[3]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3196_ (.D(FrameData[28]),
    .E(FrameStrobe[3]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3197_ (.D(FrameData[29]),
    .E(FrameStrobe[3]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3198_ (.D(FrameData[30]),
    .E(FrameStrobe[3]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3199_ (.D(FrameData[31]),
    .E(FrameStrobe[3]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame3_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3200_ (.D(FrameData[0]),
    .E(FrameStrobe[2]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3201_ (.D(FrameData[1]),
    .E(FrameStrobe[2]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3202_ (.D(FrameData[2]),
    .E(FrameStrobe[2]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3203_ (.D(FrameData[3]),
    .E(FrameStrobe[2]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3204_ (.D(FrameData[4]),
    .E(FrameStrobe[2]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3205_ (.D(FrameData[5]),
    .E(FrameStrobe[2]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3206_ (.D(FrameData[6]),
    .E(FrameStrobe[2]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3207_ (.D(FrameData[7]),
    .E(FrameStrobe[2]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3208_ (.D(FrameData[8]),
    .E(FrameStrobe[2]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3209_ (.D(FrameData[9]),
    .E(FrameStrobe[2]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3210_ (.D(FrameData[10]),
    .E(FrameStrobe[2]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3211_ (.D(FrameData[11]),
    .E(FrameStrobe[2]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3212_ (.D(FrameData[12]),
    .E(FrameStrobe[2]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3213_ (.D(FrameData[13]),
    .E(FrameStrobe[2]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3214_ (.D(FrameData[14]),
    .E(FrameStrobe[2]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3215_ (.D(FrameData[15]),
    .E(FrameStrobe[2]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3216_ (.D(FrameData[16]),
    .E(FrameStrobe[2]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3217_ (.D(FrameData[17]),
    .E(FrameStrobe[2]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3218_ (.D(FrameData[18]),
    .E(FrameStrobe[2]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3219_ (.D(FrameData[19]),
    .E(FrameStrobe[2]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3220_ (.D(FrameData[20]),
    .E(FrameStrobe[2]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3221_ (.D(FrameData[21]),
    .E(FrameStrobe[2]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3222_ (.D(FrameData[22]),
    .E(FrameStrobe[2]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3223_ (.D(FrameData[23]),
    .E(FrameStrobe[2]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3224_ (.D(FrameData[24]),
    .E(FrameStrobe[2]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3225_ (.D(FrameData[25]),
    .E(FrameStrobe[2]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3226_ (.D(FrameData[26]),
    .E(FrameStrobe[2]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3227_ (.D(FrameData[27]),
    .E(FrameStrobe[2]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3228_ (.D(FrameData[28]),
    .E(FrameStrobe[2]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3229_ (.D(FrameData[29]),
    .E(FrameStrobe[2]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3230_ (.D(FrameData[30]),
    .E(FrameStrobe[2]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3231_ (.D(FrameData[31]),
    .E(FrameStrobe[2]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame2_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3232_ (.D(FrameData[0]),
    .E(FrameStrobe[1]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3233_ (.D(FrameData[1]),
    .E(FrameStrobe[1]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3234_ (.D(FrameData[2]),
    .E(FrameStrobe[1]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3235_ (.D(FrameData[3]),
    .E(FrameStrobe[1]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3236_ (.D(FrameData[4]),
    .E(FrameStrobe[1]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3237_ (.D(FrameData[5]),
    .E(FrameStrobe[1]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3238_ (.D(FrameData[6]),
    .E(FrameStrobe[1]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3239_ (.D(FrameData[7]),
    .E(FrameStrobe[1]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3240_ (.D(FrameData[8]),
    .E(FrameStrobe[1]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3241_ (.D(FrameData[9]),
    .E(FrameStrobe[1]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3242_ (.D(FrameData[10]),
    .E(FrameStrobe[1]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3243_ (.D(FrameData[11]),
    .E(FrameStrobe[1]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3244_ (.D(FrameData[12]),
    .E(FrameStrobe[1]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3245_ (.D(FrameData[13]),
    .E(FrameStrobe[1]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3246_ (.D(FrameData[14]),
    .E(FrameStrobe[1]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3247_ (.D(FrameData[15]),
    .E(FrameStrobe[1]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3248_ (.D(FrameData[16]),
    .E(FrameStrobe[1]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3249_ (.D(FrameData[17]),
    .E(FrameStrobe[1]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3250_ (.D(FrameData[18]),
    .E(FrameStrobe[1]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3251_ (.D(FrameData[19]),
    .E(FrameStrobe[1]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3252_ (.D(FrameData[20]),
    .E(FrameStrobe[1]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3253_ (.D(FrameData[21]),
    .E(FrameStrobe[1]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3254_ (.D(FrameData[22]),
    .E(FrameStrobe[1]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3255_ (.D(FrameData[23]),
    .E(FrameStrobe[1]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3256_ (.D(FrameData[24]),
    .E(FrameStrobe[1]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3257_ (.D(FrameData[25]),
    .E(FrameStrobe[1]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3258_ (.D(FrameData[26]),
    .E(FrameStrobe[1]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3259_ (.D(FrameData[27]),
    .E(FrameStrobe[1]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3260_ (.D(FrameData[28]),
    .E(FrameStrobe[1]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3261_ (.D(FrameData[29]),
    .E(FrameStrobe[1]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3262_ (.D(FrameData[30]),
    .E(FrameStrobe[1]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3263_ (.D(FrameData[31]),
    .E(FrameStrobe[1]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame1_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3264_ (.D(FrameData[0]),
    .E(FrameStrobe[0]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3265_ (.D(FrameData[1]),
    .E(FrameStrobe[0]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3266_ (.D(FrameData[2]),
    .E(FrameStrobe[0]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3267_ (.D(FrameData[3]),
    .E(FrameStrobe[0]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3268_ (.D(FrameData[4]),
    .E(FrameStrobe[0]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3269_ (.D(FrameData[5]),
    .E(FrameStrobe[0]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3270_ (.D(FrameData[6]),
    .E(FrameStrobe[0]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3271_ (.D(FrameData[7]),
    .E(FrameStrobe[0]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3272_ (.D(FrameData[8]),
    .E(FrameStrobe[0]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3273_ (.D(FrameData[9]),
    .E(FrameStrobe[0]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3274_ (.D(FrameData[10]),
    .E(FrameStrobe[0]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3275_ (.D(FrameData[11]),
    .E(FrameStrobe[0]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3276_ (.D(FrameData[12]),
    .E(FrameStrobe[0]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3277_ (.D(FrameData[13]),
    .E(FrameStrobe[0]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3278_ (.D(FrameData[14]),
    .E(FrameStrobe[0]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3279_ (.D(FrameData[15]),
    .E(FrameStrobe[0]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3280_ (.D(FrameData[16]),
    .E(FrameStrobe[0]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3281_ (.D(FrameData[17]),
    .E(FrameStrobe[0]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3282_ (.D(FrameData[18]),
    .E(FrameStrobe[0]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3283_ (.D(FrameData[19]),
    .E(FrameStrobe[0]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3284_ (.D(FrameData[20]),
    .E(FrameStrobe[0]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3285_ (.D(FrameData[21]),
    .E(FrameStrobe[0]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3286_ (.D(FrameData[22]),
    .E(FrameStrobe[0]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3287_ (.D(FrameData[23]),
    .E(FrameStrobe[0]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3288_ (.D(FrameData[24]),
    .E(FrameStrobe[0]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3289_ (.D(FrameData[25]),
    .E(FrameStrobe[0]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3290_ (.D(FrameData[26]),
    .E(FrameStrobe[0]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3291_ (.D(FrameData[27]),
    .E(FrameStrobe[0]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3292_ (.D(FrameData[28]),
    .E(FrameStrobe[0]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3293_ (.D(FrameData[29]),
    .E(FrameStrobe[0]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3294_ (.D(FrameData[30]),
    .E(FrameStrobe[0]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _3295_ (.D(FrameData[31]),
    .E(FrameStrobe[0]),
    .Q(\Inst_RegFile_ConfigMem.Inst_frame0_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3296_ (.D(\Inst_RegFile_32x4.BD_comb[0] ),
    .CLK(clknet_4_15_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.BD_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3297_ (.D(\Inst_RegFile_32x4.BD_comb[1] ),
    .CLK(clknet_4_15_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.BD_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3298_ (.D(\Inst_RegFile_32x4.BD_comb[2] ),
    .CLK(clknet_4_14_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.BD_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3299_ (.D(\Inst_RegFile_32x4.BD_comb[3] ),
    .CLK(clknet_4_15_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.BD_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3300_ (.D(\Inst_RegFile_32x4.AD_comb[0] ),
    .CLK(clknet_4_6_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.AD_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3301_ (.D(\Inst_RegFile_32x4.AD_comb[1] ),
    .CLK(clknet_4_6_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.AD_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3302_ (.D(\Inst_RegFile_32x4.AD_comb[2] ),
    .CLK(clknet_4_3_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.AD_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3303_ (.D(\Inst_RegFile_32x4.AD_comb[3] ),
    .CLK(clknet_4_3_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.AD_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3304_ (.D(_0076_),
    .CLK(clknet_4_14_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[19][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3305_ (.D(_0077_),
    .CLK(clknet_4_11_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[19][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3306_ (.D(_0078_),
    .CLK(clknet_4_10_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[19][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3307_ (.D(_0079_),
    .CLK(clknet_4_14_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[19][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3308_ (.D(_0080_),
    .CLK(clknet_4_13_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[29][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3309_ (.D(_0081_),
    .CLK(clknet_4_9_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[29][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3310_ (.D(_0082_),
    .CLK(clknet_4_3_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[29][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3311_ (.D(_0083_),
    .CLK(clknet_4_13_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[29][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3312_ (.D(_0084_),
    .CLK(clknet_4_12_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[31][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3313_ (.D(_0085_),
    .CLK(clknet_4_9_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[31][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3314_ (.D(_0086_),
    .CLK(clknet_4_6_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[31][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3315_ (.D(_0087_),
    .CLK(clknet_4_7_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[31][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3316_ (.D(_0088_),
    .CLK(clknet_4_0_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3317_ (.D(_0089_),
    .CLK(clknet_4_1_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3318_ (.D(_0090_),
    .CLK(clknet_4_2_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3319_ (.D(_0091_),
    .CLK(clknet_4_3_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3320_ (.D(_0092_),
    .CLK(clknet_4_1_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3321_ (.D(_0093_),
    .CLK(clknet_4_1_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3322_ (.D(_0094_),
    .CLK(clknet_4_1_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3323_ (.D(_0095_),
    .CLK(clknet_4_1_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3324_ (.D(_0096_),
    .CLK(clknet_4_1_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3325_ (.D(_0097_),
    .CLK(clknet_4_1_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3326_ (.D(_0098_),
    .CLK(clknet_4_0_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3327_ (.D(_0099_),
    .CLK(clknet_4_1_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3328_ (.D(_0100_),
    .CLK(clknet_4_0_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3329_ (.D(_0101_),
    .CLK(clknet_4_1_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3330_ (.D(_0102_),
    .CLK(clknet_4_0_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3331_ (.D(_0103_),
    .CLK(clknet_4_1_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3332_ (.D(_0104_),
    .CLK(clknet_4_0_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3333_ (.D(_0105_),
    .CLK(clknet_4_4_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3334_ (.D(_0106_),
    .CLK(clknet_4_0_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3335_ (.D(_0107_),
    .CLK(clknet_4_4_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3336_ (.D(_0108_),
    .CLK(clknet_4_7_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3337_ (.D(_0109_),
    .CLK(clknet_4_7_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3338_ (.D(_0110_),
    .CLK(clknet_4_4_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3339_ (.D(_0111_),
    .CLK(clknet_4_7_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3340_ (.D(_0112_),
    .CLK(clknet_4_2_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3341_ (.D(_0113_),
    .CLK(clknet_4_2_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3342_ (.D(_0114_),
    .CLK(clknet_4_2_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3343_ (.D(_0115_),
    .CLK(clknet_4_3_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3344_ (.D(_0116_),
    .CLK(clknet_4_6_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3345_ (.D(_0117_),
    .CLK(clknet_4_7_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3346_ (.D(_0118_),
    .CLK(clknet_4_6_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3347_ (.D(_0119_),
    .CLK(clknet_4_7_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3348_ (.D(_0120_),
    .CLK(clknet_4_6_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3349_ (.D(_0121_),
    .CLK(clknet_4_6_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3350_ (.D(_0122_),
    .CLK(clknet_4_6_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3351_ (.D(_0123_),
    .CLK(clknet_4_6_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3352_ (.D(_0124_),
    .CLK(clknet_4_5_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3353_ (.D(_0125_),
    .CLK(clknet_4_5_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3354_ (.D(_0126_),
    .CLK(clknet_4_4_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _3355_ (.D(_0127_),
    .CLK(clknet_4_5_0_UserCLK_regs),
    .Q(\Inst_RegFile_32x4.mem[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3356_ (.I(\Inst_RegFile_switch_matrix.E1BEG0 ),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3357_ (.I(\Inst_RegFile_switch_matrix.E1BEG1 ),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3358_ (.I(\Inst_RegFile_switch_matrix.E1BEG2 ),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3359_ (.I(\Inst_RegFile_switch_matrix.E1BEG3 ),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3360_ (.I(\Inst_RegFile_switch_matrix.E2BEG0 ),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3361_ (.I(\Inst_RegFile_switch_matrix.E2BEG1 ),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3362_ (.I(\Inst_RegFile_switch_matrix.E2BEG2 ),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3363_ (.I(\Inst_RegFile_switch_matrix.E2BEG3 ),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3364_ (.I(\Inst_RegFile_switch_matrix.E2BEG4 ),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3365_ (.I(\Inst_RegFile_switch_matrix.E2BEG5 ),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3366_ (.I(\Inst_RegFile_switch_matrix.E2BEG6 ),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3367_ (.I(\Inst_RegFile_switch_matrix.E2BEG7 ),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3368_ (.I(E2MID[0]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3369_ (.I(E2MID[1]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3370_ (.I(E2MID[2]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3371_ (.I(E2MID[3]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3372_ (.I(E2MID[4]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3373_ (.I(E2MID[5]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3374_ (.I(E2MID[6]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3375_ (.I(E2MID[7]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3376_ (.I(E6END[2]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3377_ (.I(E6END[3]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3378_ (.I(E6END[4]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3379_ (.I(E6END[5]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3380_ (.I(E6END[6]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3381_ (.I(E6END[7]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3382_ (.I(E6END[8]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3383_ (.I(E6END[9]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3384_ (.I(E6END[10]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3385_ (.I(E6END[11]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3386_ (.I(\Inst_RegFile_switch_matrix.E6BEG0 ),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3387_ (.I(\Inst_RegFile_switch_matrix.E6BEG1 ),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3388_ (.I(EE4END[4]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3389_ (.I(EE4END[5]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3390_ (.I(EE4END[6]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3391_ (.I(EE4END[7]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3392_ (.I(EE4END[8]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3393_ (.I(EE4END[9]),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3394_ (.I(EE4END[10]),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3395_ (.I(EE4END[11]),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3396_ (.I(EE4END[12]),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3397_ (.I(EE4END[13]),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3398_ (.I(EE4END[14]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3399_ (.I(EE4END[15]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3400_ (.I(\Inst_RegFile_switch_matrix.EE4BEG0 ),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3401_ (.I(\Inst_RegFile_switch_matrix.EE4BEG1 ),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3402_ (.I(\Inst_RegFile_switch_matrix.EE4BEG2 ),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3403_ (.I(\Inst_RegFile_switch_matrix.EE4BEG3 ),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3404_ (.I(FrameData[0]),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3405_ (.I(FrameData[1]),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3406_ (.I(FrameData[2]),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3407_ (.I(FrameData[3]),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3408_ (.I(FrameData[4]),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3409_ (.I(FrameData[5]),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3410_ (.I(FrameData[6]),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3411_ (.I(FrameData[7]),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3412_ (.I(FrameData[8]),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3413_ (.I(FrameData[9]),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3414_ (.I(FrameData[10]),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3415_ (.I(FrameData[11]),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3416_ (.I(FrameData[12]),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3417_ (.I(FrameData[13]),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3418_ (.I(FrameData[14]),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3419_ (.I(FrameData[15]),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3420_ (.I(FrameData[16]),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3421_ (.I(FrameData[17]),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3422_ (.I(FrameData[18]),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3423_ (.I(FrameData[19]),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3424_ (.I(FrameData[20]),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3425_ (.I(FrameData[21]),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3426_ (.I(FrameData[22]),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3427_ (.I(FrameData[23]),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3428_ (.I(FrameData[24]),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3429_ (.I(FrameData[25]),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3430_ (.I(FrameData[26]),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3431_ (.I(FrameData[27]),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3432_ (.I(FrameData[28]),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3433_ (.I(FrameData[29]),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3434_ (.I(FrameData[30]),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3435_ (.I(FrameData[31]),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3436_ (.I(FrameStrobe[0]),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3437_ (.I(FrameStrobe[1]),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3438_ (.I(FrameStrobe[2]),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3439_ (.I(FrameStrobe[3]),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3440_ (.I(FrameStrobe[4]),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3441_ (.I(FrameStrobe[5]),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3442_ (.I(FrameStrobe[6]),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3443_ (.I(FrameStrobe[7]),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3444_ (.I(FrameStrobe[8]),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3445_ (.I(FrameStrobe[9]),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3446_ (.I(FrameStrobe[10]),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3447_ (.I(FrameStrobe[11]),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3448_ (.I(FrameStrobe[12]),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3449_ (.I(FrameStrobe[13]),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3450_ (.I(FrameStrobe[14]),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3451_ (.I(FrameStrobe[15]),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3452_ (.I(FrameStrobe[16]),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3453_ (.I(FrameStrobe[17]),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3454_ (.I(FrameStrobe[18]),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3455_ (.I(FrameStrobe[19]),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3456_ (.I(\Inst_RegFile_switch_matrix.N1BEG0 ),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3457_ (.I(\Inst_RegFile_switch_matrix.N1BEG1 ),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3458_ (.I(\Inst_RegFile_switch_matrix.N1BEG2 ),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3459_ (.I(\Inst_RegFile_switch_matrix.N1BEG3 ),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3460_ (.I(\Inst_RegFile_switch_matrix.JN2BEG0 ),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3461_ (.I(\Inst_RegFile_switch_matrix.JN2BEG1 ),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3462_ (.I(\Inst_RegFile_switch_matrix.JN2BEG2 ),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3463_ (.I(\Inst_RegFile_switch_matrix.JN2BEG3 ),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3464_ (.I(\Inst_RegFile_switch_matrix.JN2BEG4 ),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3465_ (.I(\Inst_RegFile_switch_matrix.JN2BEG5 ),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3466_ (.I(\Inst_RegFile_switch_matrix.JN2BEG6 ),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3467_ (.I(\Inst_RegFile_switch_matrix.JN2BEG7 ),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3468_ (.I(N2MID[0]),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3469_ (.I(N2MID[1]),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3470_ (.I(N2MID[2]),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3471_ (.I(N2MID[3]),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3472_ (.I(N2MID[4]),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3473_ (.I(N2MID[5]),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3474_ (.I(N2MID[6]),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3475_ (.I(N2MID[7]),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3476_ (.I(N4END[4]),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3477_ (.I(N4END[5]),
    .Z(net128));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3478_ (.I(N4END[6]),
    .Z(net129));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3479_ (.I(N4END[7]),
    .Z(net130));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3480_ (.I(N4END[8]),
    .Z(net131));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3481_ (.I(N4END[9]),
    .Z(net132));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3482_ (.I(N4END[10]),
    .Z(net133));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3483_ (.I(N4END[11]),
    .Z(net134));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3484_ (.I(N4END[12]),
    .Z(net135));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3485_ (.I(N4END[13]),
    .Z(net136));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3486_ (.I(N4END[14]),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3487_ (.I(N4END[15]),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3488_ (.I(\Inst_RegFile_switch_matrix.N4BEG0 ),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3489_ (.I(\Inst_RegFile_switch_matrix.N4BEG1 ),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3490_ (.I(\Inst_RegFile_switch_matrix.N4BEG2 ),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3491_ (.I(\Inst_RegFile_switch_matrix.N4BEG3 ),
    .Z(net127));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3492_ (.I(NN4END[4]),
    .Z(net137));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3493_ (.I(NN4END[5]),
    .Z(net144));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3494_ (.I(NN4END[6]),
    .Z(net145));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3495_ (.I(NN4END[7]),
    .Z(net146));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3496_ (.I(NN4END[8]),
    .Z(net147));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3497_ (.I(NN4END[9]),
    .Z(net148));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3498_ (.I(NN4END[10]),
    .Z(net149));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3499_ (.I(NN4END[11]),
    .Z(net150));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3500_ (.I(NN4END[12]),
    .Z(net151));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3501_ (.I(NN4END[13]),
    .Z(net152));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3502_ (.I(NN4END[14]),
    .Z(net138));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3503_ (.I(NN4END[15]),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3504_ (.I(\Inst_RegFile_switch_matrix.NN4BEG0 ),
    .Z(net140));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3505_ (.I(\Inst_RegFile_switch_matrix.NN4BEG1 ),
    .Z(net141));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3506_ (.I(\Inst_RegFile_switch_matrix.NN4BEG2 ),
    .Z(net142));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3507_ (.I(\Inst_RegFile_switch_matrix.NN4BEG3 ),
    .Z(net143));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3508_ (.I(\Inst_RegFile_switch_matrix.S1BEG0 ),
    .Z(net153));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3509_ (.I(\Inst_RegFile_switch_matrix.S1BEG1 ),
    .Z(net154));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3510_ (.I(\Inst_RegFile_switch_matrix.S1BEG2 ),
    .Z(net155));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3511_ (.I(\Inst_RegFile_switch_matrix.S1BEG3 ),
    .Z(net156));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3512_ (.I(\Inst_RegFile_switch_matrix.JS2BEG0 ),
    .Z(net157));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3513_ (.I(\Inst_RegFile_switch_matrix.JS2BEG1 ),
    .Z(net158));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3514_ (.I(\Inst_RegFile_switch_matrix.JS2BEG2 ),
    .Z(net159));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3515_ (.I(\Inst_RegFile_switch_matrix.JS2BEG3 ),
    .Z(net160));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3516_ (.I(\Inst_RegFile_switch_matrix.JS2BEG4 ),
    .Z(net161));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3517_ (.I(\Inst_RegFile_switch_matrix.JS2BEG5 ),
    .Z(net162));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3518_ (.I(\Inst_RegFile_switch_matrix.JS2BEG6 ),
    .Z(net163));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3519_ (.I(\Inst_RegFile_switch_matrix.JS2BEG7 ),
    .Z(net164));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3520_ (.I(S2MID[0]),
    .Z(net165));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3521_ (.I(S2MID[1]),
    .Z(net166));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3522_ (.I(S2MID[2]),
    .Z(net167));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3523_ (.I(S2MID[3]),
    .Z(net168));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3524_ (.I(S2MID[4]),
    .Z(net169));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3525_ (.I(S2MID[5]),
    .Z(net170));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3526_ (.I(S2MID[6]),
    .Z(net171));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3527_ (.I(S2MID[7]),
    .Z(net172));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3528_ (.I(S4END[4]),
    .Z(net173));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3529_ (.I(S4END[5]),
    .Z(net180));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3530_ (.I(S4END[6]),
    .Z(net181));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3531_ (.I(S4END[7]),
    .Z(net182));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3532_ (.I(S4END[8]),
    .Z(net183));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3533_ (.I(S4END[9]),
    .Z(net184));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3534_ (.I(S4END[10]),
    .Z(net185));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3535_ (.I(S4END[11]),
    .Z(net186));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3536_ (.I(S4END[12]),
    .Z(net187));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3537_ (.I(S4END[13]),
    .Z(net188));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3538_ (.I(S4END[14]),
    .Z(net174));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3539_ (.I(S4END[15]),
    .Z(net175));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3540_ (.I(\Inst_RegFile_switch_matrix.S4BEG0 ),
    .Z(net176));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3541_ (.I(\Inst_RegFile_switch_matrix.S4BEG1 ),
    .Z(net177));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3542_ (.I(\Inst_RegFile_switch_matrix.S4BEG2 ),
    .Z(net178));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3543_ (.I(\Inst_RegFile_switch_matrix.S4BEG3 ),
    .Z(net179));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3544_ (.I(SS4END[4]),
    .Z(net189));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3545_ (.I(SS4END[5]),
    .Z(net196));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3546_ (.I(SS4END[6]),
    .Z(net197));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3547_ (.I(SS4END[7]),
    .Z(net198));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3548_ (.I(SS4END[8]),
    .Z(net199));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3549_ (.I(SS4END[9]),
    .Z(net200));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3550_ (.I(SS4END[10]),
    .Z(net201));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3551_ (.I(SS4END[11]),
    .Z(net202));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3552_ (.I(SS4END[12]),
    .Z(net203));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3553_ (.I(SS4END[13]),
    .Z(net204));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3554_ (.I(SS4END[14]),
    .Z(net190));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3555_ (.I(SS4END[15]),
    .Z(net191));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3556_ (.I(\Inst_RegFile_switch_matrix.SS4BEG0 ),
    .Z(net192));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3557_ (.I(\Inst_RegFile_switch_matrix.SS4BEG1 ),
    .Z(net193));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3558_ (.I(\Inst_RegFile_switch_matrix.SS4BEG2 ),
    .Z(net194));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3559_ (.I(\Inst_RegFile_switch_matrix.SS4BEG3 ),
    .Z(net195));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3560_ (.I(clknet_1_0__leaf_UserCLK),
    .Z(net205));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3561_ (.I(\Inst_RegFile_switch_matrix.W1BEG0 ),
    .Z(net206));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3562_ (.I(\Inst_RegFile_switch_matrix.W1BEG1 ),
    .Z(net207));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3563_ (.I(\Inst_RegFile_switch_matrix.W1BEG2 ),
    .Z(net208));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3564_ (.I(\Inst_RegFile_switch_matrix.W1BEG3 ),
    .Z(net209));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3565_ (.I(\Inst_RegFile_switch_matrix.JW2BEG0 ),
    .Z(net210));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3566_ (.I(\Inst_RegFile_switch_matrix.JW2BEG1 ),
    .Z(net211));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3567_ (.I(\Inst_RegFile_switch_matrix.JW2BEG2 ),
    .Z(net212));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3568_ (.I(\Inst_RegFile_switch_matrix.JW2BEG3 ),
    .Z(net213));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3569_ (.I(\Inst_RegFile_switch_matrix.JW2BEG4 ),
    .Z(net214));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3570_ (.I(\Inst_RegFile_switch_matrix.JW2BEG5 ),
    .Z(net215));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3571_ (.I(\Inst_RegFile_switch_matrix.JW2BEG6 ),
    .Z(net216));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3572_ (.I(\Inst_RegFile_switch_matrix.JW2BEG7 ),
    .Z(net217));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3573_ (.I(W2MID[0]),
    .Z(net218));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3574_ (.I(W2MID[1]),
    .Z(net219));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3575_ (.I(W2MID[2]),
    .Z(net220));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3576_ (.I(W2MID[3]),
    .Z(net221));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3577_ (.I(W2MID[4]),
    .Z(net222));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3578_ (.I(W2MID[5]),
    .Z(net223));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3579_ (.I(W2MID[6]),
    .Z(net224));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3580_ (.I(W2MID[7]),
    .Z(net225));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3581_ (.I(W6END[2]),
    .Z(net226));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3582_ (.I(W6END[3]),
    .Z(net229));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3583_ (.I(W6END[4]),
    .Z(net230));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3584_ (.I(W6END[5]),
    .Z(net231));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3585_ (.I(W6END[6]),
    .Z(net232));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3586_ (.I(W6END[7]),
    .Z(net233));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3587_ (.I(W6END[8]),
    .Z(net234));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3588_ (.I(W6END[9]),
    .Z(net235));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3589_ (.I(W6END[10]),
    .Z(net236));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3590_ (.I(W6END[11]),
    .Z(net237));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3591_ (.I(\Inst_RegFile_switch_matrix.W6BEG0 ),
    .Z(net227));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3592_ (.I(\Inst_RegFile_switch_matrix.W6BEG1 ),
    .Z(net228));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3593_ (.I(WW4END[4]),
    .Z(net238));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3594_ (.I(WW4END[5]),
    .Z(net245));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3595_ (.I(WW4END[6]),
    .Z(net246));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3596_ (.I(WW4END[7]),
    .Z(net247));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3597_ (.I(WW4END[8]),
    .Z(net248));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3598_ (.I(WW4END[9]),
    .Z(net249));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3599_ (.I(WW4END[10]),
    .Z(net250));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3600_ (.I(WW4END[11]),
    .Z(net251));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3601_ (.I(WW4END[12]),
    .Z(net252));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3602_ (.I(WW4END[13]),
    .Z(net253));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3603_ (.I(WW4END[14]),
    .Z(net239));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3604_ (.I(WW4END[15]),
    .Z(net240));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3605_ (.I(\Inst_RegFile_switch_matrix.WW4BEG0 ),
    .Z(net241));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3606_ (.I(\Inst_RegFile_switch_matrix.WW4BEG1 ),
    .Z(net242));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3607_ (.I(\Inst_RegFile_switch_matrix.WW4BEG2 ),
    .Z(net243));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3608_ (.I(\Inst_RegFile_switch_matrix.WW4BEG3 ),
    .Z(net244));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Left_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Left_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Left_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Left_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Left_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Left_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Left_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Left_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Left_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_725 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output1 (.I(net1),
    .Z(E1BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output2 (.I(net2),
    .Z(E1BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output3 (.I(net3),
    .Z(E1BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output4 (.I(net4),
    .Z(E1BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output5 (.I(net5),
    .Z(E2BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output6 (.I(net6),
    .Z(E2BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output7 (.I(net7),
    .Z(E2BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output8 (.I(net8),
    .Z(E2BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output9 (.I(net9),
    .Z(E2BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output10 (.I(net10),
    .Z(E2BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output11 (.I(net11),
    .Z(E2BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output12 (.I(net12),
    .Z(E2BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output13 (.I(net13),
    .Z(E2BEGb[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output14 (.I(net14),
    .Z(E2BEGb[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output15 (.I(net15),
    .Z(E2BEGb[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output16 (.I(net16),
    .Z(E2BEGb[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output17 (.I(net17),
    .Z(E2BEGb[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output18 (.I(net18),
    .Z(E2BEGb[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output19 (.I(net19),
    .Z(E2BEGb[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output20 (.I(net20),
    .Z(E2BEGb[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output21 (.I(net21),
    .Z(E6BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output22 (.I(net22),
    .Z(E6BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output23 (.I(net23),
    .Z(E6BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output24 (.I(net24),
    .Z(E6BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output25 (.I(net25),
    .Z(E6BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output26 (.I(net26),
    .Z(E6BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output27 (.I(net27),
    .Z(E6BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output28 (.I(net28),
    .Z(E6BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output29 (.I(net29),
    .Z(E6BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output30 (.I(net30),
    .Z(E6BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output31 (.I(net31),
    .Z(E6BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output32 (.I(net32),
    .Z(E6BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output33 (.I(net33),
    .Z(EE4BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output34 (.I(net34),
    .Z(EE4BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output35 (.I(net35),
    .Z(EE4BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output36 (.I(net36),
    .Z(EE4BEG[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output37 (.I(net37),
    .Z(EE4BEG[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output38 (.I(net38),
    .Z(EE4BEG[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output39 (.I(net39),
    .Z(EE4BEG[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output40 (.I(net40),
    .Z(EE4BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output41 (.I(net41),
    .Z(EE4BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output42 (.I(net42),
    .Z(EE4BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output43 (.I(net43),
    .Z(EE4BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output44 (.I(net44),
    .Z(EE4BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output45 (.I(net45),
    .Z(EE4BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output46 (.I(net46),
    .Z(EE4BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output47 (.I(net47),
    .Z(EE4BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output48 (.I(net48),
    .Z(EE4BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output49 (.I(net49),
    .Z(FrameData_O[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output50 (.I(net50),
    .Z(FrameData_O[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output51 (.I(net51),
    .Z(FrameData_O[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output52 (.I(net52),
    .Z(FrameData_O[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output53 (.I(net53),
    .Z(FrameData_O[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output54 (.I(net54),
    .Z(FrameData_O[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output55 (.I(net55),
    .Z(FrameData_O[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output56 (.I(net56),
    .Z(FrameData_O[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output57 (.I(net57),
    .Z(FrameData_O[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output58 (.I(net58),
    .Z(FrameData_O[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output59 (.I(net59),
    .Z(FrameData_O[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output60 (.I(net60),
    .Z(FrameData_O[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output61 (.I(net61),
    .Z(FrameData_O[20]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output62 (.I(net62),
    .Z(FrameData_O[21]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output63 (.I(net63),
    .Z(FrameData_O[22]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output64 (.I(net64),
    .Z(FrameData_O[23]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output65 (.I(net65),
    .Z(FrameData_O[24]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output66 (.I(net66),
    .Z(FrameData_O[25]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output67 (.I(net67),
    .Z(FrameData_O[26]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output68 (.I(net68),
    .Z(FrameData_O[27]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output69 (.I(net69),
    .Z(FrameData_O[28]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output70 (.I(net70),
    .Z(FrameData_O[29]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output71 (.I(net71),
    .Z(FrameData_O[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output72 (.I(net72),
    .Z(FrameData_O[30]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output73 (.I(net73),
    .Z(FrameData_O[31]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output74 (.I(net74),
    .Z(FrameData_O[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output75 (.I(net75),
    .Z(FrameData_O[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output76 (.I(net76),
    .Z(FrameData_O[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output77 (.I(net77),
    .Z(FrameData_O[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output78 (.I(net78),
    .Z(FrameData_O[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output79 (.I(net79),
    .Z(FrameData_O[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output80 (.I(net80),
    .Z(FrameData_O[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output81 (.I(net81),
    .Z(FrameStrobe_O[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output82 (.I(net82),
    .Z(FrameStrobe_O[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output83 (.I(net83),
    .Z(FrameStrobe_O[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output84 (.I(net84),
    .Z(FrameStrobe_O[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output85 (.I(net85),
    .Z(FrameStrobe_O[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output86 (.I(net86),
    .Z(FrameStrobe_O[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output87 (.I(net87),
    .Z(FrameStrobe_O[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output88 (.I(net88),
    .Z(FrameStrobe_O[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output89 (.I(net89),
    .Z(FrameStrobe_O[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output90 (.I(net90),
    .Z(FrameStrobe_O[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output91 (.I(net91),
    .Z(FrameStrobe_O[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output92 (.I(net92),
    .Z(FrameStrobe_O[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output93 (.I(net93),
    .Z(FrameStrobe_O[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output94 (.I(net94),
    .Z(FrameStrobe_O[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output95 (.I(net95),
    .Z(FrameStrobe_O[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output96 (.I(net96),
    .Z(FrameStrobe_O[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output97 (.I(net97),
    .Z(FrameStrobe_O[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output98 (.I(net98),
    .Z(FrameStrobe_O[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output99 (.I(net99),
    .Z(FrameStrobe_O[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output100 (.I(net100),
    .Z(FrameStrobe_O[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output101 (.I(net101),
    .Z(N1BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output102 (.I(net102),
    .Z(N1BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output103 (.I(net103),
    .Z(N1BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output104 (.I(net104),
    .Z(N1BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output105 (.I(net105),
    .Z(N2BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output106 (.I(net106),
    .Z(N2BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output107 (.I(net107),
    .Z(N2BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output108 (.I(net108),
    .Z(N2BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output109 (.I(net109),
    .Z(N2BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output110 (.I(net110),
    .Z(N2BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output111 (.I(net111),
    .Z(N2BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output112 (.I(net112),
    .Z(N2BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output113 (.I(net113),
    .Z(N2BEGb[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output114 (.I(net114),
    .Z(N2BEGb[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output115 (.I(net115),
    .Z(N2BEGb[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output116 (.I(net116),
    .Z(N2BEGb[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output117 (.I(net117),
    .Z(N2BEGb[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output118 (.I(net118),
    .Z(N2BEGb[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output119 (.I(net119),
    .Z(N2BEGb[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output120 (.I(net120),
    .Z(N2BEGb[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output121 (.I(net121),
    .Z(N4BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output122 (.I(net122),
    .Z(N4BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output123 (.I(net123),
    .Z(N4BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output124 (.I(net124),
    .Z(N4BEG[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output125 (.I(net125),
    .Z(N4BEG[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output126 (.I(net126),
    .Z(N4BEG[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output127 (.I(net127),
    .Z(N4BEG[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output128 (.I(net128),
    .Z(N4BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output129 (.I(net129),
    .Z(N4BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output130 (.I(net130),
    .Z(N4BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output131 (.I(net131),
    .Z(N4BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output132 (.I(net132),
    .Z(N4BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output133 (.I(net133),
    .Z(N4BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output134 (.I(net134),
    .Z(N4BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output135 (.I(net135),
    .Z(N4BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output136 (.I(net136),
    .Z(N4BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output137 (.I(net137),
    .Z(NN4BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output138 (.I(net138),
    .Z(NN4BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output139 (.I(net139),
    .Z(NN4BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output140 (.I(net140),
    .Z(NN4BEG[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output141 (.I(net141),
    .Z(NN4BEG[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output142 (.I(net142),
    .Z(NN4BEG[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output143 (.I(net143),
    .Z(NN4BEG[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output144 (.I(net144),
    .Z(NN4BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output145 (.I(net145),
    .Z(NN4BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output146 (.I(net146),
    .Z(NN4BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output147 (.I(net147),
    .Z(NN4BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output148 (.I(net148),
    .Z(NN4BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output149 (.I(net149),
    .Z(NN4BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output150 (.I(net150),
    .Z(NN4BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output151 (.I(net151),
    .Z(NN4BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output152 (.I(net152),
    .Z(NN4BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output153 (.I(net153),
    .Z(S1BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output154 (.I(net154),
    .Z(S1BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output155 (.I(net155),
    .Z(S1BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output156 (.I(net156),
    .Z(S1BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output157 (.I(net157),
    .Z(S2BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output158 (.I(net158),
    .Z(S2BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output159 (.I(net159),
    .Z(S2BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output160 (.I(net160),
    .Z(S2BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output161 (.I(net161),
    .Z(S2BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output162 (.I(net162),
    .Z(S2BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output163 (.I(net163),
    .Z(S2BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output164 (.I(net164),
    .Z(S2BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output165 (.I(net165),
    .Z(S2BEGb[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output166 (.I(net166),
    .Z(S2BEGb[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output167 (.I(net167),
    .Z(S2BEGb[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output168 (.I(net168),
    .Z(S2BEGb[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output169 (.I(net169),
    .Z(S2BEGb[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output170 (.I(net170),
    .Z(S2BEGb[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output171 (.I(net171),
    .Z(S2BEGb[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output172 (.I(net172),
    .Z(S2BEGb[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output173 (.I(net173),
    .Z(S4BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output174 (.I(net174),
    .Z(S4BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output175 (.I(net175),
    .Z(S4BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output176 (.I(net176),
    .Z(S4BEG[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output177 (.I(net177),
    .Z(S4BEG[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output178 (.I(net178),
    .Z(S4BEG[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output179 (.I(net179),
    .Z(S4BEG[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output180 (.I(net180),
    .Z(S4BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output181 (.I(net181),
    .Z(S4BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output182 (.I(net182),
    .Z(S4BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output183 (.I(net183),
    .Z(S4BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output184 (.I(net184),
    .Z(S4BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output185 (.I(net185),
    .Z(S4BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output186 (.I(net186),
    .Z(S4BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output187 (.I(net187),
    .Z(S4BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output188 (.I(net188),
    .Z(S4BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output189 (.I(net189),
    .Z(SS4BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output190 (.I(net190),
    .Z(SS4BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output191 (.I(net191),
    .Z(SS4BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output192 (.I(net192),
    .Z(SS4BEG[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output193 (.I(net193),
    .Z(SS4BEG[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output194 (.I(net194),
    .Z(SS4BEG[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output195 (.I(net195),
    .Z(SS4BEG[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output196 (.I(net196),
    .Z(SS4BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output197 (.I(net197),
    .Z(SS4BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output198 (.I(net198),
    .Z(SS4BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output199 (.I(net199),
    .Z(SS4BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output200 (.I(net200),
    .Z(SS4BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output201 (.I(net201),
    .Z(SS4BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output202 (.I(net202),
    .Z(SS4BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output203 (.I(net203),
    .Z(SS4BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output204 (.I(net204),
    .Z(SS4BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output205 (.I(net205),
    .Z(UserCLKo));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output206 (.I(net206),
    .Z(W1BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output207 (.I(net207),
    .Z(W1BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output208 (.I(net208),
    .Z(W1BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output209 (.I(net209),
    .Z(W1BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output210 (.I(net210),
    .Z(W2BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output211 (.I(net211),
    .Z(W2BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output212 (.I(net212),
    .Z(W2BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output213 (.I(net213),
    .Z(W2BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output214 (.I(net214),
    .Z(W2BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output215 (.I(net215),
    .Z(W2BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output216 (.I(net216),
    .Z(W2BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output217 (.I(net217),
    .Z(W2BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output218 (.I(net218),
    .Z(W2BEGb[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output219 (.I(net219),
    .Z(W2BEGb[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output220 (.I(net220),
    .Z(W2BEGb[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output221 (.I(net221),
    .Z(W2BEGb[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output222 (.I(net222),
    .Z(W2BEGb[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output223 (.I(net223),
    .Z(W2BEGb[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output224 (.I(net224),
    .Z(W2BEGb[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output225 (.I(net225),
    .Z(W2BEGb[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output226 (.I(net226),
    .Z(W6BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output227 (.I(net227),
    .Z(W6BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output228 (.I(net228),
    .Z(W6BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output229 (.I(net229),
    .Z(W6BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output230 (.I(net230),
    .Z(W6BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output231 (.I(net231),
    .Z(W6BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output232 (.I(net232),
    .Z(W6BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output233 (.I(net233),
    .Z(W6BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output234 (.I(net234),
    .Z(W6BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output235 (.I(net235),
    .Z(W6BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output236 (.I(net236),
    .Z(W6BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output237 (.I(net237),
    .Z(W6BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output238 (.I(net238),
    .Z(WW4BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output239 (.I(net239),
    .Z(WW4BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output240 (.I(net240),
    .Z(WW4BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output241 (.I(net241),
    .Z(WW4BEG[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output242 (.I(net242),
    .Z(WW4BEG[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output243 (.I(net243),
    .Z(WW4BEG[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output244 (.I(net244),
    .Z(WW4BEG[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output245 (.I(net245),
    .Z(WW4BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output246 (.I(net246),
    .Z(WW4BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output247 (.I(net247),
    .Z(WW4BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output248 (.I(net248),
    .Z(WW4BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output249 (.I(net249),
    .Z(WW4BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output250 (.I(net250),
    .Z(WW4BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output251 (.I(net251),
    .Z(WW4BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output252 (.I(net252),
    .Z(WW4BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output253 (.I(net253),
    .Z(WW4BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_regs_0_UserCLK (.I(UserCLK),
    .Z(UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_UserCLK (.I(UserCLK),
    .Z(clknet_0_UserCLK));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_0__f_UserCLK (.I(clknet_0_UserCLK),
    .Z(clknet_1_0__leaf_UserCLK));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_UserCLK_regs (.I(UserCLK_regs),
    .Z(clknet_0_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_0_0_UserCLK_regs (.I(clknet_0_UserCLK_regs),
    .Z(clknet_4_0_0_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_1_0_UserCLK_regs (.I(clknet_0_UserCLK_regs),
    .Z(clknet_4_1_0_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_2_0_UserCLK_regs (.I(clknet_0_UserCLK_regs),
    .Z(clknet_4_2_0_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_3_0_UserCLK_regs (.I(clknet_0_UserCLK_regs),
    .Z(clknet_4_3_0_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_4_0_UserCLK_regs (.I(clknet_0_UserCLK_regs),
    .Z(clknet_4_4_0_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_5_0_UserCLK_regs (.I(clknet_0_UserCLK_regs),
    .Z(clknet_4_5_0_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_6_0_UserCLK_regs (.I(clknet_0_UserCLK_regs),
    .Z(clknet_4_6_0_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_7_0_UserCLK_regs (.I(clknet_0_UserCLK_regs),
    .Z(clknet_4_7_0_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_8_0_UserCLK_regs (.I(clknet_0_UserCLK_regs),
    .Z(clknet_4_8_0_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_9_0_UserCLK_regs (.I(clknet_0_UserCLK_regs),
    .Z(clknet_4_9_0_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_10_0_UserCLK_regs (.I(clknet_0_UserCLK_regs),
    .Z(clknet_4_10_0_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_11_0_UserCLK_regs (.I(clknet_0_UserCLK_regs),
    .Z(clknet_4_11_0_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_12_0_UserCLK_regs (.I(clknet_0_UserCLK_regs),
    .Z(clknet_4_12_0_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_13_0_UserCLK_regs (.I(clknet_0_UserCLK_regs),
    .Z(clknet_4_13_0_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_14_0_UserCLK_regs (.I(clknet_0_UserCLK_regs),
    .Z(clknet_4_14_0_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_15_0_UserCLK_regs (.I(clknet_0_UserCLK_regs),
    .Z(clknet_4_15_0_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 clkload0 (.I(clknet_4_0_0_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 clkload1 (.I(clknet_4_1_0_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 clkload2 (.I(clknet_4_2_0_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 clkload3 (.I(clknet_4_3_0_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 clkload4 (.I(clknet_4_4_0_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 clkload5 (.I(clknet_4_7_0_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 clkload6 (.I(clknet_4_8_0_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 clkload7 (.I(clknet_4_9_0_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 clkload8 (.I(clknet_4_10_0_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 clkload9 (.I(clknet_4_11_0_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 clkload10 (.I(clknet_4_12_0_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 clkload11 (.I(clknet_4_13_0_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 clkload12 (.I(clknet_4_14_0_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 clkload13 (.I(clknet_4_15_0_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_1 (.I(E6END[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_2 (.I(FrameStrobe[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_3 (.I(FrameStrobe[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_4 (.I(FrameStrobe[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_5 (.I(FrameStrobe[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_6 (.I(FrameStrobe[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_7 (.I(FrameStrobe[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_8 (.I(FrameStrobe[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_9 (.I(N2MID[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_10 (.I(W6END[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_11 (.I(W6END[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_12 (.I(W6END[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_13 (.I(W6END[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_14 (.I(W6END[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_15 (.I(WW4END[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_16 (.I(WW4END[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_17 (.I(WW4END[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_18 (.I(EE4END[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_19 (.I(FrameStrobe[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_20 (.I(W6END[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_21 (.I(WW4END[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_22 (.I(WW4END[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_23 (.I(E6END[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_24 (.I(E6END[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_25 (.I(EE4END[13]));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_560 ();
endmodule
