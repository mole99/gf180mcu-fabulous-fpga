module S_term_SRAM (UserCLK,
    UserCLKo,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N2BEG,
    N2BEGb,
    N4BEG,
    S1END,
    S2END,
    S2MID,
    S4END);
 input UserCLK;
 output UserCLKo;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 output [15:0] N4BEG;
 input [3:0] S1END;
 input [7:0] S2END;
 input [7:0] S2MID;
 input [15:0] S4END;

 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;

 gf180mcu_fd_sc_mcu7t5v0__buf_2 _00_ (.I(FrameData[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _01_ (.I(FrameData[1]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _02_ (.I(FrameData[2]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _03_ (.I(FrameData[3]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _04_ (.I(FrameData[4]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05_ (.I(FrameData[5]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06_ (.I(FrameData[6]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07_ (.I(FrameData[7]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08_ (.I(FrameData[8]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09_ (.I(FrameData[9]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10_ (.I(FrameData[10]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11_ (.I(FrameData[11]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _12_ (.I(FrameData[12]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _13_ (.I(FrameData[13]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _14_ (.I(FrameData[14]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _15_ (.I(FrameData[15]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _16_ (.I(FrameData[16]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _17_ (.I(FrameData[17]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _18_ (.I(FrameData[18]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _19_ (.I(FrameData[19]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _20_ (.I(FrameData[20]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _21_ (.I(FrameData[21]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _22_ (.I(FrameData[22]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _23_ (.I(FrameData[23]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _24_ (.I(FrameData[24]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _25_ (.I(FrameData[25]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _26_ (.I(FrameData[26]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _27_ (.I(FrameData[27]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _28_ (.I(FrameData[28]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _29_ (.I(FrameData[29]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _30_ (.I(FrameData[30]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _31_ (.I(FrameData[31]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _32_ (.I(FrameStrobe[0]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _33_ (.I(FrameStrobe[1]),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _34_ (.I(FrameStrobe[2]),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _35_ (.I(FrameStrobe[3]),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _36_ (.I(FrameStrobe[4]),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _37_ (.I(FrameStrobe[5]),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _38_ (.I(FrameStrobe[6]),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _39_ (.I(FrameStrobe[7]),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _40_ (.I(FrameStrobe[8]),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _41_ (.I(FrameStrobe[9]),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _42_ (.I(FrameStrobe[10]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _43_ (.I(FrameStrobe[11]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _44_ (.I(FrameStrobe[12]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _45_ (.I(FrameStrobe[13]),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _46_ (.I(FrameStrobe[14]),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _47_ (.I(FrameStrobe[15]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _48_ (.I(FrameStrobe[16]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _49_ (.I(FrameStrobe[17]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _50_ (.I(FrameStrobe[18]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _51_ (.I(FrameStrobe[19]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _52_ (.I(S1END[3]),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _53_ (.I(S1END[2]),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _54_ (.I(S1END[1]),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _55_ (.I(S1END[0]),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _56_ (.I(S2MID[7]),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _57_ (.I(S2MID[6]),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _58_ (.I(S2MID[5]),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _59_ (.I(S2MID[4]),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _60_ (.I(S2MID[3]),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _61_ (.I(S2MID[2]),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _62_ (.I(S2MID[1]),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _63_ (.I(S2MID[0]),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _64_ (.I(S2END[7]),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _65_ (.I(S2END[6]),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _66_ (.I(S2END[5]),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _67_ (.I(S2END[4]),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _68_ (.I(S2END[3]),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _69_ (.I(S2END[2]),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _70_ (.I(S2END[1]),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _71_ (.I(S2END[0]),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _72_ (.I(S4END[15]),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _73_ (.I(S4END[14]),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _74_ (.I(S4END[13]),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _75_ (.I(S4END[12]),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _76_ (.I(S4END[11]),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _77_ (.I(S4END[10]),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _78_ (.I(S4END[9]),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _79_ (.I(S4END[8]),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _80_ (.I(S4END[7]),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _81_ (.I(S4END[6]),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _82_ (.I(S4END[5]),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _83_ (.I(S4END[4]),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _84_ (.I(S4END[3]),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _85_ (.I(S4END[2]),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _86_ (.I(S4END[1]),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _87_ (.I(S4END[0]),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _88_ (.I(UserCLK),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_56 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_58 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_59 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_60 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_61 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_62 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_63 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_64 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_65 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_66 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_67 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_68 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_69 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_70 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_71 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_72 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_73 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_74 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_75 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_76 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_77 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_78 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_79 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_80 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_81 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_82 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_83 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_84 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_85 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_86 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_87 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_88 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_89 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_90 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_91 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_92 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_93 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_94 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output1 (.I(net1),
    .Z(FrameData_O[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output2 (.I(net2),
    .Z(FrameData_O[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output3 (.I(net3),
    .Z(FrameData_O[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output4 (.I(net4),
    .Z(FrameData_O[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output5 (.I(net5),
    .Z(FrameData_O[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output6 (.I(net6),
    .Z(FrameData_O[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output7 (.I(net7),
    .Z(FrameData_O[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output8 (.I(net8),
    .Z(FrameData_O[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output9 (.I(net9),
    .Z(FrameData_O[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output10 (.I(net10),
    .Z(FrameData_O[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output11 (.I(net11),
    .Z(FrameData_O[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output12 (.I(net12),
    .Z(FrameData_O[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output13 (.I(net13),
    .Z(FrameData_O[20]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output14 (.I(net14),
    .Z(FrameData_O[21]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output15 (.I(net15),
    .Z(FrameData_O[22]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output16 (.I(net16),
    .Z(FrameData_O[23]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output17 (.I(net17),
    .Z(FrameData_O[24]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output18 (.I(net18),
    .Z(FrameData_O[25]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output19 (.I(net19),
    .Z(FrameData_O[26]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output20 (.I(net20),
    .Z(FrameData_O[27]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output21 (.I(net21),
    .Z(FrameData_O[28]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output22 (.I(net22),
    .Z(FrameData_O[29]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output23 (.I(net23),
    .Z(FrameData_O[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output24 (.I(net24),
    .Z(FrameData_O[30]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output25 (.I(net25),
    .Z(FrameData_O[31]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output26 (.I(net26),
    .Z(FrameData_O[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output27 (.I(net27),
    .Z(FrameData_O[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output28 (.I(net28),
    .Z(FrameData_O[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output29 (.I(net29),
    .Z(FrameData_O[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output30 (.I(net30),
    .Z(FrameData_O[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output31 (.I(net31),
    .Z(FrameData_O[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output32 (.I(net32),
    .Z(FrameData_O[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output33 (.I(net33),
    .Z(FrameStrobe_O[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output34 (.I(net34),
    .Z(FrameStrobe_O[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output35 (.I(net35),
    .Z(FrameStrobe_O[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output36 (.I(net36),
    .Z(FrameStrobe_O[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output37 (.I(net37),
    .Z(FrameStrobe_O[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output38 (.I(net38),
    .Z(FrameStrobe_O[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output39 (.I(net39),
    .Z(FrameStrobe_O[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output40 (.I(net40),
    .Z(FrameStrobe_O[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output41 (.I(net41),
    .Z(FrameStrobe_O[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output42 (.I(net42),
    .Z(FrameStrobe_O[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output43 (.I(net43),
    .Z(FrameStrobe_O[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output44 (.I(net44),
    .Z(FrameStrobe_O[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output45 (.I(net45),
    .Z(FrameStrobe_O[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output46 (.I(net46),
    .Z(FrameStrobe_O[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output47 (.I(net47),
    .Z(FrameStrobe_O[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output48 (.I(net48),
    .Z(FrameStrobe_O[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output49 (.I(net49),
    .Z(FrameStrobe_O[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output50 (.I(net50),
    .Z(FrameStrobe_O[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output51 (.I(net51),
    .Z(FrameStrobe_O[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output52 (.I(net52),
    .Z(FrameStrobe_O[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output53 (.I(net53),
    .Z(N1BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output54 (.I(net54),
    .Z(N1BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output55 (.I(net55),
    .Z(N1BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output56 (.I(net56),
    .Z(N1BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output57 (.I(net57),
    .Z(N2BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output58 (.I(net58),
    .Z(N2BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output59 (.I(net59),
    .Z(N2BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output60 (.I(net60),
    .Z(N2BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output61 (.I(net61),
    .Z(N2BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output62 (.I(net62),
    .Z(N2BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output63 (.I(net63),
    .Z(N2BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output64 (.I(net64),
    .Z(N2BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output65 (.I(net65),
    .Z(N2BEGb[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output66 (.I(net66),
    .Z(N2BEGb[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output67 (.I(net67),
    .Z(N2BEGb[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output68 (.I(net68),
    .Z(N2BEGb[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output69 (.I(net69),
    .Z(N2BEGb[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output70 (.I(net70),
    .Z(N2BEGb[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output71 (.I(net71),
    .Z(N2BEGb[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output72 (.I(net72),
    .Z(N2BEGb[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output73 (.I(net73),
    .Z(N4BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output74 (.I(net74),
    .Z(N4BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output75 (.I(net75),
    .Z(N4BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output76 (.I(net76),
    .Z(N4BEG[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output77 (.I(net77),
    .Z(N4BEG[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output78 (.I(net78),
    .Z(N4BEG[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output79 (.I(net79),
    .Z(N4BEG[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output80 (.I(net80),
    .Z(N4BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output81 (.I(net81),
    .Z(N4BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output82 (.I(net82),
    .Z(N4BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output83 (.I(net83),
    .Z(N4BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output84 (.I(net84),
    .Z(N4BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output85 (.I(net85),
    .Z(N4BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output86 (.I(net86),
    .Z(N4BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output87 (.I(net87),
    .Z(N4BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output88 (.I(net88),
    .Z(N4BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output89 (.I(net89),
    .Z(UserCLKo));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__00__I (.I(FrameData[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10__I (.I(FrameData[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11__I (.I(FrameData[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12__I (.I(FrameData[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__13__I (.I(FrameData[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__14__I (.I(FrameData[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__15__I (.I(FrameData[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__16__I (.I(FrameData[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__17__I (.I(FrameData[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__18__I (.I(FrameData[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__19__I (.I(FrameData[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__01__I (.I(FrameData[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__20__I (.I(FrameData[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__21__I (.I(FrameData[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__22__I (.I(FrameData[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__23__I (.I(FrameData[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__24__I (.I(FrameData[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__25__I (.I(FrameData[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__26__I (.I(FrameData[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__27__I (.I(FrameData[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__28__I (.I(FrameData[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__29__I (.I(FrameData[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__02__I (.I(FrameData[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__30__I (.I(FrameData[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__31__I (.I(FrameData[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__03__I (.I(FrameData[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04__I (.I(FrameData[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05__I (.I(FrameData[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06__I (.I(FrameData[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07__I (.I(FrameData[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08__I (.I(FrameData[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09__I (.I(FrameData[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__32__I (.I(FrameStrobe[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__42__I (.I(FrameStrobe[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__43__I (.I(FrameStrobe[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__44__I (.I(FrameStrobe[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__45__I (.I(FrameStrobe[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__46__I (.I(FrameStrobe[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__47__I (.I(FrameStrobe[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__48__I (.I(FrameStrobe[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__49__I (.I(FrameStrobe[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__50__I (.I(FrameStrobe[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__51__I (.I(FrameStrobe[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__33__I (.I(FrameStrobe[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__34__I (.I(FrameStrobe[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__35__I (.I(FrameStrobe[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__36__I (.I(FrameStrobe[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__37__I (.I(FrameStrobe[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__38__I (.I(FrameStrobe[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__39__I (.I(FrameStrobe[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__40__I (.I(FrameStrobe[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__41__I (.I(FrameStrobe[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__55__I (.I(S1END[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__54__I (.I(S1END[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__53__I (.I(S1END[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__52__I (.I(S1END[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__71__I (.I(S2END[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__70__I (.I(S2END[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__69__I (.I(S2END[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__68__I (.I(S2END[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__67__I (.I(S2END[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__66__I (.I(S2END[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__65__I (.I(S2END[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__64__I (.I(S2END[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__63__I (.I(S2MID[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__62__I (.I(S2MID[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__61__I (.I(S2MID[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__60__I (.I(S2MID[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__59__I (.I(S2MID[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__58__I (.I(S2MID[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__57__I (.I(S2MID[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__56__I (.I(S2MID[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__87__I (.I(S4END[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__77__I (.I(S4END[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__76__I (.I(S4END[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__75__I (.I(S4END[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__74__I (.I(S4END[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__73__I (.I(S4END[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__72__I (.I(S4END[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__86__I (.I(S4END[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__85__I (.I(S4END[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__84__I (.I(S4END[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__83__I (.I(S4END[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__82__I (.I(S4END[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__81__I (.I(S4END[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__80__I (.I(S4END[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__79__I (.I(S4END[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__78__I (.I(S4END[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__88__I (.I(UserCLK));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_268 ();
endmodule
