module \$_DLATCH_P_ (input E, input D, output Q);
    gf180mcu_fd_sc_mcu7t5v0__latq_1 _TECHMAP_DLATCH_P (
        .E  (E),
        .D  (D),
        .Q  (Q)
    );
endmodule








//gf180mcu_fd_sc_mcu7t5v0__latrnq_1( E, D, RN, Q

//gf180mcu_fd_sc_mcu7t5v0__latrsnq_1 ( E, D, RN, SETN, Q

//gf180mcu_fd_sc_mcu7t5v0__latsnq_1 ( E, D, SETN, Q,
