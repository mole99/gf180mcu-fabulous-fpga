magic
tech gf180mcuD
magscale 1 10
timestamp 1764971401
<< metal1 >>
rect 672 56474 27888 56508
rect 672 56422 3806 56474
rect 3858 56422 3910 56474
rect 3962 56422 4014 56474
rect 4066 56422 23806 56474
rect 23858 56422 23910 56474
rect 23962 56422 24014 56474
rect 24066 56422 27888 56474
rect 672 56388 27888 56422
rect 3614 56306 3666 56318
rect 3614 56242 3666 56254
rect 5182 56306 5234 56318
rect 5182 56242 5234 56254
rect 8990 56306 9042 56318
rect 8990 56242 9042 56254
rect 10558 56306 10610 56318
rect 10558 56242 10610 56254
rect 13022 56306 13074 56318
rect 13022 56242 13074 56254
rect 14590 56306 14642 56318
rect 14590 56242 14642 56254
rect 16494 56306 16546 56318
rect 16494 56242 16546 56254
rect 18510 56306 18562 56318
rect 18510 56242 18562 56254
rect 20302 56306 20354 56318
rect 20302 56242 20354 56254
rect 22206 56306 22258 56318
rect 22206 56242 22258 56254
rect 24446 56306 24498 56318
rect 24446 56242 24498 56254
rect 26014 56306 26066 56318
rect 26014 56242 26066 56254
rect 7410 56142 7422 56194
rect 7474 56142 7486 56194
rect 7858 56030 7870 56082
rect 7922 56030 7934 56082
rect 21746 56030 21758 56082
rect 21810 56030 21822 56082
rect 1026 55918 1038 55970
rect 1090 55918 1102 55970
rect 3042 55918 3054 55970
rect 3106 55918 3118 55970
rect 6178 55918 6190 55970
rect 6242 55918 6254 55970
rect 9986 55918 9998 55970
rect 10050 55918 10062 55970
rect 11554 55918 11566 55970
rect 11618 55918 11630 55970
rect 14018 55918 14030 55970
rect 14082 55918 14094 55970
rect 15586 55918 15598 55970
rect 15650 55918 15662 55970
rect 17490 55918 17502 55970
rect 17554 55918 17566 55970
rect 19506 55918 19518 55970
rect 19570 55918 19582 55970
rect 21298 55918 21310 55970
rect 21362 55918 21374 55970
rect 23874 55918 23886 55970
rect 23938 55918 23950 55970
rect 25442 55918 25454 55970
rect 25506 55918 25518 55970
rect 1374 55858 1426 55870
rect 1374 55794 1426 55806
rect 672 55690 27888 55724
rect 672 55638 4466 55690
rect 4518 55638 4570 55690
rect 4622 55638 4674 55690
rect 4726 55638 24466 55690
rect 24518 55638 24570 55690
rect 24622 55638 24674 55690
rect 24726 55638 27888 55690
rect 672 55604 27888 55638
rect 22990 55522 23042 55534
rect 22990 55458 23042 55470
rect 21634 55358 21646 55410
rect 21698 55358 21710 55410
rect 20526 55298 20578 55310
rect 3490 55246 3502 55298
rect 3554 55246 3566 55298
rect 6290 55246 6302 55298
rect 6354 55246 6366 55298
rect 12898 55246 12910 55298
rect 12962 55246 12974 55298
rect 18274 55246 18286 55298
rect 18338 55246 18350 55298
rect 20066 55246 20078 55298
rect 20130 55246 20142 55298
rect 20850 55246 20862 55298
rect 20914 55246 20926 55298
rect 22418 55246 22430 55298
rect 22482 55246 22494 55298
rect 24658 55246 24670 55298
rect 24722 55246 24734 55298
rect 26450 55246 26462 55298
rect 26514 55246 26526 55298
rect 20526 55234 20578 55246
rect 2494 55186 2546 55198
rect 2494 55122 2546 55134
rect 6862 55186 6914 55198
rect 6862 55122 6914 55134
rect 11902 55186 11954 55198
rect 11902 55122 11954 55134
rect 17278 55186 17330 55198
rect 17278 55122 17330 55134
rect 25678 55074 25730 55086
rect 25678 55010 25730 55022
rect 27246 55074 27298 55086
rect 27246 55010 27298 55022
rect 672 54906 27888 54940
rect 672 54854 3806 54906
rect 3858 54854 3910 54906
rect 3962 54854 4014 54906
rect 4066 54854 23806 54906
rect 23858 54854 23910 54906
rect 23962 54854 24014 54906
rect 24066 54854 27888 54906
rect 672 54820 27888 54854
rect 22542 54738 22594 54750
rect 22542 54674 22594 54686
rect 23774 54738 23826 54750
rect 23774 54674 23826 54686
rect 19506 54574 19518 54626
rect 19570 54574 19582 54626
rect 25554 54574 25566 54626
rect 25618 54574 25630 54626
rect 21198 54514 21250 54526
rect 24098 54462 24110 54514
rect 24162 54462 24174 54514
rect 21198 54450 21250 54462
rect 21522 54350 21534 54402
rect 21586 54350 21598 54402
rect 24658 54350 24670 54402
rect 24722 54350 24734 54402
rect 26226 54350 26238 54402
rect 26290 54350 26302 54402
rect 27010 54350 27022 54402
rect 27074 54350 27086 54402
rect 19070 54290 19122 54302
rect 19070 54226 19122 54238
rect 20638 54290 20690 54302
rect 20638 54226 20690 54238
rect 672 54122 27888 54156
rect 672 54070 4466 54122
rect 4518 54070 4570 54122
rect 4622 54070 4674 54122
rect 4726 54070 24466 54122
rect 24518 54070 24570 54122
rect 24622 54070 24674 54122
rect 24726 54070 27888 54122
rect 672 54036 27888 54070
rect 21870 53842 21922 53854
rect 21870 53778 21922 53790
rect 22306 53678 22318 53730
rect 22370 53678 22382 53730
rect 22754 53678 22766 53730
rect 22818 53678 22830 53730
rect 24658 53678 24670 53730
rect 24722 53678 24734 53730
rect 26226 53678 26238 53730
rect 26290 53678 26302 53730
rect 23774 53618 23826 53630
rect 23774 53554 23826 53566
rect 25678 53618 25730 53630
rect 25678 53554 25730 53566
rect 27246 53506 27298 53518
rect 27246 53442 27298 53454
rect 672 53338 27888 53372
rect 672 53286 3806 53338
rect 3858 53286 3910 53338
rect 3962 53286 4014 53338
rect 4066 53286 23806 53338
rect 23858 53286 23910 53338
rect 23962 53286 24014 53338
rect 24066 53286 27888 53338
rect 672 53252 27888 53286
rect 24110 53170 24162 53182
rect 24110 53106 24162 53118
rect 27122 53006 27134 53058
rect 27186 53006 27198 53058
rect 23090 52782 23102 52834
rect 23154 52782 23166 52834
rect 24658 52782 24670 52834
rect 24722 52782 24734 52834
rect 25442 52782 25454 52834
rect 25506 52782 25518 52834
rect 26226 52782 26238 52834
rect 26290 52782 26302 52834
rect 672 52554 27888 52588
rect 672 52502 4466 52554
rect 4518 52502 4570 52554
rect 4622 52502 4674 52554
rect 4726 52502 24466 52554
rect 24518 52502 24570 52554
rect 24622 52502 24674 52554
rect 24726 52502 27888 52554
rect 672 52468 27888 52502
rect 21422 52386 21474 52398
rect 21422 52322 21474 52334
rect 21982 52274 22034 52286
rect 24658 52222 24670 52274
rect 24722 52222 24734 52274
rect 21982 52210 22034 52222
rect 22754 52110 22766 52162
rect 22818 52110 22830 52162
rect 26226 52110 26238 52162
rect 26290 52110 26302 52162
rect 23650 51998 23662 52050
rect 23714 51998 23726 52050
rect 25678 51938 25730 51950
rect 25678 51874 25730 51886
rect 27246 51938 27298 51950
rect 27246 51874 27298 51886
rect 672 51770 27888 51804
rect 672 51718 3806 51770
rect 3858 51718 3910 51770
rect 3962 51718 4014 51770
rect 4066 51718 23806 51770
rect 23858 51718 23910 51770
rect 23962 51718 24014 51770
rect 24066 51718 27888 51770
rect 672 51684 27888 51718
rect 25678 51602 25730 51614
rect 25678 51538 25730 51550
rect 26338 51326 26350 51378
rect 26402 51326 26414 51378
rect 24658 51214 24670 51266
rect 24722 51214 24734 51266
rect 27010 51214 27022 51266
rect 27074 51214 27086 51266
rect 672 50986 27888 51020
rect 672 50934 4466 50986
rect 4518 50934 4570 50986
rect 4622 50934 4674 50986
rect 4726 50934 24466 50986
rect 24518 50934 24570 50986
rect 24622 50934 24674 50986
rect 24726 50934 27888 50986
rect 672 50900 27888 50934
rect 23998 50594 24050 50606
rect 24658 50542 24670 50594
rect 24722 50542 24734 50594
rect 26226 50542 26238 50594
rect 26290 50542 26302 50594
rect 23998 50530 24050 50542
rect 25678 50482 25730 50494
rect 23538 50430 23550 50482
rect 23602 50430 23614 50482
rect 25678 50418 25730 50430
rect 27246 50370 27298 50382
rect 27246 50306 27298 50318
rect 672 50202 27888 50236
rect 672 50150 3806 50202
rect 3858 50150 3910 50202
rect 3962 50150 4014 50202
rect 4066 50150 23806 50202
rect 23858 50150 23910 50202
rect 23962 50150 24014 50202
rect 24066 50150 27888 50202
rect 672 50116 27888 50150
rect 25678 49922 25730 49934
rect 27122 49870 27134 49922
rect 27186 49870 27198 49922
rect 25678 49858 25730 49870
rect 26450 49758 26462 49810
rect 26514 49758 26526 49810
rect 24658 49646 24670 49698
rect 24722 49646 24734 49698
rect 672 49418 27888 49452
rect 672 49366 4466 49418
rect 4518 49366 4570 49418
rect 4622 49366 4674 49418
rect 4726 49366 24466 49418
rect 24518 49366 24570 49418
rect 24622 49366 24674 49418
rect 24726 49366 27888 49418
rect 672 49332 27888 49366
rect 24658 48974 24670 49026
rect 24722 48974 24734 49026
rect 26226 48974 26238 49026
rect 26290 48974 26302 49026
rect 25678 48802 25730 48814
rect 25678 48738 25730 48750
rect 27246 48802 27298 48814
rect 27246 48738 27298 48750
rect 672 48634 27888 48668
rect 672 48582 3806 48634
rect 3858 48582 3910 48634
rect 3962 48582 4014 48634
rect 4066 48582 23806 48634
rect 23858 48582 23910 48634
rect 23962 48582 24014 48634
rect 24066 48582 27888 48634
rect 672 48548 27888 48582
rect 26226 48078 26238 48130
rect 26290 48078 26302 48130
rect 27010 48078 27022 48130
rect 27074 48078 27086 48130
rect 672 47850 27888 47884
rect 672 47798 4466 47850
rect 4518 47798 4570 47850
rect 4622 47798 4674 47850
rect 4726 47798 24466 47850
rect 24518 47798 24570 47850
rect 24622 47798 24674 47850
rect 24726 47798 27888 47850
rect 672 47764 27888 47798
rect 24658 47406 24670 47458
rect 24722 47406 24734 47458
rect 26226 47406 26238 47458
rect 26290 47406 26302 47458
rect 25678 47346 25730 47358
rect 25678 47282 25730 47294
rect 27246 47234 27298 47246
rect 27246 47170 27298 47182
rect 672 47066 27888 47100
rect 672 47014 3806 47066
rect 3858 47014 3910 47066
rect 3962 47014 4014 47066
rect 4066 47014 23806 47066
rect 23858 47014 23910 47066
rect 23962 47014 24014 47066
rect 24066 47014 27888 47066
rect 672 46980 27888 47014
rect 25678 46786 25730 46798
rect 27122 46734 27134 46786
rect 27186 46734 27198 46786
rect 25678 46722 25730 46734
rect 24658 46510 24670 46562
rect 24722 46510 24734 46562
rect 26226 46510 26238 46562
rect 26290 46510 26302 46562
rect 672 46282 27888 46316
rect 672 46230 4466 46282
rect 4518 46230 4570 46282
rect 4622 46230 4674 46282
rect 4726 46230 24466 46282
rect 24518 46230 24570 46282
rect 24622 46230 24674 46282
rect 24726 46230 27888 46282
rect 672 46196 27888 46230
rect 24882 45838 24894 45890
rect 24946 45838 24958 45890
rect 26226 45838 26238 45890
rect 26290 45838 26302 45890
rect 25678 45666 25730 45678
rect 25678 45602 25730 45614
rect 27246 45666 27298 45678
rect 27246 45602 27298 45614
rect 672 45498 27888 45532
rect 672 45446 3806 45498
rect 3858 45446 3910 45498
rect 3962 45446 4014 45498
rect 4066 45446 23806 45498
rect 23858 45446 23910 45498
rect 23962 45446 24014 45498
rect 24066 45446 27888 45498
rect 672 45412 27888 45446
rect 26450 45054 26462 45106
rect 26514 45054 26526 45106
rect 27010 44942 27022 44994
rect 27074 44942 27086 44994
rect 672 44714 27888 44748
rect 672 44662 4466 44714
rect 4518 44662 4570 44714
rect 4622 44662 4674 44714
rect 4726 44662 24466 44714
rect 24518 44662 24570 44714
rect 24622 44662 24674 44714
rect 24726 44662 27888 44714
rect 672 44628 27888 44662
rect 24882 44270 24894 44322
rect 24946 44270 24958 44322
rect 26338 44270 26350 44322
rect 26402 44270 26414 44322
rect 25678 44210 25730 44222
rect 25678 44146 25730 44158
rect 27246 44098 27298 44110
rect 27246 44034 27298 44046
rect 672 43930 27888 43964
rect 672 43878 3806 43930
rect 3858 43878 3910 43930
rect 3962 43878 4014 43930
rect 4066 43878 23806 43930
rect 23858 43878 23910 43930
rect 23962 43878 24014 43930
rect 24066 43878 27888 43930
rect 672 43844 27888 43878
rect 25678 43650 25730 43662
rect 27122 43598 27134 43650
rect 27186 43598 27198 43650
rect 25678 43586 25730 43598
rect 24882 43486 24894 43538
rect 24946 43486 24958 43538
rect 26226 43374 26238 43426
rect 26290 43374 26302 43426
rect 672 43146 27888 43180
rect 672 43094 4466 43146
rect 4518 43094 4570 43146
rect 4622 43094 4674 43146
rect 4726 43094 24466 43146
rect 24518 43094 24570 43146
rect 24622 43094 24674 43146
rect 24726 43094 27888 43146
rect 672 43060 27888 43094
rect 24658 42702 24670 42754
rect 24722 42702 24734 42754
rect 26226 42702 26238 42754
rect 26290 42702 26302 42754
rect 25678 42530 25730 42542
rect 25678 42466 25730 42478
rect 27246 42530 27298 42542
rect 27246 42466 27298 42478
rect 672 42362 27888 42396
rect 672 42310 3806 42362
rect 3858 42310 3910 42362
rect 3962 42310 4014 42362
rect 4066 42310 23806 42362
rect 23858 42310 23910 42362
rect 23962 42310 24014 42362
rect 24066 42310 27888 42362
rect 672 42276 27888 42310
rect 14242 42030 14254 42082
rect 14306 42030 14318 42082
rect 14578 41806 14590 41858
rect 14642 41806 14654 41858
rect 26226 41806 26238 41858
rect 26290 41806 26302 41858
rect 27010 41806 27022 41858
rect 27074 41806 27086 41858
rect 15822 41746 15874 41758
rect 15822 41682 15874 41694
rect 672 41578 27888 41612
rect 672 41526 4466 41578
rect 4518 41526 4570 41578
rect 4622 41526 4674 41578
rect 4726 41526 24466 41578
rect 24518 41526 24570 41578
rect 24622 41526 24674 41578
rect 24726 41526 27888 41578
rect 672 41492 27888 41526
rect 14354 41358 14366 41410
rect 14418 41358 14430 41410
rect 10098 41246 10110 41298
rect 10162 41246 10174 41298
rect 11778 41134 11790 41186
rect 11842 41134 11854 41186
rect 13794 41134 13806 41186
rect 13858 41134 13870 41186
rect 24770 41134 24782 41186
rect 24834 41134 24846 41186
rect 26226 41134 26238 41186
rect 26290 41134 26302 41186
rect 25678 41074 25730 41086
rect 10546 41022 10558 41074
rect 10610 41022 10622 41074
rect 12114 41022 12126 41074
rect 12178 41022 12190 41074
rect 25678 41010 25730 41022
rect 8990 40962 9042 40974
rect 8990 40898 9042 40910
rect 15486 40962 15538 40974
rect 15486 40898 15538 40910
rect 27246 40962 27298 40974
rect 27246 40898 27298 40910
rect 672 40794 27888 40828
rect 672 40742 3806 40794
rect 3858 40742 3910 40794
rect 3962 40742 4014 40794
rect 4066 40742 23806 40794
rect 23858 40742 23910 40794
rect 23962 40742 24014 40794
rect 24066 40742 27888 40794
rect 672 40708 27888 40742
rect 25678 40514 25730 40526
rect 12898 40462 12910 40514
rect 12962 40462 12974 40514
rect 14466 40462 14478 40514
rect 14530 40462 14542 40514
rect 27122 40462 27134 40514
rect 27186 40462 27198 40514
rect 25678 40450 25730 40462
rect 6078 40402 6130 40414
rect 6514 40350 6526 40402
rect 6578 40350 6590 40402
rect 6850 40350 6862 40402
rect 6914 40350 6926 40402
rect 8306 40350 8318 40402
rect 8370 40350 8382 40402
rect 9202 40350 9214 40402
rect 9266 40350 9278 40402
rect 10434 40350 10446 40402
rect 10498 40350 10510 40402
rect 24658 40350 24670 40402
rect 24722 40350 24734 40402
rect 26226 40350 26238 40402
rect 26290 40350 26302 40402
rect 6078 40338 6130 40350
rect 7534 40290 7586 40302
rect 10882 40238 10894 40290
rect 10946 40238 10958 40290
rect 7534 40226 7586 40238
rect 12126 40178 12178 40190
rect 7074 40126 7086 40178
rect 7138 40126 7150 40178
rect 12126 40114 12178 40126
rect 13358 40178 13410 40190
rect 16046 40178 16098 40190
rect 14914 40126 14926 40178
rect 14978 40126 14990 40178
rect 13358 40114 13410 40126
rect 16046 40114 16098 40126
rect 672 40010 27888 40044
rect 672 39958 4466 40010
rect 4518 39958 4570 40010
rect 4622 39958 4674 40010
rect 4726 39958 24466 40010
rect 24518 39958 24570 40010
rect 24622 39958 24674 40010
rect 24726 39958 27888 40010
rect 672 39924 27888 39958
rect 6974 39842 7026 39854
rect 6974 39778 7026 39790
rect 3054 39730 3106 39742
rect 3054 39666 3106 39678
rect 7310 39730 7362 39742
rect 7310 39666 7362 39678
rect 8990 39618 9042 39630
rect 2594 39566 2606 39618
rect 2658 39566 2670 39618
rect 3826 39566 3838 39618
rect 3890 39566 3902 39618
rect 7746 39566 7758 39618
rect 7810 39566 7822 39618
rect 14018 39566 14030 39618
rect 14082 39566 14094 39618
rect 24882 39566 24894 39618
rect 24946 39566 24958 39618
rect 26226 39566 26238 39618
rect 26290 39566 26302 39618
rect 8990 39554 9042 39566
rect 6414 39506 6466 39518
rect 3490 39454 3502 39506
rect 3554 39454 3566 39506
rect 6414 39442 6466 39454
rect 9550 39506 9602 39518
rect 10546 39454 10558 39506
rect 10610 39454 10622 39506
rect 9550 39442 9602 39454
rect 25678 39394 25730 39406
rect 25678 39330 25730 39342
rect 27246 39394 27298 39406
rect 27246 39330 27298 39342
rect 672 39226 27888 39260
rect 672 39174 3806 39226
rect 3858 39174 3910 39226
rect 3962 39174 4014 39226
rect 4066 39174 23806 39226
rect 23858 39174 23910 39226
rect 23962 39174 24014 39226
rect 24066 39174 27888 39226
rect 672 39140 27888 39174
rect 6974 39058 7026 39070
rect 6974 38994 7026 39006
rect 7982 38946 8034 38958
rect 1586 38894 1598 38946
rect 1650 38894 1662 38946
rect 5394 38894 5406 38946
rect 5458 38894 5470 38946
rect 7982 38882 8034 38894
rect 12238 38946 12290 38958
rect 12238 38882 12290 38894
rect 16942 38946 16994 38958
rect 16942 38882 16994 38894
rect 2258 38782 2270 38834
rect 2322 38782 2334 38834
rect 8306 38782 8318 38834
rect 8370 38782 8382 38834
rect 8866 38794 8878 38846
rect 8930 38794 8942 38846
rect 9438 38834 9490 38846
rect 12798 38834 12850 38846
rect 14254 38834 14306 38846
rect 10098 38782 10110 38834
rect 10162 38782 10174 38834
rect 10994 38782 11006 38834
rect 11058 38782 11070 38834
rect 11778 38782 11790 38834
rect 11842 38782 11854 38834
rect 13122 38782 13134 38834
rect 13186 38782 13198 38834
rect 13570 38782 13582 38834
rect 13634 38782 13646 38834
rect 14802 38782 14814 38834
rect 14866 38782 14878 38834
rect 15810 38782 15822 38834
rect 15874 38782 15886 38834
rect 9438 38770 9490 38782
rect 12798 38770 12850 38782
rect 14254 38770 14306 38782
rect 1150 38722 1202 38734
rect 2706 38670 2718 38722
rect 2770 38670 2782 38722
rect 5842 38670 5854 38722
rect 5906 38670 5918 38722
rect 8978 38670 8990 38722
rect 9042 38670 9054 38722
rect 13794 38670 13806 38722
rect 13858 38670 13870 38722
rect 26226 38670 26238 38722
rect 26290 38670 26302 38722
rect 27010 38670 27022 38722
rect 27074 38670 27086 38722
rect 1150 38658 1202 38670
rect 3838 38610 3890 38622
rect 3838 38546 3890 38558
rect 16382 38610 16434 38622
rect 16382 38546 16434 38558
rect 672 38442 27888 38476
rect 672 38390 4466 38442
rect 4518 38390 4570 38442
rect 4622 38390 4674 38442
rect 4726 38390 24466 38442
rect 24518 38390 24570 38442
rect 24622 38390 24674 38442
rect 24726 38390 27888 38442
rect 672 38356 27888 38390
rect 5966 38274 6018 38286
rect 4834 38222 4846 38274
rect 4898 38222 4910 38274
rect 5966 38210 6018 38222
rect 8206 38274 8258 38286
rect 8206 38210 8258 38222
rect 15710 38162 15762 38174
rect 1810 38110 1822 38162
rect 1874 38110 1886 38162
rect 6962 38110 6974 38162
rect 7026 38110 7038 38162
rect 15710 38098 15762 38110
rect 15150 38050 15202 38062
rect 6626 37998 6638 38050
rect 6690 37998 6702 38050
rect 14690 37998 14702 38050
rect 14754 37998 14766 38050
rect 24658 37998 24670 38050
rect 24722 37998 24734 38050
rect 26226 37998 26238 38050
rect 26290 37998 26302 38050
rect 15150 37986 15202 37998
rect 25678 37938 25730 37950
rect 1362 37886 1374 37938
rect 1426 37886 1438 37938
rect 4386 37886 4398 37938
rect 4450 37886 4462 37938
rect 9650 37886 9662 37938
rect 9714 37886 9726 37938
rect 25678 37874 25730 37886
rect 2942 37826 2994 37838
rect 2942 37762 2994 37774
rect 27246 37826 27298 37838
rect 27246 37762 27298 37774
rect 672 37658 27888 37692
rect 672 37606 3806 37658
rect 3858 37606 3910 37658
rect 3962 37606 4014 37658
rect 4066 37606 23806 37658
rect 23858 37606 23910 37658
rect 23962 37606 24014 37658
rect 24066 37606 27888 37658
rect 672 37572 27888 37606
rect 8094 37490 8146 37502
rect 8094 37426 8146 37438
rect 2158 37378 2210 37390
rect 6514 37326 6526 37378
rect 6578 37326 6590 37378
rect 12002 37326 12014 37378
rect 12066 37326 12078 37378
rect 27122 37326 27134 37378
rect 27186 37326 27198 37378
rect 2158 37314 2210 37326
rect 16606 37266 16658 37278
rect 1698 37214 1710 37266
rect 1762 37214 1774 37266
rect 2706 37214 2718 37266
rect 2770 37214 2782 37266
rect 8642 37214 8654 37266
rect 8706 37214 8718 37266
rect 13122 37214 13134 37266
rect 13186 37214 13198 37266
rect 15474 37214 15486 37266
rect 15538 37214 15550 37266
rect 15922 37214 15934 37266
rect 15986 37214 15998 37266
rect 17154 37214 17166 37266
rect 17218 37214 17230 37266
rect 18162 37214 18174 37266
rect 18226 37214 18238 37266
rect 16606 37202 16658 37214
rect 15150 37154 15202 37166
rect 6962 37102 6974 37154
rect 7026 37102 7038 37154
rect 9314 37102 9326 37154
rect 9378 37102 9390 37154
rect 13458 37102 13470 37154
rect 13522 37102 13534 37154
rect 24658 37102 24670 37154
rect 24722 37102 24734 37154
rect 25442 37102 25454 37154
rect 25506 37102 25518 37154
rect 26226 37102 26238 37154
rect 26290 37102 26302 37154
rect 15150 37090 15202 37102
rect 4286 37042 4338 37054
rect 3154 36990 3166 37042
rect 3218 36990 3230 37042
rect 4286 36978 4338 36990
rect 14702 37042 14754 37054
rect 16146 36990 16158 37042
rect 16210 36990 16222 37042
rect 14702 36978 14754 36990
rect 672 36874 27888 36908
rect 672 36822 4466 36874
rect 4518 36822 4570 36874
rect 4622 36822 4674 36874
rect 4726 36822 24466 36874
rect 24518 36822 24570 36874
rect 24622 36822 24674 36874
rect 24726 36822 27888 36874
rect 672 36788 27888 36822
rect 10558 36706 10610 36718
rect 6402 36654 6414 36706
rect 6466 36654 6478 36706
rect 10210 36654 10222 36706
rect 10274 36654 10286 36706
rect 10558 36642 10610 36654
rect 16718 36706 16770 36718
rect 16718 36642 16770 36654
rect 17278 36594 17330 36606
rect 19854 36594 19906 36606
rect 4162 36542 4174 36594
rect 4226 36542 4238 36594
rect 18274 36542 18286 36594
rect 18338 36542 18350 36594
rect 24658 36542 24670 36594
rect 24722 36542 24734 36594
rect 17278 36530 17330 36542
rect 19854 36530 19906 36542
rect 2606 36482 2658 36494
rect 20414 36482 20466 36494
rect 4722 36430 4734 36482
rect 4786 36430 4798 36482
rect 7858 36430 7870 36482
rect 7922 36430 7934 36482
rect 10882 36430 10894 36482
rect 10946 36430 10958 36482
rect 17714 36430 17726 36482
rect 17778 36430 17790 36482
rect 26338 36430 26350 36482
rect 26402 36430 26414 36482
rect 2606 36418 2658 36430
rect 20414 36418 20466 36430
rect 2046 36370 2098 36382
rect 7422 36370 7474 36382
rect 6850 36318 6862 36370
rect 6914 36318 6926 36370
rect 13570 36318 13582 36370
rect 13634 36318 13646 36370
rect 2046 36306 2098 36318
rect 7422 36306 7474 36318
rect 3054 36258 3106 36270
rect 3054 36194 3106 36206
rect 5294 36258 5346 36270
rect 5294 36194 5346 36206
rect 19406 36258 19458 36270
rect 19406 36194 19458 36206
rect 25678 36258 25730 36270
rect 25678 36194 25730 36206
rect 27246 36258 27298 36270
rect 27246 36194 27298 36206
rect 672 36090 27888 36124
rect 672 36038 3806 36090
rect 3858 36038 3910 36090
rect 3962 36038 4014 36090
rect 4066 36038 23806 36090
rect 23858 36038 23910 36090
rect 23962 36038 24014 36090
rect 24066 36038 27888 36090
rect 672 36004 27888 36038
rect 4398 35810 4450 35822
rect 2706 35758 2718 35810
rect 2770 35758 2782 35810
rect 4398 35746 4450 35758
rect 5966 35810 6018 35822
rect 6514 35758 6526 35810
rect 6578 35758 6590 35810
rect 12002 35758 12014 35810
rect 12066 35758 12078 35810
rect 5966 35746 6018 35758
rect 5506 35646 5518 35698
rect 5570 35646 5582 35698
rect 8642 35646 8654 35698
rect 8706 35646 8718 35698
rect 13570 35646 13582 35698
rect 13634 35646 13646 35698
rect 2370 35534 2382 35586
rect 2434 35534 2446 35586
rect 9314 35534 9326 35586
rect 9378 35534 9390 35586
rect 14802 35534 14814 35586
rect 14866 35534 14878 35586
rect 26226 35534 26238 35586
rect 26290 35534 26302 35586
rect 27010 35534 27022 35586
rect 27074 35534 27086 35586
rect 1150 35474 1202 35486
rect 3838 35474 3890 35486
rect 8094 35474 8146 35486
rect 2258 35422 2270 35474
rect 2322 35422 2334 35474
rect 6962 35422 6974 35474
rect 7026 35422 7038 35474
rect 1150 35410 1202 35422
rect 3838 35410 3890 35422
rect 8094 35410 8146 35422
rect 672 35306 27888 35340
rect 672 35254 4466 35306
rect 4518 35254 4570 35306
rect 4622 35254 4674 35306
rect 4726 35254 24466 35306
rect 24518 35254 24570 35306
rect 24622 35254 24674 35306
rect 24726 35254 27888 35306
rect 672 35220 27888 35254
rect 3826 35086 3838 35138
rect 3890 35086 3902 35138
rect 4286 35026 4338 35038
rect 17950 35026 18002 35038
rect 7074 34974 7086 35026
rect 7138 34974 7150 35026
rect 14018 34974 14030 35026
rect 14082 34974 14094 35026
rect 4286 34962 4338 34974
rect 17950 34962 18002 34974
rect 18286 35026 18338 35038
rect 19282 34974 19294 35026
rect 19346 34974 19358 35026
rect 18286 34962 18338 34974
rect 2034 34862 2046 34914
rect 2098 34862 2110 34914
rect 3154 34862 3166 34914
rect 3218 34862 3230 34914
rect 3714 34862 3726 34914
rect 3778 34862 3790 34914
rect 4946 34862 4958 34914
rect 5010 34862 5022 34914
rect 5842 34862 5854 34914
rect 5906 34862 5918 34914
rect 6514 34862 6526 34914
rect 6578 34862 6590 34914
rect 9650 34862 9662 34914
rect 9714 34862 9726 34914
rect 10882 34862 10894 34914
rect 10946 34862 10958 34914
rect 17490 34862 17502 34914
rect 17554 34862 17566 34914
rect 18722 34862 18734 34914
rect 18786 34862 18798 34914
rect 19058 34862 19070 34914
rect 19122 34862 19134 34914
rect 19842 34862 19854 34914
rect 19906 34862 19918 34914
rect 20290 34862 20302 34914
rect 20354 34862 20366 34914
rect 21298 34862 21310 34914
rect 21362 34862 21374 34914
rect 24658 34862 24670 34914
rect 24722 34862 24734 34914
rect 26226 34862 26238 34914
rect 26290 34862 26302 34914
rect 2494 34802 2546 34814
rect 2494 34738 2546 34750
rect 2830 34802 2882 34814
rect 25678 34802 25730 34814
rect 9986 34750 9998 34802
rect 10050 34750 10062 34802
rect 2830 34738 2882 34750
rect 25678 34738 25730 34750
rect 8206 34690 8258 34702
rect 8206 34626 8258 34638
rect 27246 34690 27298 34702
rect 27246 34626 27298 34638
rect 672 34522 27888 34556
rect 672 34470 3806 34522
rect 3858 34470 3910 34522
rect 3962 34470 4014 34522
rect 4066 34470 23806 34522
rect 23858 34470 23910 34522
rect 23962 34470 24014 34522
rect 24066 34470 27888 34522
rect 672 34436 27888 34470
rect 18958 34354 19010 34366
rect 18958 34290 19010 34302
rect 25678 34242 25730 34254
rect 27122 34190 27134 34242
rect 27186 34190 27198 34242
rect 25678 34178 25730 34190
rect 2830 34130 2882 34142
rect 10222 34130 10274 34142
rect 19518 34130 19570 34142
rect 1474 34078 1486 34130
rect 1538 34078 1550 34130
rect 1922 34078 1934 34130
rect 1986 34078 1998 34130
rect 3154 34078 3166 34130
rect 3218 34078 3230 34130
rect 4162 34078 4174 34130
rect 4226 34078 4238 34130
rect 5058 34078 5070 34130
rect 5122 34078 5134 34130
rect 8194 34078 8206 34130
rect 8258 34078 8270 34130
rect 9090 34078 9102 34130
rect 9154 34078 9166 34130
rect 9538 34078 9550 34130
rect 9602 34078 9614 34130
rect 10882 34078 10894 34130
rect 10946 34078 10958 34130
rect 11778 34078 11790 34130
rect 11842 34078 11854 34130
rect 12674 34078 12686 34130
rect 12738 34078 12750 34130
rect 17266 34078 17278 34130
rect 17330 34078 17342 34130
rect 2830 34066 2882 34078
rect 10222 34066 10274 34078
rect 19518 34066 19570 34078
rect 1150 34018 1202 34030
rect 8766 34018 8818 34030
rect 20078 34018 20130 34030
rect 2146 33966 2158 34018
rect 2210 33966 2222 34018
rect 9762 33966 9774 34018
rect 9826 33966 9838 34018
rect 13570 33966 13582 34018
rect 13634 33966 13646 34018
rect 24658 33966 24670 34018
rect 24722 33966 24734 34018
rect 26226 33966 26238 34018
rect 26290 33966 26302 34018
rect 1150 33954 1202 33966
rect 8766 33954 8818 33966
rect 20078 33954 20130 33966
rect 5518 33906 5570 33918
rect 5518 33842 5570 33854
rect 6638 33906 6690 33918
rect 7746 33854 7758 33906
rect 7810 33854 7822 33906
rect 16258 33854 16270 33906
rect 16322 33854 16334 33906
rect 17826 33854 17838 33906
rect 17890 33854 17902 33906
rect 6638 33842 6690 33854
rect 672 33738 27888 33772
rect 672 33686 4466 33738
rect 4518 33686 4570 33738
rect 4622 33686 4674 33738
rect 4726 33686 24466 33738
rect 24518 33686 24570 33738
rect 24622 33686 24674 33738
rect 24726 33686 27888 33738
rect 672 33652 27888 33686
rect 3266 33406 3278 33458
rect 3330 33406 3342 33458
rect 7634 33406 7646 33458
rect 7698 33406 7710 33458
rect 10882 33406 10894 33458
rect 10946 33406 10958 33458
rect 18722 33406 18734 33458
rect 18786 33406 18798 33458
rect 3726 33346 3778 33358
rect 8878 33346 8930 33358
rect 2706 33294 2718 33346
rect 2770 33294 2782 33346
rect 3154 33294 3166 33346
rect 3218 33294 3230 33346
rect 4498 33294 4510 33346
rect 4562 33294 4574 33346
rect 5394 33294 5406 33346
rect 5458 33294 5470 33346
rect 12562 33294 12574 33346
rect 12626 33294 12638 33346
rect 18274 33294 18286 33346
rect 18338 33294 18350 33346
rect 24658 33294 24670 33346
rect 24722 33294 24734 33346
rect 26226 33294 26238 33346
rect 26290 33294 26302 33346
rect 3726 33282 3778 33294
rect 8878 33282 8930 33294
rect 2270 33234 2322 33246
rect 8082 33182 8094 33234
rect 8146 33182 8158 33234
rect 9314 33182 9326 33234
rect 9378 33182 9390 33234
rect 10434 33182 10446 33234
rect 10498 33182 10510 33234
rect 13234 33182 13246 33234
rect 13298 33182 13310 33234
rect 15586 33182 15598 33234
rect 15650 33182 15662 33234
rect 2270 33170 2322 33182
rect 6526 33122 6578 33134
rect 6526 33058 6578 33070
rect 12014 33122 12066 33134
rect 12014 33058 12066 33070
rect 19966 33122 20018 33134
rect 19966 33058 20018 33070
rect 25678 33122 25730 33134
rect 25678 33058 25730 33070
rect 27246 33122 27298 33134
rect 27246 33058 27298 33070
rect 672 32954 27888 32988
rect 672 32902 3806 32954
rect 3858 32902 3910 32954
rect 3962 32902 4014 32954
rect 4066 32902 23806 32954
rect 23858 32902 23910 32954
rect 23962 32902 24014 32954
rect 24066 32902 27888 32954
rect 672 32868 27888 32902
rect 2830 32786 2882 32798
rect 2830 32722 2882 32734
rect 19742 32674 19794 32686
rect 22094 32674 22146 32686
rect 5842 32622 5854 32674
rect 5906 32622 5918 32674
rect 15586 32622 15598 32674
rect 15650 32622 15662 32674
rect 20738 32622 20750 32674
rect 20802 32622 20814 32674
rect 19742 32610 19794 32622
rect 22094 32610 22146 32622
rect 19182 32562 19234 32574
rect 1138 32510 1150 32562
rect 1202 32510 1214 32562
rect 3378 32510 3390 32562
rect 3442 32510 3454 32562
rect 5170 32510 5182 32562
rect 5234 32510 5246 32562
rect 7186 32510 7198 32562
rect 7250 32510 7262 32562
rect 9874 32510 9886 32562
rect 9938 32510 9950 32562
rect 14802 32510 14814 32562
rect 14866 32510 14878 32562
rect 26338 32510 26350 32562
rect 26402 32510 26414 32562
rect 19182 32498 19234 32510
rect 3838 32450 3890 32462
rect 1586 32398 1598 32450
rect 1650 32398 1662 32450
rect 7634 32398 7646 32450
rect 7698 32398 7710 32450
rect 10322 32398 10334 32450
rect 10386 32398 10398 32450
rect 27010 32398 27022 32450
rect 27074 32398 27086 32450
rect 3838 32386 3890 32398
rect 8878 32338 8930 32350
rect 8878 32274 8930 32286
rect 11454 32338 11506 32350
rect 11454 32274 11506 32286
rect 21198 32338 21250 32350
rect 21198 32274 21250 32286
rect 21534 32338 21586 32350
rect 21534 32274 21586 32286
rect 672 32170 27888 32204
rect 672 32118 4466 32170
rect 4518 32118 4570 32170
rect 4622 32118 4674 32170
rect 4726 32118 24466 32170
rect 24518 32118 24570 32170
rect 24622 32118 24674 32170
rect 24726 32118 27888 32170
rect 672 32084 27888 32118
rect 12450 31950 12462 32002
rect 12514 31950 12526 32002
rect 21186 31950 21198 32002
rect 21250 31950 21262 32002
rect 3278 31890 3330 31902
rect 9662 31890 9714 31902
rect 2146 31838 2158 31890
rect 2210 31838 2222 31890
rect 6066 31838 6078 31890
rect 6130 31838 6142 31890
rect 3278 31826 3330 31838
rect 9662 31826 9714 31838
rect 11118 31890 11170 31902
rect 11118 31826 11170 31838
rect 12910 31890 12962 31902
rect 18610 31838 18622 31890
rect 18674 31838 18686 31890
rect 12910 31826 12962 31838
rect 10222 31778 10274 31790
rect 16718 31778 16770 31790
rect 1698 31726 1710 31778
rect 1762 31726 1774 31778
rect 5394 31726 5406 31778
rect 5458 31726 5470 31778
rect 5842 31726 5854 31778
rect 5906 31726 5918 31778
rect 6626 31726 6638 31778
rect 6690 31726 6702 31778
rect 7074 31726 7086 31778
rect 7138 31726 7150 31778
rect 8194 31726 8206 31778
rect 8258 31726 8270 31778
rect 11778 31726 11790 31778
rect 11842 31726 11854 31778
rect 10222 31714 10274 31726
rect 12338 31714 12350 31766
rect 12402 31714 12414 31766
rect 13458 31726 13470 31778
rect 13522 31726 13534 31778
rect 14466 31726 14478 31778
rect 14530 31726 14542 31778
rect 18050 31726 18062 31778
rect 18114 31726 18126 31778
rect 20626 31726 20638 31778
rect 20690 31726 20702 31778
rect 20962 31726 20974 31778
rect 21026 31726 21038 31778
rect 21746 31726 21758 31778
rect 21810 31726 21822 31778
rect 22418 31726 22430 31778
rect 22482 31726 22494 31778
rect 23202 31726 23214 31778
rect 23266 31726 23278 31778
rect 24882 31726 24894 31778
rect 24946 31726 24958 31778
rect 26450 31726 26462 31778
rect 26514 31726 26526 31778
rect 16718 31714 16770 31726
rect 5070 31666 5122 31678
rect 11454 31666 11506 31678
rect 20190 31666 20242 31678
rect 10658 31614 10670 31666
rect 10722 31614 10734 31666
rect 17154 31614 17166 31666
rect 17218 31614 17230 31666
rect 5070 31602 5122 31614
rect 11454 31602 11506 31614
rect 20190 31602 20242 31614
rect 25678 31666 25730 31678
rect 25678 31602 25730 31614
rect 19742 31554 19794 31566
rect 19742 31490 19794 31502
rect 27246 31554 27298 31566
rect 27246 31490 27298 31502
rect 672 31386 27888 31420
rect 672 31334 3806 31386
rect 3858 31334 3910 31386
rect 3962 31334 4014 31386
rect 4066 31334 23806 31386
rect 23858 31334 23910 31386
rect 23962 31334 24014 31386
rect 24066 31334 27888 31386
rect 672 31300 27888 31334
rect 4286 31218 4338 31230
rect 4286 31154 4338 31166
rect 5518 31106 5570 31118
rect 5518 31042 5570 31054
rect 6414 31106 6466 31118
rect 6414 31042 6466 31054
rect 10558 30994 10610 31006
rect 22094 30994 22146 31006
rect 2706 30942 2718 30994
rect 2770 30942 2782 30994
rect 5954 30942 5966 30994
rect 6018 30942 6030 30994
rect 6962 30942 6974 30994
rect 7026 30942 7038 30994
rect 9090 30942 9102 30994
rect 9154 30942 9166 30994
rect 9986 30942 9998 30994
rect 10050 30942 10062 30994
rect 11330 30942 11342 30994
rect 11394 30942 11406 30994
rect 11778 30942 11790 30994
rect 11842 30942 11854 30994
rect 13458 30942 13470 30994
rect 13522 30942 13534 30994
rect 15810 30942 15822 30994
rect 15874 30942 15886 30994
rect 16370 30942 16382 30994
rect 16434 30942 16446 30994
rect 17490 30942 17502 30994
rect 17554 30942 17566 30994
rect 18498 30942 18510 30994
rect 18562 30942 18574 30994
rect 20962 30942 20974 30994
rect 21026 30942 21038 30994
rect 21410 30942 21422 30994
rect 21474 30942 21486 30994
rect 22642 30942 22654 30994
rect 22706 30942 22718 30994
rect 22866 30942 22878 30994
rect 22930 30942 22942 30994
rect 23650 30942 23662 30994
rect 23714 30942 23726 30994
rect 24882 30942 24894 30994
rect 24946 30942 24958 30994
rect 26338 30942 26350 30994
rect 26402 30942 26414 30994
rect 10558 30930 10610 30942
rect 22094 30930 22146 30942
rect 12238 30882 12290 30894
rect 15038 30882 15090 30894
rect 7298 30830 7310 30882
rect 7362 30830 7374 30882
rect 11218 30830 11230 30882
rect 11282 30830 11294 30882
rect 13794 30830 13806 30882
rect 13858 30830 13870 30882
rect 12238 30818 12290 30830
rect 15038 30818 15090 30830
rect 15486 30882 15538 30894
rect 16942 30882 16994 30894
rect 16482 30830 16494 30882
rect 16546 30830 16558 30882
rect 15486 30818 15538 30830
rect 16942 30818 16994 30830
rect 20638 30882 20690 30894
rect 21634 30830 21646 30882
rect 21698 30830 21710 30882
rect 25442 30830 25454 30882
rect 25506 30830 25518 30882
rect 27010 30830 27022 30882
rect 27074 30830 27086 30882
rect 20638 30818 20690 30830
rect 4958 30770 5010 30782
rect 3154 30718 3166 30770
rect 3218 30718 3230 30770
rect 4958 30706 5010 30718
rect 8542 30770 8594 30782
rect 8542 30706 8594 30718
rect 672 30602 27888 30636
rect 672 30550 4466 30602
rect 4518 30550 4570 30602
rect 4622 30550 4674 30602
rect 4726 30550 24466 30602
rect 24518 30550 24570 30602
rect 24622 30550 24674 30602
rect 24726 30550 27888 30602
rect 672 30516 27888 30550
rect 20862 30434 20914 30446
rect 4498 30382 4510 30434
rect 4562 30382 4574 30434
rect 20862 30370 20914 30382
rect 10882 30270 10894 30322
rect 10946 30270 10958 30322
rect 13570 30270 13582 30322
rect 13634 30270 13646 30322
rect 17378 30270 17390 30322
rect 17442 30270 17454 30322
rect 19618 30270 19630 30322
rect 19682 30270 19694 30322
rect 21858 30270 21870 30322
rect 21922 30270 21934 30322
rect 4958 30210 5010 30222
rect 8878 30210 8930 30222
rect 2258 30158 2270 30210
rect 2322 30158 2334 30210
rect 2706 30158 2718 30210
rect 2770 30158 2782 30210
rect 3826 30158 3838 30210
rect 3890 30158 3902 30210
rect 4274 30158 4286 30210
rect 4338 30158 4350 30210
rect 5618 30158 5630 30210
rect 5682 30158 5694 30210
rect 6514 30158 6526 30210
rect 6578 30158 6590 30210
rect 7074 30158 7086 30210
rect 7138 30158 7150 30210
rect 4958 30146 5010 30158
rect 8878 30146 8930 30158
rect 9438 30210 9490 30222
rect 12574 30210 12626 30222
rect 14254 30210 14306 30222
rect 23102 30210 23154 30222
rect 10434 30158 10446 30210
rect 10498 30158 10510 30210
rect 12898 30158 12910 30210
rect 12962 30158 12974 30210
rect 13346 30158 13358 30210
rect 13410 30158 13422 30210
rect 14578 30158 14590 30210
rect 14642 30158 14654 30210
rect 15698 30158 15710 30210
rect 15762 30158 15774 30210
rect 26226 30158 26238 30210
rect 26290 30158 26302 30210
rect 9438 30146 9490 30158
rect 12574 30146 12626 30158
rect 14254 30146 14306 30158
rect 23102 30146 23154 30158
rect 3502 30098 3554 30110
rect 1586 30046 1598 30098
rect 1650 30046 1662 30098
rect 3042 30046 3054 30098
rect 3106 30046 3118 30098
rect 17042 30046 17054 30098
rect 17106 30046 17118 30098
rect 19282 30046 19294 30098
rect 19346 30046 19358 30098
rect 21522 30046 21534 30098
rect 21586 30046 21598 30098
rect 27122 30046 27134 30098
rect 27186 30046 27198 30098
rect 3502 30034 3554 30046
rect 7646 29986 7698 29998
rect 7646 29922 7698 29934
rect 12126 29986 12178 29998
rect 12126 29922 12178 29934
rect 18622 29986 18674 29998
rect 18622 29922 18674 29934
rect 672 29818 27888 29852
rect 672 29766 3806 29818
rect 3858 29766 3910 29818
rect 3962 29766 4014 29818
rect 4066 29766 23806 29818
rect 23858 29766 23910 29818
rect 23962 29766 24014 29818
rect 24066 29766 27888 29818
rect 672 29732 27888 29766
rect 4286 29650 4338 29662
rect 4286 29586 4338 29598
rect 7198 29650 7250 29662
rect 7198 29586 7250 29598
rect 10110 29650 10162 29662
rect 10110 29586 10162 29598
rect 14030 29538 14082 29550
rect 1138 29486 1150 29538
rect 1202 29486 1214 29538
rect 2706 29486 2718 29538
rect 2770 29486 2782 29538
rect 8530 29486 8542 29538
rect 8594 29486 8606 29538
rect 11778 29486 11790 29538
rect 11842 29486 11854 29538
rect 14030 29474 14082 29486
rect 27246 29538 27298 29550
rect 27246 29474 27298 29486
rect 16046 29426 16098 29438
rect 1474 29374 1486 29426
rect 1538 29374 1550 29426
rect 5618 29374 5630 29426
rect 5682 29374 5694 29426
rect 13570 29374 13582 29426
rect 13634 29374 13646 29426
rect 14690 29374 14702 29426
rect 14754 29374 14766 29426
rect 15138 29374 15150 29426
rect 15202 29374 15214 29426
rect 16482 29374 16494 29426
rect 16546 29374 16558 29426
rect 17490 29374 17502 29426
rect 17554 29374 17566 29426
rect 18162 29374 18174 29426
rect 18226 29374 18238 29426
rect 26226 29374 26238 29426
rect 26290 29374 26302 29426
rect 16046 29362 16098 29374
rect 14366 29314 14418 29326
rect 6066 29262 6078 29314
rect 6130 29262 6142 29314
rect 18610 29262 18622 29314
rect 18674 29262 18686 29314
rect 14366 29250 14418 29262
rect 12238 29202 12290 29214
rect 19742 29202 19794 29214
rect 3154 29150 3166 29202
rect 3218 29150 3230 29202
rect 8978 29150 8990 29202
rect 9042 29150 9054 29202
rect 15362 29150 15374 29202
rect 15426 29150 15438 29202
rect 12238 29138 12290 29150
rect 19742 29138 19794 29150
rect 672 29034 27888 29068
rect 672 28982 4466 29034
rect 4518 28982 4570 29034
rect 4622 28982 4674 29034
rect 4726 28982 24466 29034
rect 24518 28982 24570 29034
rect 24622 28982 24674 29034
rect 24726 28982 27888 29034
rect 672 28948 27888 28982
rect 3614 28866 3666 28878
rect 15486 28866 15538 28878
rect 9986 28814 9998 28866
rect 10050 28814 10062 28866
rect 12562 28814 12574 28866
rect 12626 28814 12638 28866
rect 3614 28802 3666 28814
rect 15486 28802 15538 28814
rect 11566 28754 11618 28766
rect 2370 28702 2382 28754
rect 2434 28702 2446 28754
rect 4498 28702 4510 28754
rect 4562 28702 4574 28754
rect 17826 28702 17838 28754
rect 17890 28702 17902 28754
rect 20402 28702 20414 28754
rect 20466 28702 20478 28754
rect 11566 28690 11618 28702
rect 11118 28642 11170 28654
rect 13022 28642 13074 28654
rect 16046 28642 16098 28654
rect 21086 28642 21138 28654
rect 5058 28590 5070 28642
rect 5122 28590 5134 28642
rect 7298 28590 7310 28642
rect 7362 28590 7374 28642
rect 11890 28590 11902 28642
rect 11954 28590 11966 28642
rect 12338 28590 12350 28642
rect 12402 28590 12414 28642
rect 13570 28590 13582 28642
rect 13634 28590 13646 28642
rect 14690 28590 14702 28642
rect 14754 28590 14766 28642
rect 19842 28590 19854 28642
rect 19906 28590 19918 28642
rect 20178 28590 20190 28642
rect 20242 28590 20254 28642
rect 21410 28590 21422 28642
rect 21474 28590 21486 28642
rect 22418 28590 22430 28642
rect 22482 28590 22494 28642
rect 26226 28590 26238 28642
rect 26290 28590 26302 28642
rect 11118 28578 11170 28590
rect 13022 28578 13074 28590
rect 16046 28578 16098 28590
rect 21086 28578 21138 28590
rect 19406 28530 19458 28542
rect 2034 28478 2046 28530
rect 2098 28478 2110 28530
rect 9538 28478 9550 28530
rect 9602 28478 9614 28530
rect 17378 28478 17390 28530
rect 17442 28478 17454 28530
rect 19406 28466 19458 28478
rect 27246 28530 27298 28542
rect 27246 28466 27298 28478
rect 4286 28418 4338 28430
rect 4286 28354 4338 28366
rect 8094 28418 8146 28430
rect 8094 28354 8146 28366
rect 18958 28418 19010 28430
rect 18958 28354 19010 28366
rect 672 28250 27888 28284
rect 672 28198 3806 28250
rect 3858 28198 3910 28250
rect 3962 28198 4014 28250
rect 4066 28198 23806 28250
rect 23858 28198 23910 28250
rect 23962 28198 24014 28250
rect 24066 28198 27888 28250
rect 672 28164 27888 28198
rect 7422 28082 7474 28094
rect 7422 28018 7474 28030
rect 9774 28082 9826 28094
rect 9774 28018 9826 28030
rect 12126 28082 12178 28094
rect 12126 28018 12178 28030
rect 27246 28082 27298 28094
rect 27246 28018 27298 28030
rect 13582 27970 13634 27982
rect 21198 27970 21250 27982
rect 8194 27918 8206 27970
rect 8258 27918 8270 27970
rect 18162 27918 18174 27970
rect 18226 27918 18238 27970
rect 13582 27906 13634 27918
rect 21198 27906 21250 27918
rect 25678 27970 25730 27982
rect 25678 27906 25730 27918
rect 15262 27858 15314 27870
rect 20638 27858 20690 27870
rect 2258 27806 2270 27858
rect 2322 27806 2334 27858
rect 6626 27806 6638 27858
rect 6690 27806 6702 27858
rect 10434 27806 10446 27858
rect 10498 27806 10510 27858
rect 13906 27806 13918 27858
rect 13970 27806 13982 27858
rect 14354 27806 14366 27858
rect 14418 27806 14430 27858
rect 15810 27806 15822 27858
rect 15874 27806 15886 27858
rect 16594 27806 16606 27858
rect 16658 27806 16670 27858
rect 15262 27794 15314 27806
rect 20638 27794 20690 27806
rect 5518 27746 5570 27758
rect 2818 27694 2830 27746
rect 2882 27694 2894 27746
rect 6402 27694 6414 27746
rect 6466 27694 6478 27746
rect 8642 27694 8654 27746
rect 8706 27694 8718 27746
rect 10882 27694 10894 27746
rect 10946 27694 10958 27746
rect 18498 27694 18510 27746
rect 18562 27694 18574 27746
rect 24658 27694 24670 27746
rect 24722 27694 24734 27746
rect 26226 27694 26238 27746
rect 26290 27694 26302 27746
rect 5518 27682 5570 27694
rect 3950 27634 4002 27646
rect 3950 27570 4002 27582
rect 4958 27634 5010 27646
rect 19742 27634 19794 27646
rect 14578 27582 14590 27634
rect 14642 27582 14654 27634
rect 4958 27570 5010 27582
rect 19742 27570 19794 27582
rect 672 27466 27888 27500
rect 672 27414 4466 27466
rect 4518 27414 4570 27466
rect 4622 27414 4674 27466
rect 4726 27414 24466 27466
rect 24518 27414 24570 27466
rect 24622 27414 24674 27466
rect 24726 27414 27888 27466
rect 672 27380 27888 27414
rect 13134 27298 13186 27310
rect 15374 27298 15426 27310
rect 1698 27246 1710 27298
rect 1762 27246 1774 27298
rect 4274 27246 4286 27298
rect 4338 27246 4350 27298
rect 10098 27246 10110 27298
rect 10162 27246 10174 27298
rect 12002 27246 12014 27298
rect 12066 27246 12078 27298
rect 14242 27246 14254 27298
rect 14306 27246 14318 27298
rect 13134 27234 13186 27246
rect 15374 27234 15426 27246
rect 8318 27186 8370 27198
rect 8318 27122 8370 27134
rect 17390 27186 17442 27198
rect 18386 27134 18398 27186
rect 18450 27134 18462 27186
rect 27010 27134 27022 27186
rect 27074 27134 27086 27186
rect 17390 27122 17442 27134
rect 4734 27074 4786 27086
rect 1250 27022 1262 27074
rect 1314 27022 1326 27074
rect 3602 27022 3614 27074
rect 3666 27022 3678 27074
rect 4050 27022 4062 27074
rect 4114 27022 4126 27074
rect 5282 27022 5294 27074
rect 5346 27022 5358 27074
rect 6402 27022 6414 27074
rect 6466 27022 6478 27074
rect 7858 27022 7870 27074
rect 7922 27022 7934 27074
rect 10546 27022 10558 27074
rect 10610 27022 10622 27074
rect 11442 27022 11454 27074
rect 11506 27022 11518 27074
rect 13794 27022 13806 27074
rect 13858 27022 13870 27074
rect 17714 27022 17726 27074
rect 17778 27022 17790 27074
rect 18162 27022 18174 27074
rect 18226 27022 18238 27074
rect 18946 27022 18958 27074
rect 19010 27022 19022 27074
rect 19394 27022 19406 27074
rect 19458 27022 19470 27074
rect 20402 27022 20414 27074
rect 20466 27022 20478 27074
rect 24658 27022 24670 27074
rect 24722 27022 24734 27074
rect 26226 27022 26238 27074
rect 26290 27022 26302 27074
rect 4734 27010 4786 27022
rect 3278 26962 3330 26974
rect 3278 26898 3330 26910
rect 25678 26962 25730 26974
rect 25678 26898 25730 26910
rect 2830 26850 2882 26862
rect 2830 26786 2882 26798
rect 8990 26850 9042 26862
rect 8990 26786 9042 26798
rect 672 26682 27888 26716
rect 672 26630 3806 26682
rect 3858 26630 3910 26682
rect 3962 26630 4014 26682
rect 4066 26630 23806 26682
rect 23858 26630 23910 26682
rect 23962 26630 24014 26682
rect 24066 26630 27888 26682
rect 672 26596 27888 26630
rect 3614 26514 3666 26526
rect 3614 26450 3666 26462
rect 19966 26514 20018 26526
rect 19966 26450 20018 26462
rect 27246 26514 27298 26526
rect 27246 26450 27298 26462
rect 17714 26350 17726 26402
rect 17778 26350 17790 26402
rect 10670 26290 10722 26302
rect 15262 26290 15314 26302
rect 2034 26238 2046 26290
rect 2098 26238 2110 26290
rect 6402 26238 6414 26290
rect 6466 26238 6478 26290
rect 9314 26238 9326 26290
rect 9378 26238 9390 26290
rect 9762 26238 9774 26290
rect 9826 26238 9838 26290
rect 11218 26238 11230 26290
rect 11282 26238 11294 26290
rect 12114 26238 12126 26290
rect 12178 26238 12190 26290
rect 13234 26238 13246 26290
rect 13298 26238 13310 26290
rect 18386 26238 18398 26290
rect 18450 26238 18462 26290
rect 20738 26238 20750 26290
rect 20802 26238 20814 26290
rect 10670 26226 10722 26238
rect 15262 26226 15314 26238
rect 5518 26178 5570 26190
rect 8990 26178 9042 26190
rect 15822 26178 15874 26190
rect 2370 26126 2382 26178
rect 2434 26126 2446 26178
rect 6738 26126 6750 26178
rect 6802 26126 6814 26178
rect 13682 26126 13694 26178
rect 13746 26126 13758 26178
rect 18722 26126 18734 26178
rect 18786 26126 18798 26178
rect 26226 26126 26238 26178
rect 26290 26126 26302 26178
rect 5518 26114 5570 26126
rect 8990 26114 9042 26126
rect 15822 26114 15874 26126
rect 4958 26066 5010 26078
rect 4958 26002 5010 26014
rect 7982 26066 8034 26078
rect 14814 26066 14866 26078
rect 9986 26014 9998 26066
rect 10050 26014 10062 26066
rect 7982 26002 8034 26014
rect 14814 26002 14866 26014
rect 17278 26066 17330 26078
rect 22430 26066 22482 26078
rect 21298 26014 21310 26066
rect 21362 26014 21374 26066
rect 17278 26002 17330 26014
rect 22430 26002 22482 26014
rect 672 25898 27888 25932
rect 672 25846 4466 25898
rect 4518 25846 4570 25898
rect 4622 25846 4674 25898
rect 4726 25846 24466 25898
rect 24518 25846 24570 25898
rect 24622 25846 24674 25898
rect 24726 25846 27888 25898
rect 672 25812 27888 25846
rect 10670 25730 10722 25742
rect 3602 25678 3614 25730
rect 3666 25678 3678 25730
rect 7074 25678 7086 25730
rect 7138 25678 7150 25730
rect 9538 25678 9550 25730
rect 9602 25678 9614 25730
rect 10670 25666 10722 25678
rect 18622 25730 18674 25742
rect 18622 25666 18674 25678
rect 21310 25730 21362 25742
rect 21310 25666 21362 25678
rect 17278 25618 17330 25630
rect 11778 25566 11790 25618
rect 11842 25566 11854 25618
rect 14914 25566 14926 25618
rect 14978 25566 14990 25618
rect 17278 25554 17330 25566
rect 19182 25618 19234 25630
rect 22318 25618 22370 25630
rect 20178 25566 20190 25618
rect 20242 25566 20254 25618
rect 19182 25554 19234 25566
rect 22318 25554 22370 25566
rect 21758 25506 21810 25518
rect 2034 25454 2046 25506
rect 2098 25454 2110 25506
rect 2930 25454 2942 25506
rect 2994 25454 3006 25506
rect 3378 25454 3390 25506
rect 3442 25454 3454 25506
rect 4162 25454 4174 25506
rect 4226 25454 4238 25506
rect 4722 25454 4734 25506
rect 4786 25454 4798 25506
rect 5618 25454 5630 25506
rect 5682 25454 5694 25506
rect 6514 25454 6526 25506
rect 6578 25454 6590 25506
rect 9090 25454 9102 25506
rect 9154 25454 9166 25506
rect 11330 25454 11342 25506
rect 11394 25454 11406 25506
rect 14466 25454 14478 25506
rect 14530 25454 14542 25506
rect 16818 25454 16830 25506
rect 16882 25454 16894 25506
rect 24658 25454 24670 25506
rect 24722 25454 24734 25506
rect 26226 25454 26238 25506
rect 26290 25454 26302 25506
rect 21758 25442 21810 25454
rect 1262 25394 1314 25406
rect 1262 25330 1314 25342
rect 2606 25394 2658 25406
rect 27246 25394 27298 25406
rect 19730 25342 19742 25394
rect 19794 25342 19806 25394
rect 2606 25330 2658 25342
rect 27246 25330 27298 25342
rect 8206 25282 8258 25294
rect 8206 25218 8258 25230
rect 12910 25282 12962 25294
rect 12910 25218 12962 25230
rect 16046 25282 16098 25294
rect 16046 25218 16098 25230
rect 25678 25282 25730 25294
rect 25678 25218 25730 25230
rect 672 25114 27888 25148
rect 672 25062 3806 25114
rect 3858 25062 3910 25114
rect 3962 25062 4014 25114
rect 4066 25062 23806 25114
rect 23858 25062 23910 25114
rect 23962 25062 24014 25114
rect 24066 25062 27888 25114
rect 672 25028 27888 25062
rect 5518 24946 5570 24958
rect 5518 24882 5570 24894
rect 3502 24834 3554 24846
rect 3502 24770 3554 24782
rect 18734 24834 18786 24846
rect 18734 24770 18786 24782
rect 20638 24834 20690 24846
rect 20638 24770 20690 24782
rect 25678 24834 25730 24846
rect 27122 24782 27134 24834
rect 27186 24782 27198 24834
rect 25678 24770 25730 24782
rect 8430 24722 8482 24734
rect 10558 24722 10610 24734
rect 1810 24670 1822 24722
rect 1874 24670 1886 24722
rect 4946 24670 4958 24722
rect 5010 24670 5022 24722
rect 7410 24670 7422 24722
rect 7474 24670 7486 24722
rect 7746 24670 7758 24722
rect 7810 24670 7822 24722
rect 9202 24670 9214 24722
rect 9266 24670 9278 24722
rect 9986 24670 9998 24722
rect 10050 24670 10062 24722
rect 8430 24658 8482 24670
rect 10558 24658 10610 24670
rect 11118 24722 11170 24734
rect 16046 24722 16098 24734
rect 22318 24722 22370 24734
rect 14914 24670 14926 24722
rect 14978 24670 14990 24722
rect 15362 24670 15374 24722
rect 15426 24670 15438 24722
rect 16594 24670 16606 24722
rect 16658 24670 16670 24722
rect 17602 24670 17614 24722
rect 17666 24670 17678 24722
rect 21074 24670 21086 24722
rect 21138 24670 21150 24722
rect 21522 24670 21534 24722
rect 21586 24670 21598 24722
rect 22866 24670 22878 24722
rect 22930 24670 22942 24722
rect 23762 24670 23774 24722
rect 23826 24670 23838 24722
rect 24882 24670 24894 24722
rect 24946 24670 24958 24722
rect 11118 24658 11170 24670
rect 16046 24658 16098 24670
rect 22318 24658 22370 24670
rect 6974 24610 7026 24622
rect 13358 24610 13410 24622
rect 2370 24558 2382 24610
rect 2434 24558 2446 24610
rect 7970 24558 7982 24610
rect 8034 24558 8046 24610
rect 6974 24546 7026 24558
rect 13358 24546 13410 24558
rect 14590 24610 14642 24622
rect 15586 24558 15598 24610
rect 15650 24558 15662 24610
rect 21634 24558 21646 24610
rect 21698 24558 21710 24610
rect 26226 24558 26238 24610
rect 26290 24558 26302 24610
rect 14590 24546 14642 24558
rect 12798 24498 12850 24510
rect 12798 24434 12850 24446
rect 18174 24498 18226 24510
rect 18174 24434 18226 24446
rect 672 24330 27888 24364
rect 672 24278 4466 24330
rect 4518 24278 4570 24330
rect 4622 24278 4674 24330
rect 4726 24278 24466 24330
rect 24518 24278 24570 24330
rect 24622 24278 24674 24330
rect 24726 24278 27888 24330
rect 672 24244 27888 24278
rect 22094 24162 22146 24174
rect 6626 24110 6638 24162
rect 6690 24110 6702 24162
rect 12226 24110 12238 24162
rect 12290 24110 12302 24162
rect 17714 24110 17726 24162
rect 17778 24110 17790 24162
rect 22094 24098 22146 24110
rect 10334 24050 10386 24062
rect 3378 23998 3390 24050
rect 3442 23998 3454 24050
rect 10334 23986 10386 23998
rect 16046 24050 16098 24062
rect 16046 23986 16098 23998
rect 16718 24050 16770 24062
rect 23102 24050 23154 24062
rect 20962 23998 20974 24050
rect 21026 23998 21038 24050
rect 24658 23998 24670 24050
rect 24722 23998 24734 24050
rect 16718 23986 16770 23998
rect 23102 23986 23154 23998
rect 4062 23938 4114 23950
rect 10894 23938 10946 23950
rect 12910 23938 12962 23950
rect 15486 23938 15538 23950
rect 18174 23938 18226 23950
rect 2818 23886 2830 23938
rect 2882 23886 2894 23938
rect 3154 23886 3166 23938
rect 3218 23886 3230 23938
rect 4610 23886 4622 23938
rect 4674 23886 4686 23938
rect 5506 23886 5518 23938
rect 5570 23886 5582 23938
rect 11554 23886 11566 23938
rect 11618 23886 11630 23938
rect 12002 23886 12014 23938
rect 12066 23886 12078 23938
rect 13458 23886 13470 23938
rect 13522 23886 13534 23938
rect 14354 23886 14366 23938
rect 14418 23886 14430 23938
rect 17042 23886 17054 23938
rect 17106 23886 17118 23938
rect 17602 23886 17614 23938
rect 17666 23886 17678 23938
rect 18946 23886 18958 23938
rect 19010 23886 19022 23938
rect 19730 23886 19742 23938
rect 19794 23886 19806 23938
rect 20402 23886 20414 23938
rect 20466 23886 20478 23938
rect 22642 23886 22654 23938
rect 22706 23886 22718 23938
rect 26226 23886 26238 23938
rect 26290 23886 26302 23938
rect 4062 23874 4114 23886
rect 10894 23874 10946 23886
rect 12910 23874 12962 23886
rect 15486 23874 15538 23886
rect 18174 23874 18226 23886
rect 2382 23826 2434 23838
rect 11230 23826 11282 23838
rect 6178 23774 6190 23826
rect 6242 23774 6254 23826
rect 2382 23762 2434 23774
rect 11230 23762 11282 23774
rect 27246 23826 27298 23838
rect 27246 23762 27298 23774
rect 7758 23714 7810 23726
rect 7758 23650 7810 23662
rect 25678 23714 25730 23726
rect 25678 23650 25730 23662
rect 672 23546 27888 23580
rect 672 23494 3806 23546
rect 3858 23494 3910 23546
rect 3962 23494 4014 23546
rect 4066 23494 23806 23546
rect 23858 23494 23910 23546
rect 23962 23494 24014 23546
rect 24066 23494 27888 23546
rect 672 23460 27888 23494
rect 3838 23378 3890 23390
rect 3838 23314 3890 23326
rect 16270 23378 16322 23390
rect 16270 23314 16322 23326
rect 27246 23378 27298 23390
rect 27246 23314 27298 23326
rect 1150 23266 1202 23278
rect 13246 23266 13298 23278
rect 2258 23214 2270 23266
rect 2322 23214 2334 23266
rect 6962 23214 6974 23266
rect 7026 23214 7038 23266
rect 9314 23214 9326 23266
rect 9378 23214 9390 23266
rect 1150 23202 1202 23214
rect 13246 23202 13298 23214
rect 19966 23154 20018 23166
rect 1586 23102 1598 23154
rect 1650 23102 1662 23154
rect 10322 23102 10334 23154
rect 10386 23102 10398 23154
rect 14690 23102 14702 23154
rect 14754 23102 14766 23154
rect 19966 23090 20018 23102
rect 5182 23042 5234 23054
rect 19630 23042 19682 23054
rect 2706 22990 2718 23042
rect 2770 22990 2782 23042
rect 6066 22990 6078 23042
rect 6130 22990 6142 23042
rect 8866 22990 8878 23042
rect 8930 22990 8942 23042
rect 15138 22990 15150 23042
rect 15202 22990 15214 23042
rect 26226 22990 26238 23042
rect 26290 22990 26302 23042
rect 5182 22978 5234 22990
rect 19630 22978 19682 22990
rect 5742 22930 5794 22942
rect 5742 22866 5794 22878
rect 7758 22930 7810 22942
rect 12014 22930 12066 22942
rect 10882 22878 10894 22930
rect 10946 22878 10958 22930
rect 7758 22866 7810 22878
rect 12014 22866 12066 22878
rect 13806 22930 13858 22942
rect 13806 22866 13858 22878
rect 19854 22930 19906 22942
rect 19854 22866 19906 22878
rect 20078 22930 20130 22942
rect 20078 22866 20130 22878
rect 672 22762 27888 22796
rect 672 22710 4466 22762
rect 4518 22710 4570 22762
rect 4622 22710 4674 22762
rect 4726 22710 24466 22762
rect 24518 22710 24570 22762
rect 24622 22710 24674 22762
rect 24726 22710 27888 22762
rect 672 22676 27888 22710
rect 2830 22594 2882 22606
rect 2830 22530 2882 22542
rect 13358 22594 13410 22606
rect 13358 22530 13410 22542
rect 23438 22482 23490 22494
rect 1586 22430 1598 22482
rect 1650 22430 1662 22482
rect 6066 22430 6078 22482
rect 6130 22430 6142 22482
rect 9986 22430 9998 22482
rect 10050 22430 10062 22482
rect 12226 22430 12238 22482
rect 12290 22430 12302 22482
rect 14802 22430 14814 22482
rect 14866 22430 14878 22482
rect 18050 22430 18062 22482
rect 18114 22430 18126 22482
rect 20290 22430 20302 22482
rect 20354 22430 20366 22482
rect 26226 22430 26238 22482
rect 26290 22430 26302 22482
rect 23438 22418 23490 22430
rect 20750 22370 20802 22382
rect 22878 22370 22930 22382
rect 1250 22318 1262 22370
rect 1314 22318 1326 22370
rect 4274 22318 4286 22370
rect 4338 22318 4350 22370
rect 5618 22318 5630 22370
rect 5682 22318 5694 22370
rect 9538 22318 9550 22370
rect 9602 22318 9614 22370
rect 11778 22318 11790 22370
rect 11842 22318 11854 22370
rect 18386 22318 18398 22370
rect 18450 22318 18462 22370
rect 19618 22318 19630 22370
rect 19682 22318 19694 22370
rect 20066 22318 20078 22370
rect 20130 22318 20142 22370
rect 21298 22318 21310 22370
rect 21362 22318 21374 22370
rect 21522 22318 21534 22370
rect 21586 22318 21598 22370
rect 22306 22318 22318 22370
rect 22370 22318 22382 22370
rect 24882 22318 24894 22370
rect 24946 22318 24958 22370
rect 20750 22306 20802 22318
rect 22878 22306 22930 22318
rect 3502 22258 3554 22270
rect 19294 22258 19346 22270
rect 14466 22206 14478 22258
rect 14530 22206 14542 22258
rect 3502 22194 3554 22206
rect 19294 22194 19346 22206
rect 27246 22258 27298 22270
rect 27246 22194 27298 22206
rect 7198 22146 7250 22158
rect 7198 22082 7250 22094
rect 11118 22146 11170 22158
rect 11118 22082 11170 22094
rect 16046 22146 16098 22158
rect 16046 22082 16098 22094
rect 16830 22146 16882 22158
rect 16830 22082 16882 22094
rect 25678 22146 25730 22158
rect 25678 22082 25730 22094
rect 672 21978 27888 22012
rect 672 21926 3806 21978
rect 3858 21926 3910 21978
rect 3962 21926 4014 21978
rect 4066 21926 23806 21978
rect 23858 21926 23910 21978
rect 23962 21926 24014 21978
rect 24066 21926 27888 21978
rect 672 21892 27888 21926
rect 22082 21758 22094 21810
rect 22146 21758 22158 21810
rect 18510 21698 18562 21710
rect 18162 21646 18174 21698
rect 18226 21646 18238 21698
rect 23874 21646 23886 21698
rect 23938 21646 23950 21698
rect 25778 21646 25790 21698
rect 25842 21646 25854 21698
rect 27122 21646 27134 21698
rect 27186 21646 27198 21698
rect 18510 21634 18562 21646
rect 7086 21586 7138 21598
rect 12126 21586 12178 21598
rect 16158 21586 16210 21598
rect 19294 21586 19346 21598
rect 20638 21586 20690 21598
rect 21982 21586 22034 21598
rect 2594 21534 2606 21586
rect 2658 21534 2670 21586
rect 5394 21534 5406 21586
rect 5458 21534 5470 21586
rect 6514 21534 6526 21586
rect 6578 21534 6590 21586
rect 7746 21534 7758 21586
rect 7810 21534 7822 21586
rect 8082 21534 8094 21586
rect 8146 21534 8158 21586
rect 10546 21534 10558 21586
rect 10610 21534 10622 21586
rect 14802 21534 14814 21586
rect 14866 21534 14878 21586
rect 15250 21534 15262 21586
rect 15314 21534 15326 21586
rect 16482 21534 16494 21586
rect 16546 21534 16558 21586
rect 17602 21534 17614 21586
rect 17666 21534 17678 21586
rect 19058 21534 19070 21586
rect 19122 21534 19134 21586
rect 19618 21534 19630 21586
rect 19682 21534 19694 21586
rect 20850 21534 20862 21586
rect 20914 21534 20926 21586
rect 21074 21534 21086 21586
rect 21138 21534 21150 21586
rect 22194 21534 22206 21586
rect 22258 21534 22270 21586
rect 23538 21534 23550 21586
rect 23602 21534 23614 21586
rect 7086 21522 7138 21534
rect 12126 21522 12178 21534
rect 16158 21522 16210 21534
rect 19294 21522 19346 21534
rect 20638 21522 20690 21534
rect 21982 21522 22034 21534
rect 8542 21474 8594 21486
rect 3154 21422 3166 21474
rect 3218 21422 3230 21474
rect 7522 21422 7534 21474
rect 7586 21422 7598 21474
rect 8542 21410 8594 21422
rect 14030 21474 14082 21486
rect 14030 21410 14082 21422
rect 14478 21474 14530 21486
rect 18846 21474 18898 21486
rect 15474 21422 15486 21474
rect 15538 21422 15550 21474
rect 14478 21410 14530 21422
rect 18846 21410 18898 21422
rect 20078 21474 20130 21486
rect 26226 21422 26238 21474
rect 26290 21422 26302 21474
rect 20078 21410 20130 21422
rect 4286 21362 4338 21374
rect 13470 21362 13522 21374
rect 10994 21310 11006 21362
rect 11058 21310 11070 21362
rect 4286 21298 4338 21310
rect 13470 21298 13522 21310
rect 18286 21362 18338 21374
rect 18286 21298 18338 21310
rect 19630 21362 19682 21374
rect 19630 21298 19682 21310
rect 19966 21362 20018 21374
rect 19966 21298 20018 21310
rect 25342 21362 25394 21374
rect 25342 21298 25394 21310
rect 672 21194 27888 21228
rect 672 21142 4466 21194
rect 4518 21142 4570 21194
rect 4622 21142 4674 21194
rect 4726 21142 24466 21194
rect 24518 21142 24570 21194
rect 24622 21142 24674 21194
rect 24726 21142 27888 21194
rect 672 21108 27888 21142
rect 17950 21026 18002 21038
rect 6962 20974 6974 21026
rect 7026 20974 7038 21026
rect 11330 20974 11342 21026
rect 11394 20974 11406 21026
rect 19730 20974 19742 21026
rect 19794 20974 19806 21026
rect 17950 20962 18002 20974
rect 1262 20914 1314 20926
rect 1262 20850 1314 20862
rect 1822 20914 1874 20926
rect 10334 20914 10386 20926
rect 26462 20914 26514 20926
rect 3154 20862 3166 20914
rect 3218 20862 3230 20914
rect 14802 20862 14814 20914
rect 14866 20862 14878 20914
rect 16930 20862 16942 20914
rect 16994 20862 17006 20914
rect 17266 20862 17278 20914
rect 17330 20862 17342 20914
rect 1822 20850 1874 20862
rect 10334 20850 10386 20862
rect 26462 20850 26514 20862
rect 27358 20914 27410 20926
rect 27358 20850 27410 20862
rect 3614 20802 3666 20814
rect 8878 20802 8930 20814
rect 12014 20802 12066 20814
rect 16046 20802 16098 20814
rect 20190 20802 20242 20814
rect 25902 20802 25954 20814
rect 2594 20750 2606 20802
rect 2658 20750 2670 20802
rect 2930 20750 2942 20802
rect 2994 20750 3006 20802
rect 4386 20750 4398 20802
rect 4450 20750 4462 20802
rect 5170 20750 5182 20802
rect 5234 20750 5246 20802
rect 10770 20750 10782 20802
rect 10834 20750 10846 20802
rect 11106 20750 11118 20802
rect 11170 20750 11182 20802
rect 12338 20750 12350 20802
rect 12402 20750 12414 20802
rect 13346 20750 13358 20802
rect 13410 20750 13422 20802
rect 14466 20750 14478 20802
rect 14530 20750 14542 20802
rect 16818 20750 16830 20802
rect 16882 20750 16894 20802
rect 17154 20750 17166 20802
rect 17218 20750 17230 20802
rect 19058 20750 19070 20802
rect 19122 20750 19134 20802
rect 19506 20750 19518 20802
rect 19570 20750 19582 20802
rect 20738 20750 20750 20802
rect 20802 20750 20814 20802
rect 21746 20750 21758 20802
rect 21810 20750 21822 20802
rect 26898 20750 26910 20802
rect 26962 20750 26974 20802
rect 3614 20738 3666 20750
rect 8878 20738 8930 20750
rect 12014 20738 12066 20750
rect 16046 20738 16098 20750
rect 20190 20738 20242 20750
rect 25902 20738 25954 20750
rect 2158 20690 2210 20702
rect 9438 20690 9490 20702
rect 7410 20638 7422 20690
rect 7474 20638 7486 20690
rect 2158 20626 2210 20638
rect 9438 20626 9490 20638
rect 18734 20690 18786 20702
rect 18734 20626 18786 20638
rect 5854 20578 5906 20590
rect 5854 20514 5906 20526
rect 17614 20578 17666 20590
rect 17614 20514 17666 20526
rect 672 20410 27888 20444
rect 672 20358 3806 20410
rect 3858 20358 3910 20410
rect 3962 20358 4014 20410
rect 4066 20358 23806 20410
rect 23858 20358 23910 20410
rect 23962 20358 24014 20410
rect 24066 20358 27888 20410
rect 672 20324 27888 20358
rect 5518 20242 5570 20254
rect 5518 20178 5570 20190
rect 3278 20130 3330 20142
rect 20638 20130 20690 20142
rect 11218 20078 11230 20130
rect 11282 20078 11294 20130
rect 20962 20078 20974 20130
rect 21026 20078 21038 20130
rect 3278 20066 3330 20078
rect 20638 20066 20690 20078
rect 8430 20018 8482 20030
rect 14478 20018 14530 20030
rect 19966 20018 20018 20030
rect 1698 19966 1710 20018
rect 1762 19966 1774 20018
rect 5170 19966 5182 20018
rect 5234 19966 5246 20018
rect 7298 19966 7310 20018
rect 7362 19966 7374 20018
rect 7858 19966 7870 20018
rect 7922 19966 7934 20018
rect 9202 19966 9214 20018
rect 9266 19966 9278 20018
rect 9986 19966 9998 20018
rect 10050 19966 10062 20018
rect 10546 19966 10558 20018
rect 10610 19966 10622 20018
rect 13122 19966 13134 20018
rect 13186 19966 13198 20018
rect 13570 19966 13582 20018
rect 13634 19966 13646 20018
rect 14802 19966 14814 20018
rect 14866 19966 14878 20018
rect 15810 19966 15822 20018
rect 15874 19966 15886 20018
rect 16482 19966 16494 20018
rect 16546 19966 16558 20018
rect 19730 19966 19742 20018
rect 19794 19966 19806 20018
rect 8430 19954 8482 19966
rect 14478 19954 14530 19966
rect 19966 19954 20018 19966
rect 6974 19906 7026 19918
rect 12798 19906 12850 19918
rect 18622 19906 18674 19918
rect 7970 19854 7982 19906
rect 8034 19854 8046 19906
rect 13794 19854 13806 19906
rect 13858 19854 13870 19906
rect 17042 19854 17054 19906
rect 17106 19854 17118 19906
rect 6974 19842 7026 19854
rect 12798 19842 12850 19854
rect 18622 19842 18674 19854
rect 20078 19906 20130 19918
rect 20078 19842 20130 19854
rect 11118 19794 11170 19806
rect 2146 19742 2158 19794
rect 2210 19742 2222 19794
rect 11118 19730 11170 19742
rect 18174 19794 18226 19806
rect 18174 19730 18226 19742
rect 18734 19794 18786 19806
rect 18734 19730 18786 19742
rect 18846 19794 18898 19806
rect 18846 19730 18898 19742
rect 20862 19794 20914 19806
rect 20862 19730 20914 19742
rect 672 19626 27888 19660
rect 672 19574 4466 19626
rect 4518 19574 4570 19626
rect 4622 19574 4674 19626
rect 4726 19574 24466 19626
rect 24518 19574 24570 19626
rect 24622 19574 24674 19626
rect 24726 19574 27888 19626
rect 672 19540 27888 19574
rect 9326 19458 9378 19470
rect 25902 19458 25954 19470
rect 10882 19406 10894 19458
rect 10946 19406 10958 19458
rect 13458 19406 13470 19458
rect 13522 19406 13534 19458
rect 17378 19406 17390 19458
rect 17442 19406 17454 19458
rect 20290 19406 20302 19458
rect 20354 19406 20366 19458
rect 9326 19394 9378 19406
rect 25902 19394 25954 19406
rect 6526 19346 6578 19358
rect 2258 19294 2270 19346
rect 2322 19294 2334 19346
rect 3490 19294 3502 19346
rect 3554 19294 3566 19346
rect 6066 19294 6078 19346
rect 6130 19294 6142 19346
rect 6526 19282 6578 19294
rect 9886 19346 9938 19358
rect 9886 19282 9938 19294
rect 12014 19346 12066 19358
rect 12014 19282 12066 19294
rect 26462 19346 26514 19358
rect 26462 19282 26514 19294
rect 4622 19234 4674 19246
rect 13918 19234 13970 19246
rect 16046 19234 16098 19246
rect 5394 19182 5406 19234
rect 5458 19182 5470 19234
rect 5842 19182 5854 19234
rect 5906 19182 5918 19234
rect 7074 19182 7086 19234
rect 7138 19182 7150 19234
rect 7298 19182 7310 19234
rect 7362 19182 7374 19234
rect 8194 19182 8206 19234
rect 8258 19182 8270 19234
rect 10322 19182 10334 19234
rect 10386 19182 10398 19234
rect 12786 19182 12798 19234
rect 12850 19182 12862 19234
rect 13234 19182 13246 19234
rect 13298 19182 13310 19234
rect 14466 19182 14478 19234
rect 14530 19182 14542 19234
rect 15474 19182 15486 19234
rect 15538 19182 15550 19234
rect 4622 19170 4674 19182
rect 13918 19170 13970 19182
rect 16046 19170 16098 19182
rect 16942 19234 16994 19246
rect 16942 19170 16994 19182
rect 17278 19234 17330 19246
rect 17278 19170 17330 19182
rect 17390 19234 17442 19246
rect 19630 19234 19682 19246
rect 17714 19182 17726 19234
rect 17778 19182 17790 19234
rect 18274 19182 18286 19234
rect 18338 19182 18350 19234
rect 19282 19182 19294 19234
rect 19346 19182 19358 19234
rect 20402 19182 20414 19234
rect 20466 19182 20478 19234
rect 20850 19182 20862 19234
rect 20914 19182 20926 19234
rect 17390 19170 17442 19182
rect 19630 19170 19682 19182
rect 5070 19122 5122 19134
rect 1362 19070 1374 19122
rect 1426 19070 1438 19122
rect 3042 19070 3054 19122
rect 3106 19070 3118 19122
rect 5070 19058 5122 19070
rect 12462 19122 12514 19134
rect 12462 19058 12514 19070
rect 16158 19122 16210 19134
rect 16158 19058 16210 19070
rect 21310 19122 21362 19134
rect 21310 19058 21362 19070
rect 672 18842 27888 18876
rect 672 18790 3806 18842
rect 3858 18790 3910 18842
rect 3962 18790 4014 18842
rect 4066 18790 23806 18842
rect 23858 18790 23910 18842
rect 23962 18790 24014 18842
rect 24066 18790 27888 18842
rect 672 18756 27888 18790
rect 12126 18674 12178 18686
rect 12126 18610 12178 18622
rect 14590 18674 14642 18686
rect 14590 18610 14642 18622
rect 2706 18510 2718 18562
rect 2770 18510 2782 18562
rect 5058 18510 5070 18562
rect 5122 18510 5134 18562
rect 6066 18510 6078 18562
rect 6130 18510 6142 18562
rect 10546 18510 10558 18562
rect 10610 18510 10622 18562
rect 13010 18510 13022 18562
rect 13074 18510 13086 18562
rect 2158 18450 2210 18462
rect 1698 18398 1710 18450
rect 1762 18398 1774 18450
rect 2158 18386 2210 18398
rect 5518 18450 5570 18462
rect 5518 18386 5570 18398
rect 7646 18450 7698 18462
rect 19070 18450 19122 18462
rect 8306 18398 8318 18450
rect 8370 18398 8382 18450
rect 15698 18398 15710 18450
rect 15762 18398 15774 18450
rect 16706 18398 16718 18450
rect 16770 18398 16782 18450
rect 17938 18398 17950 18450
rect 18002 18398 18014 18450
rect 18498 18398 18510 18450
rect 18562 18398 18574 18450
rect 20962 18398 20974 18450
rect 21026 18398 21038 18450
rect 21410 18398 21422 18450
rect 21474 18398 21486 18450
rect 22642 18398 22654 18450
rect 22706 18398 22718 18450
rect 23650 18398 23662 18450
rect 23714 18398 23726 18450
rect 7646 18386 7698 18398
rect 19070 18386 19122 18398
rect 17390 18338 17442 18350
rect 18846 18338 18898 18350
rect 6514 18286 6526 18338
rect 6578 18286 6590 18338
rect 8754 18286 8766 18338
rect 8818 18286 8830 18338
rect 10994 18286 11006 18338
rect 11058 18286 11070 18338
rect 13346 18286 13358 18338
rect 13410 18286 13422 18338
rect 17826 18286 17838 18338
rect 17890 18286 17902 18338
rect 17390 18274 17442 18286
rect 18846 18274 18898 18286
rect 20638 18338 20690 18350
rect 20638 18274 20690 18286
rect 22094 18338 22146 18350
rect 22094 18274 22146 18286
rect 4286 18226 4338 18238
rect 3154 18174 3166 18226
rect 3218 18174 3230 18226
rect 4286 18162 4338 18174
rect 9886 18226 9938 18238
rect 9886 18162 9938 18174
rect 19518 18226 19570 18238
rect 19518 18162 19570 18174
rect 19630 18226 19682 18238
rect 19630 18162 19682 18174
rect 19742 18226 19794 18238
rect 21634 18174 21646 18226
rect 21698 18174 21710 18226
rect 19742 18162 19794 18174
rect 672 18058 27888 18092
rect 672 18006 4466 18058
rect 4518 18006 4570 18058
rect 4622 18006 4674 18058
rect 4726 18006 24466 18058
rect 24518 18006 24570 18058
rect 24622 18006 24674 18058
rect 24726 18006 27888 18058
rect 672 17972 27888 18006
rect 13806 17890 13858 17902
rect 3714 17838 3726 17890
rect 3778 17838 3790 17890
rect 12674 17838 12686 17890
rect 12738 17838 12750 17890
rect 13806 17826 13858 17838
rect 16830 17890 16882 17902
rect 16830 17826 16882 17838
rect 6526 17778 6578 17790
rect 6066 17726 6078 17778
rect 6130 17726 6142 17778
rect 6526 17714 6578 17726
rect 8878 17778 8930 17790
rect 8878 17714 8930 17726
rect 9438 17778 9490 17790
rect 15150 17778 15202 17790
rect 10434 17726 10446 17778
rect 10498 17726 10510 17778
rect 9438 17714 9490 17726
rect 15150 17714 15202 17726
rect 17502 17778 17554 17790
rect 17502 17714 17554 17726
rect 17838 17778 17890 17790
rect 24558 17778 24610 17790
rect 18834 17726 18846 17778
rect 18898 17726 18910 17778
rect 22642 17726 22654 17778
rect 22706 17726 22718 17778
rect 17838 17714 17890 17726
rect 24558 17714 24610 17726
rect 1822 17671 1874 17683
rect 3278 17666 3330 17678
rect 4734 17666 4786 17678
rect 15710 17666 15762 17678
rect 1822 17607 1874 17619
rect 2706 17614 2718 17666
rect 2770 17614 2782 17666
rect 3826 17614 3838 17666
rect 3890 17614 3902 17666
rect 4274 17614 4286 17666
rect 4338 17614 4350 17666
rect 5394 17614 5406 17666
rect 5458 17614 5470 17666
rect 5954 17614 5966 17666
rect 6018 17614 6030 17666
rect 7298 17614 7310 17666
rect 7362 17614 7374 17666
rect 8194 17614 8206 17666
rect 8258 17614 8270 17666
rect 12114 17614 12126 17666
rect 12178 17614 12190 17666
rect 3278 17602 3330 17614
rect 4734 17602 4786 17614
rect 15710 17602 15762 17614
rect 16718 17666 16770 17678
rect 19294 17666 19346 17678
rect 21534 17666 21586 17678
rect 17154 17614 17166 17666
rect 17218 17614 17230 17666
rect 18162 17614 18174 17666
rect 18226 17614 18238 17666
rect 18610 17614 18622 17666
rect 18674 17614 18686 17666
rect 19842 17614 19854 17666
rect 19906 17614 19918 17666
rect 20066 17614 20078 17666
rect 20130 17614 20142 17666
rect 20962 17614 20974 17666
rect 21026 17614 21038 17666
rect 24994 17614 25006 17666
rect 25058 17614 25070 17666
rect 16718 17602 16770 17614
rect 19294 17602 19346 17614
rect 21534 17602 21586 17614
rect 5070 17554 5122 17566
rect 17390 17554 17442 17566
rect 9986 17502 9998 17554
rect 10050 17502 10062 17554
rect 23090 17502 23102 17554
rect 23154 17502 23166 17554
rect 5070 17490 5122 17502
rect 17390 17490 17442 17502
rect 11566 17442 11618 17454
rect 11566 17378 11618 17390
rect 672 17274 27888 17308
rect 672 17222 3806 17274
rect 3858 17222 3910 17274
rect 3962 17222 4014 17274
rect 4066 17222 23806 17274
rect 23858 17222 23910 17274
rect 23962 17222 24014 17274
rect 24066 17222 27888 17274
rect 672 17188 27888 17222
rect 2830 17106 2882 17118
rect 2830 17042 2882 17054
rect 5518 17106 5570 17118
rect 5518 17042 5570 17054
rect 18286 17106 18338 17118
rect 18286 17042 18338 17054
rect 18510 17106 18562 17118
rect 18510 17042 18562 17054
rect 19966 17106 20018 17118
rect 19966 17042 20018 17054
rect 20974 17106 21026 17118
rect 20974 17042 21026 17054
rect 1250 16942 1262 16994
rect 1314 16942 1326 16994
rect 3714 16942 3726 16994
rect 3778 16942 3790 16994
rect 19058 16942 19070 16994
rect 19122 16942 19134 16994
rect 19618 16942 19630 16994
rect 19682 16942 19694 16994
rect 10446 16882 10498 16894
rect 16158 16882 16210 16894
rect 3378 16830 3390 16882
rect 3442 16830 3454 16882
rect 4946 16830 4958 16882
rect 5010 16830 5022 16882
rect 8418 16830 8430 16882
rect 8482 16830 8494 16882
rect 9314 16830 9326 16882
rect 9378 16830 9390 16882
rect 9762 16830 9774 16882
rect 9826 16830 9838 16882
rect 10994 16830 11006 16882
rect 11058 16830 11070 16882
rect 12002 16830 12014 16882
rect 12066 16830 12078 16882
rect 15026 16830 15038 16882
rect 15090 16830 15102 16882
rect 15474 16830 15486 16882
rect 15538 16830 15550 16882
rect 16930 16830 16942 16882
rect 16994 16830 17006 16882
rect 17614 16877 17666 16889
rect 10446 16818 10498 16830
rect 16158 16818 16210 16830
rect 17614 16813 17666 16825
rect 18734 16882 18786 16894
rect 18734 16818 18786 16830
rect 19182 16882 19234 16894
rect 23762 16830 23774 16882
rect 23826 16830 23838 16882
rect 19182 16818 19234 16830
rect 8990 16770 9042 16782
rect 1586 16718 1598 16770
rect 1650 16718 1662 16770
rect 7970 16718 7982 16770
rect 8034 16718 8046 16770
rect 8990 16706 9042 16718
rect 14702 16770 14754 16782
rect 15698 16718 15710 16770
rect 15762 16718 15774 16770
rect 23314 16718 23326 16770
rect 23378 16718 23390 16770
rect 14702 16706 14754 16718
rect 6862 16658 6914 16670
rect 18958 16658 19010 16670
rect 9986 16606 9998 16658
rect 10050 16606 10062 16658
rect 6862 16594 6914 16606
rect 18958 16594 19010 16606
rect 19742 16658 19794 16670
rect 19742 16594 19794 16606
rect 20750 16658 20802 16670
rect 20750 16594 20802 16606
rect 20862 16658 20914 16670
rect 20862 16594 20914 16606
rect 22206 16658 22258 16670
rect 22206 16594 22258 16606
rect 672 16490 27888 16524
rect 672 16438 4466 16490
rect 4518 16438 4570 16490
rect 4622 16438 4674 16490
rect 4726 16438 24466 16490
rect 24518 16438 24570 16490
rect 24622 16438 24674 16490
rect 24726 16438 27888 16490
rect 672 16404 27888 16438
rect 2942 16322 2994 16334
rect 1810 16270 1822 16322
rect 1874 16270 1886 16322
rect 2942 16258 2994 16270
rect 5182 16322 5234 16334
rect 8206 16322 8258 16334
rect 7074 16270 7086 16322
rect 7138 16270 7150 16322
rect 5182 16258 5234 16270
rect 8206 16258 8258 16270
rect 9102 16322 9154 16334
rect 12798 16322 12850 16334
rect 11666 16270 11678 16322
rect 11730 16270 11742 16322
rect 17042 16270 17054 16322
rect 17106 16270 17118 16322
rect 18274 16270 18286 16322
rect 18338 16270 18350 16322
rect 19954 16270 19966 16322
rect 20018 16270 20030 16322
rect 9102 16258 9154 16270
rect 12798 16258 12850 16270
rect 5966 16210 6018 16222
rect 4050 16158 4062 16210
rect 4114 16158 4126 16210
rect 5966 16146 6018 16158
rect 10446 16210 10498 16222
rect 16046 16210 16098 16222
rect 13794 16158 13806 16210
rect 13858 16158 13870 16210
rect 10446 16146 10498 16158
rect 16046 16146 16098 16158
rect 18958 16210 19010 16222
rect 18958 16146 19010 16158
rect 20414 16210 20466 16222
rect 20414 16146 20466 16158
rect 5854 16098 5906 16110
rect 1362 16046 1374 16098
rect 1426 16046 1438 16098
rect 3602 16046 3614 16098
rect 3666 16046 3678 16098
rect 5854 16034 5906 16046
rect 6190 16098 6242 16110
rect 16718 16098 16770 16110
rect 17838 16098 17890 16110
rect 18286 16098 18338 16110
rect 9986 16046 9998 16098
rect 10050 16046 10062 16098
rect 11106 16046 11118 16098
rect 11170 16046 11182 16098
rect 13458 16046 13470 16098
rect 13522 16046 13534 16098
rect 15586 16046 15598 16098
rect 15650 16046 15662 16098
rect 16930 16046 16942 16098
rect 16994 16046 17006 16098
rect 17490 16046 17502 16098
rect 17554 16046 17566 16098
rect 18050 16046 18062 16098
rect 18114 16046 18126 16098
rect 18610 16046 18622 16098
rect 18674 16046 18686 16098
rect 19394 16046 19406 16098
rect 19458 16046 19470 16098
rect 19730 16046 19742 16098
rect 19794 16046 19806 16098
rect 21186 16046 21198 16098
rect 21250 16046 21262 16098
rect 21970 16046 21982 16098
rect 22034 16046 22046 16098
rect 6190 16034 6242 16046
rect 16718 16034 16770 16046
rect 17838 16034 17890 16046
rect 18286 16034 18338 16046
rect 6626 15934 6638 15986
rect 6690 15934 6702 15986
rect 9090 15934 9102 15986
rect 9154 15934 9166 15986
rect 8878 15874 8930 15886
rect 8878 15810 8930 15822
rect 15038 15874 15090 15886
rect 17266 15822 17278 15874
rect 17330 15822 17342 15874
rect 15038 15810 15090 15822
rect 672 15706 27888 15740
rect 672 15654 3806 15706
rect 3858 15654 3910 15706
rect 3962 15654 4014 15706
rect 4066 15654 23806 15706
rect 23858 15654 23910 15706
rect 23962 15654 24014 15706
rect 24066 15654 27888 15706
rect 672 15620 27888 15654
rect 9886 15538 9938 15550
rect 9886 15474 9938 15486
rect 12126 15538 12178 15550
rect 18610 15486 18622 15538
rect 18674 15486 18686 15538
rect 12126 15474 12178 15486
rect 2158 15426 2210 15438
rect 20638 15426 20690 15438
rect 5170 15374 5182 15426
rect 5234 15374 5246 15426
rect 10546 15374 10558 15426
rect 10610 15374 10622 15426
rect 19730 15374 19742 15426
rect 19794 15374 19806 15426
rect 2158 15362 2210 15374
rect 20638 15362 20690 15374
rect 6750 15314 6802 15326
rect 1698 15262 1710 15314
rect 1762 15262 1774 15314
rect 4274 15262 4286 15314
rect 4338 15262 4350 15314
rect 6750 15250 6802 15262
rect 7086 15314 7138 15326
rect 7086 15250 7138 15262
rect 7534 15314 7586 15326
rect 7534 15250 7586 15262
rect 7758 15314 7810 15326
rect 14366 15314 14418 15326
rect 16158 15314 16210 15326
rect 18846 15314 18898 15326
rect 8194 15262 8206 15314
rect 8258 15262 8270 15314
rect 15138 15262 15150 15314
rect 15202 15262 15214 15314
rect 15474 15262 15486 15314
rect 15538 15262 15550 15314
rect 16818 15262 16830 15314
rect 16882 15262 16894 15314
rect 17714 15262 17726 15314
rect 17778 15262 17790 15314
rect 18498 15262 18510 15314
rect 18562 15262 18574 15314
rect 7758 15250 7810 15262
rect 14366 15250 14418 15262
rect 16158 15250 16210 15262
rect 18846 15250 18898 15262
rect 19182 15314 19234 15326
rect 20962 15262 20974 15314
rect 21026 15262 21038 15314
rect 21410 15262 21422 15314
rect 21474 15262 21486 15314
rect 22866 15262 22878 15314
rect 22930 15262 22942 15314
rect 23650 15262 23662 15314
rect 23714 15262 23726 15314
rect 19182 15250 19234 15262
rect 2606 15202 2658 15214
rect 14702 15202 14754 15214
rect 20078 15202 20130 15214
rect 22094 15202 22146 15214
rect 3826 15150 3838 15202
rect 3890 15150 3902 15202
rect 5618 15150 5630 15202
rect 5682 15150 5694 15202
rect 8754 15150 8766 15202
rect 8818 15150 8830 15202
rect 10994 15150 11006 15202
rect 11058 15150 11070 15202
rect 15698 15150 15710 15202
rect 15762 15150 15774 15202
rect 21634 15150 21646 15202
rect 21698 15150 21710 15202
rect 2606 15138 2658 15150
rect 14702 15138 14754 15150
rect 20078 15138 20130 15150
rect 22094 15138 22146 15150
rect 7646 15090 7698 15102
rect 7646 15026 7698 15038
rect 14030 15090 14082 15102
rect 14030 15026 14082 15038
rect 18398 15090 18450 15102
rect 18398 15026 18450 15038
rect 19854 15090 19906 15102
rect 19854 15026 19906 15038
rect 672 14922 27888 14956
rect 672 14870 4466 14922
rect 4518 14870 4570 14922
rect 4622 14870 4674 14922
rect 4726 14870 24466 14922
rect 24518 14870 24570 14922
rect 24622 14870 24674 14922
rect 24726 14870 27888 14922
rect 672 14836 27888 14870
rect 3278 14754 3330 14766
rect 9102 14754 9154 14766
rect 5730 14702 5742 14754
rect 5794 14702 5806 14754
rect 3278 14690 3330 14702
rect 9102 14690 9154 14702
rect 12462 14754 12514 14766
rect 16830 14754 16882 14766
rect 13570 14702 13582 14754
rect 13634 14702 13646 14754
rect 22530 14702 22542 14754
rect 22594 14702 22606 14754
rect 12462 14690 12514 14702
rect 16830 14690 16882 14702
rect 4286 14642 4338 14654
rect 2146 14590 2158 14642
rect 2210 14590 2222 14642
rect 4286 14578 4338 14590
rect 6862 14642 6914 14654
rect 6862 14578 6914 14590
rect 8878 14642 8930 14654
rect 8878 14578 8930 14590
rect 9326 14642 9378 14654
rect 9326 14578 9378 14590
rect 10334 14642 10386 14654
rect 14702 14642 14754 14654
rect 11330 14590 11342 14642
rect 11394 14590 11406 14642
rect 10334 14578 10386 14590
rect 14702 14578 14754 14590
rect 15710 14642 15762 14654
rect 15710 14578 15762 14590
rect 16942 14642 16994 14654
rect 16942 14578 16994 14590
rect 17726 14642 17778 14654
rect 19182 14642 19234 14654
rect 18722 14590 18734 14642
rect 18786 14590 18798 14642
rect 25218 14590 25230 14642
rect 25282 14590 25294 14642
rect 17726 14578 17778 14590
rect 19182 14578 19234 14590
rect 4174 14530 4226 14542
rect 7982 14530 8034 14542
rect 1586 14478 1598 14530
rect 1650 14478 1662 14530
rect 3938 14478 3950 14530
rect 4002 14478 4014 14530
rect 5170 14478 5182 14530
rect 5234 14478 5246 14530
rect 7858 14478 7870 14530
rect 7922 14478 7934 14530
rect 4174 14466 4226 14478
rect 7982 14466 8034 14478
rect 8206 14530 8258 14542
rect 8206 14466 8258 14478
rect 8766 14530 8818 14542
rect 15150 14530 15202 14542
rect 9874 14478 9886 14530
rect 9938 14478 9950 14530
rect 8766 14466 8818 14478
rect 15150 14466 15202 14478
rect 16046 14530 16098 14542
rect 16046 14466 16098 14478
rect 16718 14530 16770 14542
rect 18050 14478 18062 14530
rect 18114 14478 18126 14530
rect 18498 14478 18510 14530
rect 18562 14478 18574 14530
rect 19954 14478 19966 14530
rect 20018 14478 20030 14530
rect 20738 14478 20750 14530
rect 20802 14478 20814 14530
rect 16718 14466 16770 14478
rect 8082 14366 8094 14418
rect 8146 14366 8158 14418
rect 10882 14366 10894 14418
rect 10946 14366 10958 14418
rect 13122 14366 13134 14418
rect 13186 14366 13198 14418
rect 22978 14366 22990 14418
rect 23042 14366 23054 14418
rect 24770 14366 24782 14418
rect 24834 14366 24846 14418
rect 7310 14306 7362 14318
rect 4722 14254 4734 14306
rect 4786 14254 4798 14306
rect 7310 14242 7362 14254
rect 7534 14306 7586 14318
rect 7534 14242 7586 14254
rect 16158 14306 16210 14318
rect 16158 14242 16210 14254
rect 21422 14306 21474 14318
rect 21422 14242 21474 14254
rect 26350 14306 26402 14318
rect 26350 14242 26402 14254
rect 672 14138 27888 14172
rect 672 14086 3806 14138
rect 3858 14086 3910 14138
rect 3962 14086 4014 14138
rect 4066 14086 23806 14138
rect 23858 14086 23910 14138
rect 23962 14086 24014 14138
rect 24066 14086 27888 14138
rect 672 14052 27888 14086
rect 5518 13970 5570 13982
rect 5518 13906 5570 13918
rect 17390 13970 17442 13982
rect 17390 13906 17442 13918
rect 17726 13970 17778 13982
rect 17726 13906 17778 13918
rect 19070 13970 19122 13982
rect 19070 13906 19122 13918
rect 19294 13970 19346 13982
rect 19294 13906 19346 13918
rect 23662 13970 23714 13982
rect 23662 13906 23714 13918
rect 4398 13858 4450 13870
rect 12786 13806 12798 13858
rect 12850 13806 12862 13858
rect 4398 13794 4450 13806
rect 8542 13746 8594 13758
rect 10670 13746 10722 13758
rect 21422 13746 21474 13758
rect 1810 13694 1822 13746
rect 1874 13694 1886 13746
rect 3938 13694 3950 13746
rect 4002 13694 4014 13746
rect 6962 13694 6974 13746
rect 7026 13694 7038 13746
rect 9314 13694 9326 13746
rect 9378 13694 9390 13746
rect 9762 13694 9774 13746
rect 9826 13694 9838 13746
rect 11218 13694 11230 13746
rect 11282 13694 11294 13746
rect 12114 13694 12126 13746
rect 12178 13694 12190 13746
rect 14130 13694 14142 13746
rect 14194 13694 14206 13746
rect 14578 13694 14590 13746
rect 14642 13694 14654 13746
rect 15810 13694 15822 13746
rect 15874 13694 15886 13746
rect 16706 13694 16718 13746
rect 16770 13694 16782 13746
rect 18162 13694 18174 13746
rect 18226 13694 18238 13746
rect 18386 13694 18398 13746
rect 18450 13694 18462 13746
rect 19618 13694 19630 13746
rect 19682 13694 19694 13746
rect 22978 13694 22990 13746
rect 23042 13694 23054 13746
rect 25330 13694 25342 13746
rect 25394 13694 25406 13746
rect 8542 13682 8594 13694
rect 10670 13682 10722 13694
rect 21422 13682 21474 13694
rect 3390 13634 3442 13646
rect 8990 13634 9042 13646
rect 13134 13634 13186 13646
rect 4946 13582 4958 13634
rect 5010 13582 5022 13634
rect 9986 13582 9998 13634
rect 10050 13582 10062 13634
rect 3390 13570 3442 13582
rect 8990 13570 9042 13582
rect 13134 13570 13186 13582
rect 13694 13634 13746 13646
rect 15150 13634 15202 13646
rect 19966 13634 20018 13646
rect 14690 13582 14702 13634
rect 14754 13582 14766 13634
rect 18274 13582 18286 13634
rect 18338 13582 18350 13634
rect 13694 13570 13746 13582
rect 15150 13570 15202 13582
rect 19966 13570 20018 13582
rect 20638 13634 20690 13646
rect 20638 13570 20690 13582
rect 20862 13634 20914 13646
rect 22642 13582 22654 13634
rect 22706 13582 22718 13634
rect 24770 13582 24782 13634
rect 24834 13582 24846 13634
rect 20862 13570 20914 13582
rect 12910 13522 12962 13534
rect 2258 13470 2270 13522
rect 2322 13470 2334 13522
rect 7410 13470 7422 13522
rect 7474 13470 7486 13522
rect 12910 13458 12962 13470
rect 19742 13522 19794 13534
rect 19742 13458 19794 13470
rect 19854 13522 19906 13534
rect 19854 13458 19906 13470
rect 20750 13522 20802 13534
rect 20750 13458 20802 13470
rect 672 13354 27888 13388
rect 672 13302 4466 13354
rect 4518 13302 4570 13354
rect 4622 13302 4674 13354
rect 4726 13302 24466 13354
rect 24518 13302 24570 13354
rect 24622 13302 24674 13354
rect 24726 13302 27888 13354
rect 672 13268 27888 13302
rect 3614 13186 3666 13198
rect 3614 13122 3666 13134
rect 7870 13186 7922 13198
rect 7870 13122 7922 13134
rect 8990 13186 9042 13198
rect 8990 13122 9042 13134
rect 13806 13186 13858 13198
rect 16046 13186 16098 13198
rect 14914 13134 14926 13186
rect 14978 13134 14990 13186
rect 13806 13122 13858 13134
rect 16046 13122 16098 13134
rect 3166 13074 3218 13086
rect 1474 13022 1486 13074
rect 1538 13022 1550 13074
rect 3166 13010 3218 13022
rect 3502 13074 3554 13086
rect 18734 13074 18786 13086
rect 4610 13022 4622 13074
rect 4674 13022 4686 13074
rect 10322 13022 10334 13074
rect 10386 13022 10398 13074
rect 12562 13022 12574 13074
rect 12626 13022 12638 13074
rect 17826 13022 17838 13074
rect 17890 13022 17902 13074
rect 3502 13010 3554 13022
rect 18734 13010 18786 13022
rect 19182 13074 19234 13086
rect 20178 13022 20190 13074
rect 20242 13022 20254 13074
rect 19182 13010 19234 13022
rect 2606 12962 2658 12974
rect 7982 12962 8034 12974
rect 17166 12962 17218 12974
rect 20862 12962 20914 12974
rect 25118 12962 25170 12974
rect 2258 12910 2270 12962
rect 2322 12910 2334 12962
rect 4162 12910 4174 12962
rect 4226 12910 4238 12962
rect 7298 12910 7310 12962
rect 7362 12910 7374 12962
rect 9874 12910 9886 12962
rect 9938 12910 9950 12962
rect 14354 12910 14366 12962
rect 14418 12910 14430 12962
rect 17938 12910 17950 12962
rect 18002 12910 18014 12962
rect 18386 12910 18398 12962
rect 18450 12910 18462 12962
rect 19506 12910 19518 12962
rect 19570 12910 19582 12962
rect 20066 12910 20078 12962
rect 20130 12910 20142 12962
rect 21186 12910 21198 12962
rect 21250 12910 21262 12962
rect 22194 12910 22206 12962
rect 22258 12910 22270 12962
rect 2606 12898 2658 12910
rect 7982 12898 8034 12910
rect 17166 12898 17218 12910
rect 20862 12898 20914 12910
rect 25118 12898 25170 12910
rect 5742 12850 5794 12862
rect 5742 12786 5794 12798
rect 6414 12850 6466 12862
rect 12226 12798 12238 12850
rect 12290 12798 12302 12850
rect 24658 12798 24670 12850
rect 24722 12798 24734 12850
rect 6414 12786 6466 12798
rect 7870 12738 7922 12750
rect 7870 12674 7922 12686
rect 8206 12738 8258 12750
rect 8206 12674 8258 12686
rect 8878 12738 8930 12750
rect 8878 12674 8930 12686
rect 9214 12738 9266 12750
rect 9214 12674 9266 12686
rect 11566 12738 11618 12750
rect 11566 12674 11618 12686
rect 16830 12738 16882 12750
rect 16830 12674 16882 12686
rect 18398 12738 18450 12750
rect 18398 12674 18450 12686
rect 672 12570 27888 12604
rect 672 12518 3806 12570
rect 3858 12518 3910 12570
rect 3962 12518 4014 12570
rect 4066 12518 23806 12570
rect 23858 12518 23910 12570
rect 23962 12518 24014 12570
rect 24066 12518 27888 12570
rect 672 12484 27888 12518
rect 3614 12402 3666 12414
rect 3614 12338 3666 12350
rect 11006 12402 11058 12414
rect 18286 12402 18338 12414
rect 17490 12350 17502 12402
rect 17554 12350 17566 12402
rect 11006 12338 11058 12350
rect 18286 12338 18338 12350
rect 21534 12402 21586 12414
rect 21534 12338 21586 12350
rect 19518 12290 19570 12302
rect 5282 12238 5294 12290
rect 5346 12238 5358 12290
rect 9426 12238 9438 12290
rect 9490 12238 9502 12290
rect 11890 12238 11902 12290
rect 11954 12238 11966 12290
rect 13234 12238 13246 12290
rect 13298 12238 13310 12290
rect 18722 12238 18734 12290
rect 18786 12238 18798 12290
rect 19518 12226 19570 12238
rect 20750 12290 20802 12302
rect 20750 12226 20802 12238
rect 8766 12178 8818 12190
rect 2034 12126 2046 12178
rect 2098 12126 2110 12178
rect 6066 12126 6078 12178
rect 6130 12126 6142 12178
rect 6626 12126 6638 12178
rect 6690 12126 6702 12178
rect 8766 12114 8818 12126
rect 11454 12178 11506 12190
rect 16494 12178 16546 12190
rect 14018 12126 14030 12178
rect 14082 12126 14094 12178
rect 14802 12126 14814 12178
rect 14866 12126 14878 12178
rect 11454 12114 11506 12126
rect 16494 12114 16546 12126
rect 16942 12178 16994 12190
rect 16942 12114 16994 12126
rect 17278 12178 17330 12190
rect 18062 12178 18114 12190
rect 17602 12126 17614 12178
rect 17666 12126 17678 12178
rect 17278 12114 17330 12126
rect 18062 12114 18114 12126
rect 18510 12178 18562 12190
rect 18510 12114 18562 12126
rect 18958 12178 19010 12190
rect 18958 12114 19010 12126
rect 19630 12178 19682 12190
rect 20638 12178 20690 12190
rect 19954 12126 19966 12178
rect 20018 12126 20030 12178
rect 19630 12114 19682 12126
rect 20638 12114 20690 12126
rect 20862 12178 20914 12190
rect 20862 12114 20914 12126
rect 21646 12178 21698 12190
rect 24098 12126 24110 12178
rect 24162 12126 24174 12178
rect 21646 12114 21698 12126
rect 8542 12066 8594 12078
rect 2482 12014 2494 12066
rect 2546 12014 2558 12066
rect 7298 12014 7310 12066
rect 7362 12014 7374 12066
rect 8542 12002 8594 12014
rect 8654 12066 8706 12078
rect 9762 12014 9774 12066
rect 9826 12014 9838 12066
rect 15250 12014 15262 12066
rect 15314 12014 15326 12066
rect 8654 12002 8706 12014
rect 17726 11954 17778 11966
rect 8082 11902 8094 11954
rect 8146 11902 8158 11954
rect 17726 11890 17778 11902
rect 18734 11954 18786 11966
rect 18734 11890 18786 11902
rect 19406 11954 19458 11966
rect 19406 11890 19458 11902
rect 21086 11954 21138 11966
rect 21086 11890 21138 11902
rect 22542 11954 22594 11966
rect 23650 11902 23662 11954
rect 23714 11902 23726 11954
rect 22542 11890 22594 11902
rect 672 11786 27888 11820
rect 672 11734 4466 11786
rect 4518 11734 4570 11786
rect 4622 11734 4674 11786
rect 4726 11734 24466 11786
rect 24518 11734 24570 11786
rect 24622 11734 24674 11786
rect 24726 11734 27888 11786
rect 672 11700 27888 11734
rect 1598 11618 1650 11630
rect 3726 11618 3778 11630
rect 8318 11618 8370 11630
rect 2706 11566 2718 11618
rect 2770 11566 2782 11618
rect 5506 11566 5518 11618
rect 5570 11566 5582 11618
rect 7522 11566 7534 11618
rect 7586 11566 7598 11618
rect 1598 11554 1650 11566
rect 3726 11554 3778 11566
rect 8318 11554 8370 11566
rect 9774 11618 9826 11630
rect 9774 11554 9826 11566
rect 14142 11618 14194 11630
rect 14142 11554 14194 11566
rect 15598 11618 15650 11630
rect 18722 11566 18734 11618
rect 18786 11566 18798 11618
rect 15598 11554 15650 11566
rect 7086 11506 7138 11518
rect 7086 11442 7138 11454
rect 8206 11506 8258 11518
rect 8206 11442 8258 11454
rect 9886 11506 9938 11518
rect 9886 11442 9938 11454
rect 11006 11506 11058 11518
rect 11006 11442 11058 11454
rect 11118 11506 11170 11518
rect 11118 11442 11170 11454
rect 11902 11506 11954 11518
rect 16718 11506 16770 11518
rect 13010 11454 13022 11506
rect 13074 11454 13086 11506
rect 11902 11442 11954 11454
rect 16718 11442 16770 11454
rect 23774 11506 23826 11518
rect 23774 11442 23826 11454
rect 4286 11394 4338 11406
rect 3266 11342 3278 11394
rect 3330 11342 3342 11394
rect 4286 11330 4338 11342
rect 6638 11394 6690 11406
rect 7534 11394 7586 11406
rect 8990 11394 9042 11406
rect 7298 11342 7310 11394
rect 7362 11342 7374 11394
rect 7858 11342 7870 11394
rect 7922 11342 7934 11394
rect 6638 11330 6690 11342
rect 7534 11330 7586 11342
rect 8990 11330 9042 11342
rect 9102 11394 9154 11406
rect 9102 11330 9154 11342
rect 9326 11394 9378 11406
rect 9326 11330 9378 11342
rect 10782 11394 10834 11406
rect 10782 11330 10834 11342
rect 11454 11394 11506 11406
rect 11454 11330 11506 11342
rect 11678 11394 11730 11406
rect 17054 11394 17106 11406
rect 19182 11394 19234 11406
rect 12450 11342 12462 11394
rect 12514 11342 12526 11394
rect 18162 11342 18174 11394
rect 18226 11342 18238 11394
rect 18610 11342 18622 11394
rect 18674 11342 18686 11394
rect 19954 11342 19966 11394
rect 20018 11342 20030 11394
rect 20850 11342 20862 11394
rect 20914 11342 20926 11394
rect 23314 11342 23326 11394
rect 23378 11342 23390 11394
rect 11678 11330 11730 11342
rect 17054 11330 17106 11342
rect 19182 11330 19234 11342
rect 11566 11282 11618 11294
rect 5058 11230 5070 11282
rect 5122 11230 5134 11282
rect 11566 11218 11618 11230
rect 17726 11282 17778 11294
rect 17726 11218 17778 11230
rect 9438 11170 9490 11182
rect 9438 11106 9490 11118
rect 15374 11170 15426 11182
rect 15374 11106 15426 11118
rect 15710 11170 15762 11182
rect 15710 11106 15762 11118
rect 672 11002 27888 11036
rect 672 10950 3806 11002
rect 3858 10950 3910 11002
rect 3962 10950 4014 11002
rect 4066 10950 23806 11002
rect 23858 10950 23910 11002
rect 23962 10950 24014 11002
rect 24066 10950 27888 11002
rect 672 10916 27888 10950
rect 3614 10834 3666 10846
rect 3614 10770 3666 10782
rect 7198 10834 7250 10846
rect 7198 10770 7250 10782
rect 11902 10834 11954 10846
rect 11902 10770 11954 10782
rect 18286 10834 18338 10846
rect 18286 10770 18338 10782
rect 13246 10722 13298 10734
rect 5170 10670 5182 10722
rect 5234 10670 5246 10722
rect 7970 10670 7982 10722
rect 8034 10670 8046 10722
rect 14690 10670 14702 10722
rect 14754 10670 14766 10722
rect 17602 10670 17614 10722
rect 17666 10670 17678 10722
rect 13246 10658 13298 10670
rect 7422 10610 7474 10622
rect 7870 10610 7922 10622
rect 2034 10558 2046 10610
rect 2098 10558 2110 10610
rect 7746 10558 7758 10610
rect 7810 10558 7822 10610
rect 7422 10546 7474 10558
rect 7870 10546 7922 10558
rect 8766 10610 8818 10622
rect 8766 10546 8818 10558
rect 10222 10610 10274 10622
rect 11454 10610 11506 10622
rect 12798 10610 12850 10622
rect 10882 10558 10894 10610
rect 10946 10558 10958 10610
rect 12002 10558 12014 10610
rect 12066 10558 12078 10610
rect 10222 10546 10274 10558
rect 11454 10546 11506 10558
rect 12798 10546 12850 10558
rect 13022 10610 13074 10622
rect 13022 10546 13074 10558
rect 13470 10610 13522 10622
rect 13470 10546 13522 10558
rect 16606 10610 16658 10622
rect 17490 10558 17502 10610
rect 17554 10558 17566 10610
rect 19954 10558 19966 10610
rect 20018 10558 20030 10610
rect 16606 10546 16658 10558
rect 6750 10498 6802 10510
rect 2482 10446 2494 10498
rect 2546 10446 2558 10498
rect 5618 10446 5630 10498
rect 5682 10446 5694 10498
rect 6750 10434 6802 10446
rect 9326 10498 9378 10510
rect 9326 10434 9378 10446
rect 9662 10498 9714 10510
rect 9662 10434 9714 10446
rect 10670 10498 10722 10510
rect 10670 10434 10722 10446
rect 11118 10498 11170 10510
rect 17278 10498 17330 10510
rect 11666 10446 11678 10498
rect 11730 10446 11742 10498
rect 15026 10446 15038 10498
rect 15090 10446 15102 10498
rect 11118 10434 11170 10446
rect 17278 10434 17330 10446
rect 17838 10498 17890 10510
rect 19394 10446 19406 10498
rect 19458 10446 19470 10498
rect 17838 10434 17890 10446
rect 8094 10386 8146 10398
rect 8094 10322 8146 10334
rect 9550 10386 9602 10398
rect 9550 10322 9602 10334
rect 9886 10386 9938 10398
rect 9886 10322 9938 10334
rect 11230 10386 11282 10398
rect 11230 10322 11282 10334
rect 12238 10386 12290 10398
rect 12238 10322 12290 10334
rect 13582 10386 13634 10398
rect 13582 10322 13634 10334
rect 13694 10386 13746 10398
rect 13694 10322 13746 10334
rect 16270 10386 16322 10398
rect 16270 10322 16322 10334
rect 16942 10386 16994 10398
rect 16942 10322 16994 10334
rect 17166 10386 17218 10398
rect 17166 10322 17218 10334
rect 672 10218 27888 10252
rect 672 10166 4466 10218
rect 4518 10166 4570 10218
rect 4622 10166 4674 10218
rect 4726 10166 24466 10218
rect 24518 10166 24570 10218
rect 24622 10166 24674 10218
rect 24726 10166 27888 10218
rect 672 10132 27888 10166
rect 13918 10050 13970 10062
rect 16046 10050 16098 10062
rect 5394 9998 5406 10050
rect 5458 9998 5470 10050
rect 7410 9998 7422 10050
rect 7474 9998 7486 10050
rect 12674 9998 12686 10050
rect 12738 9998 12750 10050
rect 15362 9998 15374 10050
rect 15426 9998 15438 10050
rect 18946 9998 18958 10050
rect 19010 9998 19022 10050
rect 13918 9986 13970 9998
rect 16046 9986 16098 9998
rect 6526 9938 6578 9950
rect 6526 9874 6578 9886
rect 7086 9938 7138 9950
rect 7086 9874 7138 9886
rect 9102 9938 9154 9950
rect 13134 9938 13186 9950
rect 16158 9938 16210 9950
rect 10098 9886 10110 9938
rect 10162 9886 10174 9938
rect 15138 9886 15150 9938
rect 15202 9886 15214 9938
rect 9102 9874 9154 9886
rect 13134 9874 13186 9886
rect 16158 9874 16210 9886
rect 17166 9938 17218 9950
rect 17166 9874 17218 9886
rect 19406 9938 19458 9950
rect 19406 9874 19458 9886
rect 7534 9826 7586 9838
rect 10782 9826 10834 9838
rect 13246 9826 13298 9838
rect 14926 9826 14978 9838
rect 16606 9826 16658 9838
rect 2034 9774 2046 9826
rect 2098 9774 2110 9826
rect 3826 9774 3838 9826
rect 3890 9774 3902 9826
rect 4946 9774 4958 9826
rect 5010 9774 5022 9826
rect 7298 9774 7310 9826
rect 7362 9774 7374 9826
rect 7858 9774 7870 9826
rect 7922 9774 7934 9826
rect 9538 9774 9550 9826
rect 9602 9774 9614 9826
rect 9986 9774 9998 9826
rect 10050 9774 10062 9826
rect 11330 9774 11342 9826
rect 11394 9774 11406 9826
rect 12226 9774 12238 9826
rect 12290 9774 12302 9826
rect 13458 9774 13470 9826
rect 13522 9774 13534 9826
rect 13794 9774 13806 9826
rect 13858 9774 13870 9826
rect 15698 9774 15710 9826
rect 15762 9774 15774 9826
rect 7534 9762 7586 9774
rect 10782 9762 10834 9774
rect 13246 9762 13298 9774
rect 14926 9762 14978 9774
rect 16606 9762 16658 9774
rect 17054 9826 17106 9838
rect 17054 9762 17106 9774
rect 17278 9826 17330 9838
rect 18386 9774 18398 9826
rect 18450 9774 18462 9826
rect 18834 9774 18846 9826
rect 18898 9774 18910 9826
rect 19954 9774 19966 9826
rect 20018 9774 20030 9826
rect 21074 9774 21086 9826
rect 21138 9774 21150 9826
rect 17278 9762 17330 9774
rect 1262 9714 1314 9726
rect 1262 9650 1314 9662
rect 2830 9714 2882 9726
rect 2830 9650 2882 9662
rect 17950 9714 18002 9726
rect 17950 9650 18002 9662
rect 14030 9602 14082 9614
rect 14030 9538 14082 9550
rect 14254 9602 14306 9614
rect 14254 9538 14306 9550
rect 15374 9602 15426 9614
rect 15374 9538 15426 9550
rect 672 9434 27888 9468
rect 672 9382 3806 9434
rect 3858 9382 3910 9434
rect 3962 9382 4014 9434
rect 4066 9382 23806 9434
rect 23858 9382 23910 9434
rect 23962 9382 24014 9434
rect 24066 9382 27888 9434
rect 672 9348 27888 9382
rect 1262 9266 1314 9278
rect 1262 9202 1314 9214
rect 9662 9266 9714 9278
rect 9662 9202 9714 9214
rect 12126 9266 12178 9278
rect 12126 9202 12178 9214
rect 13806 9266 13858 9278
rect 13806 9202 13858 9214
rect 16494 9266 16546 9278
rect 16494 9202 16546 9214
rect 17054 9266 17106 9278
rect 17054 9202 17106 9214
rect 5518 9154 5570 9166
rect 2930 9102 2942 9154
rect 2994 9102 3006 9154
rect 5518 9090 5570 9102
rect 6414 9154 6466 9166
rect 6414 9090 6466 9102
rect 7422 9154 7474 9166
rect 10546 9102 10558 9154
rect 10610 9102 10622 9154
rect 18610 9102 18622 9154
rect 18674 9102 18686 9154
rect 7422 9090 7474 9102
rect 4958 9042 5010 9054
rect 7534 9042 7586 9054
rect 2258 8990 2270 9042
rect 2322 8990 2334 9042
rect 3826 8990 3838 9042
rect 3890 8990 3902 9042
rect 5954 8990 5966 9042
rect 6018 8990 6030 9042
rect 6962 8990 6974 9042
rect 7026 8990 7038 9042
rect 8082 8990 8094 9042
rect 8146 8990 8158 9042
rect 12786 8990 12798 9042
rect 12850 8990 12862 9042
rect 13010 8990 13022 9042
rect 13074 8990 13086 9042
rect 14802 8990 14814 9042
rect 14866 8990 14878 9042
rect 4958 8978 5010 8990
rect 7534 8978 7586 8990
rect 7310 8930 7362 8942
rect 10882 8878 10894 8930
rect 10946 8878 10958 8930
rect 18162 8878 18174 8930
rect 18226 8878 18238 8930
rect 7310 8866 7362 8878
rect 8530 8766 8542 8818
rect 8594 8766 8606 8818
rect 15362 8766 15374 8818
rect 15426 8766 15438 8818
rect 672 8650 27888 8684
rect 672 8598 4466 8650
rect 4518 8598 4570 8650
rect 4622 8598 4674 8650
rect 4726 8598 24466 8650
rect 24518 8598 24570 8650
rect 24622 8598 24674 8650
rect 24726 8598 27888 8650
rect 672 8564 27888 8598
rect 8430 8482 8482 8494
rect 8430 8418 8482 8430
rect 12238 8482 12290 8494
rect 12238 8418 12290 8430
rect 7198 8370 7250 8382
rect 3042 8318 3054 8370
rect 3106 8318 3118 8370
rect 6290 8318 6302 8370
rect 6354 8318 6366 8370
rect 7198 8306 7250 8318
rect 8094 8370 8146 8382
rect 8094 8306 8146 8318
rect 8206 8370 8258 8382
rect 14926 8370 14978 8382
rect 11106 8318 11118 8370
rect 11170 8318 11182 8370
rect 13346 8318 13358 8370
rect 13410 8318 13422 8370
rect 8206 8306 8258 8318
rect 14926 8306 14978 8318
rect 15710 8370 15762 8382
rect 15710 8306 15762 8318
rect 17614 8370 17666 8382
rect 20974 8370 21026 8382
rect 20514 8318 20526 8370
rect 20578 8318 20590 8370
rect 17614 8306 17666 8318
rect 20974 8306 21026 8318
rect 15038 8258 15090 8270
rect 15598 8258 15650 8270
rect 2258 8206 2270 8258
rect 2322 8206 2334 8258
rect 3826 8206 3838 8258
rect 3890 8206 3902 8258
rect 6626 8206 6638 8258
rect 6690 8206 6702 8258
rect 10546 8206 10558 8258
rect 10610 8206 10622 8258
rect 12786 8206 12798 8258
rect 12850 8206 12862 8258
rect 15362 8206 15374 8258
rect 15426 8206 15438 8258
rect 15038 8194 15090 8206
rect 15598 8194 15650 8206
rect 16942 8258 16994 8270
rect 17390 8258 17442 8270
rect 17266 8206 17278 8258
rect 17330 8206 17342 8258
rect 19842 8206 19854 8258
rect 19906 8206 19918 8258
rect 20290 8206 20302 8258
rect 20354 8206 20366 8258
rect 21746 8206 21758 8258
rect 21810 8206 21822 8258
rect 22530 8206 22542 8258
rect 22594 8206 22606 8258
rect 16942 8194 16994 8206
rect 17390 8194 17442 8206
rect 1262 8146 1314 8158
rect 1262 8082 1314 8094
rect 7758 8146 7810 8158
rect 19518 8146 19570 8158
rect 17490 8094 17502 8146
rect 17554 8094 17566 8146
rect 7758 8082 7810 8094
rect 19518 8082 19570 8094
rect 5070 8034 5122 8046
rect 5070 7970 5122 7982
rect 14478 8034 14530 8046
rect 16718 8034 16770 8046
rect 16146 7982 16158 8034
rect 16210 7982 16222 8034
rect 14478 7970 14530 7982
rect 16718 7970 16770 7982
rect 672 7866 27888 7900
rect 672 7814 3806 7866
rect 3858 7814 3910 7866
rect 3962 7814 4014 7866
rect 4066 7814 23806 7866
rect 23858 7814 23910 7866
rect 23962 7814 24014 7866
rect 24066 7814 27888 7866
rect 672 7780 27888 7814
rect 2830 7698 2882 7710
rect 2830 7634 2882 7646
rect 10894 7698 10946 7710
rect 10894 7634 10946 7646
rect 12238 7698 12290 7710
rect 12238 7634 12290 7646
rect 16606 7698 16658 7710
rect 16606 7634 16658 7646
rect 16718 7698 16770 7710
rect 16718 7634 16770 7646
rect 7310 7586 7362 7598
rect 16382 7586 16434 7598
rect 1362 7534 1374 7586
rect 1426 7534 1438 7586
rect 9314 7534 9326 7586
rect 9378 7534 9390 7586
rect 13010 7534 13022 7586
rect 13074 7534 13086 7586
rect 17042 7534 17054 7586
rect 17106 7534 17118 7586
rect 7310 7522 7362 7534
rect 16382 7522 16434 7534
rect 6750 7474 6802 7486
rect 2258 7422 2270 7474
rect 2322 7422 2334 7474
rect 3826 7422 3838 7474
rect 3890 7422 3902 7474
rect 6750 7410 6802 7422
rect 12126 7474 12178 7486
rect 12126 7410 12178 7422
rect 14590 7474 14642 7486
rect 14590 7410 14642 7422
rect 15598 7474 15650 7486
rect 15598 7410 15650 7422
rect 15934 7474 15986 7486
rect 17390 7474 17442 7486
rect 16146 7422 16158 7474
rect 16210 7422 16222 7474
rect 15934 7410 15986 7422
rect 17390 7410 17442 7422
rect 9762 7310 9774 7362
rect 9826 7310 9838 7362
rect 13346 7310 13358 7362
rect 13410 7310 13422 7362
rect 15710 7250 15762 7262
rect 15710 7186 15762 7198
rect 672 7082 27888 7116
rect 672 7030 4466 7082
rect 4518 7030 4570 7082
rect 4622 7030 4674 7082
rect 4726 7030 24466 7082
rect 24518 7030 24570 7082
rect 24622 7030 24674 7082
rect 24726 7030 27888 7082
rect 672 6996 27888 7030
rect 13918 6914 13970 6926
rect 13918 6850 13970 6862
rect 12674 6750 12686 6802
rect 12738 6750 12750 6802
rect 11006 6690 11058 6702
rect 2146 6638 2158 6690
rect 2210 6638 2222 6690
rect 3602 6638 3614 6690
rect 3666 6638 3678 6690
rect 10098 6638 10110 6690
rect 10162 6638 10174 6690
rect 11006 6626 11058 6638
rect 11566 6690 11618 6702
rect 12338 6638 12350 6690
rect 12402 6638 12414 6690
rect 11566 6626 11618 6638
rect 1262 6578 1314 6590
rect 9762 6526 9774 6578
rect 9826 6526 9838 6578
rect 1262 6514 1314 6526
rect 2830 6466 2882 6478
rect 2830 6402 2882 6414
rect 672 6298 27888 6332
rect 672 6246 3806 6298
rect 3858 6246 3910 6298
rect 3962 6246 4014 6298
rect 4066 6246 23806 6298
rect 23858 6246 23910 6298
rect 23962 6246 24014 6298
rect 24066 6246 27888 6298
rect 672 6212 27888 6246
rect 7758 6130 7810 6142
rect 7758 6066 7810 6078
rect 3166 6018 3218 6030
rect 13806 6018 13858 6030
rect 1586 5966 1598 6018
rect 1650 5966 1662 6018
rect 9314 5966 9326 6018
rect 9378 5966 9390 6018
rect 3166 5954 3218 5966
rect 13806 5954 13858 5966
rect 2606 5906 2658 5918
rect 2258 5854 2270 5906
rect 2322 5854 2334 5906
rect 11666 5854 11678 5906
rect 11730 5854 11742 5906
rect 14242 5854 14254 5906
rect 14306 5854 14318 5906
rect 14690 5854 14702 5906
rect 14754 5854 14766 5906
rect 16034 5854 16046 5906
rect 16098 5854 16110 5906
rect 16930 5854 16942 5906
rect 16994 5854 17006 5906
rect 2606 5842 2658 5854
rect 12126 5794 12178 5806
rect 12126 5730 12178 5742
rect 15262 5794 15314 5806
rect 15262 5730 15314 5742
rect 8866 5630 8878 5682
rect 8930 5630 8942 5682
rect 14802 5630 14814 5682
rect 14866 5630 14878 5682
rect 672 5514 27888 5548
rect 672 5462 4466 5514
rect 4518 5462 4570 5514
rect 4622 5462 4674 5514
rect 4726 5462 24466 5514
rect 24518 5462 24570 5514
rect 24622 5462 24674 5514
rect 24726 5462 27888 5514
rect 672 5428 27888 5462
rect 3614 5346 3666 5358
rect 3614 5282 3666 5294
rect 7758 5346 7810 5358
rect 7758 5282 7810 5294
rect 12238 5346 12290 5358
rect 12238 5282 12290 5294
rect 14926 5346 14978 5358
rect 14926 5282 14978 5294
rect 15374 5346 15426 5358
rect 15374 5282 15426 5294
rect 3054 5234 3106 5246
rect 1474 5182 1486 5234
rect 1538 5182 1550 5234
rect 2258 5182 2270 5234
rect 2322 5182 2334 5234
rect 3054 5170 3106 5182
rect 8318 5234 8370 5246
rect 8318 5170 8370 5182
rect 12798 5234 12850 5246
rect 15934 5234 15986 5246
rect 13682 5182 13694 5234
rect 13746 5182 13758 5234
rect 12798 5170 12850 5182
rect 15934 5170 15986 5182
rect 13234 5070 13246 5122
rect 13298 5070 13310 5122
rect 672 4730 27888 4764
rect 672 4678 3806 4730
rect 3858 4678 3910 4730
rect 3962 4678 4014 4730
rect 4066 4678 23806 4730
rect 23858 4678 23910 4730
rect 23962 4678 24014 4730
rect 24066 4678 27888 4730
rect 672 4644 27888 4678
rect 1474 4174 1486 4226
rect 1538 4174 1550 4226
rect 2258 4174 2270 4226
rect 2322 4174 2334 4226
rect 672 3946 27888 3980
rect 672 3894 4466 3946
rect 4518 3894 4570 3946
rect 4622 3894 4674 3946
rect 4726 3894 24466 3946
rect 24518 3894 24570 3946
rect 24622 3894 24674 3946
rect 24726 3894 27888 3946
rect 672 3860 27888 3894
rect 2258 3502 2270 3554
rect 2322 3502 2334 3554
rect 1262 3330 1314 3342
rect 1262 3266 1314 3278
rect 672 3162 27888 3196
rect 672 3110 3806 3162
rect 3858 3110 3910 3162
rect 3962 3110 4014 3162
rect 4066 3110 23806 3162
rect 23858 3110 23910 3162
rect 23962 3110 24014 3162
rect 24066 3110 27888 3162
rect 672 3076 27888 3110
rect 672 2378 27888 2412
rect 672 2326 4466 2378
rect 4518 2326 4570 2378
rect 4622 2326 4674 2378
rect 4726 2326 24466 2378
rect 24518 2326 24570 2378
rect 24622 2326 24674 2378
rect 24726 2326 27888 2378
rect 672 2292 27888 2326
rect 11454 2098 11506 2110
rect 11454 2034 11506 2046
rect 13246 2098 13298 2110
rect 13246 2034 13298 2046
rect 26574 2098 26626 2110
rect 26574 2034 26626 2046
rect 27470 2098 27522 2110
rect 27470 2034 27522 2046
rect 12014 1986 12066 1998
rect 12014 1922 12066 1934
rect 13806 1986 13858 1998
rect 13806 1922 13858 1934
rect 26014 1986 26066 1998
rect 26014 1922 26066 1934
rect 26910 1986 26962 1998
rect 26910 1922 26962 1934
rect 672 1594 27888 1628
rect 672 1542 3806 1594
rect 3858 1542 3910 1594
rect 3962 1542 4014 1594
rect 4066 1542 23806 1594
rect 23858 1542 23910 1594
rect 23962 1542 24014 1594
rect 24066 1542 27888 1594
rect 672 1508 27888 1542
rect 672 810 27888 844
rect 672 758 4466 810
rect 4518 758 4570 810
rect 4622 758 4674 810
rect 4726 758 24466 810
rect 24518 758 24570 810
rect 24622 758 24674 810
rect 24726 758 27888 810
rect 672 724 27888 758
<< via1 >>
rect 3806 56422 3858 56474
rect 3910 56422 3962 56474
rect 4014 56422 4066 56474
rect 23806 56422 23858 56474
rect 23910 56422 23962 56474
rect 24014 56422 24066 56474
rect 3614 56254 3666 56306
rect 5182 56254 5234 56306
rect 8990 56254 9042 56306
rect 10558 56254 10610 56306
rect 13022 56254 13074 56306
rect 14590 56254 14642 56306
rect 16494 56254 16546 56306
rect 18510 56254 18562 56306
rect 20302 56254 20354 56306
rect 22206 56254 22258 56306
rect 24446 56254 24498 56306
rect 26014 56254 26066 56306
rect 7422 56142 7474 56194
rect 7870 56030 7922 56082
rect 21758 56030 21810 56082
rect 1038 55918 1090 55970
rect 3054 55918 3106 55970
rect 6190 55918 6242 55970
rect 9998 55918 10050 55970
rect 11566 55918 11618 55970
rect 14030 55918 14082 55970
rect 15598 55918 15650 55970
rect 17502 55918 17554 55970
rect 19518 55918 19570 55970
rect 21310 55918 21362 55970
rect 23886 55918 23938 55970
rect 25454 55918 25506 55970
rect 1374 55806 1426 55858
rect 4466 55638 4518 55690
rect 4570 55638 4622 55690
rect 4674 55638 4726 55690
rect 24466 55638 24518 55690
rect 24570 55638 24622 55690
rect 24674 55638 24726 55690
rect 22990 55470 23042 55522
rect 21646 55358 21698 55410
rect 3502 55246 3554 55298
rect 6302 55246 6354 55298
rect 12910 55246 12962 55298
rect 18286 55246 18338 55298
rect 20078 55246 20130 55298
rect 20526 55246 20578 55298
rect 20862 55246 20914 55298
rect 22430 55246 22482 55298
rect 24670 55246 24722 55298
rect 26462 55246 26514 55298
rect 2494 55134 2546 55186
rect 6862 55134 6914 55186
rect 11902 55134 11954 55186
rect 17278 55134 17330 55186
rect 25678 55022 25730 55074
rect 27246 55022 27298 55074
rect 3806 54854 3858 54906
rect 3910 54854 3962 54906
rect 4014 54854 4066 54906
rect 23806 54854 23858 54906
rect 23910 54854 23962 54906
rect 24014 54854 24066 54906
rect 22542 54686 22594 54738
rect 23774 54686 23826 54738
rect 19518 54574 19570 54626
rect 25566 54574 25618 54626
rect 21198 54462 21250 54514
rect 24110 54462 24162 54514
rect 21534 54350 21586 54402
rect 24670 54350 24722 54402
rect 26238 54350 26290 54402
rect 27022 54350 27074 54402
rect 19070 54238 19122 54290
rect 20638 54238 20690 54290
rect 4466 54070 4518 54122
rect 4570 54070 4622 54122
rect 4674 54070 4726 54122
rect 24466 54070 24518 54122
rect 24570 54070 24622 54122
rect 24674 54070 24726 54122
rect 21870 53790 21922 53842
rect 22318 53678 22370 53730
rect 22766 53678 22818 53730
rect 24670 53678 24722 53730
rect 26238 53678 26290 53730
rect 23774 53566 23826 53618
rect 25678 53566 25730 53618
rect 27246 53454 27298 53506
rect 3806 53286 3858 53338
rect 3910 53286 3962 53338
rect 4014 53286 4066 53338
rect 23806 53286 23858 53338
rect 23910 53286 23962 53338
rect 24014 53286 24066 53338
rect 24110 53118 24162 53170
rect 27134 53006 27186 53058
rect 23102 52782 23154 52834
rect 24670 52782 24722 52834
rect 25454 52782 25506 52834
rect 26238 52782 26290 52834
rect 4466 52502 4518 52554
rect 4570 52502 4622 52554
rect 4674 52502 4726 52554
rect 24466 52502 24518 52554
rect 24570 52502 24622 52554
rect 24674 52502 24726 52554
rect 21422 52334 21474 52386
rect 21982 52222 22034 52274
rect 24670 52222 24722 52274
rect 22766 52110 22818 52162
rect 26238 52110 26290 52162
rect 23662 51998 23714 52050
rect 25678 51886 25730 51938
rect 27246 51886 27298 51938
rect 3806 51718 3858 51770
rect 3910 51718 3962 51770
rect 4014 51718 4066 51770
rect 23806 51718 23858 51770
rect 23910 51718 23962 51770
rect 24014 51718 24066 51770
rect 25678 51550 25730 51602
rect 26350 51326 26402 51378
rect 24670 51214 24722 51266
rect 27022 51214 27074 51266
rect 4466 50934 4518 50986
rect 4570 50934 4622 50986
rect 4674 50934 4726 50986
rect 24466 50934 24518 50986
rect 24570 50934 24622 50986
rect 24674 50934 24726 50986
rect 23998 50542 24050 50594
rect 24670 50542 24722 50594
rect 26238 50542 26290 50594
rect 23550 50430 23602 50482
rect 25678 50430 25730 50482
rect 27246 50318 27298 50370
rect 3806 50150 3858 50202
rect 3910 50150 3962 50202
rect 4014 50150 4066 50202
rect 23806 50150 23858 50202
rect 23910 50150 23962 50202
rect 24014 50150 24066 50202
rect 25678 49870 25730 49922
rect 27134 49870 27186 49922
rect 26462 49758 26514 49810
rect 24670 49646 24722 49698
rect 4466 49366 4518 49418
rect 4570 49366 4622 49418
rect 4674 49366 4726 49418
rect 24466 49366 24518 49418
rect 24570 49366 24622 49418
rect 24674 49366 24726 49418
rect 24670 48974 24722 49026
rect 26238 48974 26290 49026
rect 25678 48750 25730 48802
rect 27246 48750 27298 48802
rect 3806 48582 3858 48634
rect 3910 48582 3962 48634
rect 4014 48582 4066 48634
rect 23806 48582 23858 48634
rect 23910 48582 23962 48634
rect 24014 48582 24066 48634
rect 26238 48078 26290 48130
rect 27022 48078 27074 48130
rect 4466 47798 4518 47850
rect 4570 47798 4622 47850
rect 4674 47798 4726 47850
rect 24466 47798 24518 47850
rect 24570 47798 24622 47850
rect 24674 47798 24726 47850
rect 24670 47406 24722 47458
rect 26238 47406 26290 47458
rect 25678 47294 25730 47346
rect 27246 47182 27298 47234
rect 3806 47014 3858 47066
rect 3910 47014 3962 47066
rect 4014 47014 4066 47066
rect 23806 47014 23858 47066
rect 23910 47014 23962 47066
rect 24014 47014 24066 47066
rect 25678 46734 25730 46786
rect 27134 46734 27186 46786
rect 24670 46510 24722 46562
rect 26238 46510 26290 46562
rect 4466 46230 4518 46282
rect 4570 46230 4622 46282
rect 4674 46230 4726 46282
rect 24466 46230 24518 46282
rect 24570 46230 24622 46282
rect 24674 46230 24726 46282
rect 24894 45838 24946 45890
rect 26238 45838 26290 45890
rect 25678 45614 25730 45666
rect 27246 45614 27298 45666
rect 3806 45446 3858 45498
rect 3910 45446 3962 45498
rect 4014 45446 4066 45498
rect 23806 45446 23858 45498
rect 23910 45446 23962 45498
rect 24014 45446 24066 45498
rect 26462 45054 26514 45106
rect 27022 44942 27074 44994
rect 4466 44662 4518 44714
rect 4570 44662 4622 44714
rect 4674 44662 4726 44714
rect 24466 44662 24518 44714
rect 24570 44662 24622 44714
rect 24674 44662 24726 44714
rect 24894 44270 24946 44322
rect 26350 44270 26402 44322
rect 25678 44158 25730 44210
rect 27246 44046 27298 44098
rect 3806 43878 3858 43930
rect 3910 43878 3962 43930
rect 4014 43878 4066 43930
rect 23806 43878 23858 43930
rect 23910 43878 23962 43930
rect 24014 43878 24066 43930
rect 25678 43598 25730 43650
rect 27134 43598 27186 43650
rect 24894 43486 24946 43538
rect 26238 43374 26290 43426
rect 4466 43094 4518 43146
rect 4570 43094 4622 43146
rect 4674 43094 4726 43146
rect 24466 43094 24518 43146
rect 24570 43094 24622 43146
rect 24674 43094 24726 43146
rect 24670 42702 24722 42754
rect 26238 42702 26290 42754
rect 25678 42478 25730 42530
rect 27246 42478 27298 42530
rect 3806 42310 3858 42362
rect 3910 42310 3962 42362
rect 4014 42310 4066 42362
rect 23806 42310 23858 42362
rect 23910 42310 23962 42362
rect 24014 42310 24066 42362
rect 14254 42030 14306 42082
rect 14590 41806 14642 41858
rect 26238 41806 26290 41858
rect 27022 41806 27074 41858
rect 15822 41694 15874 41746
rect 4466 41526 4518 41578
rect 4570 41526 4622 41578
rect 4674 41526 4726 41578
rect 24466 41526 24518 41578
rect 24570 41526 24622 41578
rect 24674 41526 24726 41578
rect 14366 41358 14418 41410
rect 10110 41246 10162 41298
rect 11790 41134 11842 41186
rect 13806 41134 13858 41186
rect 24782 41134 24834 41186
rect 26238 41134 26290 41186
rect 10558 41022 10610 41074
rect 12126 41022 12178 41074
rect 25678 41022 25730 41074
rect 8990 40910 9042 40962
rect 15486 40910 15538 40962
rect 27246 40910 27298 40962
rect 3806 40742 3858 40794
rect 3910 40742 3962 40794
rect 4014 40742 4066 40794
rect 23806 40742 23858 40794
rect 23910 40742 23962 40794
rect 24014 40742 24066 40794
rect 12910 40462 12962 40514
rect 14478 40462 14530 40514
rect 25678 40462 25730 40514
rect 27134 40462 27186 40514
rect 6078 40350 6130 40402
rect 6526 40350 6578 40402
rect 6862 40350 6914 40402
rect 8318 40350 8370 40402
rect 9214 40350 9266 40402
rect 10446 40350 10498 40402
rect 24670 40350 24722 40402
rect 26238 40350 26290 40402
rect 7534 40238 7586 40290
rect 10894 40238 10946 40290
rect 7086 40126 7138 40178
rect 12126 40126 12178 40178
rect 13358 40126 13410 40178
rect 14926 40126 14978 40178
rect 16046 40126 16098 40178
rect 4466 39958 4518 40010
rect 4570 39958 4622 40010
rect 4674 39958 4726 40010
rect 24466 39958 24518 40010
rect 24570 39958 24622 40010
rect 24674 39958 24726 40010
rect 6974 39790 7026 39842
rect 3054 39678 3106 39730
rect 7310 39678 7362 39730
rect 2606 39566 2658 39618
rect 3838 39566 3890 39618
rect 7758 39566 7810 39618
rect 8990 39566 9042 39618
rect 14030 39566 14082 39618
rect 24894 39566 24946 39618
rect 26238 39566 26290 39618
rect 3502 39454 3554 39506
rect 6414 39454 6466 39506
rect 9550 39454 9602 39506
rect 10558 39454 10610 39506
rect 25678 39342 25730 39394
rect 27246 39342 27298 39394
rect 3806 39174 3858 39226
rect 3910 39174 3962 39226
rect 4014 39174 4066 39226
rect 23806 39174 23858 39226
rect 23910 39174 23962 39226
rect 24014 39174 24066 39226
rect 6974 39006 7026 39058
rect 1598 38894 1650 38946
rect 5406 38894 5458 38946
rect 7982 38894 8034 38946
rect 12238 38894 12290 38946
rect 16942 38894 16994 38946
rect 2270 38782 2322 38834
rect 8318 38782 8370 38834
rect 8878 38794 8930 38846
rect 9438 38782 9490 38834
rect 10110 38782 10162 38834
rect 11006 38782 11058 38834
rect 11790 38782 11842 38834
rect 12798 38782 12850 38834
rect 13134 38782 13186 38834
rect 13582 38782 13634 38834
rect 14254 38782 14306 38834
rect 14814 38782 14866 38834
rect 15822 38782 15874 38834
rect 1150 38670 1202 38722
rect 2718 38670 2770 38722
rect 5854 38670 5906 38722
rect 8990 38670 9042 38722
rect 13806 38670 13858 38722
rect 26238 38670 26290 38722
rect 27022 38670 27074 38722
rect 3838 38558 3890 38610
rect 16382 38558 16434 38610
rect 4466 38390 4518 38442
rect 4570 38390 4622 38442
rect 4674 38390 4726 38442
rect 24466 38390 24518 38442
rect 24570 38390 24622 38442
rect 24674 38390 24726 38442
rect 4846 38222 4898 38274
rect 5966 38222 6018 38274
rect 8206 38222 8258 38274
rect 1822 38110 1874 38162
rect 6974 38110 7026 38162
rect 15710 38110 15762 38162
rect 6638 37998 6690 38050
rect 14702 37998 14754 38050
rect 15150 37998 15202 38050
rect 24670 37998 24722 38050
rect 26238 37998 26290 38050
rect 1374 37886 1426 37938
rect 4398 37886 4450 37938
rect 9662 37886 9714 37938
rect 25678 37886 25730 37938
rect 2942 37774 2994 37826
rect 27246 37774 27298 37826
rect 3806 37606 3858 37658
rect 3910 37606 3962 37658
rect 4014 37606 4066 37658
rect 23806 37606 23858 37658
rect 23910 37606 23962 37658
rect 24014 37606 24066 37658
rect 8094 37438 8146 37490
rect 2158 37326 2210 37378
rect 6526 37326 6578 37378
rect 12014 37326 12066 37378
rect 27134 37326 27186 37378
rect 1710 37214 1762 37266
rect 2718 37214 2770 37266
rect 8654 37214 8706 37266
rect 13134 37214 13186 37266
rect 15486 37214 15538 37266
rect 15934 37214 15986 37266
rect 16606 37214 16658 37266
rect 17166 37214 17218 37266
rect 18174 37214 18226 37266
rect 6974 37102 7026 37154
rect 9326 37102 9378 37154
rect 13470 37102 13522 37154
rect 15150 37102 15202 37154
rect 24670 37102 24722 37154
rect 25454 37102 25506 37154
rect 26238 37102 26290 37154
rect 3166 36990 3218 37042
rect 4286 36990 4338 37042
rect 14702 36990 14754 37042
rect 16158 36990 16210 37042
rect 4466 36822 4518 36874
rect 4570 36822 4622 36874
rect 4674 36822 4726 36874
rect 24466 36822 24518 36874
rect 24570 36822 24622 36874
rect 24674 36822 24726 36874
rect 6414 36654 6466 36706
rect 10222 36654 10274 36706
rect 10558 36654 10610 36706
rect 16718 36654 16770 36706
rect 4174 36542 4226 36594
rect 17278 36542 17330 36594
rect 18286 36542 18338 36594
rect 19854 36542 19906 36594
rect 24670 36542 24722 36594
rect 2606 36430 2658 36482
rect 4734 36430 4786 36482
rect 7870 36430 7922 36482
rect 10894 36430 10946 36482
rect 17726 36430 17778 36482
rect 20414 36430 20466 36482
rect 26350 36430 26402 36482
rect 2046 36318 2098 36370
rect 6862 36318 6914 36370
rect 7422 36318 7474 36370
rect 13582 36318 13634 36370
rect 3054 36206 3106 36258
rect 5294 36206 5346 36258
rect 19406 36206 19458 36258
rect 25678 36206 25730 36258
rect 27246 36206 27298 36258
rect 3806 36038 3858 36090
rect 3910 36038 3962 36090
rect 4014 36038 4066 36090
rect 23806 36038 23858 36090
rect 23910 36038 23962 36090
rect 24014 36038 24066 36090
rect 2718 35758 2770 35810
rect 4398 35758 4450 35810
rect 5966 35758 6018 35810
rect 6526 35758 6578 35810
rect 12014 35758 12066 35810
rect 5518 35646 5570 35698
rect 8654 35646 8706 35698
rect 13582 35646 13634 35698
rect 2382 35534 2434 35586
rect 9326 35534 9378 35586
rect 14814 35534 14866 35586
rect 26238 35534 26290 35586
rect 27022 35534 27074 35586
rect 1150 35422 1202 35474
rect 2270 35422 2322 35474
rect 3838 35422 3890 35474
rect 6974 35422 7026 35474
rect 8094 35422 8146 35474
rect 4466 35254 4518 35306
rect 4570 35254 4622 35306
rect 4674 35254 4726 35306
rect 24466 35254 24518 35306
rect 24570 35254 24622 35306
rect 24674 35254 24726 35306
rect 3838 35086 3890 35138
rect 4286 34974 4338 35026
rect 7086 34974 7138 35026
rect 14030 34974 14082 35026
rect 17950 34974 18002 35026
rect 18286 34974 18338 35026
rect 19294 34974 19346 35026
rect 2046 34862 2098 34914
rect 3166 34862 3218 34914
rect 3726 34862 3778 34914
rect 4958 34862 5010 34914
rect 5854 34862 5906 34914
rect 6526 34862 6578 34914
rect 9662 34862 9714 34914
rect 10894 34862 10946 34914
rect 17502 34862 17554 34914
rect 18734 34862 18786 34914
rect 19070 34862 19122 34914
rect 19854 34862 19906 34914
rect 20302 34862 20354 34914
rect 21310 34862 21362 34914
rect 24670 34862 24722 34914
rect 26238 34862 26290 34914
rect 2494 34750 2546 34802
rect 2830 34750 2882 34802
rect 9998 34750 10050 34802
rect 25678 34750 25730 34802
rect 8206 34638 8258 34690
rect 27246 34638 27298 34690
rect 3806 34470 3858 34522
rect 3910 34470 3962 34522
rect 4014 34470 4066 34522
rect 23806 34470 23858 34522
rect 23910 34470 23962 34522
rect 24014 34470 24066 34522
rect 18958 34302 19010 34354
rect 25678 34190 25730 34242
rect 27134 34190 27186 34242
rect 1486 34078 1538 34130
rect 1934 34078 1986 34130
rect 2830 34078 2882 34130
rect 3166 34078 3218 34130
rect 4174 34078 4226 34130
rect 5070 34078 5122 34130
rect 8206 34078 8258 34130
rect 9102 34078 9154 34130
rect 9550 34078 9602 34130
rect 10222 34078 10274 34130
rect 10894 34078 10946 34130
rect 11790 34078 11842 34130
rect 12686 34078 12738 34130
rect 17278 34078 17330 34130
rect 19518 34078 19570 34130
rect 1150 33966 1202 34018
rect 2158 33966 2210 34018
rect 8766 33966 8818 34018
rect 9774 33966 9826 34018
rect 13582 33966 13634 34018
rect 20078 33966 20130 34018
rect 24670 33966 24722 34018
rect 26238 33966 26290 34018
rect 5518 33854 5570 33906
rect 6638 33854 6690 33906
rect 7758 33854 7810 33906
rect 16270 33854 16322 33906
rect 17838 33854 17890 33906
rect 4466 33686 4518 33738
rect 4570 33686 4622 33738
rect 4674 33686 4726 33738
rect 24466 33686 24518 33738
rect 24570 33686 24622 33738
rect 24674 33686 24726 33738
rect 3278 33406 3330 33458
rect 7646 33406 7698 33458
rect 10894 33406 10946 33458
rect 18734 33406 18786 33458
rect 2718 33294 2770 33346
rect 3166 33294 3218 33346
rect 3726 33294 3778 33346
rect 4510 33294 4562 33346
rect 5406 33294 5458 33346
rect 8878 33294 8930 33346
rect 12574 33294 12626 33346
rect 18286 33294 18338 33346
rect 24670 33294 24722 33346
rect 26238 33294 26290 33346
rect 2270 33182 2322 33234
rect 8094 33182 8146 33234
rect 9326 33182 9378 33234
rect 10446 33182 10498 33234
rect 13246 33182 13298 33234
rect 15598 33182 15650 33234
rect 6526 33070 6578 33122
rect 12014 33070 12066 33122
rect 19966 33070 20018 33122
rect 25678 33070 25730 33122
rect 27246 33070 27298 33122
rect 3806 32902 3858 32954
rect 3910 32902 3962 32954
rect 4014 32902 4066 32954
rect 23806 32902 23858 32954
rect 23910 32902 23962 32954
rect 24014 32902 24066 32954
rect 2830 32734 2882 32786
rect 5854 32622 5906 32674
rect 15598 32622 15650 32674
rect 19742 32622 19794 32674
rect 20750 32622 20802 32674
rect 22094 32622 22146 32674
rect 1150 32510 1202 32562
rect 3390 32510 3442 32562
rect 5182 32510 5234 32562
rect 7198 32510 7250 32562
rect 9886 32510 9938 32562
rect 14814 32510 14866 32562
rect 19182 32510 19234 32562
rect 26350 32510 26402 32562
rect 1598 32398 1650 32450
rect 3838 32398 3890 32450
rect 7646 32398 7698 32450
rect 10334 32398 10386 32450
rect 27022 32398 27074 32450
rect 8878 32286 8930 32338
rect 11454 32286 11506 32338
rect 21198 32286 21250 32338
rect 21534 32286 21586 32338
rect 4466 32118 4518 32170
rect 4570 32118 4622 32170
rect 4674 32118 4726 32170
rect 24466 32118 24518 32170
rect 24570 32118 24622 32170
rect 24674 32118 24726 32170
rect 12462 31950 12514 32002
rect 21198 31950 21250 32002
rect 2158 31838 2210 31890
rect 3278 31838 3330 31890
rect 6078 31838 6130 31890
rect 9662 31838 9714 31890
rect 11118 31838 11170 31890
rect 12910 31838 12962 31890
rect 18622 31838 18674 31890
rect 1710 31726 1762 31778
rect 5406 31726 5458 31778
rect 5854 31726 5906 31778
rect 6638 31726 6690 31778
rect 7086 31726 7138 31778
rect 8206 31726 8258 31778
rect 10222 31726 10274 31778
rect 11790 31726 11842 31778
rect 12350 31714 12402 31766
rect 13470 31726 13522 31778
rect 14478 31726 14530 31778
rect 16718 31726 16770 31778
rect 18062 31726 18114 31778
rect 20638 31726 20690 31778
rect 20974 31726 21026 31778
rect 21758 31726 21810 31778
rect 22430 31726 22482 31778
rect 23214 31726 23266 31778
rect 24894 31726 24946 31778
rect 26462 31726 26514 31778
rect 5070 31614 5122 31666
rect 10670 31614 10722 31666
rect 11454 31614 11506 31666
rect 17166 31614 17218 31666
rect 20190 31614 20242 31666
rect 25678 31614 25730 31666
rect 19742 31502 19794 31554
rect 27246 31502 27298 31554
rect 3806 31334 3858 31386
rect 3910 31334 3962 31386
rect 4014 31334 4066 31386
rect 23806 31334 23858 31386
rect 23910 31334 23962 31386
rect 24014 31334 24066 31386
rect 4286 31166 4338 31218
rect 5518 31054 5570 31106
rect 6414 31054 6466 31106
rect 2718 30942 2770 30994
rect 5966 30942 6018 30994
rect 6974 30942 7026 30994
rect 9102 30942 9154 30994
rect 9998 30942 10050 30994
rect 10558 30942 10610 30994
rect 11342 30942 11394 30994
rect 11790 30942 11842 30994
rect 13470 30942 13522 30994
rect 15822 30942 15874 30994
rect 16382 30942 16434 30994
rect 17502 30942 17554 30994
rect 18510 30942 18562 30994
rect 20974 30942 21026 30994
rect 21422 30942 21474 30994
rect 22094 30942 22146 30994
rect 22654 30942 22706 30994
rect 22878 30942 22930 30994
rect 23662 30942 23714 30994
rect 24894 30942 24946 30994
rect 26350 30942 26402 30994
rect 7310 30830 7362 30882
rect 11230 30830 11282 30882
rect 12238 30830 12290 30882
rect 13806 30830 13858 30882
rect 15038 30830 15090 30882
rect 15486 30830 15538 30882
rect 16494 30830 16546 30882
rect 16942 30830 16994 30882
rect 20638 30830 20690 30882
rect 21646 30830 21698 30882
rect 25454 30830 25506 30882
rect 27022 30830 27074 30882
rect 3166 30718 3218 30770
rect 4958 30718 5010 30770
rect 8542 30718 8594 30770
rect 4466 30550 4518 30602
rect 4570 30550 4622 30602
rect 4674 30550 4726 30602
rect 24466 30550 24518 30602
rect 24570 30550 24622 30602
rect 24674 30550 24726 30602
rect 4510 30382 4562 30434
rect 20862 30382 20914 30434
rect 10894 30270 10946 30322
rect 13582 30270 13634 30322
rect 17390 30270 17442 30322
rect 19630 30270 19682 30322
rect 21870 30270 21922 30322
rect 2270 30158 2322 30210
rect 2718 30158 2770 30210
rect 3838 30158 3890 30210
rect 4286 30158 4338 30210
rect 4958 30158 5010 30210
rect 5630 30158 5682 30210
rect 6526 30158 6578 30210
rect 7086 30158 7138 30210
rect 8878 30158 8930 30210
rect 9438 30158 9490 30210
rect 10446 30158 10498 30210
rect 12574 30158 12626 30210
rect 12910 30158 12962 30210
rect 13358 30158 13410 30210
rect 14254 30158 14306 30210
rect 14590 30158 14642 30210
rect 15710 30158 15762 30210
rect 23102 30158 23154 30210
rect 26238 30158 26290 30210
rect 1598 30046 1650 30098
rect 3054 30046 3106 30098
rect 3502 30046 3554 30098
rect 17054 30046 17106 30098
rect 19294 30046 19346 30098
rect 21534 30046 21586 30098
rect 27134 30046 27186 30098
rect 7646 29934 7698 29986
rect 12126 29934 12178 29986
rect 18622 29934 18674 29986
rect 3806 29766 3858 29818
rect 3910 29766 3962 29818
rect 4014 29766 4066 29818
rect 23806 29766 23858 29818
rect 23910 29766 23962 29818
rect 24014 29766 24066 29818
rect 4286 29598 4338 29650
rect 7198 29598 7250 29650
rect 10110 29598 10162 29650
rect 1150 29486 1202 29538
rect 2718 29486 2770 29538
rect 8542 29486 8594 29538
rect 11790 29486 11842 29538
rect 14030 29486 14082 29538
rect 27246 29486 27298 29538
rect 1486 29374 1538 29426
rect 5630 29374 5682 29426
rect 13582 29374 13634 29426
rect 14702 29374 14754 29426
rect 15150 29374 15202 29426
rect 16046 29374 16098 29426
rect 16494 29374 16546 29426
rect 17502 29374 17554 29426
rect 18174 29374 18226 29426
rect 26238 29374 26290 29426
rect 6078 29262 6130 29314
rect 14366 29262 14418 29314
rect 18622 29262 18674 29314
rect 3166 29150 3218 29202
rect 8990 29150 9042 29202
rect 12238 29150 12290 29202
rect 15374 29150 15426 29202
rect 19742 29150 19794 29202
rect 4466 28982 4518 29034
rect 4570 28982 4622 29034
rect 4674 28982 4726 29034
rect 24466 28982 24518 29034
rect 24570 28982 24622 29034
rect 24674 28982 24726 29034
rect 3614 28814 3666 28866
rect 9998 28814 10050 28866
rect 12574 28814 12626 28866
rect 15486 28814 15538 28866
rect 2382 28702 2434 28754
rect 4510 28702 4562 28754
rect 11566 28702 11618 28754
rect 17838 28702 17890 28754
rect 20414 28702 20466 28754
rect 5070 28590 5122 28642
rect 7310 28590 7362 28642
rect 11118 28590 11170 28642
rect 11902 28590 11954 28642
rect 12350 28590 12402 28642
rect 13022 28590 13074 28642
rect 13582 28590 13634 28642
rect 14702 28590 14754 28642
rect 16046 28590 16098 28642
rect 19854 28590 19906 28642
rect 20190 28590 20242 28642
rect 21086 28590 21138 28642
rect 21422 28590 21474 28642
rect 22430 28590 22482 28642
rect 26238 28590 26290 28642
rect 2046 28478 2098 28530
rect 9550 28478 9602 28530
rect 17390 28478 17442 28530
rect 19406 28478 19458 28530
rect 27246 28478 27298 28530
rect 4286 28366 4338 28418
rect 8094 28366 8146 28418
rect 18958 28366 19010 28418
rect 3806 28198 3858 28250
rect 3910 28198 3962 28250
rect 4014 28198 4066 28250
rect 23806 28198 23858 28250
rect 23910 28198 23962 28250
rect 24014 28198 24066 28250
rect 7422 28030 7474 28082
rect 9774 28030 9826 28082
rect 12126 28030 12178 28082
rect 27246 28030 27298 28082
rect 8206 27918 8258 27970
rect 13582 27918 13634 27970
rect 18174 27918 18226 27970
rect 21198 27918 21250 27970
rect 25678 27918 25730 27970
rect 2270 27806 2322 27858
rect 6638 27806 6690 27858
rect 10446 27806 10498 27858
rect 13918 27806 13970 27858
rect 14366 27806 14418 27858
rect 15262 27806 15314 27858
rect 15822 27806 15874 27858
rect 16606 27806 16658 27858
rect 20638 27806 20690 27858
rect 2830 27694 2882 27746
rect 5518 27694 5570 27746
rect 6414 27694 6466 27746
rect 8654 27694 8706 27746
rect 10894 27694 10946 27746
rect 18510 27694 18562 27746
rect 24670 27694 24722 27746
rect 26238 27694 26290 27746
rect 3950 27582 4002 27634
rect 4958 27582 5010 27634
rect 14590 27582 14642 27634
rect 19742 27582 19794 27634
rect 4466 27414 4518 27466
rect 4570 27414 4622 27466
rect 4674 27414 4726 27466
rect 24466 27414 24518 27466
rect 24570 27414 24622 27466
rect 24674 27414 24726 27466
rect 1710 27246 1762 27298
rect 4286 27246 4338 27298
rect 10110 27246 10162 27298
rect 12014 27246 12066 27298
rect 13134 27246 13186 27298
rect 14254 27246 14306 27298
rect 15374 27246 15426 27298
rect 8318 27134 8370 27186
rect 17390 27134 17442 27186
rect 18398 27134 18450 27186
rect 27022 27134 27074 27186
rect 1262 27022 1314 27074
rect 3614 27022 3666 27074
rect 4062 27022 4114 27074
rect 4734 27022 4786 27074
rect 5294 27022 5346 27074
rect 6414 27022 6466 27074
rect 7870 27022 7922 27074
rect 10558 27022 10610 27074
rect 11454 27022 11506 27074
rect 13806 27022 13858 27074
rect 17726 27022 17778 27074
rect 18174 27022 18226 27074
rect 18958 27022 19010 27074
rect 19406 27022 19458 27074
rect 20414 27022 20466 27074
rect 24670 27022 24722 27074
rect 26238 27022 26290 27074
rect 3278 26910 3330 26962
rect 25678 26910 25730 26962
rect 2830 26798 2882 26850
rect 8990 26798 9042 26850
rect 3806 26630 3858 26682
rect 3910 26630 3962 26682
rect 4014 26630 4066 26682
rect 23806 26630 23858 26682
rect 23910 26630 23962 26682
rect 24014 26630 24066 26682
rect 3614 26462 3666 26514
rect 19966 26462 20018 26514
rect 27246 26462 27298 26514
rect 17726 26350 17778 26402
rect 2046 26238 2098 26290
rect 6414 26238 6466 26290
rect 9326 26238 9378 26290
rect 9774 26238 9826 26290
rect 10670 26238 10722 26290
rect 11230 26238 11282 26290
rect 12126 26238 12178 26290
rect 13246 26238 13298 26290
rect 15262 26238 15314 26290
rect 18398 26238 18450 26290
rect 20750 26238 20802 26290
rect 2382 26126 2434 26178
rect 5518 26126 5570 26178
rect 6750 26126 6802 26178
rect 8990 26126 9042 26178
rect 13694 26126 13746 26178
rect 15822 26126 15874 26178
rect 18734 26126 18786 26178
rect 26238 26126 26290 26178
rect 4958 26014 5010 26066
rect 7982 26014 8034 26066
rect 9998 26014 10050 26066
rect 14814 26014 14866 26066
rect 17278 26014 17330 26066
rect 21310 26014 21362 26066
rect 22430 26014 22482 26066
rect 4466 25846 4518 25898
rect 4570 25846 4622 25898
rect 4674 25846 4726 25898
rect 24466 25846 24518 25898
rect 24570 25846 24622 25898
rect 24674 25846 24726 25898
rect 3614 25678 3666 25730
rect 7086 25678 7138 25730
rect 9550 25678 9602 25730
rect 10670 25678 10722 25730
rect 18622 25678 18674 25730
rect 21310 25678 21362 25730
rect 11790 25566 11842 25618
rect 14926 25566 14978 25618
rect 17278 25566 17330 25618
rect 19182 25566 19234 25618
rect 20190 25566 20242 25618
rect 22318 25566 22370 25618
rect 2046 25454 2098 25506
rect 2942 25454 2994 25506
rect 3390 25454 3442 25506
rect 4174 25454 4226 25506
rect 4734 25454 4786 25506
rect 5630 25454 5682 25506
rect 6526 25454 6578 25506
rect 9102 25454 9154 25506
rect 11342 25454 11394 25506
rect 14478 25454 14530 25506
rect 16830 25454 16882 25506
rect 21758 25454 21810 25506
rect 24670 25454 24722 25506
rect 26238 25454 26290 25506
rect 1262 25342 1314 25394
rect 2606 25342 2658 25394
rect 19742 25342 19794 25394
rect 27246 25342 27298 25394
rect 8206 25230 8258 25282
rect 12910 25230 12962 25282
rect 16046 25230 16098 25282
rect 25678 25230 25730 25282
rect 3806 25062 3858 25114
rect 3910 25062 3962 25114
rect 4014 25062 4066 25114
rect 23806 25062 23858 25114
rect 23910 25062 23962 25114
rect 24014 25062 24066 25114
rect 5518 24894 5570 24946
rect 3502 24782 3554 24834
rect 18734 24782 18786 24834
rect 20638 24782 20690 24834
rect 25678 24782 25730 24834
rect 27134 24782 27186 24834
rect 1822 24670 1874 24722
rect 4958 24670 5010 24722
rect 7422 24670 7474 24722
rect 7758 24670 7810 24722
rect 8430 24670 8482 24722
rect 9214 24670 9266 24722
rect 9998 24670 10050 24722
rect 10558 24670 10610 24722
rect 11118 24670 11170 24722
rect 14926 24670 14978 24722
rect 15374 24670 15426 24722
rect 16046 24670 16098 24722
rect 16606 24670 16658 24722
rect 17614 24670 17666 24722
rect 21086 24670 21138 24722
rect 21534 24670 21586 24722
rect 22318 24670 22370 24722
rect 22878 24670 22930 24722
rect 23774 24670 23826 24722
rect 24894 24670 24946 24722
rect 2382 24558 2434 24610
rect 6974 24558 7026 24610
rect 7982 24558 8034 24610
rect 13358 24558 13410 24610
rect 14590 24558 14642 24610
rect 15598 24558 15650 24610
rect 21646 24558 21698 24610
rect 26238 24558 26290 24610
rect 12798 24446 12850 24498
rect 18174 24446 18226 24498
rect 4466 24278 4518 24330
rect 4570 24278 4622 24330
rect 4674 24278 4726 24330
rect 24466 24278 24518 24330
rect 24570 24278 24622 24330
rect 24674 24278 24726 24330
rect 6638 24110 6690 24162
rect 12238 24110 12290 24162
rect 17726 24110 17778 24162
rect 22094 24110 22146 24162
rect 3390 23998 3442 24050
rect 10334 23998 10386 24050
rect 16046 23998 16098 24050
rect 16718 23998 16770 24050
rect 20974 23998 21026 24050
rect 23102 23998 23154 24050
rect 24670 23998 24722 24050
rect 2830 23886 2882 23938
rect 3166 23886 3218 23938
rect 4062 23886 4114 23938
rect 4622 23886 4674 23938
rect 5518 23886 5570 23938
rect 10894 23886 10946 23938
rect 11566 23886 11618 23938
rect 12014 23886 12066 23938
rect 12910 23886 12962 23938
rect 13470 23886 13522 23938
rect 14366 23886 14418 23938
rect 15486 23886 15538 23938
rect 17054 23886 17106 23938
rect 17614 23886 17666 23938
rect 18174 23886 18226 23938
rect 18958 23886 19010 23938
rect 19742 23886 19794 23938
rect 20414 23886 20466 23938
rect 22654 23886 22706 23938
rect 26238 23886 26290 23938
rect 2382 23774 2434 23826
rect 6190 23774 6242 23826
rect 11230 23774 11282 23826
rect 27246 23774 27298 23826
rect 7758 23662 7810 23714
rect 25678 23662 25730 23714
rect 3806 23494 3858 23546
rect 3910 23494 3962 23546
rect 4014 23494 4066 23546
rect 23806 23494 23858 23546
rect 23910 23494 23962 23546
rect 24014 23494 24066 23546
rect 3838 23326 3890 23378
rect 16270 23326 16322 23378
rect 27246 23326 27298 23378
rect 1150 23214 1202 23266
rect 2270 23214 2322 23266
rect 6974 23214 7026 23266
rect 9326 23214 9378 23266
rect 13246 23214 13298 23266
rect 1598 23102 1650 23154
rect 10334 23102 10386 23154
rect 14702 23102 14754 23154
rect 19966 23102 20018 23154
rect 2718 22990 2770 23042
rect 5182 22990 5234 23042
rect 6078 22990 6130 23042
rect 8878 22990 8930 23042
rect 15150 22990 15202 23042
rect 19630 22990 19682 23042
rect 26238 22990 26290 23042
rect 5742 22878 5794 22930
rect 7758 22878 7810 22930
rect 10894 22878 10946 22930
rect 12014 22878 12066 22930
rect 13806 22878 13858 22930
rect 19854 22878 19906 22930
rect 20078 22878 20130 22930
rect 4466 22710 4518 22762
rect 4570 22710 4622 22762
rect 4674 22710 4726 22762
rect 24466 22710 24518 22762
rect 24570 22710 24622 22762
rect 24674 22710 24726 22762
rect 2830 22542 2882 22594
rect 13358 22542 13410 22594
rect 1598 22430 1650 22482
rect 6078 22430 6130 22482
rect 9998 22430 10050 22482
rect 12238 22430 12290 22482
rect 14814 22430 14866 22482
rect 18062 22430 18114 22482
rect 20302 22430 20354 22482
rect 23438 22430 23490 22482
rect 26238 22430 26290 22482
rect 1262 22318 1314 22370
rect 4286 22318 4338 22370
rect 5630 22318 5682 22370
rect 9550 22318 9602 22370
rect 11790 22318 11842 22370
rect 18398 22318 18450 22370
rect 19630 22318 19682 22370
rect 20078 22318 20130 22370
rect 20750 22318 20802 22370
rect 21310 22318 21362 22370
rect 21534 22318 21586 22370
rect 22318 22318 22370 22370
rect 22878 22318 22930 22370
rect 24894 22318 24946 22370
rect 3502 22206 3554 22258
rect 14478 22206 14530 22258
rect 19294 22206 19346 22258
rect 27246 22206 27298 22258
rect 7198 22094 7250 22146
rect 11118 22094 11170 22146
rect 16046 22094 16098 22146
rect 16830 22094 16882 22146
rect 25678 22094 25730 22146
rect 3806 21926 3858 21978
rect 3910 21926 3962 21978
rect 4014 21926 4066 21978
rect 23806 21926 23858 21978
rect 23910 21926 23962 21978
rect 24014 21926 24066 21978
rect 22094 21758 22146 21810
rect 18174 21646 18226 21698
rect 18510 21646 18562 21698
rect 23886 21646 23938 21698
rect 25790 21646 25842 21698
rect 27134 21646 27186 21698
rect 2606 21534 2658 21586
rect 5406 21534 5458 21586
rect 6526 21534 6578 21586
rect 7086 21534 7138 21586
rect 7758 21534 7810 21586
rect 8094 21534 8146 21586
rect 10558 21534 10610 21586
rect 12126 21534 12178 21586
rect 14814 21534 14866 21586
rect 15262 21534 15314 21586
rect 16158 21534 16210 21586
rect 16494 21534 16546 21586
rect 17614 21534 17666 21586
rect 19070 21534 19122 21586
rect 19294 21534 19346 21586
rect 19630 21534 19682 21586
rect 20638 21534 20690 21586
rect 20862 21534 20914 21586
rect 21086 21534 21138 21586
rect 21982 21534 22034 21586
rect 22206 21534 22258 21586
rect 23550 21534 23602 21586
rect 3166 21422 3218 21474
rect 7534 21422 7586 21474
rect 8542 21422 8594 21474
rect 14030 21422 14082 21474
rect 14478 21422 14530 21474
rect 15486 21422 15538 21474
rect 18846 21422 18898 21474
rect 20078 21422 20130 21474
rect 26238 21422 26290 21474
rect 4286 21310 4338 21362
rect 11006 21310 11058 21362
rect 13470 21310 13522 21362
rect 18286 21310 18338 21362
rect 19630 21310 19682 21362
rect 19966 21310 20018 21362
rect 25342 21310 25394 21362
rect 4466 21142 4518 21194
rect 4570 21142 4622 21194
rect 4674 21142 4726 21194
rect 24466 21142 24518 21194
rect 24570 21142 24622 21194
rect 24674 21142 24726 21194
rect 6974 20974 7026 21026
rect 11342 20974 11394 21026
rect 17950 20974 18002 21026
rect 19742 20974 19794 21026
rect 1262 20862 1314 20914
rect 1822 20862 1874 20914
rect 3166 20862 3218 20914
rect 10334 20862 10386 20914
rect 14814 20862 14866 20914
rect 16942 20862 16994 20914
rect 17278 20862 17330 20914
rect 26462 20862 26514 20914
rect 27358 20862 27410 20914
rect 2606 20750 2658 20802
rect 2942 20750 2994 20802
rect 3614 20750 3666 20802
rect 4398 20750 4450 20802
rect 5182 20750 5234 20802
rect 8878 20750 8930 20802
rect 10782 20750 10834 20802
rect 11118 20750 11170 20802
rect 12014 20750 12066 20802
rect 12350 20750 12402 20802
rect 13358 20750 13410 20802
rect 14478 20750 14530 20802
rect 16046 20750 16098 20802
rect 16830 20750 16882 20802
rect 17166 20750 17218 20802
rect 19070 20750 19122 20802
rect 19518 20750 19570 20802
rect 20190 20750 20242 20802
rect 20750 20750 20802 20802
rect 21758 20750 21810 20802
rect 25902 20750 25954 20802
rect 26910 20750 26962 20802
rect 2158 20638 2210 20690
rect 7422 20638 7474 20690
rect 9438 20638 9490 20690
rect 18734 20638 18786 20690
rect 5854 20526 5906 20578
rect 17614 20526 17666 20578
rect 3806 20358 3858 20410
rect 3910 20358 3962 20410
rect 4014 20358 4066 20410
rect 23806 20358 23858 20410
rect 23910 20358 23962 20410
rect 24014 20358 24066 20410
rect 5518 20190 5570 20242
rect 3278 20078 3330 20130
rect 11230 20078 11282 20130
rect 20638 20078 20690 20130
rect 20974 20078 21026 20130
rect 1710 19966 1762 20018
rect 5182 19966 5234 20018
rect 7310 19966 7362 20018
rect 7870 19966 7922 20018
rect 8430 19966 8482 20018
rect 9214 19966 9266 20018
rect 9998 19966 10050 20018
rect 10558 19966 10610 20018
rect 13134 19966 13186 20018
rect 13582 19966 13634 20018
rect 14478 19966 14530 20018
rect 14814 19966 14866 20018
rect 15822 19966 15874 20018
rect 16494 19966 16546 20018
rect 19742 19966 19794 20018
rect 19966 19966 20018 20018
rect 6974 19854 7026 19906
rect 7982 19854 8034 19906
rect 12798 19854 12850 19906
rect 13806 19854 13858 19906
rect 17054 19854 17106 19906
rect 18622 19854 18674 19906
rect 20078 19854 20130 19906
rect 2158 19742 2210 19794
rect 11118 19742 11170 19794
rect 18174 19742 18226 19794
rect 18734 19742 18786 19794
rect 18846 19742 18898 19794
rect 20862 19742 20914 19794
rect 4466 19574 4518 19626
rect 4570 19574 4622 19626
rect 4674 19574 4726 19626
rect 24466 19574 24518 19626
rect 24570 19574 24622 19626
rect 24674 19574 24726 19626
rect 9326 19406 9378 19458
rect 10894 19406 10946 19458
rect 13470 19406 13522 19458
rect 17390 19406 17442 19458
rect 20302 19406 20354 19458
rect 25902 19406 25954 19458
rect 2270 19294 2322 19346
rect 3502 19294 3554 19346
rect 6078 19294 6130 19346
rect 6526 19294 6578 19346
rect 9886 19294 9938 19346
rect 12014 19294 12066 19346
rect 26462 19294 26514 19346
rect 4622 19182 4674 19234
rect 5406 19182 5458 19234
rect 5854 19182 5906 19234
rect 7086 19182 7138 19234
rect 7310 19182 7362 19234
rect 8206 19182 8258 19234
rect 10334 19182 10386 19234
rect 12798 19182 12850 19234
rect 13246 19182 13298 19234
rect 13918 19182 13970 19234
rect 14478 19182 14530 19234
rect 15486 19182 15538 19234
rect 16046 19182 16098 19234
rect 16942 19182 16994 19234
rect 17278 19182 17330 19234
rect 17390 19182 17442 19234
rect 17726 19182 17778 19234
rect 18286 19182 18338 19234
rect 19294 19182 19346 19234
rect 19630 19182 19682 19234
rect 20414 19182 20466 19234
rect 20862 19182 20914 19234
rect 1374 19070 1426 19122
rect 3054 19070 3106 19122
rect 5070 19070 5122 19122
rect 12462 19070 12514 19122
rect 16158 19070 16210 19122
rect 21310 19070 21362 19122
rect 3806 18790 3858 18842
rect 3910 18790 3962 18842
rect 4014 18790 4066 18842
rect 23806 18790 23858 18842
rect 23910 18790 23962 18842
rect 24014 18790 24066 18842
rect 12126 18622 12178 18674
rect 14590 18622 14642 18674
rect 2718 18510 2770 18562
rect 5070 18510 5122 18562
rect 6078 18510 6130 18562
rect 10558 18510 10610 18562
rect 13022 18510 13074 18562
rect 1710 18398 1762 18450
rect 2158 18398 2210 18450
rect 5518 18398 5570 18450
rect 7646 18398 7698 18450
rect 8318 18398 8370 18450
rect 15710 18398 15762 18450
rect 16718 18398 16770 18450
rect 17950 18398 18002 18450
rect 18510 18398 18562 18450
rect 19070 18398 19122 18450
rect 20974 18398 21026 18450
rect 21422 18398 21474 18450
rect 22654 18398 22706 18450
rect 23662 18398 23714 18450
rect 6526 18286 6578 18338
rect 8766 18286 8818 18338
rect 11006 18286 11058 18338
rect 13358 18286 13410 18338
rect 17390 18286 17442 18338
rect 17838 18286 17890 18338
rect 18846 18286 18898 18338
rect 20638 18286 20690 18338
rect 22094 18286 22146 18338
rect 3166 18174 3218 18226
rect 4286 18174 4338 18226
rect 9886 18174 9938 18226
rect 19518 18174 19570 18226
rect 19630 18174 19682 18226
rect 19742 18174 19794 18226
rect 21646 18174 21698 18226
rect 4466 18006 4518 18058
rect 4570 18006 4622 18058
rect 4674 18006 4726 18058
rect 24466 18006 24518 18058
rect 24570 18006 24622 18058
rect 24674 18006 24726 18058
rect 3726 17838 3778 17890
rect 12686 17838 12738 17890
rect 13806 17838 13858 17890
rect 16830 17838 16882 17890
rect 6078 17726 6130 17778
rect 6526 17726 6578 17778
rect 8878 17726 8930 17778
rect 9438 17726 9490 17778
rect 10446 17726 10498 17778
rect 15150 17726 15202 17778
rect 17502 17726 17554 17778
rect 17838 17726 17890 17778
rect 18846 17726 18898 17778
rect 22654 17726 22706 17778
rect 24558 17726 24610 17778
rect 1822 17619 1874 17671
rect 2718 17614 2770 17666
rect 3278 17614 3330 17666
rect 3838 17614 3890 17666
rect 4286 17614 4338 17666
rect 4734 17614 4786 17666
rect 5406 17614 5458 17666
rect 5966 17614 6018 17666
rect 7310 17614 7362 17666
rect 8206 17614 8258 17666
rect 12126 17614 12178 17666
rect 15710 17614 15762 17666
rect 16718 17614 16770 17666
rect 17166 17614 17218 17666
rect 18174 17614 18226 17666
rect 18622 17614 18674 17666
rect 19294 17614 19346 17666
rect 19854 17614 19906 17666
rect 20078 17614 20130 17666
rect 20974 17614 21026 17666
rect 21534 17614 21586 17666
rect 25006 17614 25058 17666
rect 5070 17502 5122 17554
rect 9998 17502 10050 17554
rect 17390 17502 17442 17554
rect 23102 17502 23154 17554
rect 11566 17390 11618 17442
rect 3806 17222 3858 17274
rect 3910 17222 3962 17274
rect 4014 17222 4066 17274
rect 23806 17222 23858 17274
rect 23910 17222 23962 17274
rect 24014 17222 24066 17274
rect 2830 17054 2882 17106
rect 5518 17054 5570 17106
rect 18286 17054 18338 17106
rect 18510 17054 18562 17106
rect 19966 17054 20018 17106
rect 20974 17054 21026 17106
rect 1262 16942 1314 16994
rect 3726 16942 3778 16994
rect 19070 16942 19122 16994
rect 19630 16942 19682 16994
rect 3390 16830 3442 16882
rect 4958 16830 5010 16882
rect 8430 16830 8482 16882
rect 9326 16830 9378 16882
rect 9774 16830 9826 16882
rect 10446 16830 10498 16882
rect 11006 16830 11058 16882
rect 12014 16830 12066 16882
rect 15038 16830 15090 16882
rect 15486 16830 15538 16882
rect 16158 16830 16210 16882
rect 16942 16830 16994 16882
rect 17614 16825 17666 16877
rect 18734 16830 18786 16882
rect 19182 16830 19234 16882
rect 23774 16830 23826 16882
rect 1598 16718 1650 16770
rect 7982 16718 8034 16770
rect 8990 16718 9042 16770
rect 14702 16718 14754 16770
rect 15710 16718 15762 16770
rect 23326 16718 23378 16770
rect 6862 16606 6914 16658
rect 9998 16606 10050 16658
rect 18958 16606 19010 16658
rect 19742 16606 19794 16658
rect 20750 16606 20802 16658
rect 20862 16606 20914 16658
rect 22206 16606 22258 16658
rect 4466 16438 4518 16490
rect 4570 16438 4622 16490
rect 4674 16438 4726 16490
rect 24466 16438 24518 16490
rect 24570 16438 24622 16490
rect 24674 16438 24726 16490
rect 1822 16270 1874 16322
rect 2942 16270 2994 16322
rect 5182 16270 5234 16322
rect 7086 16270 7138 16322
rect 8206 16270 8258 16322
rect 9102 16270 9154 16322
rect 11678 16270 11730 16322
rect 12798 16270 12850 16322
rect 17054 16270 17106 16322
rect 18286 16270 18338 16322
rect 19966 16270 20018 16322
rect 4062 16158 4114 16210
rect 5966 16158 6018 16210
rect 10446 16158 10498 16210
rect 13806 16158 13858 16210
rect 16046 16158 16098 16210
rect 18958 16158 19010 16210
rect 20414 16158 20466 16210
rect 1374 16046 1426 16098
rect 3614 16046 3666 16098
rect 5854 16046 5906 16098
rect 6190 16046 6242 16098
rect 9998 16046 10050 16098
rect 11118 16046 11170 16098
rect 13470 16046 13522 16098
rect 15598 16046 15650 16098
rect 16718 16046 16770 16098
rect 16942 16046 16994 16098
rect 17502 16046 17554 16098
rect 17838 16046 17890 16098
rect 18062 16046 18114 16098
rect 18286 16046 18338 16098
rect 18622 16046 18674 16098
rect 19406 16046 19458 16098
rect 19742 16046 19794 16098
rect 21198 16046 21250 16098
rect 21982 16046 22034 16098
rect 6638 15934 6690 15986
rect 9102 15934 9154 15986
rect 8878 15822 8930 15874
rect 15038 15822 15090 15874
rect 17278 15822 17330 15874
rect 3806 15654 3858 15706
rect 3910 15654 3962 15706
rect 4014 15654 4066 15706
rect 23806 15654 23858 15706
rect 23910 15654 23962 15706
rect 24014 15654 24066 15706
rect 9886 15486 9938 15538
rect 12126 15486 12178 15538
rect 18622 15486 18674 15538
rect 2158 15374 2210 15426
rect 5182 15374 5234 15426
rect 10558 15374 10610 15426
rect 19742 15374 19794 15426
rect 20638 15374 20690 15426
rect 1710 15262 1762 15314
rect 4286 15262 4338 15314
rect 6750 15262 6802 15314
rect 7086 15262 7138 15314
rect 7534 15262 7586 15314
rect 7758 15262 7810 15314
rect 8206 15262 8258 15314
rect 14366 15262 14418 15314
rect 15150 15262 15202 15314
rect 15486 15262 15538 15314
rect 16158 15262 16210 15314
rect 16830 15262 16882 15314
rect 17726 15262 17778 15314
rect 18510 15262 18562 15314
rect 18846 15262 18898 15314
rect 19182 15262 19234 15314
rect 20974 15262 21026 15314
rect 21422 15262 21474 15314
rect 22878 15262 22930 15314
rect 23662 15262 23714 15314
rect 2606 15150 2658 15202
rect 3838 15150 3890 15202
rect 5630 15150 5682 15202
rect 8766 15150 8818 15202
rect 11006 15150 11058 15202
rect 14702 15150 14754 15202
rect 15710 15150 15762 15202
rect 20078 15150 20130 15202
rect 21646 15150 21698 15202
rect 22094 15150 22146 15202
rect 7646 15038 7698 15090
rect 14030 15038 14082 15090
rect 18398 15038 18450 15090
rect 19854 15038 19906 15090
rect 4466 14870 4518 14922
rect 4570 14870 4622 14922
rect 4674 14870 4726 14922
rect 24466 14870 24518 14922
rect 24570 14870 24622 14922
rect 24674 14870 24726 14922
rect 3278 14702 3330 14754
rect 5742 14702 5794 14754
rect 9102 14702 9154 14754
rect 12462 14702 12514 14754
rect 13582 14702 13634 14754
rect 16830 14702 16882 14754
rect 22542 14702 22594 14754
rect 2158 14590 2210 14642
rect 4286 14590 4338 14642
rect 6862 14590 6914 14642
rect 8878 14590 8930 14642
rect 9326 14590 9378 14642
rect 10334 14590 10386 14642
rect 11342 14590 11394 14642
rect 14702 14590 14754 14642
rect 15710 14590 15762 14642
rect 16942 14590 16994 14642
rect 17726 14590 17778 14642
rect 18734 14590 18786 14642
rect 19182 14590 19234 14642
rect 25230 14590 25282 14642
rect 1598 14478 1650 14530
rect 3950 14478 4002 14530
rect 4174 14478 4226 14530
rect 5182 14478 5234 14530
rect 7870 14478 7922 14530
rect 7982 14478 8034 14530
rect 8206 14478 8258 14530
rect 8766 14478 8818 14530
rect 9886 14478 9938 14530
rect 15150 14478 15202 14530
rect 16046 14478 16098 14530
rect 16718 14478 16770 14530
rect 18062 14478 18114 14530
rect 18510 14478 18562 14530
rect 19966 14478 20018 14530
rect 20750 14478 20802 14530
rect 8094 14366 8146 14418
rect 10894 14366 10946 14418
rect 13134 14366 13186 14418
rect 22990 14366 23042 14418
rect 24782 14366 24834 14418
rect 4734 14254 4786 14306
rect 7310 14254 7362 14306
rect 7534 14254 7586 14306
rect 16158 14254 16210 14306
rect 21422 14254 21474 14306
rect 26350 14254 26402 14306
rect 3806 14086 3858 14138
rect 3910 14086 3962 14138
rect 4014 14086 4066 14138
rect 23806 14086 23858 14138
rect 23910 14086 23962 14138
rect 24014 14086 24066 14138
rect 5518 13918 5570 13970
rect 17390 13918 17442 13970
rect 17726 13918 17778 13970
rect 19070 13918 19122 13970
rect 19294 13918 19346 13970
rect 23662 13918 23714 13970
rect 4398 13806 4450 13858
rect 12798 13806 12850 13858
rect 1822 13694 1874 13746
rect 3950 13694 4002 13746
rect 6974 13694 7026 13746
rect 8542 13694 8594 13746
rect 9326 13694 9378 13746
rect 9774 13694 9826 13746
rect 10670 13694 10722 13746
rect 11230 13694 11282 13746
rect 12126 13694 12178 13746
rect 14142 13694 14194 13746
rect 14590 13694 14642 13746
rect 15822 13694 15874 13746
rect 16718 13694 16770 13746
rect 18174 13694 18226 13746
rect 18398 13694 18450 13746
rect 19630 13694 19682 13746
rect 21422 13694 21474 13746
rect 22990 13694 23042 13746
rect 25342 13694 25394 13746
rect 3390 13582 3442 13634
rect 4958 13582 5010 13634
rect 8990 13582 9042 13634
rect 9998 13582 10050 13634
rect 13134 13582 13186 13634
rect 13694 13582 13746 13634
rect 14702 13582 14754 13634
rect 15150 13582 15202 13634
rect 18286 13582 18338 13634
rect 19966 13582 20018 13634
rect 20638 13582 20690 13634
rect 20862 13582 20914 13634
rect 22654 13582 22706 13634
rect 24782 13582 24834 13634
rect 2270 13470 2322 13522
rect 7422 13470 7474 13522
rect 12910 13470 12962 13522
rect 19742 13470 19794 13522
rect 19854 13470 19906 13522
rect 20750 13470 20802 13522
rect 4466 13302 4518 13354
rect 4570 13302 4622 13354
rect 4674 13302 4726 13354
rect 24466 13302 24518 13354
rect 24570 13302 24622 13354
rect 24674 13302 24726 13354
rect 3614 13134 3666 13186
rect 7870 13134 7922 13186
rect 8990 13134 9042 13186
rect 13806 13134 13858 13186
rect 14926 13134 14978 13186
rect 16046 13134 16098 13186
rect 1486 13022 1538 13074
rect 3166 13022 3218 13074
rect 3502 13022 3554 13074
rect 4622 13022 4674 13074
rect 10334 13022 10386 13074
rect 12574 13022 12626 13074
rect 17838 13022 17890 13074
rect 18734 13022 18786 13074
rect 19182 13022 19234 13074
rect 20190 13022 20242 13074
rect 2270 12910 2322 12962
rect 2606 12910 2658 12962
rect 4174 12910 4226 12962
rect 7310 12910 7362 12962
rect 7982 12910 8034 12962
rect 9886 12910 9938 12962
rect 14366 12910 14418 12962
rect 17166 12910 17218 12962
rect 17950 12910 18002 12962
rect 18398 12910 18450 12962
rect 19518 12910 19570 12962
rect 20078 12910 20130 12962
rect 20862 12910 20914 12962
rect 21198 12910 21250 12962
rect 22206 12910 22258 12962
rect 25118 12910 25170 12962
rect 5742 12798 5794 12850
rect 6414 12798 6466 12850
rect 12238 12798 12290 12850
rect 24670 12798 24722 12850
rect 7870 12686 7922 12738
rect 8206 12686 8258 12738
rect 8878 12686 8930 12738
rect 9214 12686 9266 12738
rect 11566 12686 11618 12738
rect 16830 12686 16882 12738
rect 18398 12686 18450 12738
rect 3806 12518 3858 12570
rect 3910 12518 3962 12570
rect 4014 12518 4066 12570
rect 23806 12518 23858 12570
rect 23910 12518 23962 12570
rect 24014 12518 24066 12570
rect 3614 12350 3666 12402
rect 11006 12350 11058 12402
rect 17502 12350 17554 12402
rect 18286 12350 18338 12402
rect 21534 12350 21586 12402
rect 5294 12238 5346 12290
rect 9438 12238 9490 12290
rect 11902 12238 11954 12290
rect 13246 12238 13298 12290
rect 18734 12238 18786 12290
rect 19518 12238 19570 12290
rect 20750 12238 20802 12290
rect 2046 12126 2098 12178
rect 6078 12126 6130 12178
rect 6638 12126 6690 12178
rect 8766 12126 8818 12178
rect 11454 12126 11506 12178
rect 14030 12126 14082 12178
rect 14814 12126 14866 12178
rect 16494 12126 16546 12178
rect 16942 12126 16994 12178
rect 17278 12126 17330 12178
rect 17614 12126 17666 12178
rect 18062 12126 18114 12178
rect 18510 12126 18562 12178
rect 18958 12126 19010 12178
rect 19630 12126 19682 12178
rect 19966 12126 20018 12178
rect 20638 12126 20690 12178
rect 20862 12126 20914 12178
rect 21646 12126 21698 12178
rect 24110 12126 24162 12178
rect 2494 12014 2546 12066
rect 7310 12014 7362 12066
rect 8542 12014 8594 12066
rect 8654 12014 8706 12066
rect 9774 12014 9826 12066
rect 15262 12014 15314 12066
rect 8094 11902 8146 11954
rect 17726 11902 17778 11954
rect 18734 11902 18786 11954
rect 19406 11902 19458 11954
rect 21086 11902 21138 11954
rect 22542 11902 22594 11954
rect 23662 11902 23714 11954
rect 4466 11734 4518 11786
rect 4570 11734 4622 11786
rect 4674 11734 4726 11786
rect 24466 11734 24518 11786
rect 24570 11734 24622 11786
rect 24674 11734 24726 11786
rect 1598 11566 1650 11618
rect 2718 11566 2770 11618
rect 3726 11566 3778 11618
rect 5518 11566 5570 11618
rect 7534 11566 7586 11618
rect 8318 11566 8370 11618
rect 9774 11566 9826 11618
rect 14142 11566 14194 11618
rect 15598 11566 15650 11618
rect 18734 11566 18786 11618
rect 7086 11454 7138 11506
rect 8206 11454 8258 11506
rect 9886 11454 9938 11506
rect 11006 11454 11058 11506
rect 11118 11454 11170 11506
rect 11902 11454 11954 11506
rect 13022 11454 13074 11506
rect 16718 11454 16770 11506
rect 23774 11454 23826 11506
rect 3278 11342 3330 11394
rect 4286 11342 4338 11394
rect 6638 11342 6690 11394
rect 7310 11342 7362 11394
rect 7534 11342 7586 11394
rect 7870 11342 7922 11394
rect 8990 11342 9042 11394
rect 9102 11342 9154 11394
rect 9326 11342 9378 11394
rect 10782 11342 10834 11394
rect 11454 11342 11506 11394
rect 11678 11342 11730 11394
rect 12462 11342 12514 11394
rect 17054 11342 17106 11394
rect 18174 11342 18226 11394
rect 18622 11342 18674 11394
rect 19182 11342 19234 11394
rect 19966 11342 20018 11394
rect 20862 11342 20914 11394
rect 23326 11342 23378 11394
rect 5070 11230 5122 11282
rect 11566 11230 11618 11282
rect 17726 11230 17778 11282
rect 9438 11118 9490 11170
rect 15374 11118 15426 11170
rect 15710 11118 15762 11170
rect 3806 10950 3858 11002
rect 3910 10950 3962 11002
rect 4014 10950 4066 11002
rect 23806 10950 23858 11002
rect 23910 10950 23962 11002
rect 24014 10950 24066 11002
rect 3614 10782 3666 10834
rect 7198 10782 7250 10834
rect 11902 10782 11954 10834
rect 18286 10782 18338 10834
rect 5182 10670 5234 10722
rect 7982 10670 8034 10722
rect 13246 10670 13298 10722
rect 14702 10670 14754 10722
rect 17614 10670 17666 10722
rect 2046 10558 2098 10610
rect 7422 10558 7474 10610
rect 7758 10558 7810 10610
rect 7870 10558 7922 10610
rect 8766 10558 8818 10610
rect 10222 10558 10274 10610
rect 10894 10558 10946 10610
rect 11454 10558 11506 10610
rect 12014 10558 12066 10610
rect 12798 10558 12850 10610
rect 13022 10558 13074 10610
rect 13470 10558 13522 10610
rect 16606 10558 16658 10610
rect 17502 10558 17554 10610
rect 19966 10558 20018 10610
rect 2494 10446 2546 10498
rect 5630 10446 5682 10498
rect 6750 10446 6802 10498
rect 9326 10446 9378 10498
rect 9662 10446 9714 10498
rect 10670 10446 10722 10498
rect 11118 10446 11170 10498
rect 11678 10446 11730 10498
rect 15038 10446 15090 10498
rect 17278 10446 17330 10498
rect 17838 10446 17890 10498
rect 19406 10446 19458 10498
rect 8094 10334 8146 10386
rect 9550 10334 9602 10386
rect 9886 10334 9938 10386
rect 11230 10334 11282 10386
rect 12238 10334 12290 10386
rect 13582 10334 13634 10386
rect 13694 10334 13746 10386
rect 16270 10334 16322 10386
rect 16942 10334 16994 10386
rect 17166 10334 17218 10386
rect 4466 10166 4518 10218
rect 4570 10166 4622 10218
rect 4674 10166 4726 10218
rect 24466 10166 24518 10218
rect 24570 10166 24622 10218
rect 24674 10166 24726 10218
rect 5406 9998 5458 10050
rect 7422 9998 7474 10050
rect 12686 9998 12738 10050
rect 13918 9998 13970 10050
rect 15374 9998 15426 10050
rect 16046 9998 16098 10050
rect 18958 9998 19010 10050
rect 6526 9886 6578 9938
rect 7086 9886 7138 9938
rect 9102 9886 9154 9938
rect 10110 9886 10162 9938
rect 13134 9886 13186 9938
rect 15150 9886 15202 9938
rect 16158 9886 16210 9938
rect 17166 9886 17218 9938
rect 19406 9886 19458 9938
rect 2046 9774 2098 9826
rect 3838 9774 3890 9826
rect 4958 9774 5010 9826
rect 7310 9774 7362 9826
rect 7534 9774 7586 9826
rect 7870 9774 7922 9826
rect 9550 9774 9602 9826
rect 9998 9774 10050 9826
rect 10782 9774 10834 9826
rect 11342 9774 11394 9826
rect 12238 9774 12290 9826
rect 13246 9774 13298 9826
rect 13470 9774 13522 9826
rect 13806 9774 13858 9826
rect 14926 9774 14978 9826
rect 15710 9774 15762 9826
rect 16606 9774 16658 9826
rect 17054 9774 17106 9826
rect 17278 9774 17330 9826
rect 18398 9774 18450 9826
rect 18846 9774 18898 9826
rect 19966 9774 20018 9826
rect 21086 9774 21138 9826
rect 1262 9662 1314 9714
rect 2830 9662 2882 9714
rect 17950 9662 18002 9714
rect 14030 9550 14082 9602
rect 14254 9550 14306 9602
rect 15374 9550 15426 9602
rect 3806 9382 3858 9434
rect 3910 9382 3962 9434
rect 4014 9382 4066 9434
rect 23806 9382 23858 9434
rect 23910 9382 23962 9434
rect 24014 9382 24066 9434
rect 1262 9214 1314 9266
rect 9662 9214 9714 9266
rect 12126 9214 12178 9266
rect 13806 9214 13858 9266
rect 16494 9214 16546 9266
rect 17054 9214 17106 9266
rect 2942 9102 2994 9154
rect 5518 9102 5570 9154
rect 6414 9102 6466 9154
rect 7422 9102 7474 9154
rect 10558 9102 10610 9154
rect 18622 9102 18674 9154
rect 2270 8990 2322 9042
rect 3838 8990 3890 9042
rect 4958 8990 5010 9042
rect 5966 8990 6018 9042
rect 6974 8990 7026 9042
rect 7534 8990 7586 9042
rect 8094 8990 8146 9042
rect 12798 8990 12850 9042
rect 13022 8990 13074 9042
rect 14814 8990 14866 9042
rect 7310 8878 7362 8930
rect 10894 8878 10946 8930
rect 18174 8878 18226 8930
rect 8542 8766 8594 8818
rect 15374 8766 15426 8818
rect 4466 8598 4518 8650
rect 4570 8598 4622 8650
rect 4674 8598 4726 8650
rect 24466 8598 24518 8650
rect 24570 8598 24622 8650
rect 24674 8598 24726 8650
rect 8430 8430 8482 8482
rect 12238 8430 12290 8482
rect 3054 8318 3106 8370
rect 6302 8318 6354 8370
rect 7198 8318 7250 8370
rect 8094 8318 8146 8370
rect 8206 8318 8258 8370
rect 11118 8318 11170 8370
rect 13358 8318 13410 8370
rect 14926 8318 14978 8370
rect 15710 8318 15762 8370
rect 17614 8318 17666 8370
rect 20526 8318 20578 8370
rect 20974 8318 21026 8370
rect 2270 8206 2322 8258
rect 3838 8206 3890 8258
rect 6638 8206 6690 8258
rect 10558 8206 10610 8258
rect 12798 8206 12850 8258
rect 15038 8206 15090 8258
rect 15374 8206 15426 8258
rect 15598 8206 15650 8258
rect 16942 8206 16994 8258
rect 17278 8206 17330 8258
rect 17390 8206 17442 8258
rect 19854 8206 19906 8258
rect 20302 8206 20354 8258
rect 21758 8206 21810 8258
rect 22542 8206 22594 8258
rect 1262 8094 1314 8146
rect 7758 8094 7810 8146
rect 17502 8094 17554 8146
rect 19518 8094 19570 8146
rect 5070 7982 5122 8034
rect 14478 7982 14530 8034
rect 16158 7982 16210 8034
rect 16718 7982 16770 8034
rect 3806 7814 3858 7866
rect 3910 7814 3962 7866
rect 4014 7814 4066 7866
rect 23806 7814 23858 7866
rect 23910 7814 23962 7866
rect 24014 7814 24066 7866
rect 2830 7646 2882 7698
rect 10894 7646 10946 7698
rect 12238 7646 12290 7698
rect 16606 7646 16658 7698
rect 16718 7646 16770 7698
rect 1374 7534 1426 7586
rect 7310 7534 7362 7586
rect 9326 7534 9378 7586
rect 13022 7534 13074 7586
rect 16382 7534 16434 7586
rect 17054 7534 17106 7586
rect 2270 7422 2322 7474
rect 3838 7422 3890 7474
rect 6750 7422 6802 7474
rect 12126 7422 12178 7474
rect 14590 7422 14642 7474
rect 15598 7422 15650 7474
rect 15934 7422 15986 7474
rect 16158 7422 16210 7474
rect 17390 7422 17442 7474
rect 9774 7310 9826 7362
rect 13358 7310 13410 7362
rect 15710 7198 15762 7250
rect 4466 7030 4518 7082
rect 4570 7030 4622 7082
rect 4674 7030 4726 7082
rect 24466 7030 24518 7082
rect 24570 7030 24622 7082
rect 24674 7030 24726 7082
rect 13918 6862 13970 6914
rect 12686 6750 12738 6802
rect 2158 6638 2210 6690
rect 3614 6638 3666 6690
rect 10110 6638 10162 6690
rect 11006 6638 11058 6690
rect 11566 6638 11618 6690
rect 12350 6638 12402 6690
rect 1262 6526 1314 6578
rect 9774 6526 9826 6578
rect 2830 6414 2882 6466
rect 3806 6246 3858 6298
rect 3910 6246 3962 6298
rect 4014 6246 4066 6298
rect 23806 6246 23858 6298
rect 23910 6246 23962 6298
rect 24014 6246 24066 6298
rect 7758 6078 7810 6130
rect 1598 5966 1650 6018
rect 3166 5966 3218 6018
rect 9326 5966 9378 6018
rect 13806 5966 13858 6018
rect 2270 5854 2322 5906
rect 2606 5854 2658 5906
rect 11678 5854 11730 5906
rect 14254 5854 14306 5906
rect 14702 5854 14754 5906
rect 16046 5854 16098 5906
rect 16942 5854 16994 5906
rect 12126 5742 12178 5794
rect 15262 5742 15314 5794
rect 8878 5630 8930 5682
rect 14814 5630 14866 5682
rect 4466 5462 4518 5514
rect 4570 5462 4622 5514
rect 4674 5462 4726 5514
rect 24466 5462 24518 5514
rect 24570 5462 24622 5514
rect 24674 5462 24726 5514
rect 3614 5294 3666 5346
rect 7758 5294 7810 5346
rect 12238 5294 12290 5346
rect 14926 5294 14978 5346
rect 15374 5294 15426 5346
rect 1486 5182 1538 5234
rect 2270 5182 2322 5234
rect 3054 5182 3106 5234
rect 8318 5182 8370 5234
rect 12798 5182 12850 5234
rect 13694 5182 13746 5234
rect 15934 5182 15986 5234
rect 13246 5070 13298 5122
rect 3806 4678 3858 4730
rect 3910 4678 3962 4730
rect 4014 4678 4066 4730
rect 23806 4678 23858 4730
rect 23910 4678 23962 4730
rect 24014 4678 24066 4730
rect 1486 4174 1538 4226
rect 2270 4174 2322 4226
rect 4466 3894 4518 3946
rect 4570 3894 4622 3946
rect 4674 3894 4726 3946
rect 24466 3894 24518 3946
rect 24570 3894 24622 3946
rect 24674 3894 24726 3946
rect 2270 3502 2322 3554
rect 1262 3278 1314 3330
rect 3806 3110 3858 3162
rect 3910 3110 3962 3162
rect 4014 3110 4066 3162
rect 23806 3110 23858 3162
rect 23910 3110 23962 3162
rect 24014 3110 24066 3162
rect 4466 2326 4518 2378
rect 4570 2326 4622 2378
rect 4674 2326 4726 2378
rect 24466 2326 24518 2378
rect 24570 2326 24622 2378
rect 24674 2326 24726 2378
rect 11454 2046 11506 2098
rect 13246 2046 13298 2098
rect 26574 2046 26626 2098
rect 27470 2046 27522 2098
rect 12014 1934 12066 1986
rect 13806 1934 13858 1986
rect 26014 1934 26066 1986
rect 26910 1934 26962 1986
rect 3806 1542 3858 1594
rect 3910 1542 3962 1594
rect 4014 1542 4066 1594
rect 23806 1542 23858 1594
rect 23910 1542 23962 1594
rect 24014 1542 24066 1594
rect 4466 758 4518 810
rect 4570 758 4622 810
rect 4674 758 4726 810
rect 24466 758 24518 810
rect 24570 758 24622 810
rect 24674 758 24726 810
<< metal2 >>
rect 672 57344 784 57456
rect 2016 57344 2128 57456
rect 3360 57344 3472 57456
rect 4704 57344 4816 57456
rect 6048 57344 6160 57456
rect 7392 57344 7504 57456
rect 8736 57344 8848 57456
rect 10080 57344 10192 57456
rect 11424 57344 11536 57456
rect 12768 57344 12880 57456
rect 14112 57344 14224 57456
rect 15456 57344 15568 57456
rect 16800 57344 16912 57456
rect 18144 57344 18256 57456
rect 19488 57344 19600 57456
rect 19852 57372 20356 57428
rect 700 55972 756 57344
rect 1036 55972 1092 55982
rect 700 55970 1092 55972
rect 700 55918 1038 55970
rect 1090 55918 1092 55970
rect 700 55916 1092 55918
rect 1036 55906 1092 55916
rect 1372 55858 1428 55870
rect 1372 55806 1374 55858
rect 1426 55806 1428 55858
rect 1372 53844 1428 55806
rect 2044 55468 2100 57344
rect 3388 56308 3444 57344
rect 4732 56644 4788 57344
rect 4732 56588 5236 56644
rect 3804 56476 4068 56486
rect 3860 56420 3908 56476
rect 3964 56420 4012 56476
rect 3804 56410 4068 56420
rect 3612 56308 3668 56318
rect 3388 56306 3668 56308
rect 3388 56254 3614 56306
rect 3666 56254 3668 56306
rect 3388 56252 3668 56254
rect 3612 56242 3668 56252
rect 5180 56306 5236 56588
rect 5180 56254 5182 56306
rect 5234 56254 5236 56306
rect 5180 56242 5236 56254
rect 3052 55970 3108 55982
rect 3052 55918 3054 55970
rect 3106 55918 3108 55970
rect 3052 55468 3108 55918
rect 4464 55692 4728 55702
rect 4520 55636 4568 55692
rect 4624 55636 4672 55692
rect 4464 55626 4728 55636
rect 2044 55412 2548 55468
rect 2492 55186 2548 55412
rect 2492 55134 2494 55186
rect 2546 55134 2548 55186
rect 2492 55122 2548 55134
rect 2716 55412 3108 55468
rect 1372 53778 1428 53788
rect 2044 53396 2100 53406
rect 1484 52500 1540 52510
rect 588 41748 644 41758
rect 252 39620 308 39630
rect 252 532 308 39564
rect 588 38612 644 41692
rect 364 37380 420 37390
rect 364 23268 420 37324
rect 364 23202 420 23212
rect 476 29428 532 29438
rect 476 1652 532 29372
rect 588 21812 644 38556
rect 924 40964 980 40974
rect 812 38164 868 38174
rect 812 28532 868 38108
rect 812 28466 868 28476
rect 588 21746 644 21756
rect 700 18452 756 18462
rect 700 9268 756 18396
rect 700 9202 756 9212
rect 812 12180 868 12190
rect 812 6580 868 12124
rect 924 6916 980 40908
rect 1148 38722 1204 38734
rect 1148 38670 1150 38722
rect 1202 38670 1204 38722
rect 1148 38612 1204 38670
rect 1484 38668 1540 52444
rect 1596 45220 1652 45230
rect 1596 38946 1652 45164
rect 1932 42644 1988 42654
rect 1820 40852 1876 40862
rect 1596 38894 1598 38946
rect 1650 38894 1652 38946
rect 1596 38882 1652 38894
rect 1708 39060 1764 39070
rect 1484 38612 1652 38668
rect 1148 38276 1204 38556
rect 1148 38210 1204 38220
rect 1372 37938 1428 37950
rect 1372 37886 1374 37938
rect 1426 37886 1428 37938
rect 1372 35812 1428 37886
rect 1036 35756 1372 35812
rect 1036 32676 1092 35756
rect 1372 35746 1428 35756
rect 1148 35476 1204 35486
rect 1148 35474 1540 35476
rect 1148 35422 1150 35474
rect 1202 35422 1540 35474
rect 1148 35420 1540 35422
rect 1148 35410 1204 35420
rect 1484 34130 1540 35420
rect 1484 34078 1486 34130
rect 1538 34078 1540 34130
rect 1484 34066 1540 34078
rect 1148 34020 1204 34030
rect 1148 33926 1204 33964
rect 1036 32564 1092 32620
rect 1484 32676 1540 32686
rect 1148 32564 1204 32574
rect 1036 32562 1204 32564
rect 1036 32510 1150 32562
rect 1202 32510 1204 32562
rect 1036 32508 1204 32510
rect 1148 32498 1204 32508
rect 1484 31780 1540 32620
rect 1484 31714 1540 31724
rect 1596 32450 1652 38612
rect 1708 37492 1764 39004
rect 1820 38162 1876 40796
rect 1932 40180 1988 42588
rect 1932 40114 1988 40124
rect 1820 38110 1822 38162
rect 1874 38110 1876 38162
rect 1820 37716 1876 38110
rect 1820 37650 1876 37660
rect 1708 37436 1876 37492
rect 1708 37266 1764 37278
rect 1708 37214 1710 37266
rect 1762 37214 1764 37266
rect 1708 36932 1764 37214
rect 1708 36484 1764 36876
rect 1708 36418 1764 36428
rect 1596 32398 1598 32450
rect 1650 32398 1652 32450
rect 1596 30324 1652 32398
rect 1708 36260 1764 36270
rect 1708 32004 1764 36204
rect 1708 31938 1764 31948
rect 1596 30258 1652 30268
rect 1708 31780 1764 31790
rect 1596 30098 1652 30110
rect 1596 30046 1598 30098
rect 1650 30046 1652 30098
rect 1036 29988 1092 29998
rect 1036 22148 1092 29932
rect 1148 29540 1204 29550
rect 1148 29446 1204 29484
rect 1484 29428 1540 29438
rect 1484 29334 1540 29372
rect 1484 28532 1540 28542
rect 1484 27300 1540 28476
rect 1484 27234 1540 27244
rect 1596 28420 1652 30046
rect 1596 27972 1652 28364
rect 1260 27076 1316 27086
rect 1260 26982 1316 27020
rect 1596 26908 1652 27916
rect 1708 27524 1764 31724
rect 1820 28756 1876 37436
rect 1932 37156 1988 37166
rect 1932 36372 1988 37100
rect 2044 36596 2100 53340
rect 2716 43708 2772 55412
rect 2380 43652 2772 43708
rect 2828 55300 2884 55310
rect 2156 39956 2212 39966
rect 2156 37716 2212 39900
rect 2268 38834 2324 38846
rect 2268 38782 2270 38834
rect 2322 38782 2324 38834
rect 2268 37828 2324 38782
rect 2380 38668 2436 43652
rect 2604 40180 2660 40190
rect 2604 39618 2660 40124
rect 2604 39566 2606 39618
rect 2658 39566 2660 39618
rect 2604 38836 2660 39566
rect 2604 38770 2660 38780
rect 2716 39844 2772 39854
rect 2716 38722 2772 39788
rect 2716 38670 2718 38722
rect 2770 38670 2772 38722
rect 2380 38612 2660 38668
rect 2716 38658 2772 38670
rect 2268 37772 2548 37828
rect 2156 37660 2436 37716
rect 2156 37492 2212 37502
rect 2156 37378 2212 37436
rect 2156 37326 2158 37378
rect 2210 37326 2212 37378
rect 2156 37314 2212 37326
rect 2044 36540 2212 36596
rect 2044 36372 2100 36382
rect 1932 36370 2100 36372
rect 1932 36318 2046 36370
rect 2098 36318 2100 36370
rect 1932 36316 2100 36318
rect 2044 36306 2100 36316
rect 1932 34916 1988 34926
rect 1932 34130 1988 34860
rect 1932 34078 1934 34130
rect 1986 34078 1988 34130
rect 1932 34066 1988 34078
rect 2044 34914 2100 34926
rect 2044 34862 2046 34914
rect 2098 34862 2100 34914
rect 2044 34020 2100 34862
rect 2156 34244 2212 36540
rect 2380 35586 2436 37660
rect 2492 36932 2548 37772
rect 2492 36866 2548 36876
rect 2604 36708 2660 38612
rect 2828 37492 2884 55244
rect 3500 55298 3556 55310
rect 3500 55246 3502 55298
rect 3554 55246 3556 55298
rect 2940 48916 2996 48926
rect 2940 40292 2996 48860
rect 2940 40226 2996 40236
rect 3052 46788 3108 46798
rect 3052 39730 3108 46732
rect 3052 39678 3054 39730
rect 3106 39678 3108 39730
rect 3052 39666 3108 39678
rect 3164 40516 3220 40526
rect 2828 37426 2884 37436
rect 2940 37826 2996 37838
rect 2940 37774 2942 37826
rect 2994 37774 2996 37826
rect 2716 37266 2772 37278
rect 2716 37214 2718 37266
rect 2770 37214 2772 37266
rect 2716 37044 2772 37214
rect 2716 36978 2772 36988
rect 2380 35534 2382 35586
rect 2434 35534 2436 35586
rect 2380 35522 2436 35534
rect 2492 36652 2660 36708
rect 2268 35474 2324 35486
rect 2268 35422 2270 35474
rect 2322 35422 2324 35474
rect 2268 34468 2324 35422
rect 2492 35028 2548 36652
rect 2828 36596 2884 36606
rect 2604 36482 2660 36494
rect 2604 36430 2606 36482
rect 2658 36430 2660 36482
rect 2604 35252 2660 36430
rect 2716 35812 2772 35822
rect 2716 35718 2772 35756
rect 2828 35476 2884 36540
rect 2604 35186 2660 35196
rect 2716 35420 2884 35476
rect 2492 34972 2660 35028
rect 2268 34402 2324 34412
rect 2380 34804 2436 34814
rect 2156 34188 2324 34244
rect 2156 34020 2212 34030
rect 2044 34018 2212 34020
rect 2044 33966 2158 34018
rect 2210 33966 2212 34018
rect 2044 33964 2212 33966
rect 2156 33954 2212 33964
rect 1820 28690 1876 28700
rect 1932 33908 1988 33918
rect 1708 27468 1876 27524
rect 1484 26852 1652 26908
rect 1708 27300 1764 27310
rect 1260 26516 1316 26526
rect 1260 25394 1316 26460
rect 1260 25342 1262 25394
rect 1314 25342 1316 25394
rect 1260 25330 1316 25342
rect 1372 23828 1428 23838
rect 1148 23268 1204 23278
rect 1148 23174 1204 23212
rect 1260 23156 1316 23166
rect 1260 22370 1316 23100
rect 1260 22318 1262 22370
rect 1314 22318 1316 22370
rect 1260 22306 1316 22318
rect 1036 22092 1316 22148
rect 1260 20914 1316 22092
rect 1260 20862 1262 20914
rect 1314 20862 1316 20914
rect 1260 20850 1316 20862
rect 1148 19348 1204 19358
rect 1036 17556 1092 17566
rect 1036 8428 1092 17500
rect 1148 9716 1204 19292
rect 1372 19122 1428 23772
rect 1484 23268 1540 26852
rect 1708 24500 1764 27244
rect 1820 27076 1876 27468
rect 1820 24722 1876 27020
rect 1932 25508 1988 33852
rect 2268 33460 2324 34188
rect 2156 33404 2324 33460
rect 2380 34020 2436 34748
rect 2492 34802 2548 34814
rect 2492 34750 2494 34802
rect 2546 34750 2548 34802
rect 2492 34356 2548 34750
rect 2492 34290 2548 34300
rect 2156 31890 2212 33404
rect 2268 33236 2324 33246
rect 2380 33236 2436 33964
rect 2268 33234 2436 33236
rect 2268 33182 2270 33234
rect 2322 33182 2436 33234
rect 2268 33180 2436 33182
rect 2492 34132 2548 34142
rect 2268 32340 2324 33180
rect 2268 32274 2324 32284
rect 2156 31838 2158 31890
rect 2210 31838 2212 31890
rect 2044 28530 2100 28542
rect 2044 28478 2046 28530
rect 2098 28478 2100 28530
rect 2044 28420 2100 28478
rect 2044 28354 2100 28364
rect 2044 26290 2100 26302
rect 2044 26238 2046 26290
rect 2098 26238 2100 26290
rect 2044 25956 2100 26238
rect 2156 26180 2212 31838
rect 2380 32004 2436 32014
rect 2268 30210 2324 30222
rect 2268 30158 2270 30210
rect 2322 30158 2324 30210
rect 2268 29540 2324 30158
rect 2380 29876 2436 31948
rect 2492 30100 2548 34076
rect 2604 30548 2660 34972
rect 2716 34132 2772 35420
rect 2828 34804 2884 34814
rect 2828 34710 2884 34748
rect 2716 34066 2772 34076
rect 2828 34132 2884 34142
rect 2940 34132 2996 37774
rect 3164 37380 3220 40460
rect 3500 39732 3556 55246
rect 6076 55188 6132 57344
rect 7420 56194 7476 57344
rect 8764 56644 8820 57344
rect 10108 56756 10164 57344
rect 10108 56700 10612 56756
rect 8764 56588 9044 56644
rect 8988 56306 9044 56588
rect 8988 56254 8990 56306
rect 9042 56254 9044 56306
rect 8988 56242 9044 56254
rect 10556 56306 10612 56700
rect 10556 56254 10558 56306
rect 10610 56254 10612 56306
rect 10556 56242 10612 56254
rect 7420 56142 7422 56194
rect 7474 56142 7476 56194
rect 7420 56130 7476 56142
rect 7868 56082 7924 56094
rect 7868 56030 7870 56082
rect 7922 56030 7924 56082
rect 6188 55972 6244 55982
rect 6188 55878 6244 55916
rect 6300 55300 6356 55310
rect 6300 55206 6356 55244
rect 6076 55122 6132 55132
rect 6860 55188 6916 55198
rect 6860 55094 6916 55132
rect 3804 54908 4068 54918
rect 3860 54852 3908 54908
rect 3964 54852 4012 54908
rect 3804 54842 4068 54852
rect 5964 54292 6020 54302
rect 4464 54124 4728 54134
rect 4520 54068 4568 54124
rect 4624 54068 4672 54124
rect 4464 54058 4728 54068
rect 3804 53340 4068 53350
rect 3860 53284 3908 53340
rect 3964 53284 4012 53340
rect 3804 53274 4068 53284
rect 4464 52556 4728 52566
rect 4520 52500 4568 52556
rect 4624 52500 4672 52556
rect 4464 52490 4728 52500
rect 3804 51772 4068 51782
rect 3860 51716 3908 51772
rect 3964 51716 4012 51772
rect 3804 51706 4068 51716
rect 4464 50988 4728 50998
rect 4520 50932 4568 50988
rect 4624 50932 4672 50988
rect 4464 50922 4728 50932
rect 5964 50428 6020 54236
rect 6748 54068 6804 54078
rect 5964 50372 6244 50428
rect 3804 50204 4068 50214
rect 3860 50148 3908 50204
rect 3964 50148 4012 50204
rect 3804 50138 4068 50148
rect 5292 49812 5348 49822
rect 4464 49420 4728 49430
rect 4520 49364 4568 49420
rect 4624 49364 4672 49420
rect 4464 49354 4728 49364
rect 3804 48636 4068 48646
rect 3860 48580 3908 48636
rect 3964 48580 4012 48636
rect 3804 48570 4068 48580
rect 4464 47852 4728 47862
rect 4520 47796 4568 47852
rect 4624 47796 4672 47852
rect 4464 47786 4728 47796
rect 3804 47068 4068 47078
rect 3860 47012 3908 47068
rect 3964 47012 4012 47068
rect 3804 47002 4068 47012
rect 4464 46284 4728 46294
rect 4520 46228 4568 46284
rect 4624 46228 4672 46284
rect 4464 46218 4728 46228
rect 3804 45500 4068 45510
rect 3860 45444 3908 45500
rect 3964 45444 4012 45500
rect 3804 45434 4068 45444
rect 4464 44716 4728 44726
rect 4520 44660 4568 44716
rect 4624 44660 4672 44716
rect 4464 44650 4728 44660
rect 3804 43932 4068 43942
rect 3860 43876 3908 43932
rect 3964 43876 4012 43932
rect 3804 43866 4068 43876
rect 4464 43148 4728 43158
rect 4520 43092 4568 43148
rect 4624 43092 4672 43148
rect 4464 43082 4728 43092
rect 3804 42364 4068 42374
rect 3860 42308 3908 42364
rect 3964 42308 4012 42364
rect 3804 42298 4068 42308
rect 4464 41580 4728 41590
rect 4520 41524 4568 41580
rect 4624 41524 4672 41580
rect 4464 41514 4728 41524
rect 3804 40796 4068 40806
rect 3860 40740 3908 40796
rect 3964 40740 4012 40796
rect 3804 40730 4068 40740
rect 5180 40180 5236 40190
rect 4464 40012 4728 40022
rect 4520 39956 4568 40012
rect 4624 39956 4672 40012
rect 4464 39946 4728 39956
rect 3500 39666 3556 39676
rect 4172 39844 4228 39854
rect 3836 39620 3892 39630
rect 3836 39526 3892 39564
rect 4172 39620 4228 39788
rect 3500 39506 3556 39518
rect 3500 39454 3502 39506
rect 3554 39454 3556 39506
rect 3500 38948 3556 39454
rect 3804 39228 4068 39238
rect 3860 39172 3908 39228
rect 3964 39172 4012 39228
rect 3804 39162 4068 39172
rect 3500 38882 3556 38892
rect 4172 38668 4228 39564
rect 5068 38948 5124 38958
rect 3836 38610 3892 38622
rect 4172 38612 4340 38668
rect 3836 38558 3838 38610
rect 3890 38558 3892 38610
rect 3836 37828 3892 38558
rect 3836 37772 4228 37828
rect 3804 37660 4068 37670
rect 3860 37604 3908 37660
rect 3964 37604 4012 37660
rect 3804 37594 4068 37604
rect 4172 37492 4228 37772
rect 3164 37314 3220 37324
rect 4060 37436 4228 37492
rect 3164 37042 3220 37054
rect 3164 36990 3166 37042
rect 3218 36990 3220 37042
rect 3164 36596 3220 36990
rect 3164 36530 3220 36540
rect 3388 37044 3444 37054
rect 3052 36258 3108 36270
rect 3052 36206 3054 36258
rect 3106 36206 3108 36258
rect 3052 34916 3108 36206
rect 3164 34916 3220 34926
rect 3052 34914 3220 34916
rect 3052 34862 3166 34914
rect 3218 34862 3220 34914
rect 3052 34860 3220 34862
rect 3164 34850 3220 34860
rect 2828 34130 2996 34132
rect 2828 34078 2830 34130
rect 2882 34078 2996 34130
rect 2828 34076 2996 34078
rect 3052 34468 3108 34478
rect 2828 34066 2884 34076
rect 2716 33346 2772 33358
rect 2716 33294 2718 33346
rect 2770 33294 2772 33346
rect 2716 32788 2772 33294
rect 2828 32788 2884 32798
rect 2716 32786 2884 32788
rect 2716 32734 2830 32786
rect 2882 32734 2884 32786
rect 2716 32732 2884 32734
rect 2828 32722 2884 32732
rect 2716 30994 2772 31006
rect 2716 30942 2718 30994
rect 2770 30942 2772 30994
rect 2716 30884 2772 30942
rect 2716 30818 2772 30828
rect 3052 30772 3108 34412
rect 3164 34130 3220 34142
rect 3164 34078 3166 34130
rect 3218 34078 3220 34130
rect 3164 33572 3220 34078
rect 3388 33796 3444 36988
rect 3612 36596 3668 36606
rect 3612 35252 3668 36540
rect 4060 36372 4116 37436
rect 4284 37380 4340 38612
rect 4464 38444 4728 38454
rect 4520 38388 4568 38444
rect 4624 38388 4672 38444
rect 4464 38378 4728 38388
rect 4844 38276 4900 38286
rect 4844 38182 4900 38220
rect 4396 37940 4452 37950
rect 4396 37846 4452 37884
rect 4172 37324 4340 37380
rect 4844 37380 4900 37390
rect 4172 36596 4228 37324
rect 4172 36502 4228 36540
rect 4284 37042 4340 37054
rect 4284 36990 4286 37042
rect 4338 36990 4340 37042
rect 4060 36316 4228 36372
rect 3804 36092 4068 36102
rect 3860 36036 3908 36092
rect 3964 36036 4012 36092
rect 3804 36026 4068 36036
rect 3836 35476 3892 35486
rect 3724 35474 3892 35476
rect 3724 35422 3838 35474
rect 3890 35422 3892 35474
rect 3724 35420 3892 35422
rect 3724 35252 3780 35420
rect 3836 35410 3892 35420
rect 3388 33730 3444 33740
rect 3500 35196 3780 35252
rect 3836 35252 3892 35262
rect 3164 33506 3220 33516
rect 3276 33460 3332 33470
rect 3276 33458 3444 33460
rect 3276 33406 3278 33458
rect 3330 33406 3444 33458
rect 3276 33404 3444 33406
rect 3276 33394 3332 33404
rect 3164 33346 3220 33358
rect 3164 33294 3166 33346
rect 3218 33294 3220 33346
rect 3164 30996 3220 33294
rect 3276 33236 3332 33246
rect 3276 31890 3332 33180
rect 3388 32562 3444 33404
rect 3388 32510 3390 32562
rect 3442 32510 3444 32562
rect 3388 32498 3444 32510
rect 3500 32340 3556 35196
rect 3836 35138 3892 35196
rect 3836 35086 3838 35138
rect 3890 35086 3892 35138
rect 3836 35074 3892 35086
rect 3724 35028 3780 35038
rect 3724 34914 3780 34972
rect 3724 34862 3726 34914
rect 3778 34862 3780 34914
rect 3724 34850 3780 34862
rect 4172 34804 4228 36316
rect 4284 35026 4340 36990
rect 4844 37044 4900 37324
rect 4464 36876 4728 36886
rect 4520 36820 4568 36876
rect 4624 36820 4672 36876
rect 4464 36810 4728 36820
rect 4732 36484 4788 36494
rect 4844 36484 4900 36988
rect 4732 36482 4900 36484
rect 4732 36430 4734 36482
rect 4786 36430 4900 36482
rect 4732 36428 4900 36430
rect 4732 36418 4788 36428
rect 4396 35812 4452 35822
rect 4396 35718 4452 35756
rect 4464 35308 4728 35318
rect 4520 35252 4568 35308
rect 4624 35252 4672 35308
rect 4464 35242 4728 35252
rect 4284 34974 4286 35026
rect 4338 34974 4340 35026
rect 4284 34962 4340 34974
rect 4956 34914 5012 34926
rect 4956 34862 4958 34914
rect 5010 34862 5012 34914
rect 4172 34748 4340 34804
rect 3804 34524 4068 34534
rect 3860 34468 3908 34524
rect 3964 34468 4012 34524
rect 3804 34458 4068 34468
rect 4172 34132 4228 34142
rect 4172 34038 4228 34076
rect 3276 31838 3278 31890
rect 3330 31838 3332 31890
rect 3276 31826 3332 31838
rect 3388 32284 3556 32340
rect 3612 33796 3668 33806
rect 4284 33796 4340 34748
rect 3164 30940 3332 30996
rect 2604 30482 2660 30492
rect 2940 30716 3108 30772
rect 3164 30772 3220 30782
rect 2940 30436 2996 30716
rect 3164 30678 3220 30716
rect 2828 30324 2884 30334
rect 2492 30034 2548 30044
rect 2716 30210 2772 30222
rect 2716 30158 2718 30210
rect 2770 30158 2772 30210
rect 2380 29820 2548 29876
rect 2268 29474 2324 29484
rect 2492 28868 2548 29820
rect 2716 29540 2772 30158
rect 2716 29446 2772 29484
rect 2492 28802 2548 28812
rect 2380 28756 2436 28766
rect 2156 26114 2212 26124
rect 2268 27858 2324 27870
rect 2268 27806 2270 27858
rect 2322 27806 2324 27858
rect 2268 25956 2324 27806
rect 2380 26908 2436 28700
rect 2828 27748 2884 30268
rect 2940 29092 2996 30380
rect 3052 30548 3108 30558
rect 3052 30098 3108 30492
rect 3052 30046 3054 30098
rect 3106 30046 3108 30098
rect 3052 30034 3108 30046
rect 3276 30212 3332 30940
rect 3276 29428 3332 30156
rect 2940 29026 2996 29036
rect 3052 29372 3332 29428
rect 2716 27746 2884 27748
rect 2716 27694 2830 27746
rect 2882 27694 2884 27746
rect 2716 27692 2884 27694
rect 2380 26852 2548 26908
rect 2380 26180 2436 26190
rect 2380 26086 2436 26124
rect 2044 25900 2324 25956
rect 2044 25508 2100 25518
rect 1932 25506 2100 25508
rect 1932 25454 2046 25506
rect 2098 25454 2100 25506
rect 1932 25452 2100 25454
rect 2044 25442 2100 25452
rect 1820 24670 1822 24722
rect 1874 24670 1876 24722
rect 1820 24658 1876 24670
rect 2044 25284 2100 25294
rect 1708 24444 1988 24500
rect 1484 23202 1540 23212
rect 1596 24052 1652 24062
rect 1596 23154 1652 23996
rect 1596 23102 1598 23154
rect 1650 23102 1652 23154
rect 1596 23090 1652 23102
rect 1708 23268 1764 23278
rect 1596 22482 1652 22494
rect 1596 22430 1598 22482
rect 1650 22430 1652 22482
rect 1372 19070 1374 19122
rect 1426 19070 1428 19122
rect 1372 19058 1428 19070
rect 1484 22036 1540 22046
rect 1372 18676 1428 18686
rect 1260 17444 1316 17454
rect 1260 16994 1316 17388
rect 1260 16942 1262 16994
rect 1314 16942 1316 16994
rect 1260 16930 1316 16942
rect 1372 16098 1428 18620
rect 1372 16046 1374 16098
rect 1426 16046 1428 16098
rect 1372 14532 1428 16046
rect 1372 14466 1428 14476
rect 1372 13972 1428 13982
rect 1260 9716 1316 9726
rect 1148 9714 1316 9716
rect 1148 9662 1262 9714
rect 1314 9662 1316 9714
rect 1148 9660 1316 9662
rect 1260 9650 1316 9660
rect 1260 9268 1316 9278
rect 1260 9174 1316 9212
rect 1036 8372 1316 8428
rect 1260 8146 1316 8372
rect 1260 8094 1262 8146
rect 1314 8094 1316 8146
rect 1260 8082 1316 8094
rect 1372 7586 1428 13916
rect 1484 13074 1540 21980
rect 1596 21812 1652 22430
rect 1596 21746 1652 21756
rect 1708 20018 1764 23212
rect 1820 20916 1876 20926
rect 1820 20822 1876 20860
rect 1932 20692 1988 24444
rect 1708 19966 1710 20018
rect 1762 19966 1764 20018
rect 1708 18676 1764 19966
rect 1596 18620 1764 18676
rect 1820 20636 1988 20692
rect 1596 18004 1652 18620
rect 1708 18452 1764 18462
rect 1820 18452 1876 20636
rect 1708 18450 1876 18452
rect 1708 18398 1710 18450
rect 1762 18398 1876 18450
rect 1708 18396 1876 18398
rect 1932 20468 1988 20478
rect 1708 18228 1764 18396
rect 1708 18162 1764 18172
rect 1596 17948 1764 18004
rect 1708 17444 1764 17948
rect 1708 17378 1764 17388
rect 1820 17671 1876 17683
rect 1820 17619 1822 17671
rect 1874 17619 1876 17671
rect 1820 17108 1876 17619
rect 1820 17042 1876 17052
rect 1596 16772 1652 16782
rect 1596 16678 1652 16716
rect 1820 16324 1876 16362
rect 1820 16258 1876 16268
rect 1708 15316 1764 15326
rect 1708 15222 1764 15260
rect 1596 14532 1652 14542
rect 1596 14438 1652 14476
rect 1932 14308 1988 20412
rect 2044 16772 2100 25228
rect 2268 24052 2324 25900
rect 2380 24612 2436 24622
rect 2492 24612 2548 26852
rect 2380 24610 2548 24612
rect 2380 24558 2382 24610
rect 2434 24558 2548 24610
rect 2380 24556 2548 24558
rect 2380 24546 2436 24556
rect 2492 24388 2548 24556
rect 2604 25394 2660 25406
rect 2604 25342 2606 25394
rect 2658 25342 2660 25394
rect 2604 24612 2660 25342
rect 2716 25284 2772 27692
rect 2828 27682 2884 27692
rect 2940 28868 2996 28878
rect 2828 26850 2884 26862
rect 2828 26798 2830 26850
rect 2882 26798 2884 26850
rect 2828 25508 2884 26798
rect 2940 26068 2996 28812
rect 3052 26908 3108 29372
rect 3388 29316 3444 32284
rect 3612 30436 3668 33740
rect 4172 33740 4340 33796
rect 4464 33740 4728 33750
rect 3724 33346 3780 33358
rect 3724 33294 3726 33346
rect 3778 33294 3780 33346
rect 3724 33236 3780 33294
rect 3724 33170 3780 33180
rect 3804 32956 4068 32966
rect 3860 32900 3908 32956
rect 3964 32900 4012 32956
rect 3804 32890 4068 32900
rect 3836 32452 3892 32462
rect 3836 32358 3892 32396
rect 3804 31388 4068 31398
rect 3860 31332 3908 31388
rect 3964 31332 4012 31388
rect 3804 31322 4068 31332
rect 3612 30380 4116 30436
rect 3836 30212 3892 30222
rect 3612 30210 3892 30212
rect 3612 30158 3838 30210
rect 3890 30158 3892 30210
rect 3612 30156 3892 30158
rect 3500 30098 3556 30110
rect 3500 30046 3502 30098
rect 3554 30046 3556 30098
rect 3500 29428 3556 30046
rect 3500 29362 3556 29372
rect 3388 29250 3444 29260
rect 3164 29202 3220 29214
rect 3164 29150 3166 29202
rect 3218 29150 3220 29202
rect 3164 28532 3220 29150
rect 3276 29092 3332 29102
rect 3332 29036 3556 29092
rect 3276 29026 3332 29036
rect 3164 28466 3220 28476
rect 3276 26964 3332 27002
rect 3052 26852 3220 26908
rect 3276 26898 3332 26908
rect 3164 26292 3220 26852
rect 2940 26012 3108 26068
rect 2940 25508 2996 25518
rect 2828 25506 2996 25508
rect 2828 25454 2942 25506
rect 2994 25454 2996 25506
rect 2828 25452 2996 25454
rect 2940 25442 2996 25452
rect 2716 25218 2772 25228
rect 2604 24546 2660 24556
rect 2492 24332 2996 24388
rect 2268 23996 2660 24052
rect 2380 23828 2436 23838
rect 2268 23268 2324 23278
rect 2268 23174 2324 23212
rect 2156 20690 2212 20702
rect 2156 20638 2158 20690
rect 2210 20638 2212 20690
rect 2156 20188 2212 20638
rect 2156 20132 2324 20188
rect 2156 19796 2212 19806
rect 2156 19702 2212 19740
rect 2268 19572 2324 20132
rect 2156 19516 2324 19572
rect 2156 18676 2212 19516
rect 2268 19348 2324 19358
rect 2268 19254 2324 19292
rect 2156 18620 2324 18676
rect 2156 18452 2212 18462
rect 2156 18358 2212 18396
rect 2268 18228 2324 18620
rect 2044 16706 2100 16716
rect 2156 18172 2324 18228
rect 2156 16996 2212 18172
rect 2156 15764 2212 16940
rect 1484 13022 1486 13074
rect 1538 13022 1540 13074
rect 1484 13010 1540 13022
rect 1708 14252 1988 14308
rect 2044 15708 2212 15764
rect 2268 16772 2324 16782
rect 1596 11620 1652 11630
rect 1596 11526 1652 11564
rect 1372 7534 1374 7586
rect 1426 7534 1428 7586
rect 1372 7522 1428 7534
rect 1596 8596 1652 8606
rect 924 6850 980 6860
rect 1484 6804 1540 6814
rect 1260 6580 1316 6590
rect 812 6578 1316 6580
rect 812 6526 1262 6578
rect 1314 6526 1316 6578
rect 812 6524 1316 6526
rect 1260 6514 1316 6524
rect 1484 5234 1540 6748
rect 1596 6018 1652 8540
rect 1708 7700 1764 14252
rect 1820 13746 1876 13758
rect 1820 13694 1822 13746
rect 1874 13694 1876 13746
rect 1820 11732 1876 13694
rect 2044 13076 2100 15708
rect 2156 15540 2212 15550
rect 2156 15426 2212 15484
rect 2156 15374 2158 15426
rect 2210 15374 2212 15426
rect 2156 15362 2212 15374
rect 1820 11666 1876 11676
rect 1932 13020 2100 13076
rect 2156 14642 2212 14654
rect 2156 14590 2158 14642
rect 2210 14590 2212 14642
rect 1708 7634 1764 7644
rect 1820 8428 1876 8438
rect 1596 5966 1598 6018
rect 1650 5966 1652 6018
rect 1596 5954 1652 5966
rect 1484 5182 1486 5234
rect 1538 5182 1540 5234
rect 1484 5170 1540 5182
rect 1484 4226 1540 4238
rect 1484 4174 1486 4226
rect 1538 4174 1540 4226
rect 1484 4116 1540 4174
rect 1484 4050 1540 4060
rect 1260 3330 1316 3342
rect 1260 3278 1262 3330
rect 1314 3278 1316 3330
rect 1260 3220 1316 3278
rect 1260 3154 1316 3164
rect 1820 2324 1876 8372
rect 1932 5012 1988 13020
rect 2044 12178 2100 12190
rect 2044 12126 2046 12178
rect 2098 12126 2100 12178
rect 2044 11732 2100 12126
rect 2156 12180 2212 14590
rect 2268 13522 2324 16716
rect 2268 13470 2270 13522
rect 2322 13470 2324 13522
rect 2268 13188 2324 13470
rect 2268 13122 2324 13132
rect 2156 12114 2212 12124
rect 2268 12962 2324 12974
rect 2268 12910 2270 12962
rect 2322 12910 2324 12962
rect 2044 11666 2100 11676
rect 2268 11620 2324 12910
rect 2268 11554 2324 11564
rect 2268 11396 2324 11406
rect 2044 10612 2100 10622
rect 2044 10518 2100 10556
rect 2044 9826 2100 9838
rect 2044 9774 2046 9826
rect 2098 9774 2100 9826
rect 2044 9044 2100 9774
rect 2044 8978 2100 8988
rect 2268 9042 2324 11340
rect 2268 8990 2270 9042
rect 2322 8990 2324 9042
rect 2268 8978 2324 8990
rect 2380 8820 2436 23772
rect 2604 22372 2660 23996
rect 2828 23938 2884 23950
rect 2828 23886 2830 23938
rect 2882 23886 2884 23938
rect 2716 23156 2772 23166
rect 2716 23042 2772 23100
rect 2716 22990 2718 23042
rect 2770 22990 2772 23042
rect 2716 22978 2772 22990
rect 2828 22594 2884 23886
rect 2828 22542 2830 22594
rect 2882 22542 2884 22594
rect 2828 22530 2884 22542
rect 2604 21588 2660 22316
rect 2828 22260 2884 22270
rect 2604 21586 2772 21588
rect 2604 21534 2606 21586
rect 2658 21534 2772 21586
rect 2604 21532 2772 21534
rect 2604 21522 2660 21532
rect 2604 20802 2660 20814
rect 2604 20750 2606 20802
rect 2658 20750 2660 20802
rect 2492 19796 2548 19806
rect 2492 12964 2548 19740
rect 2604 18340 2660 20750
rect 2716 18562 2772 21532
rect 2828 20468 2884 22204
rect 2940 21700 2996 24332
rect 2940 21634 2996 21644
rect 2828 20402 2884 20412
rect 2940 20802 2996 20814
rect 2940 20750 2942 20802
rect 2994 20750 2996 20802
rect 2716 18510 2718 18562
rect 2770 18510 2772 18562
rect 2716 18498 2772 18510
rect 2940 20244 2996 20750
rect 2604 18284 2884 18340
rect 2716 17666 2772 17678
rect 2716 17614 2718 17666
rect 2770 17614 2772 17666
rect 2716 17556 2772 17614
rect 2716 17490 2772 17500
rect 2828 17106 2884 18284
rect 2940 17892 2996 20188
rect 3052 20188 3108 26012
rect 3164 23938 3220 26236
rect 3388 25506 3444 25518
rect 3388 25454 3390 25506
rect 3442 25454 3444 25506
rect 3388 24948 3444 25454
rect 3500 25060 3556 29036
rect 3612 28866 3668 30156
rect 3836 30146 3892 30156
rect 4060 30100 4116 30380
rect 4172 30324 4228 33740
rect 4520 33684 4568 33740
rect 4624 33684 4672 33740
rect 4464 33674 4728 33684
rect 4844 33684 4900 33694
rect 4508 33572 4564 33582
rect 4508 33346 4564 33516
rect 4508 33294 4510 33346
rect 4562 33294 4564 33346
rect 4508 32564 4564 33294
rect 4508 32498 4564 32508
rect 4464 32172 4728 32182
rect 4520 32116 4568 32172
rect 4624 32116 4672 32172
rect 4464 32106 4728 32116
rect 4284 31220 4340 31230
rect 4284 31126 4340 31164
rect 4844 30884 4900 33628
rect 4956 33572 5012 34862
rect 5068 34130 5124 38892
rect 5068 34078 5070 34130
rect 5122 34078 5124 34130
rect 5068 34020 5124 34078
rect 5068 33954 5124 33964
rect 4956 33506 5012 33516
rect 5180 32788 5236 40124
rect 5292 38724 5348 49756
rect 5292 38658 5348 38668
rect 5404 42084 5460 42094
rect 5404 38946 5460 42028
rect 6076 40402 6132 40414
rect 6076 40350 6078 40402
rect 6130 40350 6132 40402
rect 6076 40180 6132 40350
rect 6076 40114 6132 40124
rect 5404 38894 5406 38946
rect 5458 38894 5460 38946
rect 5404 37940 5460 38894
rect 5852 38836 5908 38846
rect 5852 38722 5908 38780
rect 5852 38670 5854 38722
rect 5906 38670 5908 38722
rect 5852 38668 5908 38670
rect 6188 38668 6244 50372
rect 6524 40402 6580 40414
rect 6524 40350 6526 40402
rect 6578 40350 6580 40402
rect 6412 39506 6468 39518
rect 6412 39454 6414 39506
rect 6466 39454 6468 39506
rect 6412 38668 6468 39454
rect 5292 36258 5348 36270
rect 5292 36206 5294 36258
rect 5346 36206 5348 36258
rect 5292 33908 5348 36206
rect 5404 35028 5460 37884
rect 5740 38612 5908 38668
rect 5964 38612 6244 38668
rect 6300 38612 6468 38668
rect 5628 37492 5684 37502
rect 5516 35698 5572 35710
rect 5516 35646 5518 35698
rect 5570 35646 5572 35698
rect 5516 35252 5572 35646
rect 5516 35186 5572 35196
rect 5404 34972 5572 35028
rect 5292 33842 5348 33852
rect 5404 34692 5460 34702
rect 5404 34132 5460 34636
rect 5068 32732 5236 32788
rect 5292 33572 5348 33582
rect 5068 31668 5124 32732
rect 5180 32564 5236 32574
rect 5292 32564 5348 33516
rect 5404 33348 5460 34076
rect 5516 33906 5572 34972
rect 5516 33854 5518 33906
rect 5570 33854 5572 33906
rect 5516 33572 5572 33854
rect 5516 33506 5572 33516
rect 5404 33346 5572 33348
rect 5404 33294 5406 33346
rect 5458 33294 5572 33346
rect 5404 33292 5572 33294
rect 5404 33282 5460 33292
rect 5180 32562 5348 32564
rect 5180 32510 5182 32562
rect 5234 32510 5348 32562
rect 5180 32508 5348 32510
rect 5180 32498 5236 32508
rect 5068 31666 5236 31668
rect 5068 31614 5070 31666
rect 5122 31614 5236 31666
rect 5068 31612 5236 31614
rect 5068 31602 5124 31612
rect 4284 30828 4900 30884
rect 4284 30436 4340 30828
rect 4956 30772 5012 30782
rect 4844 30770 5012 30772
rect 4844 30718 4958 30770
rect 5010 30718 5012 30770
rect 4844 30716 5012 30718
rect 4464 30604 4728 30614
rect 4520 30548 4568 30604
rect 4624 30548 4672 30604
rect 4464 30538 4728 30548
rect 4508 30436 4564 30446
rect 4844 30436 4900 30716
rect 4956 30706 5012 30716
rect 4284 30380 4452 30436
rect 4172 30258 4228 30268
rect 4284 30212 4340 30222
rect 4284 30118 4340 30156
rect 4060 30044 4228 30100
rect 3804 29820 4068 29830
rect 3860 29764 3908 29820
rect 3964 29764 4012 29820
rect 3804 29754 4068 29764
rect 4172 29316 4228 30044
rect 4284 29652 4340 29662
rect 4284 29558 4340 29596
rect 3612 28814 3614 28866
rect 3666 28814 3668 28866
rect 3612 28802 3668 28814
rect 4060 29260 4228 29316
rect 4060 28756 4116 29260
rect 4396 29204 4452 30380
rect 4508 30434 4900 30436
rect 4508 30382 4510 30434
rect 4562 30382 4900 30434
rect 4508 30380 4900 30382
rect 4508 30370 4564 30380
rect 4060 28690 4116 28700
rect 4172 29148 4452 29204
rect 4844 30212 4900 30222
rect 3804 28252 4068 28262
rect 3860 28196 3908 28252
rect 3964 28196 4012 28252
rect 3804 28186 4068 28196
rect 4172 28084 4228 29148
rect 4464 29036 4728 29046
rect 4520 28980 4568 29036
rect 4624 28980 4672 29036
rect 4464 28970 4728 28980
rect 4508 28756 4564 28766
rect 4508 28662 4564 28700
rect 3836 28028 4228 28084
rect 4284 28418 4340 28430
rect 4284 28366 4286 28418
rect 4338 28366 4340 28418
rect 3612 27074 3668 27086
rect 3612 27022 3614 27074
rect 3666 27022 3668 27074
rect 3612 26514 3668 27022
rect 3836 26852 3892 28028
rect 3948 27634 4004 27646
rect 3948 27582 3950 27634
rect 4002 27582 4004 27634
rect 3948 27076 4004 27582
rect 4284 27524 4340 28366
rect 4172 27468 4340 27524
rect 4464 27468 4728 27478
rect 3948 27010 4004 27020
rect 4060 27412 4116 27422
rect 4060 27074 4116 27356
rect 4060 27022 4062 27074
rect 4114 27022 4116 27074
rect 4060 27010 4116 27022
rect 4172 27076 4228 27468
rect 4520 27412 4568 27468
rect 4624 27412 4672 27468
rect 4464 27402 4728 27412
rect 4284 27300 4340 27310
rect 4284 27206 4340 27244
rect 4732 27076 4788 27086
rect 4172 27020 4452 27076
rect 3836 26796 4340 26852
rect 3804 26684 4068 26694
rect 3860 26628 3908 26684
rect 3964 26628 4012 26684
rect 3804 26618 4068 26628
rect 3612 26462 3614 26514
rect 3666 26462 3668 26514
rect 3612 26450 3668 26462
rect 3612 25732 3668 25742
rect 3612 25638 3668 25676
rect 4172 25506 4228 25518
rect 4172 25454 4174 25506
rect 4226 25454 4228 25506
rect 3804 25116 4068 25126
rect 3860 25060 3908 25116
rect 3964 25060 4012 25116
rect 3500 25004 3668 25060
rect 3804 25050 4068 25060
rect 3388 24836 3444 24892
rect 3164 23886 3166 23938
rect 3218 23886 3220 23938
rect 3164 22260 3220 23886
rect 3276 24780 3444 24836
rect 3500 24836 3556 24846
rect 3276 23828 3332 24780
rect 3500 24742 3556 24780
rect 3500 24388 3556 24398
rect 3388 24052 3444 24062
rect 3388 23958 3444 23996
rect 3276 23762 3332 23772
rect 3164 22194 3220 22204
rect 3500 22258 3556 24332
rect 3500 22206 3502 22258
rect 3554 22206 3556 22258
rect 3500 22194 3556 22206
rect 3164 21812 3220 21822
rect 3164 21474 3220 21756
rect 3164 21422 3166 21474
rect 3218 21422 3220 21474
rect 3164 21410 3220 21422
rect 3612 21140 3668 25004
rect 4172 24836 4228 25454
rect 4172 24770 4228 24780
rect 4060 23940 4116 23950
rect 4060 23938 4228 23940
rect 4060 23886 4062 23938
rect 4114 23886 4228 23938
rect 4060 23884 4228 23886
rect 4060 23874 4116 23884
rect 3804 23548 4068 23558
rect 3860 23492 3908 23548
rect 3964 23492 4012 23548
rect 3804 23482 4068 23492
rect 3836 23380 3892 23390
rect 4172 23380 4228 23884
rect 3836 23378 4228 23380
rect 3836 23326 3838 23378
rect 3890 23326 4228 23378
rect 3836 23324 4228 23326
rect 3836 23314 3892 23324
rect 4284 22370 4340 26796
rect 4396 26068 4452 27020
rect 4732 26982 4788 27020
rect 4396 26002 4452 26012
rect 4464 25900 4728 25910
rect 4520 25844 4568 25900
rect 4624 25844 4672 25900
rect 4464 25834 4728 25844
rect 4732 25506 4788 25518
rect 4732 25454 4734 25506
rect 4786 25454 4788 25506
rect 4732 24836 4788 25454
rect 4732 24770 4788 24780
rect 4844 24724 4900 30156
rect 4956 30210 5012 30222
rect 4956 30158 4958 30210
rect 5010 30158 5012 30210
rect 4956 29652 5012 30158
rect 4956 29586 5012 29596
rect 5068 29540 5124 29550
rect 5068 28642 5124 29484
rect 5068 28590 5070 28642
rect 5122 28590 5124 28642
rect 5068 28578 5124 28590
rect 5180 28420 5236 31612
rect 5292 30884 5348 32508
rect 5404 31778 5460 31790
rect 5404 31726 5406 31778
rect 5458 31726 5460 31778
rect 5404 31220 5460 31726
rect 5516 31556 5572 33292
rect 5516 31490 5572 31500
rect 5404 31154 5460 31164
rect 5516 31108 5572 31118
rect 5628 31108 5684 37436
rect 5516 31106 5684 31108
rect 5516 31054 5518 31106
rect 5570 31054 5684 31106
rect 5516 31052 5684 31054
rect 5516 31042 5572 31052
rect 5292 29428 5348 30828
rect 5628 30210 5684 30222
rect 5628 30158 5630 30210
rect 5682 30158 5684 30210
rect 5628 30100 5684 30158
rect 5628 30034 5684 30044
rect 5292 29362 5348 29372
rect 5628 29428 5684 29438
rect 5628 29334 5684 29372
rect 5180 28354 5236 28364
rect 5516 27746 5572 27758
rect 5516 27694 5518 27746
rect 5570 27694 5572 27746
rect 4956 27634 5012 27646
rect 4956 27582 4958 27634
rect 5010 27582 5012 27634
rect 4956 27300 5012 27582
rect 5516 27412 5572 27694
rect 5516 27346 5572 27356
rect 4956 27234 5012 27244
rect 5292 27076 5348 27086
rect 5292 26982 5348 27020
rect 5404 26964 5460 26974
rect 4956 26066 5012 26078
rect 4956 26014 4958 26066
rect 5010 26014 5012 26066
rect 4956 25732 5012 26014
rect 4956 25666 5012 25676
rect 5292 26068 5348 26078
rect 4956 24724 5012 24734
rect 4844 24722 5012 24724
rect 4844 24670 4958 24722
rect 5010 24670 5012 24722
rect 4844 24668 5012 24670
rect 4956 24658 5012 24668
rect 4464 24332 4728 24342
rect 4520 24276 4568 24332
rect 4624 24276 4672 24332
rect 4464 24266 4728 24276
rect 4620 23940 4676 23950
rect 4620 23846 4676 23884
rect 5068 23940 5124 23950
rect 4844 23604 4900 23614
rect 4464 22764 4728 22774
rect 4520 22708 4568 22764
rect 4624 22708 4672 22764
rect 4464 22698 4728 22708
rect 4284 22318 4286 22370
rect 4338 22318 4340 22370
rect 4284 22306 4340 22318
rect 3804 21980 4068 21990
rect 3860 21924 3908 21980
rect 3964 21924 4012 21980
rect 3804 21914 4068 21924
rect 3612 21074 3668 21084
rect 4172 21812 4228 21822
rect 3164 20916 3220 20926
rect 3164 20822 3220 20860
rect 3612 20802 3668 20814
rect 3612 20750 3614 20802
rect 3666 20750 3668 20802
rect 3612 20188 3668 20750
rect 3804 20412 4068 20422
rect 3860 20356 3908 20412
rect 3964 20356 4012 20412
rect 3804 20346 4068 20356
rect 3052 20132 3220 20188
rect 3052 19124 3108 19134
rect 3052 19030 3108 19068
rect 3164 18226 3220 20132
rect 3276 20132 3668 20188
rect 3276 20130 3332 20132
rect 3276 20078 3278 20130
rect 3330 20078 3332 20130
rect 3276 20066 3332 20078
rect 3164 18174 3166 18226
rect 3218 18174 3220 18226
rect 2940 17836 3108 17892
rect 2828 17054 2830 17106
rect 2882 17054 2884 17106
rect 2828 17042 2884 17054
rect 2940 17668 2996 17678
rect 2940 16322 2996 17612
rect 2940 16270 2942 16322
rect 2994 16270 2996 16322
rect 2940 16258 2996 16270
rect 2716 16212 2772 16222
rect 2604 15204 2660 15214
rect 2604 15110 2660 15148
rect 2604 12964 2660 12974
rect 2492 12962 2660 12964
rect 2492 12910 2606 12962
rect 2658 12910 2660 12962
rect 2492 12908 2660 12910
rect 2492 12068 2548 12908
rect 2604 12898 2660 12908
rect 2492 11974 2548 12012
rect 2604 12180 2660 12190
rect 2380 8754 2436 8764
rect 2492 11844 2548 11854
rect 2492 10498 2548 11788
rect 2604 11620 2660 12124
rect 2716 11956 2772 16156
rect 2716 11890 2772 11900
rect 2828 15764 2884 15774
rect 2716 11620 2772 11630
rect 2604 11618 2772 11620
rect 2604 11566 2718 11618
rect 2770 11566 2772 11618
rect 2604 11564 2772 11566
rect 2716 11554 2772 11564
rect 2492 10446 2494 10498
rect 2546 10446 2548 10498
rect 2492 10052 2548 10446
rect 2156 8428 2212 8438
rect 2492 8428 2548 9996
rect 2604 10724 2660 10734
rect 2604 8708 2660 10668
rect 2828 9714 2884 15708
rect 2828 9662 2830 9714
rect 2882 9662 2884 9714
rect 2828 9650 2884 9662
rect 2940 13076 2996 13086
rect 2604 8642 2660 8652
rect 2716 9492 2772 9502
rect 2492 8372 2660 8428
rect 1932 4946 1988 4956
rect 2044 6916 2100 6926
rect 1820 2258 1876 2268
rect 476 1586 532 1596
rect 252 466 308 476
rect 700 644 756 654
rect 700 112 756 588
rect 2044 112 2100 6860
rect 2156 6690 2212 8372
rect 2268 8260 2324 8270
rect 2268 8258 2436 8260
rect 2268 8206 2270 8258
rect 2322 8206 2436 8258
rect 2268 8204 2436 8206
rect 2268 8194 2324 8204
rect 2268 8036 2324 8046
rect 2268 7474 2324 7980
rect 2268 7422 2270 7474
rect 2322 7422 2324 7474
rect 2268 7410 2324 7422
rect 2380 6916 2436 8204
rect 2380 6850 2436 6860
rect 2156 6638 2158 6690
rect 2210 6638 2212 6690
rect 2156 6626 2212 6638
rect 2268 6132 2324 6142
rect 2268 5906 2324 6076
rect 2268 5854 2270 5906
rect 2322 5854 2324 5906
rect 2268 5842 2324 5854
rect 2604 5906 2660 8372
rect 2716 7700 2772 9436
rect 2940 9154 2996 13020
rect 3052 11508 3108 17836
rect 3164 15316 3220 18174
rect 3500 19346 3556 19358
rect 3500 19294 3502 19346
rect 3554 19294 3556 19346
rect 3500 18228 3556 19294
rect 3804 18844 4068 18854
rect 3860 18788 3908 18844
rect 3964 18788 4012 18844
rect 3804 18778 4068 18788
rect 3500 18162 3556 18172
rect 3948 18452 4004 18462
rect 3724 17892 3780 17902
rect 3724 17798 3780 17836
rect 3836 17780 3892 17790
rect 3164 15250 3220 15260
rect 3276 17666 3332 17678
rect 3276 17614 3278 17666
rect 3330 17614 3332 17666
rect 3276 14754 3332 17614
rect 3836 17666 3892 17724
rect 3836 17614 3838 17666
rect 3890 17614 3892 17666
rect 3836 17602 3892 17614
rect 3948 17444 4004 18396
rect 3612 17388 4004 17444
rect 3612 16996 3668 17388
rect 3804 17276 4068 17286
rect 3860 17220 3908 17276
rect 3964 17220 4012 17276
rect 3804 17210 4068 17220
rect 3724 16996 3780 17006
rect 3612 16994 3780 16996
rect 3612 16942 3726 16994
rect 3778 16942 3780 16994
rect 3612 16940 3780 16942
rect 3724 16930 3780 16940
rect 3388 16884 3444 16894
rect 3388 16790 3444 16828
rect 3836 16884 3892 16894
rect 3612 16212 3668 16222
rect 3612 16098 3668 16156
rect 3612 16046 3614 16098
rect 3666 16046 3668 16098
rect 3612 16034 3668 16046
rect 3276 14702 3278 14754
rect 3330 14702 3332 14754
rect 3276 14690 3332 14702
rect 3388 15876 3444 15886
rect 3836 15876 3892 16828
rect 4060 16212 4116 16222
rect 4060 16118 4116 16156
rect 3388 15204 3444 15820
rect 3388 14084 3444 15148
rect 3500 15820 3892 15876
rect 3500 14308 3556 15820
rect 3804 15708 4068 15718
rect 3860 15652 3908 15708
rect 3964 15652 4012 15708
rect 3804 15642 4068 15652
rect 4172 15540 4228 21756
rect 4284 21364 4340 21374
rect 4284 21270 4340 21308
rect 4464 21196 4728 21206
rect 4520 21140 4568 21196
rect 4624 21140 4672 21196
rect 4464 21130 4728 21140
rect 4396 20804 4452 20814
rect 4396 20710 4452 20748
rect 4464 19628 4728 19638
rect 4520 19572 4568 19628
rect 4624 19572 4672 19628
rect 4464 19562 4728 19572
rect 4620 19236 4676 19246
rect 4620 19142 4676 19180
rect 4844 18452 4900 23548
rect 4844 18386 4900 18396
rect 4956 21700 5012 21710
rect 4284 18226 4340 18238
rect 4284 18174 4286 18226
rect 4338 18174 4340 18226
rect 4284 17892 4340 18174
rect 4464 18060 4728 18070
rect 4520 18004 4568 18060
rect 4624 18004 4672 18060
rect 4464 17994 4728 18004
rect 4956 17892 5012 21644
rect 5068 19122 5124 23884
rect 5292 23828 5348 26012
rect 5404 23940 5460 26908
rect 5516 26180 5572 26190
rect 5516 26086 5572 26124
rect 5516 25620 5572 25630
rect 5516 24946 5572 25564
rect 5516 24894 5518 24946
rect 5570 24894 5572 24946
rect 5516 24882 5572 24894
rect 5628 25506 5684 25518
rect 5628 25454 5630 25506
rect 5682 25454 5684 25506
rect 5516 23940 5572 23950
rect 5404 23884 5516 23940
rect 5516 23846 5572 23884
rect 5292 23772 5460 23828
rect 5292 23156 5348 23166
rect 5180 23044 5236 23054
rect 5180 22950 5236 22988
rect 5292 22820 5348 23100
rect 5180 22764 5348 22820
rect 5180 22148 5236 22764
rect 5404 22260 5460 23772
rect 5628 23380 5684 25454
rect 5628 23314 5684 23324
rect 5740 23156 5796 38612
rect 5964 38500 6020 38612
rect 5852 38444 6020 38500
rect 5852 35140 5908 38444
rect 5964 38276 6020 38286
rect 5964 38182 6020 38220
rect 5964 36372 6020 36382
rect 5964 35810 6020 36316
rect 5964 35758 5966 35810
rect 6018 35758 6020 35810
rect 5964 35746 6020 35758
rect 5852 35084 6020 35140
rect 5852 34914 5908 34926
rect 5852 34862 5854 34914
rect 5906 34862 5908 34914
rect 5852 34692 5908 34862
rect 5852 34626 5908 34636
rect 5852 32900 5908 32910
rect 5852 32676 5908 32844
rect 5852 32582 5908 32620
rect 5852 31780 5908 31818
rect 5852 31714 5908 31724
rect 5740 23090 5796 23100
rect 5852 31556 5908 31566
rect 5180 22082 5236 22092
rect 5292 22204 5460 22260
rect 5516 22932 5572 22942
rect 5180 21476 5236 21486
rect 5180 20802 5236 21420
rect 5292 21364 5348 22204
rect 5404 21588 5460 21598
rect 5404 21494 5460 21532
rect 5292 21308 5460 21364
rect 5180 20750 5182 20802
rect 5234 20750 5236 20802
rect 5180 20738 5236 20750
rect 5292 21028 5348 21038
rect 5068 19070 5070 19122
rect 5122 19070 5124 19122
rect 5068 18788 5124 19070
rect 5068 18722 5124 18732
rect 5180 20018 5236 20030
rect 5180 19966 5182 20018
rect 5234 19966 5236 20018
rect 5068 18564 5124 18574
rect 5068 18470 5124 18508
rect 4284 17826 4340 17836
rect 4620 17836 5012 17892
rect 4284 17668 4340 17678
rect 4284 17574 4340 17612
rect 4620 16772 4676 17836
rect 5180 17780 5236 19966
rect 5292 18228 5348 20972
rect 5404 20020 5460 21308
rect 5516 20242 5572 22876
rect 5740 22930 5796 22942
rect 5740 22878 5742 22930
rect 5794 22878 5796 22930
rect 5628 22596 5684 22606
rect 5628 22372 5684 22540
rect 5628 22306 5684 22316
rect 5516 20190 5518 20242
rect 5570 20190 5572 20242
rect 5516 20178 5572 20190
rect 5628 22148 5684 22158
rect 5404 19964 5572 20020
rect 5404 19236 5460 19246
rect 5404 19142 5460 19180
rect 5516 19012 5572 19964
rect 5404 18956 5572 19012
rect 5404 18452 5460 18956
rect 5404 18386 5460 18396
rect 5516 18788 5572 18798
rect 5516 18450 5572 18732
rect 5516 18398 5518 18450
rect 5570 18398 5572 18450
rect 5516 18386 5572 18398
rect 5292 18172 5572 18228
rect 4956 17724 5236 17780
rect 4732 17668 4788 17678
rect 4732 17574 4788 17612
rect 4956 17332 5012 17724
rect 5404 17668 5460 17678
rect 5180 17666 5460 17668
rect 5180 17614 5406 17666
rect 5458 17614 5460 17666
rect 5180 17612 5460 17614
rect 5068 17556 5124 17566
rect 5068 17462 5124 17500
rect 4956 17276 5124 17332
rect 4956 16884 5012 16894
rect 4956 16790 5012 16828
rect 4620 16716 4788 16772
rect 4732 16660 4788 16716
rect 4732 16604 5012 16660
rect 4464 16492 4728 16502
rect 4520 16436 4568 16492
rect 4624 16436 4672 16492
rect 4464 16426 4728 16436
rect 3836 15484 4228 15540
rect 3836 15202 3892 15484
rect 4284 15428 4340 15438
rect 4284 15316 4340 15372
rect 3836 15150 3838 15202
rect 3890 15150 3892 15202
rect 3836 15138 3892 15150
rect 4060 15314 4340 15316
rect 4060 15262 4286 15314
rect 4338 15262 4340 15314
rect 4060 15260 4340 15262
rect 3948 14532 4004 14542
rect 3500 14242 3556 14252
rect 3612 14530 4004 14532
rect 3612 14478 3950 14530
rect 4002 14478 4004 14530
rect 3612 14476 4004 14478
rect 3388 14028 3556 14084
rect 3388 13636 3444 13646
rect 3388 13542 3444 13580
rect 3164 13076 3220 13086
rect 3164 12982 3220 13020
rect 3500 13074 3556 14028
rect 3612 13186 3668 14476
rect 3948 14466 4004 14476
rect 4060 14308 4116 15260
rect 4284 15250 4340 15260
rect 4284 15092 4340 15102
rect 4284 14642 4340 15036
rect 4464 14924 4728 14934
rect 4520 14868 4568 14924
rect 4624 14868 4672 14924
rect 4464 14858 4728 14868
rect 4284 14590 4286 14642
rect 4338 14590 4340 14642
rect 4284 14578 4340 14590
rect 4172 14532 4228 14542
rect 4172 14438 4228 14476
rect 4732 14308 4788 14318
rect 4060 14252 4228 14308
rect 3804 14140 4068 14150
rect 3860 14084 3908 14140
rect 3964 14084 4012 14140
rect 3804 14074 4068 14084
rect 3612 13134 3614 13186
rect 3666 13134 3668 13186
rect 3612 13122 3668 13134
rect 3724 13972 3780 13982
rect 3500 13022 3502 13074
rect 3554 13022 3556 13074
rect 3500 13010 3556 13022
rect 3724 12964 3780 13916
rect 3948 13972 4004 13982
rect 3948 13746 4004 13916
rect 3948 13694 3950 13746
rect 4002 13694 4004 13746
rect 3948 13682 4004 13694
rect 3612 12908 3780 12964
rect 4172 12962 4228 14252
rect 4732 14214 4788 14252
rect 4396 13972 4452 13982
rect 4396 13858 4452 13916
rect 4956 13860 5012 16604
rect 4396 13806 4398 13858
rect 4450 13806 4452 13858
rect 4396 13794 4452 13806
rect 4844 13804 5012 13860
rect 4464 13356 4728 13366
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4464 13290 4728 13300
rect 4620 13188 4676 13198
rect 4844 13188 4900 13804
rect 4956 13636 5012 13646
rect 4956 13542 5012 13580
rect 4956 13188 5012 13198
rect 4844 13132 4956 13188
rect 4620 13076 4676 13132
rect 4620 13074 4900 13076
rect 4620 13022 4622 13074
rect 4674 13022 4900 13074
rect 4620 13020 4900 13022
rect 4620 13010 4676 13020
rect 4172 12910 4174 12962
rect 4226 12910 4228 12962
rect 3612 12402 3668 12908
rect 4172 12898 4228 12910
rect 3804 12572 4068 12582
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 3804 12506 4068 12516
rect 3612 12350 3614 12402
rect 3666 12350 3668 12402
rect 3612 12338 3668 12350
rect 3724 12292 3780 12302
rect 3276 11732 3332 11742
rect 3052 11452 3220 11508
rect 2940 9102 2942 9154
rect 2994 9102 2996 9154
rect 2940 9090 2996 9102
rect 3052 11284 3108 11294
rect 3052 8370 3108 11228
rect 3164 10388 3220 11452
rect 3276 11394 3332 11676
rect 3724 11618 3780 12236
rect 3724 11566 3726 11618
rect 3778 11566 3780 11618
rect 3724 11554 3780 11566
rect 4172 11956 4228 11966
rect 3276 11342 3278 11394
rect 3330 11342 3332 11394
rect 3276 11284 3332 11342
rect 3276 11218 3332 11228
rect 3612 11508 3668 11518
rect 3164 10322 3220 10332
rect 3276 11060 3332 11070
rect 3276 8428 3332 11004
rect 3612 10834 3668 11452
rect 3804 11004 4068 11014
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 3804 10938 4068 10948
rect 3612 10782 3614 10834
rect 3666 10782 3668 10834
rect 3612 10770 3668 10782
rect 3836 9826 3892 9838
rect 3836 9774 3838 9826
rect 3890 9774 3892 9826
rect 3836 9716 3892 9774
rect 3836 9650 3892 9660
rect 3804 9436 4068 9446
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 3804 9370 4068 9380
rect 3836 9044 3892 9054
rect 4172 9044 4228 11900
rect 4464 11788 4728 11798
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4464 11722 4728 11732
rect 4284 11396 4340 11406
rect 4284 11302 4340 11340
rect 4464 10220 4728 10230
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4464 10154 4728 10164
rect 3836 9042 4228 9044
rect 3836 8990 3838 9042
rect 3890 8990 4228 9042
rect 3836 8988 4228 8990
rect 4844 9044 4900 13020
rect 4956 12292 5012 13132
rect 4956 12226 5012 12236
rect 5068 11508 5124 17276
rect 5180 16322 5236 17612
rect 5404 17602 5460 17612
rect 5404 17444 5460 17454
rect 5180 16270 5182 16322
rect 5234 16270 5236 16322
rect 5180 16258 5236 16270
rect 5292 16660 5348 16670
rect 5180 15428 5236 15438
rect 5180 14530 5236 15372
rect 5180 14478 5182 14530
rect 5234 14478 5236 14530
rect 5180 14466 5236 14478
rect 5292 12290 5348 16604
rect 5292 12238 5294 12290
rect 5346 12238 5348 12290
rect 5292 12226 5348 12238
rect 5068 11442 5124 11452
rect 5068 11284 5124 11294
rect 5068 11282 5236 11284
rect 5068 11230 5070 11282
rect 5122 11230 5236 11282
rect 5068 11228 5236 11230
rect 5068 11218 5124 11228
rect 5180 10836 5236 11228
rect 5180 10724 5236 10780
rect 4956 10722 5236 10724
rect 4956 10670 5182 10722
rect 5234 10670 5236 10722
rect 4956 10668 5236 10670
rect 4956 9826 5012 10668
rect 5180 10658 5236 10668
rect 5404 10276 5460 17388
rect 5516 17106 5572 18172
rect 5516 17054 5518 17106
rect 5570 17054 5572 17106
rect 5516 17042 5572 17054
rect 5516 16324 5572 16334
rect 5516 13970 5572 16268
rect 5628 15202 5684 22092
rect 5740 22036 5796 22878
rect 5740 21970 5796 21980
rect 5852 20804 5908 31500
rect 5964 31220 6020 35084
rect 6188 34020 6244 34030
rect 5964 31154 6020 31164
rect 6076 31890 6132 31902
rect 6076 31838 6078 31890
rect 6130 31838 6132 31890
rect 5964 30996 6020 31006
rect 6076 30996 6132 31838
rect 5964 30994 6132 30996
rect 5964 30942 5966 30994
rect 6018 30942 6132 30994
rect 5964 30940 6132 30942
rect 5964 30930 6020 30940
rect 5740 20748 5908 20804
rect 5964 30548 6020 30558
rect 5964 27636 6020 30492
rect 5740 19012 5796 20748
rect 5852 20580 5908 20590
rect 5852 20486 5908 20524
rect 5964 20356 6020 27580
rect 6076 30324 6132 30334
rect 6076 29314 6132 30268
rect 6076 29262 6078 29314
rect 6130 29262 6132 29314
rect 6076 23268 6132 29262
rect 6188 23826 6244 33964
rect 6300 33572 6356 38612
rect 6524 38276 6580 40350
rect 6524 38210 6580 38220
rect 6636 39508 6692 39518
rect 6636 38948 6692 39452
rect 6636 38050 6692 38892
rect 6636 37998 6638 38050
rect 6690 37998 6692 38050
rect 6636 37986 6692 37998
rect 6524 37380 6580 37390
rect 6524 37286 6580 37324
rect 6412 36708 6468 36718
rect 6412 36614 6468 36652
rect 6524 36484 6580 36494
rect 6524 35810 6580 36428
rect 6524 35758 6526 35810
rect 6578 35758 6580 35810
rect 6524 34914 6580 35758
rect 6524 34862 6526 34914
rect 6578 34862 6580 34914
rect 6524 34850 6580 34862
rect 6636 33906 6692 33918
rect 6636 33854 6638 33906
rect 6690 33854 6692 33906
rect 6636 33684 6692 33854
rect 6636 33618 6692 33628
rect 6300 33506 6356 33516
rect 6524 33122 6580 33134
rect 6524 33070 6526 33122
rect 6578 33070 6580 33122
rect 6524 31668 6580 33070
rect 6524 31602 6580 31612
rect 6636 31778 6692 31790
rect 6636 31726 6638 31778
rect 6690 31726 6692 31778
rect 6412 31556 6468 31566
rect 6300 31220 6356 31230
rect 6300 30324 6356 31164
rect 6412 31106 6468 31500
rect 6412 31054 6414 31106
rect 6466 31054 6468 31106
rect 6412 31042 6468 31054
rect 6300 30258 6356 30268
rect 6524 30884 6580 30894
rect 6524 30210 6580 30828
rect 6524 30158 6526 30210
rect 6578 30158 6580 30210
rect 6524 30146 6580 30158
rect 6524 29876 6580 29886
rect 6412 27748 6468 27758
rect 6188 23774 6190 23826
rect 6242 23774 6244 23826
rect 6188 23492 6244 23774
rect 6188 23426 6244 23436
rect 6300 27746 6468 27748
rect 6300 27694 6414 27746
rect 6466 27694 6468 27746
rect 6300 27692 6468 27694
rect 6076 23212 6244 23268
rect 6076 23042 6132 23054
rect 6076 22990 6078 23042
rect 6130 22990 6132 23042
rect 6076 22820 6132 22990
rect 6076 22754 6132 22764
rect 6076 22482 6132 22494
rect 6076 22430 6078 22482
rect 6130 22430 6132 22482
rect 6076 22148 6132 22430
rect 6076 22082 6132 22092
rect 6188 21028 6244 23212
rect 6300 21812 6356 27692
rect 6412 27682 6468 27692
rect 6412 27076 6468 27086
rect 6412 26982 6468 27020
rect 6412 26292 6468 26302
rect 6524 26292 6580 29820
rect 6636 29652 6692 31726
rect 6636 29586 6692 29596
rect 6636 28644 6692 28654
rect 6636 27858 6692 28588
rect 6636 27806 6638 27858
rect 6690 27806 6692 27858
rect 6636 27794 6692 27806
rect 6748 26908 6804 54012
rect 6860 50484 6916 50494
rect 6860 45220 6916 50428
rect 6860 45154 6916 45164
rect 7644 47236 7700 47246
rect 6860 40402 6916 40414
rect 6860 40350 6862 40402
rect 6914 40350 6916 40402
rect 6860 39060 6916 40350
rect 7532 40292 7588 40302
rect 7196 40290 7588 40292
rect 7196 40238 7534 40290
rect 7586 40238 7588 40290
rect 7196 40236 7588 40238
rect 7084 40180 7140 40190
rect 6972 40178 7140 40180
rect 6972 40126 7086 40178
rect 7138 40126 7140 40178
rect 6972 40124 7140 40126
rect 6972 39842 7028 40124
rect 7084 40114 7140 40124
rect 6972 39790 6974 39842
rect 7026 39790 7028 39842
rect 6972 39778 7028 39790
rect 7196 39508 7252 40236
rect 7532 40226 7588 40236
rect 7644 40068 7700 47180
rect 7420 40012 7700 40068
rect 7756 40852 7812 40862
rect 7308 39732 7364 39742
rect 7308 39638 7364 39676
rect 6860 38994 6916 39004
rect 6972 39452 7252 39508
rect 6972 39058 7028 39452
rect 6972 39006 6974 39058
rect 7026 39006 7028 39058
rect 6972 38994 7028 39006
rect 6860 38724 6916 38734
rect 6860 36596 6916 38668
rect 7420 38668 7476 40012
rect 7756 39618 7812 40796
rect 7756 39566 7758 39618
rect 7810 39566 7812 39618
rect 7756 39508 7812 39566
rect 7644 39452 7812 39508
rect 7420 38612 7588 38668
rect 6972 38162 7028 38174
rect 6972 38110 6974 38162
rect 7026 38110 7028 38162
rect 6972 37716 7028 38110
rect 6972 37154 7028 37660
rect 6972 37102 6974 37154
rect 7026 37102 7028 37154
rect 6972 37090 7028 37102
rect 6860 36540 7028 36596
rect 6860 36370 6916 36382
rect 6860 36318 6862 36370
rect 6914 36318 6916 36370
rect 6860 36260 6916 36318
rect 6860 36194 6916 36204
rect 6972 36036 7028 36540
rect 6860 35980 7028 36036
rect 7420 36370 7476 36382
rect 7420 36318 7422 36370
rect 7474 36318 7476 36370
rect 6860 28420 6916 35980
rect 6972 35474 7028 35486
rect 6972 35422 6974 35474
rect 7026 35422 7028 35474
rect 6972 33460 7028 35422
rect 7084 35252 7140 35262
rect 7084 35028 7140 35196
rect 7084 34934 7140 34972
rect 6972 33394 7028 33404
rect 7196 32562 7252 32574
rect 7196 32510 7198 32562
rect 7250 32510 7252 32562
rect 7084 31778 7140 31790
rect 7084 31726 7086 31778
rect 7138 31726 7140 31778
rect 7084 31332 7140 31726
rect 7084 31266 7140 31276
rect 6972 30996 7028 31006
rect 7196 30996 7252 32510
rect 7420 31556 7476 36318
rect 7532 32676 7588 38612
rect 7644 36820 7700 39452
rect 7756 39172 7812 39182
rect 7756 36932 7812 39116
rect 7868 37828 7924 56030
rect 9212 55972 9268 55982
rect 8540 46116 8596 46126
rect 8316 42756 8372 42766
rect 8316 40628 8372 42700
rect 8316 40572 8484 40628
rect 8316 40402 8372 40414
rect 8316 40350 8318 40402
rect 8370 40350 8372 40402
rect 7980 40180 8036 40190
rect 7980 38946 8036 40124
rect 8316 39172 8372 40350
rect 8316 39106 8372 39116
rect 7980 38894 7982 38946
rect 8034 38894 8036 38946
rect 7980 38882 8036 38894
rect 8092 38892 8260 38948
rect 7868 37762 7924 37772
rect 8092 37490 8148 38892
rect 8204 38836 8260 38892
rect 8316 38836 8372 38846
rect 8204 38834 8372 38836
rect 8204 38782 8318 38834
rect 8370 38782 8372 38834
rect 8204 38780 8372 38782
rect 8316 38770 8372 38780
rect 8428 38668 8484 40572
rect 8204 38612 8260 38622
rect 8204 38274 8260 38556
rect 8204 38222 8206 38274
rect 8258 38222 8260 38274
rect 8204 38210 8260 38222
rect 8316 38612 8484 38668
rect 8092 37438 8094 37490
rect 8146 37438 8148 37490
rect 8092 37426 8148 37438
rect 7756 36876 8036 36932
rect 7644 36764 7924 36820
rect 7868 36484 7924 36764
rect 7868 36390 7924 36428
rect 7868 36260 7924 36270
rect 7756 35028 7812 35038
rect 7756 33906 7812 34972
rect 7868 34020 7924 36204
rect 7868 33954 7924 33964
rect 7756 33854 7758 33906
rect 7810 33854 7812 33906
rect 7644 33460 7700 33470
rect 7644 33366 7700 33404
rect 7532 32610 7588 32620
rect 7644 32450 7700 32462
rect 7644 32398 7646 32450
rect 7698 32398 7700 32450
rect 7644 32004 7700 32398
rect 7644 31938 7700 31948
rect 7420 31500 7588 31556
rect 7420 31332 7476 31342
rect 6972 30994 7252 30996
rect 6972 30942 6974 30994
rect 7026 30942 7252 30994
rect 6972 30940 7252 30942
rect 7308 31220 7364 31230
rect 6972 29876 7028 30940
rect 7308 30882 7364 31164
rect 7308 30830 7310 30882
rect 7362 30830 7364 30882
rect 7308 30818 7364 30830
rect 7420 30548 7476 31276
rect 7420 30482 7476 30492
rect 6972 29810 7028 29820
rect 7084 30210 7140 30222
rect 7084 30158 7086 30210
rect 7138 30158 7140 30210
rect 7084 29540 7140 30158
rect 7308 30212 7364 30222
rect 7196 29652 7252 29662
rect 7196 29558 7252 29596
rect 7084 29474 7140 29484
rect 7308 28644 7364 30156
rect 7532 29764 7588 31500
rect 7644 29986 7700 29998
rect 7644 29934 7646 29986
rect 7698 29934 7700 29986
rect 7644 29876 7700 29934
rect 7644 29810 7700 29820
rect 7532 29698 7588 29708
rect 7308 28550 7364 28588
rect 7420 28532 7476 28542
rect 6860 28364 7364 28420
rect 7084 28084 7140 28094
rect 6748 26852 6916 26908
rect 6412 26290 6580 26292
rect 6412 26238 6414 26290
rect 6466 26238 6580 26290
rect 6412 26236 6580 26238
rect 6412 26226 6468 26236
rect 6524 25506 6580 26236
rect 6748 26404 6804 26414
rect 6748 26180 6804 26348
rect 6524 25454 6526 25506
rect 6578 25454 6580 25506
rect 6524 25442 6580 25454
rect 6636 26178 6804 26180
rect 6636 26126 6750 26178
rect 6802 26126 6804 26178
rect 6636 26124 6804 26126
rect 6636 24162 6692 26124
rect 6748 26114 6804 26124
rect 6636 24110 6638 24162
rect 6690 24110 6692 24162
rect 6636 24098 6692 24110
rect 6748 23940 6804 23950
rect 6412 23492 6468 23502
rect 6412 22820 6468 23436
rect 6412 22754 6468 22764
rect 6300 21756 6468 21812
rect 6188 20972 6356 21028
rect 5852 20300 6020 20356
rect 5852 19234 5908 20300
rect 6188 20132 6244 20142
rect 6076 19348 6132 19358
rect 5852 19182 5854 19234
rect 5906 19182 5908 19234
rect 5852 19170 5908 19182
rect 5964 19346 6132 19348
rect 5964 19294 6078 19346
rect 6130 19294 6132 19346
rect 5964 19292 6132 19294
rect 5740 18946 5796 18956
rect 5964 18788 6020 19292
rect 6076 19282 6132 19292
rect 5964 18722 6020 18732
rect 6076 18676 6132 18686
rect 6188 18676 6244 20076
rect 6132 18620 6244 18676
rect 6076 18562 6132 18620
rect 6076 18510 6078 18562
rect 6130 18510 6132 18562
rect 6076 18498 6132 18510
rect 6188 18452 6244 18462
rect 5964 18116 6020 18126
rect 5852 17780 5908 17790
rect 5964 17780 6020 18060
rect 5908 17724 6020 17780
rect 5852 17714 5908 17724
rect 5964 17666 6020 17724
rect 6076 17780 6132 17790
rect 6076 17686 6132 17724
rect 5964 17614 5966 17666
rect 6018 17614 6020 17666
rect 5964 17602 6020 17614
rect 5852 17556 5908 17566
rect 5852 17220 5908 17500
rect 5852 17154 5908 17164
rect 6188 16548 6244 18396
rect 6188 16482 6244 16492
rect 5964 16212 6020 16222
rect 5964 16210 6132 16212
rect 5964 16158 5966 16210
rect 6018 16158 6132 16210
rect 5964 16156 6132 16158
rect 5964 16146 6020 16156
rect 5852 16098 5908 16110
rect 5852 16046 5854 16098
rect 5906 16046 5908 16098
rect 5852 15876 5908 16046
rect 5852 15810 5908 15820
rect 5628 15150 5630 15202
rect 5682 15150 5684 15202
rect 5628 15138 5684 15150
rect 5740 15316 5796 15326
rect 5740 14754 5796 15260
rect 5740 14702 5742 14754
rect 5794 14702 5796 14754
rect 5740 14690 5796 14702
rect 5516 13918 5518 13970
rect 5570 13918 5572 13970
rect 5516 13906 5572 13918
rect 5852 13524 5908 13534
rect 5740 12852 5796 12862
rect 5740 12758 5796 12796
rect 5516 12180 5572 12190
rect 5516 11844 5572 12124
rect 5516 11618 5572 11788
rect 5516 11566 5518 11618
rect 5570 11566 5572 11618
rect 5516 11554 5572 11566
rect 5628 12068 5684 12078
rect 5628 10498 5684 12012
rect 5628 10446 5630 10498
rect 5682 10446 5684 10498
rect 5628 10434 5684 10446
rect 5852 10276 5908 13468
rect 6076 12404 6132 16156
rect 6188 16098 6244 16110
rect 6188 16046 6190 16098
rect 6242 16046 6244 16098
rect 6188 14868 6244 16046
rect 6188 14802 6244 14812
rect 6076 12348 6244 12404
rect 6076 12178 6132 12190
rect 6076 12126 6078 12178
rect 6130 12126 6132 12178
rect 4956 9774 4958 9826
rect 5010 9774 5012 9826
rect 4956 9762 5012 9774
rect 5292 10220 5460 10276
rect 5516 10220 5908 10276
rect 5964 11844 6020 11854
rect 4956 9044 5012 9054
rect 4844 9042 5012 9044
rect 4844 8990 4958 9042
rect 5010 8990 5012 9042
rect 4844 8988 5012 8990
rect 3836 8978 3892 8988
rect 4956 8978 5012 8988
rect 4464 8652 4728 8662
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4464 8586 4728 8596
rect 3052 8318 3054 8370
rect 3106 8318 3108 8370
rect 3052 8306 3108 8318
rect 3164 8372 3332 8428
rect 2828 7700 2884 7710
rect 2716 7698 2884 7700
rect 2716 7646 2830 7698
rect 2882 7646 2884 7698
rect 2716 7644 2884 7646
rect 2828 7634 2884 7644
rect 3164 6804 3220 8372
rect 2940 6748 3220 6804
rect 3612 8260 3668 8270
rect 2604 5854 2606 5906
rect 2658 5854 2660 5906
rect 2604 5842 2660 5854
rect 2828 6466 2884 6478
rect 2828 6414 2830 6466
rect 2882 6414 2884 6466
rect 2828 5908 2884 6414
rect 2828 5842 2884 5852
rect 2268 5236 2324 5246
rect 2940 5236 2996 6748
rect 3612 6690 3668 8204
rect 3836 8258 3892 8270
rect 3836 8206 3838 8258
rect 3890 8206 3892 8258
rect 3836 8148 3892 8206
rect 3836 8082 3892 8092
rect 5068 8036 5124 8046
rect 5068 7942 5124 7980
rect 3804 7868 4068 7878
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 3804 7802 4068 7812
rect 3836 7476 3892 7486
rect 3836 7382 3892 7420
rect 4464 7084 4728 7094
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4464 7018 4728 7028
rect 3612 6638 3614 6690
rect 3666 6638 3668 6690
rect 3612 6626 3668 6638
rect 2268 5234 2996 5236
rect 2268 5182 2270 5234
rect 2322 5182 2996 5234
rect 2268 5180 2996 5182
rect 3052 6468 3108 6478
rect 3052 5234 3108 6412
rect 3804 6300 4068 6310
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 3804 6234 4068 6244
rect 3164 6020 3220 6030
rect 3164 5926 3220 5964
rect 4464 5516 4728 5526
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4464 5450 4728 5460
rect 3612 5348 3668 5358
rect 3612 5254 3668 5292
rect 3052 5182 3054 5234
rect 3106 5182 3108 5234
rect 2268 5170 2324 5180
rect 3052 5170 3108 5182
rect 3804 4732 4068 4742
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 3804 4666 4068 4676
rect 2268 4228 2324 4238
rect 2268 4134 2324 4172
rect 4464 3948 4728 3958
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4464 3882 4728 3892
rect 2268 3556 2324 3566
rect 2268 3462 2324 3500
rect 3804 3164 4068 3174
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 3804 3098 4068 3108
rect 4464 2380 4728 2390
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4464 2314 4728 2324
rect 3388 1652 3444 1662
rect 3388 112 3444 1596
rect 3804 1596 4068 1606
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 3804 1530 4068 1540
rect 4464 812 4728 822
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4464 746 4728 756
rect 4732 532 4788 542
rect 4732 112 4788 476
rect 672 0 784 112
rect 2016 0 2128 112
rect 3360 0 3472 112
rect 4704 0 4816 112
rect 5292 84 5348 10220
rect 5404 10052 5460 10062
rect 5404 9958 5460 9996
rect 5516 9154 5572 10220
rect 5516 9102 5518 9154
rect 5570 9102 5572 9154
rect 5516 9090 5572 9102
rect 5964 9042 6020 11788
rect 5964 8990 5966 9042
rect 6018 8990 6020 9042
rect 5964 8978 6020 8990
rect 6076 6804 6132 12126
rect 6188 10276 6244 12348
rect 6300 11844 6356 20972
rect 6412 17444 6468 21756
rect 6524 21586 6580 21598
rect 6524 21534 6526 21586
rect 6578 21534 6580 21586
rect 6524 20804 6580 21534
rect 6748 21252 6804 23884
rect 6748 21186 6804 21196
rect 6580 20748 6804 20804
rect 6524 20738 6580 20748
rect 6524 20580 6580 20590
rect 6524 19346 6580 20524
rect 6748 19684 6804 20748
rect 6748 19618 6804 19628
rect 6524 19294 6526 19346
rect 6578 19294 6580 19346
rect 6524 19282 6580 19294
rect 6524 18340 6580 18350
rect 6580 18284 6692 18340
rect 6524 18246 6580 18284
rect 6524 17892 6580 17902
rect 6524 17778 6580 17836
rect 6524 17726 6526 17778
rect 6578 17726 6580 17778
rect 6524 17714 6580 17726
rect 6412 17378 6468 17388
rect 6412 16772 6468 16782
rect 6412 15652 6468 16716
rect 6636 16772 6692 18284
rect 6860 16884 6916 26852
rect 7084 25732 7140 28028
rect 7084 25638 7140 25676
rect 6972 24612 7028 24622
rect 6972 24276 7028 24556
rect 6972 24210 7028 24220
rect 7196 24164 7252 24174
rect 7084 23716 7140 23726
rect 6972 23268 7028 23278
rect 6972 23174 7028 23212
rect 6972 21700 7028 21710
rect 6972 21026 7028 21644
rect 7084 21586 7140 23660
rect 7196 23492 7252 24108
rect 7196 23426 7252 23436
rect 7084 21534 7086 21586
rect 7138 21534 7140 21586
rect 7084 21522 7140 21534
rect 7196 22146 7252 22158
rect 7196 22094 7198 22146
rect 7250 22094 7252 22146
rect 6972 20974 6974 21026
rect 7026 20974 7028 21026
rect 6972 20962 7028 20974
rect 7084 21252 7140 21262
rect 6972 19906 7028 19918
rect 6972 19854 6974 19906
rect 7026 19854 7028 19906
rect 6972 19684 7028 19854
rect 6972 19618 7028 19628
rect 7084 19234 7140 21196
rect 7196 20692 7252 22094
rect 7308 21588 7364 28364
rect 7420 28082 7476 28476
rect 7420 28030 7422 28082
rect 7474 28030 7476 28082
rect 7420 28018 7476 28030
rect 7532 28420 7588 28430
rect 7420 27860 7476 27870
rect 7420 27188 7476 27804
rect 7420 26404 7476 27132
rect 7420 26338 7476 26348
rect 7420 26068 7476 26078
rect 7420 24722 7476 26012
rect 7420 24670 7422 24722
rect 7474 24670 7476 24722
rect 7420 24658 7476 24670
rect 7532 23156 7588 28364
rect 7756 28084 7812 33854
rect 7980 33684 8036 36876
rect 8092 35474 8148 35486
rect 8092 35422 8094 35474
rect 8146 35422 8148 35474
rect 8092 34132 8148 35422
rect 8204 34692 8260 34702
rect 8204 34598 8260 34636
rect 8092 34066 8148 34076
rect 8204 34130 8260 34142
rect 8204 34078 8206 34130
rect 8258 34078 8260 34130
rect 8204 34020 8260 34078
rect 8204 33954 8260 33964
rect 7980 33628 8260 33684
rect 7980 33460 8036 33470
rect 7756 28018 7812 28028
rect 7868 31108 7924 31118
rect 7868 30100 7924 31052
rect 7868 27860 7924 30044
rect 7756 27804 7924 27860
rect 7980 27860 8036 33404
rect 7756 26908 7812 27804
rect 7980 27794 8036 27804
rect 8092 33236 8148 33246
rect 8092 32228 8148 33180
rect 8092 28418 8148 32172
rect 8092 28366 8094 28418
rect 8146 28366 8148 28418
rect 7868 27188 7924 27198
rect 7868 27074 7924 27132
rect 7868 27022 7870 27074
rect 7922 27022 7924 27074
rect 7868 27010 7924 27022
rect 8092 27188 8148 28366
rect 8204 31778 8260 33628
rect 8204 31726 8206 31778
rect 8258 31726 8260 31778
rect 8204 28308 8260 31726
rect 8316 29988 8372 38612
rect 8316 29922 8372 29932
rect 8428 34916 8484 34926
rect 8204 28242 8260 28252
rect 8316 29652 8372 29662
rect 8204 27972 8260 27982
rect 8204 27878 8260 27916
rect 7644 26852 7812 26908
rect 7644 24948 7700 26852
rect 7980 26068 8036 26078
rect 7980 25974 8036 26012
rect 7644 24724 7700 24892
rect 7756 24724 7812 24734
rect 7644 24722 7812 24724
rect 7644 24670 7758 24722
rect 7810 24670 7812 24722
rect 7644 24668 7812 24670
rect 7756 24658 7812 24668
rect 7980 24612 8036 24622
rect 7980 24518 8036 24556
rect 7756 23716 7812 23726
rect 7756 23622 7812 23660
rect 8092 23548 8148 27132
rect 8316 27186 8372 29596
rect 8428 29316 8484 34860
rect 8540 31108 8596 46060
rect 8764 45332 8820 45342
rect 8764 38724 8820 45276
rect 9212 41188 9268 55916
rect 9996 55970 10052 55982
rect 9996 55918 9998 55970
rect 10050 55918 10052 55970
rect 9212 41122 9268 41132
rect 9884 41748 9940 41758
rect 9772 41076 9828 41086
rect 8988 40964 9044 40974
rect 8988 40962 9492 40964
rect 8988 40910 8990 40962
rect 9042 40910 9492 40962
rect 8988 40908 9492 40910
rect 8988 40898 9044 40908
rect 9212 40402 9268 40414
rect 9212 40350 9214 40402
rect 9266 40350 9268 40402
rect 9100 40292 9156 40302
rect 8988 39618 9044 39630
rect 8988 39566 8990 39618
rect 9042 39566 9044 39618
rect 8876 39060 8932 39070
rect 8876 38846 8932 39004
rect 8876 38794 8878 38846
rect 8930 38794 8932 38846
rect 8876 38782 8932 38794
rect 8764 38668 8932 38724
rect 8652 37268 8708 37278
rect 8652 35698 8708 37212
rect 8652 35646 8654 35698
rect 8706 35646 8708 35698
rect 8652 35634 8708 35646
rect 8764 34018 8820 34030
rect 8764 33966 8766 34018
rect 8818 33966 8820 34018
rect 8652 33460 8708 33470
rect 8652 32900 8708 33404
rect 8652 32834 8708 32844
rect 8540 31052 8708 31108
rect 8540 30770 8596 30782
rect 8540 30718 8542 30770
rect 8594 30718 8596 30770
rect 8540 30100 8596 30718
rect 8540 30034 8596 30044
rect 8540 29540 8596 29550
rect 8540 29446 8596 29484
rect 8428 29260 8596 29316
rect 8316 27134 8318 27186
rect 8370 27134 8372 27186
rect 8316 27122 8372 27134
rect 8204 25284 8260 25294
rect 8204 25282 8372 25284
rect 8204 25230 8206 25282
rect 8258 25230 8372 25282
rect 8204 25228 8372 25230
rect 8204 25218 8260 25228
rect 8316 24724 8372 25228
rect 8428 24724 8484 24734
rect 8316 24722 8484 24724
rect 8316 24670 8430 24722
rect 8482 24670 8484 24722
rect 8316 24668 8484 24670
rect 8428 24658 8484 24668
rect 7980 23492 8148 23548
rect 8204 23940 8260 23950
rect 7532 23100 7700 23156
rect 7532 22036 7588 22046
rect 7308 21532 7476 21588
rect 7196 20626 7252 20636
rect 7308 21364 7364 21374
rect 7308 20018 7364 21308
rect 7420 20916 7476 21532
rect 7532 21474 7588 21980
rect 7644 21588 7700 23100
rect 7756 22932 7812 22942
rect 7756 22838 7812 22876
rect 7756 21588 7812 21598
rect 7644 21586 7924 21588
rect 7644 21534 7758 21586
rect 7810 21534 7924 21586
rect 7644 21532 7924 21534
rect 7756 21522 7812 21532
rect 7532 21422 7534 21474
rect 7586 21422 7588 21474
rect 7532 21410 7588 21422
rect 7420 20860 7588 20916
rect 7308 19966 7310 20018
rect 7362 19966 7364 20018
rect 7308 19954 7364 19966
rect 7420 20690 7476 20702
rect 7420 20638 7422 20690
rect 7474 20638 7476 20690
rect 7084 19182 7086 19234
rect 7138 19182 7140 19234
rect 7084 19170 7140 19182
rect 7308 19236 7364 19246
rect 7308 19142 7364 19180
rect 7420 19124 7476 20638
rect 7420 19058 7476 19068
rect 7532 18228 7588 20860
rect 7868 20020 7924 21532
rect 7980 20132 8036 23492
rect 8092 22932 8148 22942
rect 8092 21586 8148 22876
rect 8092 21534 8094 21586
rect 8146 21534 8148 21586
rect 8092 21522 8148 21534
rect 7980 20066 8036 20076
rect 7868 19926 7924 19964
rect 7980 19908 8036 19918
rect 7980 19814 8036 19852
rect 8204 19796 8260 23884
rect 8540 21700 8596 29260
rect 8652 27746 8708 31052
rect 8652 27694 8654 27746
rect 8706 27694 8708 27746
rect 8652 25732 8708 27694
rect 8652 25666 8708 25676
rect 8540 21644 8708 21700
rect 8540 21476 8596 21486
rect 8540 21382 8596 21420
rect 8092 19740 8260 19796
rect 8316 21140 8372 21150
rect 8092 19684 8148 19740
rect 7644 19628 8148 19684
rect 7644 18450 7700 19628
rect 8204 19572 8260 19582
rect 7644 18398 7646 18450
rect 7698 18398 7700 18450
rect 7644 18386 7700 18398
rect 7868 19236 7924 19246
rect 6636 16706 6692 16716
rect 6748 16828 6916 16884
rect 7084 18172 7588 18228
rect 6636 16548 6692 16558
rect 6636 15988 6692 16492
rect 6636 15894 6692 15932
rect 6412 15586 6468 15596
rect 6748 15540 6804 16828
rect 6636 15484 6804 15540
rect 6860 16658 6916 16670
rect 6860 16606 6862 16658
rect 6914 16606 6916 16658
rect 6412 14756 6468 14766
rect 6412 12850 6468 14700
rect 6636 13524 6692 15484
rect 6748 15316 6804 15354
rect 6748 15250 6804 15260
rect 6860 15148 6916 16606
rect 7084 16324 7140 18172
rect 7308 18004 7364 18014
rect 7308 17668 7364 17948
rect 7308 17574 7364 17612
rect 7532 17444 7588 17454
rect 7532 16996 7588 17388
rect 7532 16930 7588 16940
rect 7756 16996 7812 17006
rect 7084 16230 7140 16268
rect 7532 15876 7588 15886
rect 7084 15316 7140 15326
rect 7084 15222 7140 15260
rect 7532 15314 7588 15820
rect 7532 15262 7534 15314
rect 7586 15262 7588 15314
rect 6636 13458 6692 13468
rect 6748 15092 6916 15148
rect 6412 12798 6414 12850
rect 6466 12798 6468 12850
rect 6412 12786 6468 12798
rect 6300 11778 6356 11788
rect 6636 12178 6692 12190
rect 6636 12126 6638 12178
rect 6690 12126 6692 12178
rect 6524 11732 6580 11742
rect 6524 10612 6580 11676
rect 6636 11620 6692 12126
rect 6748 11956 6804 15092
rect 7084 14980 7140 14990
rect 6860 14644 6916 14654
rect 6860 14550 6916 14588
rect 6972 13748 7028 13758
rect 6972 12404 7028 13692
rect 6972 12338 7028 12348
rect 7084 12180 7140 14924
rect 7532 14532 7588 15262
rect 7756 15314 7812 16940
rect 7756 15262 7758 15314
rect 7810 15262 7812 15314
rect 7756 15204 7812 15262
rect 7756 15138 7812 15148
rect 7868 15148 7924 19180
rect 8204 19234 8260 19516
rect 8204 19182 8206 19234
rect 8258 19182 8260 19234
rect 8204 19170 8260 19182
rect 8316 18676 8372 21084
rect 8428 20692 8484 20702
rect 8428 20018 8484 20636
rect 8428 19966 8430 20018
rect 8482 19966 8484 20018
rect 8428 19954 8484 19966
rect 8092 18620 8372 18676
rect 7980 18340 8036 18350
rect 7980 16770 8036 18284
rect 7980 16718 7982 16770
rect 8034 16718 8036 16770
rect 7980 16706 8036 16718
rect 8092 15540 8148 18620
rect 8316 18450 8372 18462
rect 8316 18398 8318 18450
rect 8370 18398 8372 18450
rect 8204 17668 8260 17678
rect 8204 17574 8260 17612
rect 8204 16884 8260 16894
rect 8204 16322 8260 16828
rect 8204 16270 8206 16322
rect 8258 16270 8260 16322
rect 8204 16258 8260 16270
rect 8092 15474 8148 15484
rect 8204 15988 8260 15998
rect 8204 15314 8260 15932
rect 8316 15540 8372 18398
rect 8652 18004 8708 21644
rect 8764 20132 8820 33966
rect 8876 33796 8932 38668
rect 8988 38722 9044 39566
rect 8988 38670 8990 38722
rect 9042 38670 9044 38722
rect 8988 38658 9044 38670
rect 9100 34916 9156 40236
rect 9212 39284 9268 40350
rect 9212 39218 9268 39228
rect 9324 39732 9380 39742
rect 9324 38668 9380 39676
rect 9436 38834 9492 40908
rect 9436 38782 9438 38834
rect 9490 38782 9492 38834
rect 9436 38770 9492 38782
rect 9548 39506 9604 39518
rect 9548 39454 9550 39506
rect 9602 39454 9604 39506
rect 9100 34850 9156 34860
rect 9212 38612 9380 38668
rect 9100 34692 9156 34702
rect 9100 34130 9156 34636
rect 9100 34078 9102 34130
rect 9154 34078 9156 34130
rect 9100 34066 9156 34078
rect 8876 33730 8932 33740
rect 8876 33348 8932 33358
rect 8876 33254 8932 33292
rect 9212 33236 9268 38612
rect 9324 37156 9380 37166
rect 9324 37154 9492 37156
rect 9324 37102 9326 37154
rect 9378 37102 9492 37154
rect 9324 37100 9492 37102
rect 9324 37090 9380 37100
rect 9324 35586 9380 35598
rect 9324 35534 9326 35586
rect 9378 35534 9380 35586
rect 9324 34468 9380 35534
rect 9436 35364 9492 37100
rect 9548 36820 9604 39454
rect 9660 37938 9716 37950
rect 9660 37886 9662 37938
rect 9714 37886 9716 37938
rect 9660 37268 9716 37886
rect 9660 37202 9716 37212
rect 9548 36754 9604 36764
rect 9772 35308 9828 41020
rect 9884 40180 9940 41692
rect 9996 41300 10052 55918
rect 11452 55188 11508 57344
rect 12796 56644 12852 57344
rect 14140 56756 14196 57344
rect 14140 56700 14644 56756
rect 12796 56588 13076 56644
rect 13020 56306 13076 56588
rect 13020 56254 13022 56306
rect 13074 56254 13076 56306
rect 13020 56242 13076 56254
rect 14588 56306 14644 56700
rect 14588 56254 14590 56306
rect 14642 56254 14644 56306
rect 14588 56242 14644 56254
rect 15484 56308 15540 57344
rect 16828 57204 16884 57344
rect 16828 57148 16996 57204
rect 15484 56242 15540 56252
rect 16492 56308 16548 56318
rect 16492 56214 16548 56252
rect 11452 55122 11508 55132
rect 11564 55970 11620 55982
rect 11564 55918 11566 55970
rect 11618 55918 11620 55970
rect 11564 54516 11620 55918
rect 14028 55970 14084 55982
rect 14028 55918 14030 55970
rect 14082 55918 14084 55970
rect 14028 55748 14084 55918
rect 14028 55682 14084 55692
rect 15596 55970 15652 55982
rect 15596 55918 15598 55970
rect 15650 55918 15652 55970
rect 12908 55298 12964 55310
rect 12908 55246 12910 55298
rect 12962 55246 12964 55298
rect 11900 55188 11956 55198
rect 11900 55094 11956 55132
rect 11564 54450 11620 54460
rect 10220 53844 10276 53854
rect 9996 41234 10052 41244
rect 10108 41298 10164 41310
rect 10108 41246 10110 41298
rect 10162 41246 10164 41298
rect 10108 40292 10164 41246
rect 10108 40226 10164 40236
rect 9884 40124 10052 40180
rect 9436 35298 9492 35308
rect 9548 35252 9828 35308
rect 9884 39284 9940 39294
rect 9884 38836 9940 39228
rect 9548 34692 9604 35252
rect 9660 34916 9716 34926
rect 9660 34914 9828 34916
rect 9660 34862 9662 34914
rect 9714 34862 9828 34914
rect 9660 34860 9828 34862
rect 9660 34850 9716 34860
rect 9548 34636 9716 34692
rect 9324 34402 9380 34412
rect 9548 34468 9604 34478
rect 9548 34130 9604 34412
rect 9548 34078 9550 34130
rect 9602 34078 9604 34130
rect 9548 34066 9604 34078
rect 9436 33460 9492 33470
rect 9324 33236 9380 33246
rect 9212 33234 9380 33236
rect 9212 33182 9326 33234
rect 9378 33182 9380 33234
rect 9212 33180 9380 33182
rect 9324 33170 9380 33180
rect 9324 32676 9380 32686
rect 8876 32338 8932 32350
rect 8876 32286 8878 32338
rect 8930 32286 8932 32338
rect 8876 30996 8932 32286
rect 8876 30930 8932 30940
rect 9100 30994 9156 31006
rect 9100 30942 9102 30994
rect 9154 30942 9156 30994
rect 9100 30884 9156 30942
rect 9100 30818 9156 30828
rect 8876 30212 8932 30222
rect 8876 30118 8932 30156
rect 8988 29202 9044 29214
rect 8988 29150 8990 29202
rect 9042 29150 9044 29202
rect 8988 28980 9044 29150
rect 8988 28914 9044 28924
rect 9324 26964 9380 32620
rect 9436 30436 9492 33404
rect 9660 31890 9716 34636
rect 9772 34018 9828 34860
rect 9772 33966 9774 34018
rect 9826 33966 9828 34018
rect 9772 33954 9828 33966
rect 9884 32788 9940 38780
rect 9996 34802 10052 40124
rect 10108 39172 10164 39182
rect 10108 38834 10164 39116
rect 10108 38782 10110 38834
rect 10162 38782 10164 38834
rect 10108 38770 10164 38782
rect 10220 36706 10276 53788
rect 10892 52612 10948 52622
rect 10780 50708 10836 50718
rect 10556 41076 10612 41086
rect 10332 41074 10612 41076
rect 10332 41022 10558 41074
rect 10610 41022 10612 41074
rect 10332 41020 10612 41022
rect 10332 37380 10388 41020
rect 10556 41010 10612 41020
rect 10444 40402 10500 40414
rect 10444 40350 10446 40402
rect 10498 40350 10500 40402
rect 10444 39508 10500 40350
rect 10444 39442 10500 39452
rect 10556 39506 10612 39518
rect 10556 39454 10558 39506
rect 10610 39454 10612 39506
rect 10332 37314 10388 37324
rect 10444 38052 10500 38062
rect 10220 36654 10222 36706
rect 10274 36654 10276 36706
rect 10220 36642 10276 36654
rect 9996 34750 9998 34802
rect 10050 34750 10052 34802
rect 9996 34738 10052 34750
rect 10220 34132 10276 34142
rect 10220 34038 10276 34076
rect 10444 33572 10500 37996
rect 10556 36706 10612 39454
rect 10556 36654 10558 36706
rect 10610 36654 10612 36706
rect 10556 36642 10612 36654
rect 10668 37716 10724 37726
rect 9772 32732 9940 32788
rect 10332 33516 10500 33572
rect 9772 32340 9828 32732
rect 9884 32564 9940 32574
rect 9884 32562 10052 32564
rect 9884 32510 9886 32562
rect 9938 32510 10052 32562
rect 9884 32508 10052 32510
rect 9884 32498 9940 32508
rect 9772 32284 9940 32340
rect 9660 31838 9662 31890
rect 9714 31838 9716 31890
rect 9660 31826 9716 31838
rect 9660 30660 9716 30670
rect 9436 30380 9604 30436
rect 9436 30212 9492 30222
rect 9436 30118 9492 30156
rect 9548 28756 9604 30380
rect 9436 28700 9604 28756
rect 9436 27524 9492 28700
rect 9548 28532 9604 28542
rect 9548 28438 9604 28476
rect 9660 28308 9716 30604
rect 9436 27458 9492 27468
rect 9548 28252 9716 28308
rect 9772 29764 9828 29774
rect 9324 26898 9380 26908
rect 9436 27300 9492 27310
rect 8988 26852 9044 26862
rect 8988 26850 9156 26852
rect 8988 26798 8990 26850
rect 9042 26798 9156 26850
rect 8988 26796 9156 26798
rect 8988 26786 9044 26796
rect 9100 26292 9156 26796
rect 9324 26292 9380 26302
rect 9100 26290 9380 26292
rect 9100 26238 9326 26290
rect 9378 26238 9380 26290
rect 9100 26236 9380 26238
rect 9324 26226 9380 26236
rect 8988 26178 9044 26190
rect 8988 26126 8990 26178
rect 9042 26126 9044 26178
rect 8988 24052 9044 26126
rect 9100 25508 9156 25518
rect 9100 25414 9156 25452
rect 9212 24836 9268 24846
rect 9212 24722 9268 24780
rect 9212 24670 9214 24722
rect 9266 24670 9268 24722
rect 9212 24658 9268 24670
rect 8988 23986 9044 23996
rect 8988 23828 9044 23838
rect 8876 23492 8932 23502
rect 8876 23042 8932 23436
rect 8876 22990 8878 23042
rect 8930 22990 8932 23042
rect 8876 22978 8932 22990
rect 8764 20066 8820 20076
rect 8876 20802 8932 20814
rect 8876 20750 8878 20802
rect 8930 20750 8932 20802
rect 8876 19908 8932 20750
rect 8876 19842 8932 19852
rect 8764 18340 8820 18350
rect 8764 18246 8820 18284
rect 8652 17948 8820 18004
rect 8316 15474 8372 15484
rect 8428 16882 8484 16894
rect 8428 16830 8430 16882
rect 8482 16830 8484 16882
rect 8204 15262 8206 15314
rect 8258 15262 8260 15314
rect 8204 15250 8260 15262
rect 7644 15090 7700 15102
rect 7868 15092 8372 15148
rect 7644 15038 7646 15090
rect 7698 15038 7700 15090
rect 7644 14756 7700 15038
rect 7644 14690 7700 14700
rect 7868 14644 7924 14654
rect 7532 14476 7812 14532
rect 7308 14308 7364 14318
rect 7308 14214 7364 14252
rect 7532 14308 7588 14318
rect 7532 14306 7700 14308
rect 7532 14254 7534 14306
rect 7586 14254 7700 14306
rect 7532 14252 7700 14254
rect 7532 14242 7588 14252
rect 7308 13860 7364 13870
rect 6748 11890 6804 11900
rect 6972 12124 7140 12180
rect 7196 12964 7252 12974
rect 6636 11564 6804 11620
rect 6636 11396 6692 11406
rect 6636 11302 6692 11340
rect 6748 11284 6804 11564
rect 6748 10724 6804 11228
rect 6748 10668 6916 10724
rect 6580 10556 6692 10612
rect 6524 10518 6580 10556
rect 6188 10210 6244 10220
rect 6524 9940 6580 9950
rect 6524 9846 6580 9884
rect 6412 9156 6468 9166
rect 6412 9062 6468 9100
rect 6300 8372 6356 8382
rect 6300 8278 6356 8316
rect 6636 8258 6692 10556
rect 6748 10500 6804 10510
rect 6748 10406 6804 10444
rect 6748 10052 6804 10062
rect 6748 8932 6804 9996
rect 6748 8866 6804 8876
rect 6636 8206 6638 8258
rect 6690 8206 6692 8258
rect 6636 8194 6692 8206
rect 6748 8372 6804 8382
rect 6748 7474 6804 8316
rect 6748 7422 6750 7474
rect 6802 7422 6804 7474
rect 6748 7410 6804 7422
rect 6076 6738 6132 6748
rect 5852 252 6132 308
rect 5852 84 5908 252
rect 6076 112 6132 252
rect 6860 196 6916 10668
rect 6972 10164 7028 12124
rect 7084 11508 7140 11518
rect 7196 11508 7252 12908
rect 7308 12962 7364 13804
rect 7420 13524 7476 13534
rect 7420 13430 7476 13468
rect 7308 12910 7310 12962
rect 7362 12910 7364 12962
rect 7308 12898 7364 12910
rect 7420 12740 7476 12750
rect 7308 12066 7364 12078
rect 7308 12014 7310 12066
rect 7362 12014 7364 12066
rect 7308 11844 7364 12014
rect 7308 11778 7364 11788
rect 7084 11506 7252 11508
rect 7084 11454 7086 11506
rect 7138 11454 7252 11506
rect 7084 11452 7252 11454
rect 7084 11442 7140 11452
rect 7308 11394 7364 11406
rect 7308 11342 7310 11394
rect 7362 11342 7364 11394
rect 6972 10098 7028 10108
rect 7084 11284 7140 11294
rect 7084 10388 7140 11228
rect 7196 10948 7252 10958
rect 7196 10834 7252 10892
rect 7196 10782 7198 10834
rect 7250 10782 7252 10834
rect 7196 10770 7252 10782
rect 6972 9940 7028 9950
rect 6972 9042 7028 9884
rect 7084 9938 7140 10332
rect 7084 9886 7086 9938
rect 7138 9886 7140 9938
rect 7084 9874 7140 9886
rect 7308 9826 7364 11342
rect 7420 11396 7476 12684
rect 7644 12628 7700 14252
rect 7756 12964 7812 14476
rect 7868 14530 7924 14588
rect 7868 14478 7870 14530
rect 7922 14478 7924 14530
rect 7868 14466 7924 14478
rect 7980 14530 8036 14542
rect 7980 14478 7982 14530
rect 8034 14478 8036 14530
rect 7868 13188 7924 13198
rect 7980 13188 8036 14478
rect 8204 14532 8260 14542
rect 8204 14438 8260 14476
rect 7868 13186 8036 13188
rect 7868 13134 7870 13186
rect 7922 13134 8036 13186
rect 7868 13132 8036 13134
rect 8092 14418 8148 14430
rect 8092 14366 8094 14418
rect 8146 14366 8148 14418
rect 7868 13122 7924 13132
rect 7980 12964 8036 12974
rect 7812 12962 8036 12964
rect 7812 12910 7982 12962
rect 8034 12910 8036 12962
rect 7812 12908 8036 12910
rect 7756 12870 7812 12908
rect 7980 12898 8036 12908
rect 7868 12740 7924 12750
rect 7868 12646 7924 12684
rect 7532 12572 7700 12628
rect 7532 11618 7588 12572
rect 8092 12180 8148 14366
rect 8204 14308 8260 14318
rect 8204 13524 8260 14252
rect 8204 13458 8260 13468
rect 8204 12740 8260 12750
rect 8204 12646 8260 12684
rect 8316 12628 8372 15092
rect 8428 14420 8484 16830
rect 8428 14354 8484 14364
rect 8540 15988 8596 15998
rect 8540 13972 8596 15932
rect 8764 15202 8820 17948
rect 8876 17780 8932 17790
rect 8876 17686 8932 17724
rect 8988 16996 9044 23772
rect 9100 23716 9156 23726
rect 9100 20244 9156 23660
rect 9324 23268 9380 23278
rect 9324 23174 9380 23212
rect 9100 20178 9156 20188
rect 9212 21476 9268 21486
rect 9212 20018 9268 21420
rect 9436 20916 9492 27244
rect 9548 26292 9604 28252
rect 9772 28082 9828 29708
rect 9772 28030 9774 28082
rect 9826 28030 9828 28082
rect 9772 28018 9828 28030
rect 9548 26226 9604 26236
rect 9660 27524 9716 27534
rect 9548 25732 9604 25742
rect 9548 25638 9604 25676
rect 9660 25508 9716 27468
rect 9772 26292 9828 26302
rect 9772 26198 9828 26236
rect 9660 25442 9716 25452
rect 9772 26068 9828 26078
rect 9660 23716 9716 23726
rect 9548 23268 9604 23278
rect 9548 22370 9604 23212
rect 9548 22318 9550 22370
rect 9602 22318 9604 22370
rect 9548 21924 9604 22318
rect 9548 21858 9604 21868
rect 9212 19966 9214 20018
rect 9266 19966 9268 20018
rect 8988 16930 9044 16940
rect 9100 17668 9156 17678
rect 9100 17108 9156 17612
rect 9212 17556 9268 19966
rect 9324 20860 9492 20916
rect 9324 19458 9380 20860
rect 9436 20692 9492 20702
rect 9660 20692 9716 23660
rect 9772 23492 9828 26012
rect 9772 23426 9828 23436
rect 9436 20690 9716 20692
rect 9436 20638 9438 20690
rect 9490 20638 9716 20690
rect 9436 20636 9716 20638
rect 9772 23268 9828 23278
rect 9436 20626 9492 20636
rect 9772 20580 9828 23212
rect 9324 19406 9326 19458
rect 9378 19406 9380 19458
rect 9324 18340 9380 19406
rect 9324 18274 9380 18284
rect 9548 20524 9828 20580
rect 9436 17780 9492 17790
rect 9548 17780 9604 20524
rect 9436 17778 9604 17780
rect 9436 17726 9438 17778
rect 9490 17726 9604 17778
rect 9436 17724 9604 17726
rect 9772 20244 9828 20254
rect 9436 17714 9492 17724
rect 9772 17668 9828 20188
rect 9884 19572 9940 32284
rect 9996 32228 10052 32508
rect 9996 32162 10052 32172
rect 10332 32450 10388 33516
rect 10668 33460 10724 37660
rect 10780 34356 10836 50652
rect 10892 41636 10948 52556
rect 10892 41570 10948 41580
rect 11228 48020 11284 48030
rect 10892 40292 10948 40302
rect 10892 38052 10948 40236
rect 11004 38836 11060 38846
rect 11004 38742 11060 38780
rect 11228 38668 11284 47964
rect 11900 47348 11956 47358
rect 11788 41186 11844 41198
rect 11788 41134 11790 41186
rect 11842 41134 11844 41186
rect 11788 40964 11844 41134
rect 11788 40898 11844 40908
rect 11788 38948 11844 38958
rect 11788 38834 11844 38892
rect 11788 38782 11790 38834
rect 11842 38782 11844 38834
rect 11228 38612 11396 38668
rect 10892 37986 10948 37996
rect 10892 36482 10948 36494
rect 10892 36430 10894 36482
rect 10946 36430 10948 36482
rect 10892 34916 10948 36430
rect 10892 34822 10948 34860
rect 11228 35252 11284 35262
rect 10780 34300 11060 34356
rect 10892 34132 10948 34142
rect 10892 34038 10948 34076
rect 10892 33460 10948 33470
rect 10668 33458 10948 33460
rect 10668 33406 10894 33458
rect 10946 33406 10948 33458
rect 10668 33404 10948 33406
rect 10444 33236 10500 33246
rect 10444 33234 10836 33236
rect 10444 33182 10446 33234
rect 10498 33182 10836 33234
rect 10444 33180 10836 33182
rect 10444 33170 10500 33180
rect 10332 32398 10334 32450
rect 10386 32398 10388 32450
rect 10332 31892 10388 32398
rect 10108 31780 10164 31790
rect 10108 31444 10164 31724
rect 10220 31778 10276 31790
rect 10220 31726 10222 31778
rect 10274 31726 10276 31778
rect 10220 31668 10276 31726
rect 10220 31602 10276 31612
rect 9996 31108 10052 31118
rect 9996 30994 10052 31052
rect 9996 30942 9998 30994
rect 10050 30942 10052 30994
rect 9996 30930 10052 30942
rect 10108 30212 10164 31388
rect 10332 30548 10388 31836
rect 9996 30156 10164 30212
rect 10220 30492 10388 30548
rect 10444 33012 10500 33022
rect 9996 29428 10052 30156
rect 10108 29988 10164 29998
rect 10108 29650 10164 29932
rect 10108 29598 10110 29650
rect 10162 29598 10164 29650
rect 10108 29586 10164 29598
rect 9996 29372 10164 29428
rect 9996 28980 10052 28990
rect 9996 28866 10052 28924
rect 9996 28814 9998 28866
rect 10050 28814 10052 28866
rect 9996 27300 10052 28814
rect 10108 27972 10164 29372
rect 10108 27906 10164 27916
rect 10220 27748 10276 30492
rect 10444 30436 10500 32956
rect 10668 31666 10724 31678
rect 10668 31614 10670 31666
rect 10722 31614 10724 31666
rect 10220 27682 10276 27692
rect 10332 30380 10500 30436
rect 10556 30994 10612 31006
rect 10556 30942 10558 30994
rect 10610 30942 10612 30994
rect 10108 27300 10164 27310
rect 10052 27298 10164 27300
rect 10052 27246 10110 27298
rect 10162 27246 10164 27298
rect 10052 27244 10164 27246
rect 9996 27206 10052 27244
rect 10108 27234 10164 27244
rect 10220 27076 10276 27086
rect 9996 26068 10052 26078
rect 9996 25974 10052 26012
rect 9996 24722 10052 24734
rect 9996 24670 9998 24722
rect 10050 24670 10052 24722
rect 9996 23716 10052 24670
rect 9996 23660 10164 23716
rect 9996 23492 10052 23502
rect 9996 23156 10052 23436
rect 10108 23380 10164 23660
rect 10108 23314 10164 23324
rect 9996 22484 10052 23100
rect 9996 22482 10164 22484
rect 9996 22430 9998 22482
rect 10050 22430 10164 22482
rect 9996 22428 10164 22430
rect 9996 22418 10052 22428
rect 10108 20804 10164 22428
rect 10220 21028 10276 27020
rect 10332 24050 10388 30380
rect 10444 30210 10500 30222
rect 10444 30158 10446 30210
rect 10498 30158 10500 30210
rect 10444 29876 10500 30158
rect 10556 29988 10612 30942
rect 10556 29922 10612 29932
rect 10444 29810 10500 29820
rect 10332 23998 10334 24050
rect 10386 23998 10388 24050
rect 10332 23986 10388 23998
rect 10444 28532 10500 28542
rect 10444 27858 10500 28476
rect 10444 27806 10446 27858
rect 10498 27806 10500 27858
rect 10332 23154 10388 23166
rect 10332 23102 10334 23154
rect 10386 23102 10388 23154
rect 10332 22820 10388 23102
rect 10332 22754 10388 22764
rect 10220 20916 10276 20972
rect 10444 22596 10500 27806
rect 10556 28420 10612 28430
rect 10556 27524 10612 28364
rect 10556 27074 10612 27468
rect 10556 27022 10558 27074
rect 10610 27022 10612 27074
rect 10556 27010 10612 27022
rect 10668 26908 10724 31614
rect 10780 30212 10836 33180
rect 10892 31780 10948 33404
rect 10892 31714 10948 31724
rect 10892 30772 10948 30782
rect 10892 30322 10948 30716
rect 10892 30270 10894 30322
rect 10946 30270 10948 30322
rect 10892 30258 10948 30270
rect 10780 30100 10836 30156
rect 10780 30044 10948 30100
rect 10892 28756 10948 30044
rect 10892 28084 10948 28700
rect 10892 28018 10948 28028
rect 11004 27860 11060 34300
rect 11228 34132 11284 35196
rect 11116 31892 11172 31902
rect 11116 31798 11172 31836
rect 11228 31668 11284 34076
rect 11116 31612 11284 31668
rect 11116 30660 11172 31612
rect 11340 31444 11396 38612
rect 11788 36708 11844 38782
rect 11788 36642 11844 36652
rect 11676 35476 11732 35486
rect 11452 32338 11508 32350
rect 11452 32286 11454 32338
rect 11506 32286 11508 32338
rect 11452 31892 11508 32286
rect 11676 32228 11732 35420
rect 11788 34132 11844 34142
rect 11788 34038 11844 34076
rect 11676 32162 11732 32172
rect 11452 31836 11620 31892
rect 11564 31780 11620 31836
rect 11788 31780 11844 31790
rect 11564 31778 11844 31780
rect 11564 31726 11790 31778
rect 11842 31726 11844 31778
rect 11564 31724 11844 31726
rect 11788 31714 11844 31724
rect 11452 31668 11508 31678
rect 11452 31574 11508 31612
rect 11340 31378 11396 31388
rect 11676 31444 11732 31454
rect 11228 31108 11284 31118
rect 11228 30882 11284 31052
rect 11228 30830 11230 30882
rect 11282 30830 11284 30882
rect 11228 30818 11284 30830
rect 11340 30994 11396 31006
rect 11340 30942 11342 30994
rect 11394 30942 11396 30994
rect 11340 30660 11396 30942
rect 11116 30604 11284 30660
rect 11116 28644 11172 28654
rect 11116 28550 11172 28588
rect 11004 27794 11060 27804
rect 11116 28420 11172 28430
rect 10892 27746 10948 27758
rect 10892 27694 10894 27746
rect 10946 27694 10948 27746
rect 10668 26852 10836 26908
rect 10668 26290 10724 26302
rect 10668 26238 10670 26290
rect 10722 26238 10724 26290
rect 10556 26068 10612 26078
rect 10556 24722 10612 26012
rect 10668 25730 10724 26238
rect 10668 25678 10670 25730
rect 10722 25678 10724 25730
rect 10668 25666 10724 25678
rect 10556 24670 10558 24722
rect 10610 24670 10612 24722
rect 10556 24658 10612 24670
rect 10668 25508 10724 25518
rect 10332 20916 10388 20926
rect 10220 20914 10388 20916
rect 10220 20862 10334 20914
rect 10386 20862 10388 20914
rect 10220 20860 10388 20862
rect 10332 20850 10388 20860
rect 10108 20748 10276 20804
rect 9996 20020 10052 20030
rect 9996 19926 10052 19964
rect 9884 19516 10052 19572
rect 9884 19348 9940 19358
rect 9884 19254 9940 19292
rect 9884 18226 9940 18238
rect 9884 18174 9886 18226
rect 9938 18174 9940 18226
rect 9884 17780 9940 18174
rect 9996 17780 10052 19516
rect 9996 17724 10164 17780
rect 9884 17714 9940 17724
rect 9716 17612 9828 17668
rect 9212 17500 9604 17556
rect 8988 16770 9044 16782
rect 8988 16718 8990 16770
rect 9042 16718 9044 16770
rect 8988 16212 9044 16718
rect 9100 16324 9156 17052
rect 9324 16884 9380 16894
rect 9324 16790 9380 16828
rect 9100 16322 9380 16324
rect 9100 16270 9102 16322
rect 9154 16270 9380 16322
rect 9100 16268 9380 16270
rect 9100 16258 9156 16268
rect 8988 16146 9044 16156
rect 9100 15988 9156 15998
rect 9100 15894 9156 15932
rect 8876 15876 8932 15886
rect 8876 15782 8932 15820
rect 8764 15150 8766 15202
rect 8818 15150 8820 15202
rect 8764 15148 8820 15150
rect 8652 15092 8820 15148
rect 9324 15148 9380 16268
rect 9324 15092 9492 15148
rect 8652 14308 8708 15092
rect 9324 14868 9380 14878
rect 9100 14756 9156 14766
rect 9100 14662 9156 14700
rect 8876 14644 8932 14654
rect 8876 14550 8932 14588
rect 9324 14642 9380 14812
rect 9324 14590 9326 14642
rect 9378 14590 9380 14642
rect 9324 14578 9380 14590
rect 8764 14532 8820 14542
rect 8764 14438 8820 14476
rect 8652 14242 8708 14252
rect 8316 12562 8372 12572
rect 8428 13916 8596 13972
rect 8428 12404 8484 13916
rect 8540 13748 8596 13758
rect 8540 13654 8596 13692
rect 9324 13748 9380 13758
rect 9324 13654 9380 13692
rect 7532 11566 7534 11618
rect 7586 11566 7588 11618
rect 7532 11554 7588 11566
rect 7644 12124 8148 12180
rect 8204 12348 8484 12404
rect 8764 13636 8820 13646
rect 7532 11396 7588 11406
rect 7420 11394 7588 11396
rect 7420 11342 7534 11394
rect 7586 11342 7588 11394
rect 7420 11340 7588 11342
rect 7532 11330 7588 11340
rect 7644 11172 7700 12124
rect 8092 11956 8148 11966
rect 7644 11106 7700 11116
rect 7756 11954 8148 11956
rect 7756 11902 8094 11954
rect 8146 11902 8148 11954
rect 7756 11900 8148 11902
rect 7756 10948 7812 11900
rect 8092 11890 8148 11900
rect 8204 11732 8260 12348
rect 8764 12178 8820 13580
rect 8988 13636 9044 13646
rect 8988 13542 9044 13580
rect 8988 13188 9044 13198
rect 9436 13188 9492 15092
rect 8988 13186 9492 13188
rect 8988 13134 8990 13186
rect 9042 13134 9492 13186
rect 8988 13132 9492 13134
rect 8988 13122 9044 13132
rect 8764 12126 8766 12178
rect 8818 12126 8820 12178
rect 8764 12114 8820 12126
rect 8876 12738 8932 12750
rect 8876 12686 8878 12738
rect 8930 12686 8932 12738
rect 8540 12068 8596 12078
rect 8540 11974 8596 12012
rect 8652 12066 8708 12078
rect 8652 12014 8654 12066
rect 8706 12014 8708 12066
rect 8652 11732 8708 12014
rect 7868 11676 8260 11732
rect 8316 11676 8708 11732
rect 8764 11844 8820 11854
rect 7868 11394 7924 11676
rect 8316 11618 8372 11676
rect 8316 11566 8318 11618
rect 8370 11566 8372 11618
rect 8316 11554 8372 11566
rect 8204 11508 8260 11518
rect 8204 11414 8260 11452
rect 7868 11342 7870 11394
rect 7922 11342 7924 11394
rect 7868 11330 7924 11342
rect 7756 10882 7812 10892
rect 8652 11172 8708 11182
rect 7980 10724 8036 10734
rect 7980 10630 8036 10668
rect 7420 10610 7476 10622
rect 7420 10558 7422 10610
rect 7474 10558 7476 10610
rect 7420 10050 7476 10558
rect 7756 10610 7812 10622
rect 7756 10558 7758 10610
rect 7810 10558 7812 10610
rect 7756 10500 7812 10558
rect 7868 10612 7924 10622
rect 7868 10518 7924 10556
rect 7756 10434 7812 10444
rect 7420 9998 7422 10050
rect 7474 9998 7476 10050
rect 7420 9986 7476 9998
rect 7644 10388 7700 10398
rect 7308 9774 7310 9826
rect 7362 9774 7364 9826
rect 7308 9716 7364 9774
rect 7532 9940 7588 9950
rect 7532 9826 7588 9884
rect 7532 9774 7534 9826
rect 7586 9774 7588 9826
rect 7532 9762 7588 9774
rect 6972 8990 6974 9042
rect 7026 8990 7028 9042
rect 6972 8978 7028 8990
rect 7084 9660 7364 9716
rect 7084 7812 7140 9660
rect 7420 9156 7476 9166
rect 7420 9062 7476 9100
rect 7532 9044 7588 9054
rect 7644 9044 7700 10332
rect 8092 10388 8148 10398
rect 8092 10294 8148 10332
rect 8204 10276 8260 10286
rect 7868 9828 7924 9838
rect 7868 9734 7924 9772
rect 7532 9042 8036 9044
rect 7532 8990 7534 9042
rect 7586 8990 8036 9042
rect 7532 8988 8036 8990
rect 7532 8978 7588 8988
rect 7308 8932 7364 8942
rect 7308 8838 7364 8876
rect 7196 8708 7252 8718
rect 7196 8370 7252 8652
rect 7196 8318 7198 8370
rect 7250 8318 7252 8370
rect 7196 8306 7252 8318
rect 7980 8372 8036 8988
rect 8092 9042 8148 9054
rect 8092 8990 8094 9042
rect 8146 8990 8148 9042
rect 8092 8596 8148 8990
rect 8092 8530 8148 8540
rect 8092 8372 8148 8382
rect 7980 8370 8148 8372
rect 7980 8318 8094 8370
rect 8146 8318 8148 8370
rect 7980 8316 8148 8318
rect 8092 8306 8148 8316
rect 8204 8370 8260 10220
rect 8540 8818 8596 8830
rect 8540 8766 8542 8818
rect 8594 8766 8596 8818
rect 8540 8708 8596 8766
rect 8540 8642 8596 8652
rect 8428 8484 8484 8494
rect 8428 8390 8484 8428
rect 8204 8318 8206 8370
rect 8258 8318 8260 8370
rect 8204 8306 8260 8318
rect 7756 8148 7812 8158
rect 7756 8054 7812 8092
rect 7084 7746 7140 7756
rect 7308 7588 7364 7598
rect 7308 7494 7364 7532
rect 7756 6804 7812 6814
rect 7756 6130 7812 6748
rect 7756 6078 7758 6130
rect 7810 6078 7812 6130
rect 7756 6066 7812 6078
rect 7756 5684 7812 5694
rect 7756 5346 7812 5628
rect 7756 5294 7758 5346
rect 7810 5294 7812 5346
rect 7756 5282 7812 5294
rect 8316 5236 8372 5246
rect 8316 5142 8372 5180
rect 8652 3388 8708 11116
rect 8764 10948 8820 11788
rect 8764 10882 8820 10892
rect 8764 10724 8820 10734
rect 8764 10610 8820 10668
rect 8764 10558 8766 10610
rect 8818 10558 8820 10610
rect 8764 10546 8820 10558
rect 8876 9828 8932 12686
rect 9212 12738 9268 12750
rect 9212 12686 9214 12738
rect 9266 12686 9268 12738
rect 8988 12068 9044 12078
rect 8988 11394 9044 12012
rect 9212 11508 9268 12686
rect 8988 11342 8990 11394
rect 9042 11342 9044 11394
rect 8988 9940 9044 11342
rect 9100 11396 9156 11406
rect 9212 11396 9268 11452
rect 9100 11394 9268 11396
rect 9100 11342 9102 11394
rect 9154 11342 9268 11394
rect 9100 11340 9268 11342
rect 9324 12740 9380 12750
rect 9324 11956 9380 12684
rect 9436 12404 9492 12414
rect 9436 12290 9492 12348
rect 9436 12238 9438 12290
rect 9490 12238 9492 12290
rect 9436 12226 9492 12238
rect 9324 11394 9380 11900
rect 9324 11342 9326 11394
rect 9378 11342 9380 11394
rect 9100 11330 9156 11340
rect 9324 11330 9380 11342
rect 9548 11284 9604 17500
rect 9716 17332 9772 17612
rect 9996 17554 10052 17566
rect 9996 17502 9998 17554
rect 10050 17502 10052 17554
rect 9996 17332 10052 17502
rect 9716 17276 9828 17332
rect 9660 16996 9716 17006
rect 9660 16660 9716 16940
rect 9772 16882 9828 17276
rect 9996 17266 10052 17276
rect 10108 17556 10164 17724
rect 10108 16996 10164 17500
rect 10108 16930 10164 16940
rect 9772 16830 9774 16882
rect 9826 16830 9828 16882
rect 9772 16818 9828 16830
rect 9884 16884 9940 16894
rect 9660 16604 9828 16660
rect 9660 16324 9716 16334
rect 9660 15204 9716 16268
rect 9660 12068 9716 15148
rect 9772 13746 9828 16604
rect 9884 15538 9940 16828
rect 10108 16772 10164 16782
rect 9996 16658 10052 16670
rect 9996 16606 9998 16658
rect 10050 16606 10052 16658
rect 9996 16098 10052 16606
rect 9996 16046 9998 16098
rect 10050 16046 10052 16098
rect 9996 16034 10052 16046
rect 10108 16436 10164 16716
rect 9884 15486 9886 15538
rect 9938 15486 9940 15538
rect 9884 15474 9940 15486
rect 9996 15540 10052 15550
rect 9996 14756 10052 15484
rect 9996 14690 10052 14700
rect 9884 14532 9940 14542
rect 9884 14530 10052 14532
rect 9884 14478 9886 14530
rect 9938 14478 10052 14530
rect 9884 14476 10052 14478
rect 9884 14466 9940 14476
rect 9772 13694 9774 13746
rect 9826 13694 9828 13746
rect 9772 12740 9828 13694
rect 9884 14308 9940 14318
rect 9884 12962 9940 14252
rect 9996 13634 10052 14476
rect 10108 13748 10164 16380
rect 10108 13682 10164 13692
rect 9996 13582 9998 13634
rect 10050 13582 10052 13634
rect 9996 13570 10052 13582
rect 9884 12910 9886 12962
rect 9938 12910 9940 12962
rect 9884 12898 9940 12910
rect 10108 13524 10164 13534
rect 10108 12852 10164 13468
rect 10220 13076 10276 20748
rect 10444 20020 10500 22540
rect 10556 21588 10612 21598
rect 10556 21494 10612 21532
rect 10556 20020 10612 20030
rect 10444 20018 10612 20020
rect 10444 19966 10558 20018
rect 10610 19966 10612 20018
rect 10444 19964 10612 19966
rect 10556 19954 10612 19964
rect 10332 19234 10388 19246
rect 10332 19182 10334 19234
rect 10386 19182 10388 19234
rect 10332 17332 10388 19182
rect 10556 18676 10612 18686
rect 10556 18562 10612 18620
rect 10556 18510 10558 18562
rect 10610 18510 10612 18562
rect 10556 18498 10612 18510
rect 10444 17780 10500 17790
rect 10668 17780 10724 25452
rect 10780 24948 10836 26852
rect 10892 25844 10948 27694
rect 11004 26740 11060 26750
rect 11004 26068 11060 26684
rect 11004 26002 11060 26012
rect 11116 25844 11172 28364
rect 11228 26740 11284 30604
rect 11340 30594 11396 30604
rect 11564 29540 11620 29550
rect 11564 29092 11620 29484
rect 11564 28754 11620 29036
rect 11564 28702 11566 28754
rect 11618 28702 11620 28754
rect 11564 28690 11620 28702
rect 11676 28420 11732 31388
rect 11788 30994 11844 31006
rect 11788 30942 11790 30994
rect 11842 30942 11844 30994
rect 11788 29764 11844 30942
rect 11900 30772 11956 47292
rect 12348 45892 12404 45902
rect 12124 41074 12180 41086
rect 12124 41022 12126 41074
rect 12178 41022 12180 41074
rect 12124 40852 12180 41022
rect 12124 40786 12180 40796
rect 12124 40178 12180 40190
rect 12124 40126 12126 40178
rect 12178 40126 12180 40178
rect 12124 38836 12180 40126
rect 12236 38948 12292 38958
rect 12348 38948 12404 45836
rect 12908 40852 12964 55246
rect 15036 53508 15092 53518
rect 14140 52388 14196 52398
rect 12908 40786 12964 40796
rect 13692 51604 13748 51614
rect 12908 40516 12964 40526
rect 12908 40514 13076 40516
rect 12908 40462 12910 40514
rect 12962 40462 13076 40514
rect 12908 40460 13076 40462
rect 12908 40450 12964 40460
rect 12236 38946 12404 38948
rect 12236 38894 12238 38946
rect 12290 38894 12404 38946
rect 12236 38892 12404 38894
rect 12236 38882 12292 38892
rect 12796 38836 12852 38846
rect 12124 38770 12180 38780
rect 12460 38834 12852 38836
rect 12460 38782 12798 38834
rect 12850 38782 12852 38834
rect 12460 38780 12852 38782
rect 12012 37380 12068 37390
rect 12012 37286 12068 37324
rect 12124 37268 12180 37278
rect 12012 35812 12068 35822
rect 12124 35812 12180 37212
rect 12012 35810 12180 35812
rect 12012 35758 12014 35810
rect 12066 35758 12180 35810
rect 12012 35756 12180 35758
rect 12012 35746 12068 35756
rect 12012 33122 12068 33134
rect 12012 33070 12014 33122
rect 12066 33070 12068 33122
rect 12012 32004 12068 33070
rect 12012 31938 12068 31948
rect 12124 31780 12180 35756
rect 12124 31714 12180 31724
rect 12236 36148 12292 36158
rect 12236 31108 12292 36092
rect 12460 32900 12516 38780
rect 12796 38770 12852 38780
rect 12796 37380 12852 37390
rect 12684 34132 12740 34142
rect 12460 32834 12516 32844
rect 12572 34130 12740 34132
rect 12572 34078 12686 34130
rect 12738 34078 12740 34130
rect 12572 34076 12740 34078
rect 12572 33346 12628 34076
rect 12684 34066 12740 34076
rect 12572 33294 12574 33346
rect 12626 33294 12628 33346
rect 12572 32676 12628 33294
rect 12572 32610 12628 32620
rect 12460 32116 12516 32126
rect 12460 32002 12516 32060
rect 12460 31950 12462 32002
rect 12514 31950 12516 32002
rect 12460 31938 12516 31950
rect 12124 31052 12292 31108
rect 12348 31766 12404 31778
rect 12348 31714 12350 31766
rect 12402 31714 12404 31766
rect 12348 31444 12404 31714
rect 12796 31556 12852 37324
rect 12908 32004 12964 32014
rect 12908 31890 12964 31948
rect 12908 31838 12910 31890
rect 12962 31838 12964 31890
rect 12908 31826 12964 31838
rect 11900 30716 12068 30772
rect 11788 29698 11844 29708
rect 11676 28354 11732 28364
rect 11788 29538 11844 29550
rect 11788 29486 11790 29538
rect 11842 29486 11844 29538
rect 11228 26674 11284 26684
rect 11340 28084 11396 28094
rect 11228 26516 11284 26526
rect 11228 26290 11284 26460
rect 11228 26238 11230 26290
rect 11282 26238 11284 26290
rect 11228 26226 11284 26238
rect 10892 25788 11060 25844
rect 10780 24882 10836 24892
rect 11004 25732 11060 25788
rect 11004 24500 11060 25676
rect 11116 25284 11172 25788
rect 11116 25218 11172 25228
rect 11228 26068 11284 26078
rect 11116 24724 11172 24734
rect 11116 24630 11172 24668
rect 11004 24444 11172 24500
rect 10892 23940 10948 23950
rect 10892 23938 11060 23940
rect 10892 23886 10894 23938
rect 10946 23886 11060 23938
rect 10892 23884 11060 23886
rect 10892 23874 10948 23884
rect 10892 23044 10948 23054
rect 10892 22930 10948 22988
rect 10892 22878 10894 22930
rect 10946 22878 10948 22930
rect 10892 22372 10948 22878
rect 11004 22820 11060 23884
rect 11004 22754 11060 22764
rect 11116 22708 11172 24444
rect 11228 23828 11284 26012
rect 11340 25506 11396 28028
rect 11564 27748 11620 27758
rect 11452 27188 11508 27198
rect 11452 27074 11508 27132
rect 11452 27022 11454 27074
rect 11506 27022 11508 27074
rect 11452 27010 11508 27022
rect 11564 26908 11620 27692
rect 11340 25454 11342 25506
rect 11394 25454 11396 25506
rect 11340 25442 11396 25454
rect 11452 26852 11620 26908
rect 11228 23734 11284 23772
rect 11340 25284 11396 25294
rect 11340 23044 11396 25228
rect 11340 22978 11396 22988
rect 11116 22642 11172 22652
rect 11340 22820 11396 22830
rect 10892 22306 10948 22316
rect 11116 22148 11172 22158
rect 10780 22146 11172 22148
rect 10780 22094 11118 22146
rect 11170 22094 11172 22146
rect 10780 22092 11172 22094
rect 10780 20802 10836 22092
rect 11116 22082 11172 22092
rect 11228 22036 11284 22046
rect 10780 20750 10782 20802
rect 10834 20750 10836 20802
rect 10780 20738 10836 20750
rect 10892 21924 10948 21934
rect 10892 20020 10948 21868
rect 11116 21812 11172 21822
rect 11004 21364 11060 21374
rect 11004 21270 11060 21308
rect 11116 20802 11172 21756
rect 11116 20750 11118 20802
rect 11170 20750 11172 20802
rect 11116 20244 11172 20750
rect 11116 20178 11172 20188
rect 11228 21588 11284 21980
rect 11228 20130 11284 21532
rect 11340 21026 11396 22764
rect 11452 22484 11508 26852
rect 11788 25844 11844 29486
rect 11900 28644 11956 28654
rect 11900 28550 11956 28588
rect 12012 28420 12068 30716
rect 12124 30324 12180 31052
rect 12236 30882 12292 30894
rect 12236 30830 12238 30882
rect 12290 30830 12292 30882
rect 12236 30548 12292 30830
rect 12348 30660 12404 31388
rect 12348 30594 12404 30604
rect 12572 31500 12852 31556
rect 12236 30482 12292 30492
rect 12124 30268 12292 30324
rect 12124 29988 12180 29998
rect 12124 29894 12180 29932
rect 12236 29428 12292 30268
rect 12572 30212 12628 31500
rect 12796 30660 12852 30670
rect 12572 30210 12740 30212
rect 12572 30158 12574 30210
rect 12626 30158 12740 30210
rect 12572 30156 12740 30158
rect 12572 30146 12628 30156
rect 11676 25788 11844 25844
rect 11900 28364 12068 28420
rect 12124 29372 12292 29428
rect 11676 25396 11732 25788
rect 11788 25620 11844 25630
rect 11788 25526 11844 25564
rect 11676 25340 11844 25396
rect 11788 24052 11844 25340
rect 11788 23986 11844 23996
rect 11564 23940 11620 23950
rect 11564 23846 11620 23884
rect 11676 23828 11732 23838
rect 11676 23716 11732 23772
rect 11452 22418 11508 22428
rect 11564 23660 11732 23716
rect 11340 20974 11342 21026
rect 11394 20974 11396 21026
rect 11340 20962 11396 20974
rect 11228 20078 11230 20130
rect 11282 20078 11284 20130
rect 11228 20066 11284 20078
rect 11340 20132 11396 20142
rect 10780 19964 10948 20020
rect 10780 18676 10836 19964
rect 10892 19796 10948 19806
rect 10892 19458 10948 19740
rect 10892 19406 10894 19458
rect 10946 19406 10948 19458
rect 10892 19394 10948 19406
rect 11116 19794 11172 19806
rect 11116 19742 11118 19794
rect 11170 19742 11172 19794
rect 11116 19124 11172 19742
rect 11116 19058 11172 19068
rect 10780 18610 10836 18620
rect 11004 18340 11060 18378
rect 11004 18274 11060 18284
rect 10444 17778 10724 17780
rect 10444 17726 10446 17778
rect 10498 17726 10724 17778
rect 10444 17724 10724 17726
rect 11004 18116 11060 18126
rect 10444 17714 10500 17724
rect 10332 17266 10388 17276
rect 10444 16884 10500 16894
rect 10444 16790 10500 16828
rect 10332 16324 10388 16334
rect 10332 14642 10388 16268
rect 10444 16212 10500 16222
rect 10444 16118 10500 16156
rect 10556 15988 10612 17724
rect 11004 17444 11060 18060
rect 11004 16882 11060 17388
rect 11004 16830 11006 16882
rect 11058 16830 11060 16882
rect 11004 16818 11060 16830
rect 11116 17332 11172 17342
rect 11116 16098 11172 17276
rect 11116 16046 11118 16098
rect 11170 16046 11172 16098
rect 11116 16034 11172 16046
rect 11228 16772 11284 16782
rect 10332 14590 10334 14642
rect 10386 14590 10388 14642
rect 10332 14578 10388 14590
rect 10444 15932 10612 15988
rect 10332 13076 10388 13086
rect 10220 13074 10388 13076
rect 10220 13022 10334 13074
rect 10386 13022 10388 13074
rect 10220 13020 10388 13022
rect 10332 13010 10388 13020
rect 10108 12796 10388 12852
rect 9772 12684 10052 12740
rect 9772 12068 9828 12078
rect 9660 12066 9828 12068
rect 9660 12014 9774 12066
rect 9826 12014 9828 12066
rect 9660 12012 9828 12014
rect 9772 12002 9828 12012
rect 9884 11956 9940 11966
rect 9884 11732 9940 11900
rect 9772 11676 9940 11732
rect 9772 11618 9828 11676
rect 9772 11566 9774 11618
rect 9826 11566 9828 11618
rect 9772 11554 9828 11566
rect 9884 11508 9940 11518
rect 9884 11414 9940 11452
rect 9548 11218 9604 11228
rect 9436 11170 9492 11182
rect 9436 11118 9438 11170
rect 9490 11118 9492 11170
rect 8988 9874 9044 9884
rect 9100 11060 9156 11070
rect 9100 9938 9156 11004
rect 9100 9886 9102 9938
rect 9154 9886 9156 9938
rect 9100 9874 9156 9886
rect 9212 10948 9268 10958
rect 8876 9762 8932 9772
rect 9212 6020 9268 10892
rect 9436 10612 9492 11118
rect 9436 10546 9492 10556
rect 9324 10498 9380 10510
rect 9324 10446 9326 10498
rect 9378 10446 9380 10498
rect 9324 9268 9380 10446
rect 9660 10500 9716 10510
rect 9660 10406 9716 10444
rect 9548 10388 9604 10398
rect 9548 10294 9604 10332
rect 9884 10386 9940 10398
rect 9884 10334 9886 10386
rect 9938 10334 9940 10386
rect 9772 10052 9828 10062
rect 9548 9826 9604 9838
rect 9548 9774 9550 9826
rect 9602 9774 9604 9826
rect 9548 9268 9604 9774
rect 9660 9268 9716 9278
rect 9548 9266 9716 9268
rect 9548 9214 9662 9266
rect 9714 9214 9716 9266
rect 9548 9212 9716 9214
rect 9324 9202 9380 9212
rect 9660 9202 9716 9212
rect 9772 8708 9828 9996
rect 9884 9156 9940 10334
rect 9996 9826 10052 12684
rect 10108 12516 10164 12526
rect 10108 10164 10164 12460
rect 10108 10098 10164 10108
rect 10220 10610 10276 10622
rect 10220 10558 10222 10610
rect 10274 10558 10276 10610
rect 9996 9774 9998 9826
rect 10050 9774 10052 9826
rect 9996 9762 10052 9774
rect 10108 9938 10164 9950
rect 10108 9886 10110 9938
rect 10162 9886 10164 9938
rect 9884 9090 9940 9100
rect 9772 8642 9828 8652
rect 9324 8596 9380 8606
rect 9324 7586 9380 8540
rect 9324 7534 9326 7586
rect 9378 7534 9380 7586
rect 9324 7522 9380 7534
rect 9772 7364 9828 7374
rect 9772 7270 9828 7308
rect 10108 6690 10164 9886
rect 10220 8484 10276 10558
rect 10220 8418 10276 8428
rect 10332 8372 10388 12796
rect 10332 8306 10388 8316
rect 10444 7364 10500 15932
rect 10556 15540 10612 15550
rect 10556 15426 10612 15484
rect 10556 15374 10558 15426
rect 10610 15374 10612 15426
rect 10556 15362 10612 15374
rect 11004 15316 11060 15326
rect 11004 15202 11060 15260
rect 11004 15150 11006 15202
rect 11058 15150 11060 15202
rect 11004 15138 11060 15150
rect 11228 15148 11284 16716
rect 11116 15092 11284 15148
rect 10892 14418 10948 14430
rect 10892 14366 10894 14418
rect 10946 14366 10948 14418
rect 10892 13860 10948 14366
rect 11116 13860 11172 15092
rect 11340 14868 11396 20076
rect 10892 13804 11172 13860
rect 10668 13748 10724 13758
rect 10668 13746 10948 13748
rect 10668 13694 10670 13746
rect 10722 13694 10948 13746
rect 10668 13692 10948 13694
rect 10668 13682 10724 13692
rect 10668 13300 10724 13310
rect 10556 12964 10612 12974
rect 10556 9492 10612 12908
rect 10668 10724 10724 13244
rect 10892 12404 10948 13692
rect 11004 12404 11060 12414
rect 10892 12402 11060 12404
rect 10892 12350 11006 12402
rect 11058 12350 11060 12402
rect 10892 12348 11060 12350
rect 11004 12338 11060 12348
rect 11116 11956 11172 13804
rect 11116 11890 11172 11900
rect 11228 14812 11396 14868
rect 11452 18340 11508 18350
rect 11228 13746 11284 14812
rect 11228 13694 11230 13746
rect 11282 13694 11284 13746
rect 11116 11732 11172 11742
rect 11004 11506 11060 11518
rect 11004 11454 11006 11506
rect 11058 11454 11060 11506
rect 10668 10658 10724 10668
rect 10780 11394 10836 11406
rect 10780 11342 10782 11394
rect 10834 11342 10836 11394
rect 10668 10500 10724 10510
rect 10780 10500 10836 11342
rect 10892 10948 10948 10958
rect 10892 10610 10948 10892
rect 10892 10558 10894 10610
rect 10946 10558 10948 10610
rect 10892 10546 10948 10558
rect 10668 10498 10836 10500
rect 10668 10446 10670 10498
rect 10722 10446 10836 10498
rect 10668 10444 10836 10446
rect 10668 10434 10724 10444
rect 10556 9426 10612 9436
rect 10780 9826 10836 9838
rect 10780 9774 10782 9826
rect 10834 9774 10836 9826
rect 10556 9268 10612 9278
rect 10556 9154 10612 9212
rect 10556 9102 10558 9154
rect 10610 9102 10612 9154
rect 10556 8258 10612 9102
rect 10556 8206 10558 8258
rect 10610 8206 10612 8258
rect 10556 8194 10612 8206
rect 10780 7700 10836 9774
rect 10892 9492 10948 9502
rect 10892 8930 10948 9436
rect 11004 9044 11060 11454
rect 11116 11506 11172 11676
rect 11116 11454 11118 11506
rect 11170 11454 11172 11506
rect 11116 11396 11172 11454
rect 11116 11330 11172 11340
rect 11116 10836 11172 10846
rect 11116 10498 11172 10780
rect 11228 10612 11284 13694
rect 11340 14642 11396 14654
rect 11340 14590 11342 14642
rect 11394 14590 11396 14642
rect 11340 13524 11396 14590
rect 11340 13458 11396 13468
rect 11452 13076 11508 18284
rect 11564 18116 11620 23660
rect 11788 22596 11844 22606
rect 11564 18050 11620 18060
rect 11676 22372 11732 22382
rect 11564 17444 11620 17454
rect 11564 17350 11620 17388
rect 11676 17220 11732 22316
rect 11788 22370 11844 22540
rect 11788 22318 11790 22370
rect 11842 22318 11844 22370
rect 11788 22306 11844 22318
rect 11900 21028 11956 28364
rect 12124 28308 12180 29372
rect 12236 29202 12292 29214
rect 12236 29150 12238 29202
rect 12290 29150 12292 29202
rect 12236 28868 12292 29150
rect 12236 28802 12292 28812
rect 12572 28868 12628 28878
rect 12572 28774 12628 28812
rect 12012 28252 12180 28308
rect 12348 28642 12404 28654
rect 12348 28590 12350 28642
rect 12402 28590 12404 28642
rect 12348 28308 12404 28590
rect 12012 27300 12068 28252
rect 12348 28242 12404 28252
rect 12684 28308 12740 30156
rect 12684 28242 12740 28252
rect 12124 28084 12180 28094
rect 12124 27990 12180 28028
rect 12796 27748 12852 30604
rect 12908 30210 12964 30222
rect 12908 30158 12910 30210
rect 12962 30158 12964 30210
rect 12908 30100 12964 30158
rect 12908 30034 12964 30044
rect 13020 29540 13076 40460
rect 13356 40178 13412 40190
rect 13356 40126 13358 40178
rect 13410 40126 13412 40178
rect 13132 38834 13188 38846
rect 13132 38782 13134 38834
rect 13186 38782 13188 38834
rect 13132 38724 13188 38782
rect 13132 38658 13188 38668
rect 13356 38724 13412 40126
rect 13356 38658 13412 38668
rect 13468 40180 13524 40190
rect 13468 39620 13524 40124
rect 13132 37268 13188 37278
rect 13132 37266 13300 37268
rect 13132 37214 13134 37266
rect 13186 37214 13300 37266
rect 13132 37212 13300 37214
rect 13132 37202 13188 37212
rect 13244 33460 13300 37212
rect 13468 37154 13524 39564
rect 13580 39172 13636 39182
rect 13580 38834 13636 39116
rect 13580 38782 13582 38834
rect 13634 38782 13636 38834
rect 13580 38770 13636 38782
rect 13468 37102 13470 37154
rect 13522 37102 13524 37154
rect 13468 37090 13524 37102
rect 13580 36370 13636 36382
rect 13580 36318 13582 36370
rect 13634 36318 13636 36370
rect 13580 35698 13636 36318
rect 13580 35646 13582 35698
rect 13634 35646 13636 35698
rect 13580 35634 13636 35646
rect 13580 34018 13636 34030
rect 13580 33966 13582 34018
rect 13634 33966 13636 34018
rect 13244 33394 13300 33404
rect 13356 33908 13412 33918
rect 13244 33234 13300 33246
rect 13244 33182 13246 33234
rect 13298 33182 13300 33234
rect 13244 33124 13300 33182
rect 13244 33058 13300 33068
rect 13244 31780 13300 31790
rect 13244 30772 13300 31724
rect 13244 30436 13300 30716
rect 13356 30660 13412 33852
rect 13468 33124 13524 33134
rect 13468 31778 13524 33068
rect 13468 31726 13470 31778
rect 13522 31726 13524 31778
rect 13468 31220 13524 31726
rect 13580 31444 13636 33966
rect 13580 31378 13636 31388
rect 13468 31154 13524 31164
rect 13468 30994 13524 31006
rect 13468 30942 13470 30994
rect 13522 30942 13524 30994
rect 13468 30772 13524 30942
rect 13468 30706 13524 30716
rect 13356 30594 13412 30604
rect 13468 30548 13524 30558
rect 13244 30380 13356 30436
rect 13300 30222 13356 30380
rect 13300 30210 13412 30222
rect 13300 30158 13358 30210
rect 13410 30158 13412 30210
rect 13300 30156 13412 30158
rect 13356 30146 13412 30156
rect 13020 29474 13076 29484
rect 13020 28642 13076 28654
rect 13020 28590 13022 28642
rect 13074 28590 13076 28642
rect 13020 28084 13076 28590
rect 13468 28644 13524 30492
rect 13580 30322 13636 30334
rect 13580 30270 13582 30322
rect 13634 30270 13636 30322
rect 13580 29426 13636 30270
rect 13580 29374 13582 29426
rect 13634 29374 13636 29426
rect 13580 29362 13636 29374
rect 13580 28644 13636 28654
rect 13468 28642 13636 28644
rect 13468 28590 13582 28642
rect 13634 28590 13636 28642
rect 13468 28588 13636 28590
rect 13580 28578 13636 28588
rect 13020 28018 13076 28028
rect 13580 28308 13636 28318
rect 13468 27972 13524 27982
rect 12796 27682 12852 27692
rect 12908 27860 12964 27870
rect 12012 27298 12404 27300
rect 12012 27246 12014 27298
rect 12066 27246 12404 27298
rect 12012 27244 12404 27246
rect 12012 27234 12068 27244
rect 12124 26852 12180 26862
rect 12124 26290 12180 26796
rect 12124 26238 12126 26290
rect 12178 26238 12180 26290
rect 12124 26226 12180 26238
rect 12236 26292 12292 26302
rect 12236 24724 12292 26236
rect 12348 25844 12404 27244
rect 12572 26964 12628 26974
rect 12572 26292 12628 26908
rect 12572 26226 12628 26236
rect 12348 25788 12740 25844
rect 12124 24668 12292 24724
rect 12572 25396 12628 25406
rect 12012 23938 12068 23950
rect 12012 23886 12014 23938
rect 12066 23886 12068 23938
rect 12012 23828 12068 23886
rect 12012 23762 12068 23772
rect 11452 12178 11508 13020
rect 11564 17164 11732 17220
rect 11788 20972 11956 21028
rect 12012 22930 12068 22942
rect 12012 22878 12014 22930
rect 12066 22878 12068 22930
rect 11564 12964 11620 17164
rect 11676 16436 11732 16446
rect 11676 16322 11732 16380
rect 11676 16270 11678 16322
rect 11730 16270 11732 16322
rect 11676 16258 11732 16270
rect 11564 12898 11620 12908
rect 11452 12126 11454 12178
rect 11506 12126 11508 12178
rect 11452 12114 11508 12126
rect 11564 12738 11620 12750
rect 11564 12686 11566 12738
rect 11618 12686 11620 12738
rect 11564 11620 11620 12686
rect 11340 11564 11620 11620
rect 11340 10836 11396 11564
rect 11340 10770 11396 10780
rect 11452 11396 11508 11406
rect 11452 10612 11508 11340
rect 11676 11394 11732 11406
rect 11676 11342 11678 11394
rect 11730 11342 11732 11394
rect 11564 11282 11620 11294
rect 11564 11230 11566 11282
rect 11618 11230 11620 11282
rect 11564 10948 11620 11230
rect 11564 10882 11620 10892
rect 11676 10724 11732 11342
rect 11228 10556 11396 10612
rect 11116 10446 11118 10498
rect 11170 10446 11172 10498
rect 11116 10434 11172 10446
rect 11228 10388 11284 10398
rect 11228 10294 11284 10332
rect 11340 9826 11396 10556
rect 11452 10518 11508 10556
rect 11564 10668 11732 10724
rect 11564 10500 11620 10668
rect 11340 9774 11342 9826
rect 11394 9774 11396 9826
rect 11340 9604 11396 9774
rect 11340 9538 11396 9548
rect 11452 10052 11508 10062
rect 11004 8988 11284 9044
rect 10892 8878 10894 8930
rect 10946 8878 10948 8930
rect 10892 8866 10948 8878
rect 11116 8372 11172 8382
rect 10892 7700 10948 7710
rect 10780 7698 10948 7700
rect 10780 7646 10894 7698
rect 10946 7646 10948 7698
rect 10780 7644 10948 7646
rect 10892 7634 10948 7644
rect 10444 7298 10500 7308
rect 11004 7364 11060 7374
rect 10108 6638 10110 6690
rect 10162 6638 10164 6690
rect 10108 6626 10164 6638
rect 11004 6804 11060 7308
rect 11004 6690 11060 6748
rect 11004 6638 11006 6690
rect 11058 6638 11060 6690
rect 11004 6626 11060 6638
rect 9772 6578 9828 6590
rect 9772 6526 9774 6578
rect 9826 6526 9828 6578
rect 9772 6244 9828 6526
rect 9772 6178 9828 6188
rect 9324 6020 9380 6030
rect 9212 6018 9380 6020
rect 9212 5966 9326 6018
rect 9378 5966 9380 6018
rect 9212 5964 9380 5966
rect 9324 5954 9380 5964
rect 8876 5684 8932 5694
rect 8876 5590 8932 5628
rect 11116 5684 11172 8316
rect 11228 7252 11284 8988
rect 11452 8596 11508 9996
rect 11564 9156 11620 10444
rect 11676 10498 11732 10510
rect 11676 10446 11678 10498
rect 11730 10446 11732 10498
rect 11676 10164 11732 10446
rect 11676 10098 11732 10108
rect 11564 9090 11620 9100
rect 11452 8530 11508 8540
rect 11228 7186 11284 7196
rect 11564 6692 11620 6702
rect 11788 6692 11844 20972
rect 12012 20802 12068 22878
rect 12124 21812 12180 24668
rect 12236 24500 12292 24510
rect 12236 24162 12292 24444
rect 12236 24110 12238 24162
rect 12290 24110 12292 24162
rect 12236 24098 12292 24110
rect 12460 23940 12516 23950
rect 12348 23828 12404 23838
rect 12236 22482 12292 22494
rect 12236 22430 12238 22482
rect 12290 22430 12292 22482
rect 12236 22372 12292 22430
rect 12236 22306 12292 22316
rect 12348 21812 12404 23772
rect 12124 21756 12292 21812
rect 12124 21588 12180 21598
rect 12124 21494 12180 21532
rect 12012 20750 12014 20802
rect 12066 20750 12068 20802
rect 12012 20738 12068 20750
rect 12236 20580 12292 21756
rect 12348 21746 12404 21756
rect 12348 20804 12404 20814
rect 12348 20710 12404 20748
rect 11900 20524 12292 20580
rect 11900 12516 11956 20524
rect 12460 19460 12516 23884
rect 12572 20580 12628 25340
rect 12572 20514 12628 20524
rect 12684 20188 12740 25788
rect 12908 25508 12964 27804
rect 13020 27748 13076 27758
rect 13020 26908 13076 27692
rect 13132 27300 13188 27310
rect 13132 27206 13188 27244
rect 13468 26908 13524 27916
rect 13580 27970 13636 28252
rect 13580 27918 13582 27970
rect 13634 27918 13636 27970
rect 13580 27524 13636 27918
rect 13580 27458 13636 27468
rect 13020 26852 13188 26908
rect 13468 26852 13636 26908
rect 12908 25442 12964 25452
rect 13020 26740 13076 26750
rect 12908 25282 12964 25294
rect 12908 25230 12910 25282
rect 12962 25230 12964 25282
rect 12796 24500 12852 24510
rect 12796 24406 12852 24444
rect 12908 23938 12964 25230
rect 12908 23886 12910 23938
rect 12962 23886 12964 23938
rect 12908 23874 12964 23886
rect 13020 23044 13076 26684
rect 13132 23268 13188 26852
rect 13244 26290 13300 26302
rect 13244 26238 13246 26290
rect 13298 26238 13300 26290
rect 13244 25956 13300 26238
rect 13244 25890 13300 25900
rect 13356 24610 13412 24622
rect 13356 24558 13358 24610
rect 13410 24558 13412 24610
rect 13244 23268 13300 23278
rect 13132 23266 13300 23268
rect 13132 23214 13246 23266
rect 13298 23214 13300 23266
rect 13132 23212 13300 23214
rect 13244 23202 13300 23212
rect 13020 22988 13300 23044
rect 12684 20132 12964 20188
rect 12124 19404 12516 19460
rect 12796 20020 12852 20030
rect 12796 19906 12852 19964
rect 12796 19854 12798 19906
rect 12850 19854 12852 19906
rect 12796 19460 12852 19854
rect 12012 19348 12068 19358
rect 12012 19254 12068 19292
rect 12124 19124 12180 19404
rect 12796 19394 12852 19404
rect 12572 19348 12628 19358
rect 11900 12450 11956 12460
rect 12012 19068 12180 19124
rect 12460 19124 12516 19134
rect 12572 19124 12628 19292
rect 12796 19234 12852 19246
rect 12796 19182 12798 19234
rect 12850 19182 12852 19234
rect 12796 19124 12852 19182
rect 12572 19068 12852 19124
rect 12012 16882 12068 19068
rect 12460 19030 12516 19068
rect 12908 19012 12964 20132
rect 13132 20020 13188 20030
rect 12684 18956 12964 19012
rect 13020 20018 13188 20020
rect 13020 19966 13134 20018
rect 13186 19966 13188 20018
rect 13020 19964 13188 19966
rect 12124 18900 12180 18910
rect 12124 18674 12180 18844
rect 12124 18622 12126 18674
rect 12178 18622 12180 18674
rect 12124 18610 12180 18622
rect 12684 17892 12740 18956
rect 13020 18900 13076 19964
rect 13132 19954 13188 19964
rect 13244 19796 13300 22988
rect 13356 22820 13412 24558
rect 13468 23940 13524 23950
rect 13468 23846 13524 23884
rect 13356 22754 13412 22764
rect 13356 22596 13412 22606
rect 13356 22502 13412 22540
rect 13356 21924 13412 21934
rect 13356 20802 13412 21868
rect 13356 20750 13358 20802
rect 13410 20750 13412 20802
rect 13356 20738 13412 20750
rect 13468 21362 13524 21374
rect 13468 21310 13470 21362
rect 13522 21310 13524 21362
rect 13020 18834 13076 18844
rect 13132 19740 13300 19796
rect 13356 20580 13412 20590
rect 12684 17798 12740 17836
rect 13020 18676 13076 18686
rect 13020 18562 13076 18620
rect 13020 18510 13022 18562
rect 13074 18510 13076 18562
rect 12124 17666 12180 17678
rect 12124 17614 12126 17666
rect 12178 17614 12180 17666
rect 12124 17332 12180 17614
rect 12124 17266 12180 17276
rect 12012 16830 12014 16882
rect 12066 16830 12068 16882
rect 11900 12292 11956 12302
rect 12012 12292 12068 16830
rect 12796 16884 12852 16894
rect 12124 16548 12180 16558
rect 12124 15538 12180 16492
rect 12796 16322 12852 16828
rect 13020 16772 13076 18510
rect 13020 16706 13076 16716
rect 12796 16270 12798 16322
rect 12850 16270 12852 16322
rect 12796 16258 12852 16270
rect 13132 16100 13188 19740
rect 13244 19236 13300 19246
rect 13244 19142 13300 19180
rect 13356 18340 13412 20524
rect 13468 19458 13524 21310
rect 13580 20916 13636 26852
rect 13692 26178 13748 51548
rect 14028 43428 14084 43438
rect 13804 41186 13860 41198
rect 13804 41134 13806 41186
rect 13858 41134 13860 41186
rect 13804 40964 13860 41134
rect 13804 40898 13860 40908
rect 14028 40852 14084 43372
rect 13916 40796 14084 40852
rect 13804 38724 13860 38762
rect 13804 38658 13860 38668
rect 13916 34020 13972 40796
rect 14028 39618 14084 39630
rect 14028 39566 14030 39618
rect 14082 39566 14084 39618
rect 14028 35026 14084 39566
rect 14028 34974 14030 35026
rect 14082 34974 14084 35026
rect 14028 34962 14084 34974
rect 13916 33964 14084 34020
rect 13916 32340 13972 32350
rect 13804 30882 13860 30894
rect 13804 30830 13806 30882
rect 13858 30830 13860 30882
rect 13804 30436 13860 30830
rect 13804 30370 13860 30380
rect 13804 29988 13860 29998
rect 13804 28756 13860 29932
rect 13916 29652 13972 32284
rect 13916 29586 13972 29596
rect 14028 29538 14084 33964
rect 14028 29486 14030 29538
rect 14082 29486 14084 29538
rect 14028 29474 14084 29486
rect 13804 27074 13860 28700
rect 13916 27858 13972 27870
rect 13916 27806 13918 27858
rect 13970 27806 13972 27858
rect 13916 27300 13972 27806
rect 13916 27234 13972 27244
rect 13804 27022 13806 27074
rect 13858 27022 13860 27074
rect 13804 27010 13860 27022
rect 13916 27076 13972 27086
rect 13916 26908 13972 27020
rect 14140 26964 14196 52332
rect 14252 42084 14308 42094
rect 14252 41990 14308 42028
rect 14588 41860 14644 41870
rect 14364 41858 14644 41860
rect 14364 41806 14590 41858
rect 14642 41806 14644 41858
rect 14364 41804 14644 41806
rect 14364 41410 14420 41804
rect 14588 41794 14644 41804
rect 14364 41358 14366 41410
rect 14418 41358 14420 41410
rect 14364 38948 14420 41358
rect 14476 40964 14532 40974
rect 14476 40514 14532 40908
rect 14476 40462 14478 40514
rect 14530 40462 14532 40514
rect 14476 40450 14532 40462
rect 14924 40180 14980 40190
rect 14924 40086 14980 40124
rect 14364 38882 14420 38892
rect 14252 38836 14308 38846
rect 14252 38742 14308 38780
rect 14812 38834 14868 38846
rect 14812 38782 14814 38834
rect 14866 38782 14868 38834
rect 14812 38668 14868 38782
rect 15036 38668 15092 53452
rect 15596 41412 15652 55918
rect 16940 55468 16996 57148
rect 18172 56308 18228 57344
rect 19516 57316 19572 57344
rect 19516 57250 19572 57260
rect 19852 57316 19908 57372
rect 19852 57250 19908 57260
rect 18508 56308 18564 56318
rect 18172 56306 18564 56308
rect 18172 56254 18510 56306
rect 18562 56254 18564 56306
rect 18172 56252 18564 56254
rect 18508 56242 18564 56252
rect 20300 56306 20356 57372
rect 20832 57344 20944 57456
rect 22176 57344 22288 57456
rect 22540 57372 23044 57428
rect 20300 56254 20302 56306
rect 20354 56254 20356 56306
rect 20300 56242 20356 56254
rect 20860 56308 20916 57344
rect 22204 57204 22260 57344
rect 22540 57204 22596 57372
rect 22204 57148 22596 57204
rect 20860 56242 20916 56252
rect 21644 56644 21700 56654
rect 17500 55970 17556 55982
rect 17500 55918 17502 55970
rect 17554 55918 17556 55970
rect 16940 55412 17332 55468
rect 17276 55186 17332 55412
rect 17276 55134 17278 55186
rect 17330 55134 17332 55186
rect 17276 55122 17332 55134
rect 16828 53620 16884 53630
rect 15596 41346 15652 41356
rect 15708 44548 15764 44558
rect 14588 38612 14868 38668
rect 14924 38612 15092 38668
rect 15484 40962 15540 40974
rect 15484 40910 15486 40962
rect 15538 40910 15540 40962
rect 14364 37044 14420 37054
rect 14252 30212 14308 30222
rect 14252 30118 14308 30156
rect 14364 29540 14420 36988
rect 14476 31780 14532 31790
rect 14476 30884 14532 31724
rect 14476 30818 14532 30828
rect 14588 30548 14644 38612
rect 14700 38052 14756 38062
rect 14700 38050 14868 38052
rect 14700 37998 14702 38050
rect 14754 37998 14868 38050
rect 14700 37996 14868 37998
rect 14700 37986 14756 37996
rect 14588 30482 14644 30492
rect 14700 37042 14756 37054
rect 14700 36990 14702 37042
rect 14754 36990 14756 37042
rect 14588 30212 14644 30222
rect 13692 26126 13694 26178
rect 13746 26126 13748 26178
rect 13692 25060 13748 26126
rect 13692 24994 13748 25004
rect 13804 26852 13972 26908
rect 14028 26908 14196 26964
rect 14252 29484 14420 29540
rect 14476 30210 14644 30212
rect 14476 30158 14590 30210
rect 14642 30158 14644 30210
rect 14476 30156 14644 30158
rect 14252 27298 14308 29484
rect 14364 29316 14420 29326
rect 14476 29316 14532 30156
rect 14588 30146 14644 30156
rect 14700 29426 14756 36990
rect 14812 35586 14868 37996
rect 14812 35534 14814 35586
rect 14866 35534 14868 35586
rect 14812 32562 14868 35534
rect 14812 32510 14814 32562
rect 14866 32510 14868 32562
rect 14812 32498 14868 32510
rect 14700 29374 14702 29426
rect 14754 29374 14756 29426
rect 14700 29362 14756 29374
rect 14364 29314 14532 29316
rect 14364 29262 14366 29314
rect 14418 29262 14532 29314
rect 14364 29260 14532 29262
rect 14364 29250 14420 29260
rect 14364 27860 14420 27870
rect 14364 27766 14420 27804
rect 14252 27246 14254 27298
rect 14306 27246 14308 27298
rect 13580 20850 13636 20860
rect 13692 24612 13748 24622
rect 13468 19406 13470 19458
rect 13522 19406 13524 19458
rect 13468 19394 13524 19406
rect 13580 20020 13636 20030
rect 13580 19236 13636 19964
rect 13580 19170 13636 19180
rect 12124 15486 12126 15538
rect 12178 15486 12180 15538
rect 12124 15474 12180 15486
rect 12796 16044 13188 16100
rect 13244 18338 13412 18340
rect 13244 18286 13358 18338
rect 13410 18286 13412 18338
rect 13244 18284 13412 18286
rect 12460 15316 12516 15326
rect 12460 14754 12516 15260
rect 12796 15092 12852 16044
rect 13244 15988 13300 18284
rect 13356 18274 13412 18284
rect 13580 18228 13636 18238
rect 12796 15026 12852 15036
rect 12908 15932 13300 15988
rect 13356 17892 13412 17902
rect 12460 14702 12462 14754
rect 12514 14702 12516 14754
rect 12460 14690 12516 14702
rect 12124 14308 12180 14318
rect 12124 13746 12180 14252
rect 12908 14084 12964 15932
rect 13244 15540 13300 15550
rect 13132 14418 13188 14430
rect 13132 14366 13134 14418
rect 13186 14366 13188 14418
rect 13132 14196 13188 14366
rect 13132 14130 13188 14140
rect 12124 13694 12126 13746
rect 12178 13694 12180 13746
rect 12124 13682 12180 13694
rect 12684 14028 12964 14084
rect 12572 13076 12628 13086
rect 12572 12982 12628 13020
rect 12236 12850 12292 12862
rect 12236 12798 12238 12850
rect 12290 12798 12292 12850
rect 12236 12404 12292 12798
rect 12572 12516 12628 12526
rect 12292 12348 12516 12404
rect 12236 12338 12292 12348
rect 12012 12236 12180 12292
rect 11900 12198 11956 12236
rect 11900 11506 11956 11518
rect 11900 11454 11902 11506
rect 11954 11454 11956 11506
rect 11900 10834 11956 11454
rect 11900 10782 11902 10834
rect 11954 10782 11956 10834
rect 11900 10052 11956 10782
rect 12012 11060 12068 11070
rect 12012 10610 12068 11004
rect 12012 10558 12014 10610
rect 12066 10558 12068 10610
rect 12012 10546 12068 10558
rect 12124 10388 12180 12236
rect 12460 11394 12516 12348
rect 12460 11342 12462 11394
rect 12514 11342 12516 11394
rect 12460 11330 12516 11342
rect 12348 10612 12404 10622
rect 11900 9986 11956 9996
rect 12012 10332 12180 10388
rect 12236 10500 12292 10510
rect 12236 10386 12292 10444
rect 12236 10334 12238 10386
rect 12290 10334 12292 10386
rect 11564 6690 11844 6692
rect 11564 6638 11566 6690
rect 11618 6638 11844 6690
rect 11564 6636 11844 6638
rect 11564 6626 11620 6636
rect 11676 5908 11732 5918
rect 11676 5814 11732 5852
rect 11116 5618 11172 5628
rect 10108 3892 10164 3902
rect 8652 3332 8820 3388
rect 6860 130 6916 140
rect 7420 196 7476 206
rect 7420 112 7476 140
rect 8764 112 8820 3332
rect 10108 112 10164 3836
rect 12012 3388 12068 10332
rect 12236 10322 12292 10334
rect 12124 10052 12180 10062
rect 12124 9604 12180 9996
rect 12236 9940 12292 9950
rect 12236 9826 12292 9884
rect 12236 9774 12238 9826
rect 12290 9774 12292 9826
rect 12236 9762 12292 9774
rect 12124 9548 12292 9604
rect 12124 9380 12180 9390
rect 12124 9266 12180 9324
rect 12124 9214 12126 9266
rect 12178 9214 12180 9266
rect 12124 7474 12180 9214
rect 12236 8482 12292 9548
rect 12348 9380 12404 10556
rect 12348 9314 12404 9324
rect 12236 8430 12238 8482
rect 12290 8430 12292 8482
rect 12236 8418 12292 8430
rect 12460 9268 12516 9278
rect 12236 7700 12292 7710
rect 12236 7606 12292 7644
rect 12124 7422 12126 7474
rect 12178 7422 12180 7474
rect 12124 7410 12180 7422
rect 12236 7364 12292 7374
rect 12124 5796 12180 5806
rect 12124 5702 12180 5740
rect 12236 5346 12292 7308
rect 12348 6692 12404 6702
rect 12460 6692 12516 9212
rect 12348 6690 12516 6692
rect 12348 6638 12350 6690
rect 12402 6638 12516 6690
rect 12348 6636 12516 6638
rect 12348 6626 12404 6636
rect 12236 5294 12238 5346
rect 12290 5294 12292 5346
rect 12236 5282 12292 5294
rect 12572 3388 12628 12460
rect 12684 11396 12740 14028
rect 12684 11330 12740 11340
rect 12796 13858 12852 13870
rect 12796 13806 12798 13858
rect 12850 13806 12852 13858
rect 12796 11060 12852 13806
rect 13132 13636 13188 13646
rect 13020 13634 13188 13636
rect 13020 13582 13134 13634
rect 13186 13582 13188 13634
rect 13020 13580 13188 13582
rect 12908 13522 12964 13534
rect 12908 13470 12910 13522
rect 12962 13470 12964 13522
rect 12908 13300 12964 13470
rect 12908 11508 12964 13244
rect 13020 11732 13076 13580
rect 13132 13570 13188 13580
rect 13244 12290 13300 15484
rect 13244 12238 13246 12290
rect 13298 12238 13300 12290
rect 13244 12226 13300 12238
rect 13020 11666 13076 11676
rect 12908 11442 12964 11452
rect 13020 11506 13076 11518
rect 13020 11454 13022 11506
rect 13074 11454 13076 11506
rect 12796 10994 12852 11004
rect 13020 11396 13076 11454
rect 13020 11060 13076 11340
rect 13020 10994 13076 11004
rect 13244 10836 13300 10846
rect 13244 10722 13300 10780
rect 13244 10670 13246 10722
rect 13298 10670 13300 10722
rect 13244 10658 13300 10670
rect 12796 10610 12852 10622
rect 12796 10558 12798 10610
rect 12850 10558 12852 10610
rect 12684 10052 12740 10062
rect 12796 10052 12852 10558
rect 13020 10610 13076 10622
rect 13020 10558 13022 10610
rect 13074 10558 13076 10610
rect 13020 10500 13076 10558
rect 13020 10434 13076 10444
rect 12684 10050 12852 10052
rect 12684 9998 12686 10050
rect 12738 9998 12852 10050
rect 12684 9996 12852 9998
rect 13132 10052 13188 10062
rect 12684 9986 12740 9996
rect 13132 9938 13188 9996
rect 13132 9886 13134 9938
rect 13186 9886 13188 9938
rect 13132 9828 13188 9886
rect 13132 9762 13188 9772
rect 13244 9826 13300 9838
rect 13244 9774 13246 9826
rect 13298 9774 13300 9826
rect 12796 9268 12852 9278
rect 12796 9042 12852 9212
rect 12796 8990 12798 9042
rect 12850 8990 12852 9042
rect 12796 8978 12852 8990
rect 13020 9042 13076 9054
rect 13020 8990 13022 9042
rect 13074 8990 13076 9042
rect 12796 8484 12852 8494
rect 12796 8258 12852 8428
rect 12796 8206 12798 8258
rect 12850 8206 12852 8258
rect 12796 8194 12852 8206
rect 13020 7586 13076 8990
rect 13020 7534 13022 7586
rect 13074 7534 13076 7586
rect 13020 7522 13076 7534
rect 13132 8484 13188 8494
rect 12684 6804 12740 6814
rect 12684 6710 12740 6748
rect 12796 5348 12852 5358
rect 12796 5234 12852 5292
rect 12796 5182 12798 5234
rect 12850 5182 12852 5234
rect 12796 5170 12852 5182
rect 13132 5124 13188 8428
rect 13244 7700 13300 9774
rect 13244 7634 13300 7644
rect 13356 8370 13412 17836
rect 13468 16772 13524 16782
rect 13468 16098 13524 16716
rect 13468 16046 13470 16098
rect 13522 16046 13524 16098
rect 13468 16034 13524 16046
rect 13580 14754 13636 18172
rect 13580 14702 13582 14754
rect 13634 14702 13636 14754
rect 13580 14690 13636 14702
rect 13468 14196 13524 14206
rect 13468 12964 13524 14140
rect 13468 12898 13524 12908
rect 13692 13634 13748 24556
rect 13804 23604 13860 26852
rect 13804 23538 13860 23548
rect 13916 26740 13972 26750
rect 13804 22930 13860 22942
rect 13804 22878 13806 22930
rect 13858 22878 13860 22930
rect 13804 19906 13860 22878
rect 13804 19854 13806 19906
rect 13858 19854 13860 19906
rect 13804 19842 13860 19854
rect 13916 19796 13972 26684
rect 14028 26516 14084 26908
rect 14252 26740 14308 27246
rect 14476 26908 14532 29260
rect 14700 28642 14756 28654
rect 14700 28590 14702 28642
rect 14754 28590 14756 28642
rect 14252 26674 14308 26684
rect 14364 26852 14532 26908
rect 14588 27634 14644 27646
rect 14588 27582 14590 27634
rect 14642 27582 14644 27634
rect 14028 26460 14196 26516
rect 14028 25060 14084 25070
rect 14028 21700 14084 25004
rect 14140 22148 14196 26460
rect 14252 26404 14308 26414
rect 14252 24388 14308 26348
rect 14252 24322 14308 24332
rect 14364 24164 14420 26852
rect 14588 26292 14644 27582
rect 14588 26226 14644 26236
rect 14476 25956 14532 25966
rect 14476 25506 14532 25900
rect 14476 25454 14478 25506
rect 14530 25454 14532 25506
rect 14476 25442 14532 25454
rect 14588 24612 14644 24622
rect 14588 24518 14644 24556
rect 14700 24388 14756 28590
rect 14924 26908 14980 38612
rect 15148 38052 15204 38062
rect 15148 37958 15204 37996
rect 15484 37266 15540 40910
rect 15484 37214 15486 37266
rect 15538 37214 15540 37266
rect 15484 37202 15540 37214
rect 15596 39060 15652 39070
rect 15148 37156 15204 37166
rect 15148 37154 15316 37156
rect 15148 37102 15150 37154
rect 15202 37102 15316 37154
rect 15148 37100 15316 37102
rect 15148 37090 15204 37100
rect 15036 30884 15092 30894
rect 15036 30790 15092 30828
rect 14812 26852 14980 26908
rect 15148 29426 15204 29438
rect 15148 29374 15150 29426
rect 15202 29374 15204 29426
rect 14812 26404 14868 26852
rect 14812 26338 14868 26348
rect 14812 26066 14868 26078
rect 14812 26014 14814 26066
rect 14866 26014 14868 26066
rect 14812 24724 14868 26014
rect 14924 25618 14980 25630
rect 14924 25566 14926 25618
rect 14978 25566 14980 25618
rect 14924 25508 14980 25566
rect 14924 25442 14980 25452
rect 14924 24724 14980 24734
rect 14812 24722 14980 24724
rect 14812 24670 14926 24722
rect 14978 24670 14980 24722
rect 14812 24668 14980 24670
rect 14924 24658 14980 24668
rect 14700 24322 14756 24332
rect 15036 24612 15092 24622
rect 14252 24108 14420 24164
rect 14252 23548 14308 24108
rect 14364 23940 14420 23950
rect 14364 23846 14420 23884
rect 14252 23492 14420 23548
rect 14140 22082 14196 22092
rect 14028 21634 14084 21644
rect 14028 21476 14084 21486
rect 14028 21382 14084 21420
rect 14364 21476 14420 23492
rect 14700 23156 14756 23166
rect 14476 22260 14532 22270
rect 14476 22258 14644 22260
rect 14476 22206 14478 22258
rect 14530 22206 14644 22258
rect 14476 22204 14644 22206
rect 14476 22194 14532 22204
rect 14476 21476 14532 21486
rect 14364 21474 14532 21476
rect 14364 21422 14478 21474
rect 14530 21422 14532 21474
rect 14364 21420 14532 21422
rect 13916 19730 13972 19740
rect 13916 19236 13972 19246
rect 13804 19234 13972 19236
rect 13804 19182 13918 19234
rect 13970 19182 13972 19234
rect 13804 19180 13972 19182
rect 13804 17890 13860 19180
rect 13916 19170 13972 19180
rect 14364 19012 14420 21420
rect 14476 21410 14532 21420
rect 14476 20804 14532 20814
rect 14588 20804 14644 22204
rect 14700 22036 14756 23100
rect 14812 22484 14868 22494
rect 14812 22390 14868 22428
rect 14700 21970 14756 21980
rect 14812 21588 14868 21598
rect 14812 21494 14868 21532
rect 14812 20916 14868 20926
rect 14812 20822 14868 20860
rect 14476 20802 14644 20804
rect 14476 20750 14478 20802
rect 14530 20750 14644 20802
rect 14476 20748 14644 20750
rect 14476 20738 14532 20748
rect 14588 20244 14644 20748
rect 15036 20188 15092 24556
rect 15148 24276 15204 29374
rect 15260 28980 15316 37100
rect 15596 35028 15652 39004
rect 15708 38162 15764 44492
rect 15820 41748 15876 41758
rect 15820 41746 15988 41748
rect 15820 41694 15822 41746
rect 15874 41694 15988 41746
rect 15820 41692 15988 41694
rect 15820 41682 15876 41692
rect 15708 38110 15710 38162
rect 15762 38110 15764 38162
rect 15708 38098 15764 38110
rect 15820 38834 15876 38846
rect 15820 38782 15822 38834
rect 15874 38782 15876 38834
rect 15596 33684 15652 34972
rect 15596 33234 15652 33628
rect 15596 33182 15598 33234
rect 15650 33182 15652 33234
rect 15596 33170 15652 33182
rect 15596 32676 15652 32686
rect 15596 32582 15652 32620
rect 15820 32228 15876 38782
rect 15932 38668 15988 41692
rect 16044 40180 16100 40190
rect 16044 40178 16660 40180
rect 16044 40126 16046 40178
rect 16098 40126 16660 40178
rect 16044 40124 16660 40126
rect 16044 40114 16100 40124
rect 15932 38612 16100 38668
rect 15932 37268 15988 37278
rect 15932 37174 15988 37212
rect 15596 32172 15876 32228
rect 15484 30882 15540 30894
rect 15484 30830 15486 30882
rect 15538 30830 15540 30882
rect 15484 29428 15540 30830
rect 15484 29362 15540 29372
rect 15372 29204 15428 29214
rect 15372 29202 15540 29204
rect 15372 29150 15374 29202
rect 15426 29150 15540 29202
rect 15372 29148 15540 29150
rect 15372 29138 15428 29148
rect 15260 28914 15316 28924
rect 15484 28866 15540 29148
rect 15484 28814 15486 28866
rect 15538 28814 15540 28866
rect 15484 28802 15540 28814
rect 15596 28084 15652 32172
rect 15932 31668 15988 31678
rect 15820 30996 15876 31006
rect 15820 30902 15876 30940
rect 15708 30212 15764 30222
rect 15708 30118 15764 30156
rect 15484 28028 15652 28084
rect 15708 28980 15764 28990
rect 15260 27858 15316 27870
rect 15260 27806 15262 27858
rect 15314 27806 15316 27858
rect 15260 27300 15316 27806
rect 15372 27300 15428 27310
rect 15260 27298 15428 27300
rect 15260 27246 15374 27298
rect 15426 27246 15428 27298
rect 15260 27244 15428 27246
rect 15372 27234 15428 27244
rect 15484 26908 15540 28028
rect 15372 26852 15540 26908
rect 15260 26292 15316 26302
rect 15260 26198 15316 26236
rect 15372 24948 15428 26852
rect 15260 24892 15428 24948
rect 15484 25284 15540 25294
rect 15260 24388 15316 24892
rect 15372 24722 15428 24734
rect 15372 24670 15374 24722
rect 15426 24670 15428 24722
rect 15372 24612 15428 24670
rect 15372 24546 15428 24556
rect 15260 24332 15428 24388
rect 15204 24220 15316 24276
rect 15148 24210 15204 24220
rect 15148 23492 15204 23502
rect 15148 23044 15204 23436
rect 15148 22950 15204 22988
rect 14588 20178 14644 20188
rect 14700 20132 15092 20188
rect 15148 21812 15204 21822
rect 14476 20020 14532 20030
rect 14700 20020 14756 20132
rect 14476 20018 14644 20020
rect 14476 19966 14478 20018
rect 14530 19966 14644 20018
rect 14476 19964 14644 19966
rect 14476 19954 14532 19964
rect 14476 19572 14532 19582
rect 14476 19234 14532 19516
rect 14476 19182 14478 19234
rect 14530 19182 14532 19234
rect 14476 19170 14532 19182
rect 14364 18956 14532 19012
rect 13804 17838 13806 17890
rect 13858 17838 13860 17890
rect 13804 17826 13860 17838
rect 14364 16996 14420 17006
rect 13804 16210 13860 16222
rect 13804 16158 13806 16210
rect 13858 16158 13860 16210
rect 13804 15204 13860 16158
rect 14364 15314 14420 16940
rect 14364 15262 14366 15314
rect 14418 15262 14420 15314
rect 14364 15250 14420 15262
rect 13804 14868 13860 15148
rect 14028 15092 14084 15102
rect 14028 15090 14308 15092
rect 14028 15038 14030 15090
rect 14082 15038 14308 15090
rect 14028 15036 14308 15038
rect 14028 15026 14084 15036
rect 13804 14802 13860 14812
rect 14140 13746 14196 13758
rect 14140 13694 14142 13746
rect 14194 13694 14196 13746
rect 13692 13582 13694 13634
rect 13746 13582 13748 13634
rect 13692 12740 13748 13582
rect 13804 13636 13860 13646
rect 13804 13186 13860 13580
rect 13804 13134 13806 13186
rect 13858 13134 13860 13186
rect 13804 13122 13860 13134
rect 13692 11844 13748 12684
rect 14028 12964 14084 12974
rect 14028 12180 14084 12908
rect 14028 12086 14084 12124
rect 13692 11788 14084 11844
rect 13468 10612 13524 10622
rect 13468 10610 13972 10612
rect 13468 10558 13470 10610
rect 13522 10558 13972 10610
rect 13468 10556 13972 10558
rect 13468 10546 13524 10556
rect 13580 10386 13636 10398
rect 13580 10334 13582 10386
rect 13634 10334 13636 10386
rect 13356 8318 13358 8370
rect 13410 8318 13412 8370
rect 13356 7364 13412 8318
rect 13468 9826 13524 9838
rect 13468 9774 13470 9826
rect 13522 9774 13524 9826
rect 13468 8036 13524 9774
rect 13468 7970 13524 7980
rect 13580 7476 13636 10334
rect 13692 10388 13748 10398
rect 13692 10294 13748 10332
rect 13580 7410 13636 7420
rect 13692 10052 13748 10062
rect 13356 7270 13412 7308
rect 13692 5908 13748 9996
rect 13916 10050 13972 10556
rect 13916 9998 13918 10050
rect 13970 9998 13972 10050
rect 13916 9986 13972 9998
rect 13804 9828 13860 9838
rect 14028 9828 14084 11788
rect 14140 11618 14196 13694
rect 14140 11566 14142 11618
rect 14194 11566 14196 11618
rect 14140 11554 14196 11566
rect 14252 9828 14308 15036
rect 14364 14980 14420 14990
rect 14364 13748 14420 14924
rect 14476 14196 14532 18956
rect 14588 18674 14644 19964
rect 14700 19954 14756 19964
rect 14812 20018 14868 20030
rect 14812 19966 14814 20018
rect 14866 19966 14868 20018
rect 14812 19908 14868 19966
rect 14812 19572 14868 19852
rect 14812 19506 14868 19516
rect 14924 20020 14980 20030
rect 14588 18622 14590 18674
rect 14642 18622 14644 18674
rect 14588 18610 14644 18622
rect 14700 18452 14756 18462
rect 14700 17108 14756 18396
rect 14700 16770 14756 17052
rect 14700 16718 14702 16770
rect 14754 16718 14756 16770
rect 14700 15204 14756 16718
rect 14924 15540 14980 19964
rect 15148 17778 15204 21756
rect 15260 21586 15316 24220
rect 15372 22372 15428 24332
rect 15484 24164 15540 25228
rect 15596 24612 15652 24622
rect 15596 24518 15652 24556
rect 15484 24108 15652 24164
rect 15372 21924 15428 22316
rect 15372 21858 15428 21868
rect 15484 23938 15540 23950
rect 15484 23886 15486 23938
rect 15538 23886 15540 23938
rect 15260 21534 15262 21586
rect 15314 21534 15316 21586
rect 15260 20692 15316 21534
rect 15260 20626 15316 20636
rect 15372 21476 15428 21486
rect 15148 17726 15150 17778
rect 15202 17726 15204 17778
rect 15148 17714 15204 17726
rect 15036 16884 15092 16894
rect 15036 16790 15092 16828
rect 15036 15876 15092 15886
rect 15036 15782 15092 15820
rect 14924 15474 14980 15484
rect 15148 15316 15204 15326
rect 15148 15222 15204 15260
rect 14700 15202 14868 15204
rect 14700 15150 14702 15202
rect 14754 15150 14868 15202
rect 14700 15148 14868 15150
rect 14700 15138 14756 15148
rect 14700 14644 14756 14654
rect 14700 14550 14756 14588
rect 14476 14130 14532 14140
rect 14700 14420 14756 14430
rect 14588 13748 14644 13758
rect 14364 13746 14644 13748
rect 14364 13694 14590 13746
rect 14642 13694 14644 13746
rect 14364 13692 14644 13694
rect 14364 12964 14420 12974
rect 14364 12870 14420 12908
rect 14588 10500 14644 13692
rect 14700 13634 14756 14364
rect 14812 13748 14868 15148
rect 15372 15148 15428 21420
rect 15484 21474 15540 23886
rect 15484 21422 15486 21474
rect 15538 21422 15540 21474
rect 15484 21410 15540 21422
rect 15484 19348 15540 19358
rect 15484 19234 15540 19292
rect 15484 19182 15486 19234
rect 15538 19182 15540 19234
rect 15484 19170 15540 19182
rect 15596 19012 15652 24108
rect 15708 19796 15764 28924
rect 15820 27860 15876 27870
rect 15932 27860 15988 31612
rect 16044 29426 16100 38612
rect 16380 38610 16436 38622
rect 16380 38558 16382 38610
rect 16434 38558 16436 38610
rect 16380 37716 16436 38558
rect 16380 37650 16436 37660
rect 16604 37266 16660 40124
rect 16604 37214 16606 37266
rect 16658 37214 16660 37266
rect 16604 37202 16660 37214
rect 16156 37042 16212 37054
rect 16156 36990 16158 37042
rect 16210 36990 16212 37042
rect 16156 36708 16212 36990
rect 16156 36642 16212 36652
rect 16268 37044 16324 37054
rect 16268 34132 16324 36988
rect 16716 36708 16772 36718
rect 16716 36614 16772 36652
rect 16044 29374 16046 29426
rect 16098 29374 16100 29426
rect 16044 29362 16100 29374
rect 16156 34076 16324 34132
rect 16380 34916 16436 34926
rect 16044 28644 16100 28654
rect 16044 28550 16100 28588
rect 15820 27858 15988 27860
rect 15820 27806 15822 27858
rect 15874 27806 15988 27858
rect 15820 27804 15988 27806
rect 15820 27794 15876 27804
rect 15820 26180 15876 26190
rect 15820 26086 15876 26124
rect 16044 25282 16100 25294
rect 16044 25230 16046 25282
rect 16098 25230 16100 25282
rect 16044 24722 16100 25230
rect 16044 24670 16046 24722
rect 16098 24670 16100 24722
rect 16044 24658 16100 24670
rect 16044 24500 16100 24510
rect 15820 24388 15876 24398
rect 15820 20020 15876 24332
rect 16044 24050 16100 24444
rect 16044 23998 16046 24050
rect 16098 23998 16100 24050
rect 16044 23986 16100 23998
rect 16044 22148 16100 22158
rect 16044 22054 16100 22092
rect 16156 21812 16212 34076
rect 16268 33908 16324 33918
rect 16380 33908 16436 34860
rect 16268 33906 16436 33908
rect 16268 33854 16270 33906
rect 16322 33854 16436 33906
rect 16268 33852 16436 33854
rect 16268 33842 16324 33852
rect 16380 30994 16436 33852
rect 16716 31780 16772 31790
rect 16380 30942 16382 30994
rect 16434 30942 16436 30994
rect 16380 26852 16436 30942
rect 16492 31778 16772 31780
rect 16492 31726 16718 31778
rect 16770 31726 16772 31778
rect 16492 31724 16772 31726
rect 16492 30882 16548 31724
rect 16716 31714 16772 31724
rect 16492 30830 16494 30882
rect 16546 30830 16548 30882
rect 16492 30818 16548 30830
rect 16268 25732 16324 25742
rect 16268 23604 16324 25676
rect 16380 25284 16436 26796
rect 16380 25218 16436 25228
rect 16492 30212 16548 30222
rect 16492 29426 16548 30156
rect 16828 29764 16884 53564
rect 16940 46564 16996 46574
rect 16940 38946 16996 46508
rect 17276 42980 17332 42990
rect 17052 41860 17108 41870
rect 17052 39284 17108 41804
rect 17052 39218 17108 39228
rect 16940 38894 16942 38946
rect 16994 38894 16996 38946
rect 16940 38882 16996 38894
rect 17164 37380 17220 37390
rect 17164 37266 17220 37324
rect 17164 37214 17166 37266
rect 17218 37214 17220 37266
rect 17164 37202 17220 37214
rect 17276 36594 17332 42924
rect 17500 37828 17556 55918
rect 19516 55972 19572 55982
rect 19516 55878 19572 55916
rect 21308 55972 21364 55982
rect 21308 55878 21364 55916
rect 19516 55748 19572 55758
rect 18284 55300 18340 55310
rect 18284 55206 18340 55244
rect 19516 54626 19572 55692
rect 21644 55410 21700 56588
rect 22204 56308 22260 56318
rect 22204 56214 22260 56252
rect 21644 55358 21646 55410
rect 21698 55358 21700 55410
rect 21644 55346 21700 55358
rect 21756 56082 21812 56094
rect 21756 56030 21758 56082
rect 21810 56030 21812 56082
rect 20076 55298 20132 55310
rect 20076 55246 20078 55298
rect 20130 55246 20132 55298
rect 20076 55188 20132 55246
rect 20524 55300 20580 55310
rect 20524 55206 20580 55244
rect 20860 55300 20916 55310
rect 20860 55206 20916 55244
rect 20076 55122 20132 55132
rect 19516 54574 19518 54626
rect 19570 54574 19572 54626
rect 19516 54562 19572 54574
rect 21196 54516 21252 54526
rect 21196 54422 21252 54460
rect 21532 54402 21588 54414
rect 21532 54350 21534 54402
rect 21586 54350 21588 54402
rect 19068 54292 19124 54302
rect 19068 54198 19124 54236
rect 20636 54290 20692 54302
rect 20636 54238 20638 54290
rect 20690 54238 20692 54290
rect 20524 54180 20580 54190
rect 20076 52836 20132 52846
rect 19740 47460 19796 47470
rect 17724 44436 17780 44446
rect 17724 43708 17780 44380
rect 17724 43652 18004 43708
rect 17500 37762 17556 37772
rect 17612 39620 17668 39630
rect 17276 36542 17278 36594
rect 17330 36542 17332 36594
rect 17276 36530 17332 36542
rect 17612 35476 17668 39564
rect 17948 38668 18004 43652
rect 19180 43540 19236 43550
rect 18284 41972 18340 41982
rect 18284 38668 18340 41916
rect 17836 38612 18004 38668
rect 18060 38612 18340 38668
rect 18396 40180 18452 40190
rect 17164 35420 17668 35476
rect 17724 36482 17780 36494
rect 17724 36430 17726 36482
rect 17778 36430 17780 36482
rect 17164 31666 17220 35420
rect 17500 35252 17556 35262
rect 17500 34914 17556 35196
rect 17500 34862 17502 34914
rect 17554 34862 17556 34914
rect 17500 34804 17556 34862
rect 17500 34738 17556 34748
rect 17164 31614 17166 31666
rect 17218 31614 17220 31666
rect 17164 31602 17220 31614
rect 17276 34132 17332 34142
rect 17724 34132 17780 36430
rect 17276 34130 17780 34132
rect 17276 34078 17278 34130
rect 17330 34078 17780 34130
rect 17276 34076 17780 34078
rect 17836 34132 17892 38612
rect 17948 35028 18004 35038
rect 18060 35028 18116 38612
rect 17948 35026 18116 35028
rect 17948 34974 17950 35026
rect 18002 34974 18116 35026
rect 17948 34972 18116 34974
rect 18172 37266 18228 37278
rect 18172 37214 18174 37266
rect 18226 37214 18228 37266
rect 17948 34962 18004 34972
rect 18060 34804 18116 34814
rect 18060 34244 18116 34748
rect 17836 34076 18004 34132
rect 16940 30884 16996 30894
rect 16940 30790 16996 30828
rect 17052 30100 17108 30110
rect 17052 30006 17108 30044
rect 17276 29988 17332 34076
rect 17836 33906 17892 33918
rect 17836 33854 17838 33906
rect 17890 33854 17892 33906
rect 17500 33684 17556 33694
rect 17388 32788 17444 32798
rect 17388 30322 17444 32732
rect 17388 30270 17390 30322
rect 17442 30270 17444 30322
rect 17388 30258 17444 30270
rect 17500 30994 17556 33628
rect 17836 33460 17892 33854
rect 17836 32788 17892 33404
rect 17836 32722 17892 32732
rect 17948 32340 18004 34076
rect 17948 32274 18004 32284
rect 18060 32228 18116 34188
rect 18060 32162 18116 32172
rect 18172 32004 18228 37214
rect 18284 36594 18340 36606
rect 18284 36542 18286 36594
rect 18338 36542 18340 36594
rect 18284 35252 18340 36542
rect 18284 35186 18340 35196
rect 18284 35028 18340 35038
rect 18284 34934 18340 34972
rect 17500 30942 17502 30994
rect 17554 30942 17556 30994
rect 17500 30212 17556 30942
rect 17724 31948 18228 32004
rect 18284 33346 18340 33358
rect 18284 33294 18286 33346
rect 18338 33294 18340 33346
rect 17724 30212 17780 31948
rect 18060 31780 18116 31790
rect 18284 31780 18340 33294
rect 17500 30146 17556 30156
rect 17612 30156 17780 30212
rect 17948 31778 18340 31780
rect 17948 31726 18062 31778
rect 18114 31726 18340 31778
rect 17948 31724 18340 31726
rect 17276 29922 17332 29932
rect 16828 29708 17108 29764
rect 16492 29374 16494 29426
rect 16546 29374 16548 29426
rect 16268 23548 16436 23604
rect 16268 23380 16324 23390
rect 16268 23286 16324 23324
rect 16156 21746 16212 21756
rect 16156 21588 16212 21598
rect 16156 21494 16212 21532
rect 16044 20804 16100 20814
rect 16044 20710 16100 20748
rect 15820 20018 15988 20020
rect 15820 19966 15822 20018
rect 15874 19966 15988 20018
rect 15820 19964 15988 19966
rect 15820 19954 15876 19964
rect 15708 19740 15876 19796
rect 15484 18956 15652 19012
rect 15484 16882 15540 18956
rect 15708 18452 15764 18462
rect 15596 18450 15764 18452
rect 15596 18398 15710 18450
rect 15762 18398 15764 18450
rect 15596 18396 15764 18398
rect 15596 17332 15652 18396
rect 15708 18386 15764 18396
rect 15596 17266 15652 17276
rect 15708 17666 15764 17678
rect 15708 17614 15710 17666
rect 15762 17614 15764 17666
rect 15484 16830 15486 16882
rect 15538 16830 15540 16882
rect 15484 15314 15540 16830
rect 15708 16770 15764 17614
rect 15708 16718 15710 16770
rect 15762 16718 15764 16770
rect 15708 16706 15764 16718
rect 15484 15262 15486 15314
rect 15538 15262 15540 15314
rect 15484 15250 15540 15262
rect 15596 16098 15652 16110
rect 15596 16046 15598 16098
rect 15650 16046 15652 16098
rect 15596 15204 15652 16046
rect 15708 15204 15764 15214
rect 15596 15202 15764 15204
rect 15596 15150 15710 15202
rect 15762 15150 15764 15202
rect 15596 15148 15764 15150
rect 15372 15092 15540 15148
rect 15708 15138 15764 15148
rect 15148 14532 15204 14542
rect 15092 14530 15204 14532
rect 15092 14478 15150 14530
rect 15202 14478 15204 14530
rect 15092 14466 15204 14478
rect 15092 14430 15148 14466
rect 15036 14420 15148 14430
rect 15092 14364 15148 14420
rect 15036 14354 15092 14364
rect 14812 13682 14868 13692
rect 15260 14084 15316 14094
rect 14700 13582 14702 13634
rect 14754 13582 14756 13634
rect 14700 13570 14756 13582
rect 15148 13636 15204 13646
rect 15148 13542 15204 13580
rect 15036 13524 15092 13534
rect 14924 13188 14980 13198
rect 14924 13094 14980 13132
rect 14812 12180 14868 12190
rect 14700 10724 14756 10734
rect 14812 10724 14868 12124
rect 14700 10722 14812 10724
rect 14700 10670 14702 10722
rect 14754 10670 14812 10722
rect 14700 10668 14812 10670
rect 14700 10658 14756 10668
rect 14588 10444 14756 10500
rect 13804 9734 13860 9772
rect 13916 9772 14084 9828
rect 14140 9772 14308 9828
rect 13804 9268 13860 9278
rect 13804 9174 13860 9212
rect 13916 9044 13972 9772
rect 14028 9602 14084 9614
rect 14028 9550 14030 9602
rect 14082 9550 14084 9602
rect 14028 9380 14084 9550
rect 14028 9314 14084 9324
rect 13804 8988 13972 9044
rect 13804 6018 13860 8988
rect 13916 8484 13972 8494
rect 13916 6914 13972 8428
rect 13916 6862 13918 6914
rect 13970 6862 13972 6914
rect 13916 6850 13972 6862
rect 14140 6132 14196 9772
rect 14252 9602 14308 9614
rect 14252 9550 14254 9602
rect 14306 9550 14308 9602
rect 14252 7812 14308 9550
rect 14252 7746 14308 7756
rect 14476 8034 14532 8046
rect 14476 7982 14478 8034
rect 14530 7982 14532 8034
rect 14140 6066 14196 6076
rect 13804 5966 13806 6018
rect 13858 5966 13860 6018
rect 13804 5954 13860 5966
rect 13692 5234 13748 5852
rect 14252 5908 14308 5918
rect 14476 5908 14532 7982
rect 14588 7476 14644 7486
rect 14588 7382 14644 7420
rect 14252 5906 14532 5908
rect 14252 5854 14254 5906
rect 14306 5854 14532 5906
rect 14252 5852 14532 5854
rect 14700 5906 14756 10444
rect 14812 9268 14868 10668
rect 15036 10498 15092 13468
rect 15260 12066 15316 14028
rect 15260 12014 15262 12066
rect 15314 12014 15316 12066
rect 15260 12002 15316 12014
rect 15372 11172 15428 11182
rect 15036 10446 15038 10498
rect 15090 10446 15092 10498
rect 15036 10052 15092 10446
rect 15260 11170 15428 11172
rect 15260 11118 15374 11170
rect 15426 11118 15428 11170
rect 15260 11116 15428 11118
rect 15036 9986 15092 9996
rect 15148 10164 15204 10174
rect 15148 9938 15204 10108
rect 15148 9886 15150 9938
rect 15202 9886 15204 9938
rect 15148 9874 15204 9886
rect 14924 9828 14980 9838
rect 15260 9828 15316 11116
rect 15372 11106 15428 11116
rect 15484 11060 15540 15092
rect 15820 14868 15876 19740
rect 15932 19348 15988 19964
rect 15932 19282 15988 19292
rect 16268 19460 16324 19470
rect 16044 19234 16100 19246
rect 16044 19182 16046 19234
rect 16098 19182 16100 19234
rect 15932 19124 15988 19134
rect 16044 19124 16100 19182
rect 15988 19068 16100 19124
rect 15932 19058 15988 19068
rect 16044 18900 16100 19068
rect 16156 19124 16212 19134
rect 16156 19030 16212 19068
rect 16044 18834 16100 18844
rect 16156 17444 16212 17454
rect 16156 16882 16212 17388
rect 16156 16830 16158 16882
rect 16210 16830 16212 16882
rect 16156 16818 16212 16830
rect 15932 16660 15988 16670
rect 15932 16324 15988 16604
rect 15932 16258 15988 16268
rect 16044 16212 16100 16222
rect 16044 16118 16100 16156
rect 15596 14812 15876 14868
rect 15932 16100 15988 16110
rect 15596 13748 15652 14812
rect 15932 14756 15988 16044
rect 16156 15876 16212 15886
rect 16156 15314 16212 15820
rect 16156 15262 16158 15314
rect 16210 15262 16212 15314
rect 16156 15250 16212 15262
rect 15708 14700 15988 14756
rect 15708 14642 15764 14700
rect 15708 14590 15710 14642
rect 15762 14590 15764 14642
rect 15708 14578 15764 14590
rect 16044 14530 16100 14542
rect 16044 14478 16046 14530
rect 16098 14478 16100 14530
rect 15820 13748 15876 13758
rect 15596 13746 15876 13748
rect 15596 13694 15822 13746
rect 15874 13694 15876 13746
rect 15596 13692 15876 13694
rect 15484 10994 15540 11004
rect 15596 11732 15652 11742
rect 15596 11618 15652 11676
rect 15596 11566 15598 11618
rect 15650 11566 15652 11618
rect 15596 10388 15652 11566
rect 15596 10322 15652 10332
rect 15708 11170 15764 11182
rect 15708 11118 15710 11170
rect 15762 11118 15764 11170
rect 15372 10052 15428 10062
rect 15372 10050 15540 10052
rect 15372 9998 15374 10050
rect 15426 9998 15540 10050
rect 15372 9996 15540 9998
rect 15372 9986 15428 9996
rect 14924 9826 15092 9828
rect 14924 9774 14926 9826
rect 14978 9774 15092 9826
rect 14924 9772 15092 9774
rect 14924 9762 14980 9772
rect 14812 9042 14868 9212
rect 14812 8990 14814 9042
rect 14866 8990 14868 9042
rect 14812 8978 14868 8990
rect 15036 9716 15092 9772
rect 15260 9716 15316 9772
rect 15036 9660 15316 9716
rect 14924 8484 14980 8494
rect 15036 8484 15092 9660
rect 15372 9602 15428 9614
rect 15372 9550 15374 9602
rect 15426 9550 15428 9602
rect 15372 9492 15428 9550
rect 15372 9426 15428 9436
rect 15372 8820 15428 8830
rect 15372 8726 15428 8764
rect 14980 8428 15092 8484
rect 14924 8370 14980 8428
rect 14924 8318 14926 8370
rect 14978 8318 14980 8370
rect 14924 7364 14980 8318
rect 15036 8260 15092 8270
rect 15372 8260 15428 8270
rect 15036 8258 15428 8260
rect 15036 8206 15038 8258
rect 15090 8206 15374 8258
rect 15426 8206 15428 8258
rect 15036 8204 15428 8206
rect 15036 8194 15092 8204
rect 15372 8194 15428 8204
rect 15484 8260 15540 9996
rect 15708 9826 15764 11118
rect 15708 9774 15710 9826
rect 15762 9774 15764 9826
rect 15708 9762 15764 9774
rect 15708 9492 15764 9502
rect 15708 8370 15764 9436
rect 15820 9156 15876 13692
rect 16044 13186 16100 14478
rect 16044 13134 16046 13186
rect 16098 13134 16100 13186
rect 16044 12964 16100 13134
rect 16044 12898 16100 12908
rect 16156 14306 16212 14318
rect 16156 14254 16158 14306
rect 16210 14254 16212 14306
rect 16156 12292 16212 14254
rect 16156 12226 16212 12236
rect 16268 11172 16324 19404
rect 16380 16100 16436 23548
rect 16492 21586 16548 29374
rect 16716 29428 16772 29438
rect 16604 27860 16660 27870
rect 16604 27766 16660 27804
rect 16604 27412 16660 27422
rect 16604 24722 16660 27356
rect 16604 24670 16606 24722
rect 16658 24670 16660 24722
rect 16604 24658 16660 24670
rect 16716 27188 16772 29372
rect 16716 24276 16772 27132
rect 16940 27860 16996 27870
rect 16828 25506 16884 25518
rect 16828 25454 16830 25506
rect 16882 25454 16884 25506
rect 16828 24612 16884 25454
rect 16828 24546 16884 24556
rect 16716 24050 16772 24220
rect 16716 23998 16718 24050
rect 16770 23998 16772 24050
rect 16716 23986 16772 23998
rect 16940 23940 16996 27804
rect 17052 26908 17108 29708
rect 17500 29426 17556 29438
rect 17500 29374 17502 29426
rect 17554 29374 17556 29426
rect 17388 28532 17444 28542
rect 17388 28438 17444 28476
rect 17388 27188 17444 27198
rect 17388 27094 17444 27132
rect 17500 26908 17556 29374
rect 17612 27860 17668 30156
rect 17612 27794 17668 27804
rect 17724 29988 17780 29998
rect 17724 27074 17780 29932
rect 17836 28756 17892 28766
rect 17836 28662 17892 28700
rect 17724 27022 17726 27074
rect 17778 27022 17780 27074
rect 17724 27010 17780 27022
rect 17052 26852 17444 26908
rect 17500 26852 17892 26908
rect 17388 26628 17444 26852
rect 17388 26572 17780 26628
rect 17724 26402 17780 26572
rect 17836 26516 17892 26852
rect 17836 26450 17892 26460
rect 17724 26350 17726 26402
rect 17778 26350 17780 26402
rect 17724 26338 17780 26350
rect 17276 26066 17332 26078
rect 17276 26014 17278 26066
rect 17330 26014 17332 26066
rect 17276 25844 17332 26014
rect 17948 25956 18004 31724
rect 18060 31714 18116 31724
rect 18396 31444 18452 40124
rect 19180 38668 19236 43484
rect 19180 38612 19684 38668
rect 19404 36260 19460 36270
rect 19404 36166 19460 36204
rect 19292 35028 19348 35038
rect 19292 35026 19572 35028
rect 19292 34974 19294 35026
rect 19346 34974 19572 35026
rect 19292 34972 19572 34974
rect 19292 34962 19348 34972
rect 18732 34916 18788 34926
rect 19068 34916 19124 34926
rect 18732 34914 19012 34916
rect 18732 34862 18734 34914
rect 18786 34862 19012 34914
rect 18732 34860 19012 34862
rect 18732 34850 18788 34860
rect 18956 34354 19012 34860
rect 19068 34822 19124 34860
rect 18956 34302 18958 34354
rect 19010 34302 19012 34354
rect 18956 34290 19012 34302
rect 19516 34130 19572 34972
rect 19516 34078 19518 34130
rect 19570 34078 19572 34130
rect 19516 34066 19572 34078
rect 18732 33460 18788 33470
rect 18620 32228 18676 32238
rect 18620 31890 18676 32172
rect 18620 31838 18622 31890
rect 18674 31838 18676 31890
rect 17948 25890 18004 25900
rect 18060 31388 18452 31444
rect 18508 31668 18564 31678
rect 17276 25778 17332 25788
rect 17276 25620 17332 25630
rect 18060 25620 18116 31388
rect 18508 30996 18564 31612
rect 18508 30902 18564 30940
rect 18620 30772 18676 31838
rect 18508 30716 18676 30772
rect 18284 29876 18340 29886
rect 18172 29426 18228 29438
rect 18172 29374 18174 29426
rect 18226 29374 18228 29426
rect 18172 29316 18228 29374
rect 18172 27970 18228 29260
rect 18172 27918 18174 27970
rect 18226 27918 18228 27970
rect 18172 27906 18228 27918
rect 17276 25618 18116 25620
rect 17276 25566 17278 25618
rect 17330 25566 18116 25618
rect 17276 25564 18116 25566
rect 18172 27074 18228 27086
rect 18172 27022 18174 27074
rect 18226 27022 18228 27074
rect 17276 25554 17332 25564
rect 18172 24836 18228 27022
rect 18284 26908 18340 29820
rect 18508 28756 18564 30716
rect 18620 29988 18676 29998
rect 18620 29894 18676 29932
rect 18620 29316 18676 29326
rect 18732 29316 18788 33404
rect 19180 33460 19236 33470
rect 19180 32562 19236 33404
rect 19180 32510 19182 32562
rect 19234 32510 19236 32562
rect 19180 32498 19236 32510
rect 19628 30324 19684 38612
rect 19740 32674 19796 47404
rect 20076 43708 20132 52780
rect 19964 43652 20132 43708
rect 19852 41188 19908 41198
rect 19852 36594 19908 41132
rect 19852 36542 19854 36594
rect 19906 36542 19908 36594
rect 19852 36530 19908 36542
rect 19852 36260 19908 36270
rect 19852 34914 19908 36204
rect 19852 34862 19854 34914
rect 19906 34862 19908 34914
rect 19852 34850 19908 34862
rect 19964 33348 20020 43652
rect 20412 36482 20468 36494
rect 20412 36430 20414 36482
rect 20466 36430 20468 36482
rect 20300 34914 20356 34926
rect 20300 34862 20302 34914
rect 20354 34862 20356 34914
rect 19740 32622 19742 32674
rect 19794 32622 19796 32674
rect 19740 32610 19796 32622
rect 19852 33292 20020 33348
rect 20076 34018 20132 34030
rect 20076 33966 20078 34018
rect 20130 33966 20132 34018
rect 19740 31554 19796 31566
rect 19740 31502 19742 31554
rect 19794 31502 19796 31554
rect 19740 30996 19796 31502
rect 19740 30930 19796 30940
rect 18620 29314 18788 29316
rect 18620 29262 18622 29314
rect 18674 29262 18788 29314
rect 18620 29260 18788 29262
rect 18844 30322 19684 30324
rect 18844 30270 19630 30322
rect 19682 30270 19684 30322
rect 18844 30268 19684 30270
rect 18620 29250 18676 29260
rect 18508 27746 18564 28700
rect 18508 27694 18510 27746
rect 18562 27694 18564 27746
rect 18508 27682 18564 27694
rect 18396 27188 18452 27198
rect 18396 27186 18676 27188
rect 18396 27134 18398 27186
rect 18450 27134 18676 27186
rect 18396 27132 18676 27134
rect 18396 27122 18452 27132
rect 18284 26852 18452 26908
rect 18396 26290 18452 26852
rect 18396 26238 18398 26290
rect 18450 26238 18452 26290
rect 18396 25396 18452 26238
rect 18620 25730 18676 27132
rect 18732 26178 18788 26190
rect 18732 26126 18734 26178
rect 18786 26126 18788 26178
rect 18732 25844 18788 26126
rect 18732 25778 18788 25788
rect 18620 25678 18622 25730
rect 18674 25678 18676 25730
rect 18620 25666 18676 25678
rect 18396 25330 18452 25340
rect 18732 25508 18788 25518
rect 17612 24722 17668 24734
rect 17612 24670 17614 24722
rect 17666 24670 17668 24722
rect 17612 24500 17668 24670
rect 18172 24724 18228 24780
rect 18732 24834 18788 25452
rect 18732 24782 18734 24834
rect 18786 24782 18788 24834
rect 18732 24770 18788 24782
rect 18172 24668 18340 24724
rect 18172 24500 18228 24510
rect 17612 24434 17668 24444
rect 17724 24498 18228 24500
rect 17724 24446 18174 24498
rect 18226 24446 18228 24498
rect 17724 24444 18228 24446
rect 17724 24162 17780 24444
rect 18172 24434 18228 24444
rect 17724 24110 17726 24162
rect 17778 24110 17780 24162
rect 17724 24098 17780 24110
rect 17164 24052 17220 24062
rect 16940 23874 16996 23884
rect 17052 23938 17108 23950
rect 17052 23886 17054 23938
rect 17106 23886 17108 23938
rect 17052 23380 17108 23886
rect 17052 23314 17108 23324
rect 16492 21534 16494 21586
rect 16546 21534 16548 21586
rect 16492 21476 16548 21534
rect 16492 21410 16548 21420
rect 16604 23044 16660 23054
rect 16492 20020 16548 20030
rect 16492 19926 16548 19964
rect 16604 18564 16660 22988
rect 16828 22146 16884 22158
rect 16828 22094 16830 22146
rect 16882 22094 16884 22146
rect 16828 21588 16884 22094
rect 16828 21522 16884 21532
rect 16828 21364 16884 21374
rect 17164 21364 17220 23996
rect 17612 23938 17668 23950
rect 17612 23886 17614 23938
rect 17666 23886 17668 23938
rect 17612 23604 17668 23886
rect 17612 23538 17668 23548
rect 18172 23938 18228 23950
rect 18172 23886 18174 23938
rect 18226 23886 18228 23938
rect 18172 22596 18228 23886
rect 18284 23604 18340 24668
rect 18844 24052 18900 30268
rect 19628 30258 19684 30268
rect 19292 30100 19348 30110
rect 19292 30006 19348 30044
rect 19852 29428 19908 33292
rect 19964 33122 20020 33134
rect 19964 33070 19966 33122
rect 20018 33070 20020 33122
rect 19964 31220 20020 33070
rect 19964 31154 20020 31164
rect 19852 29362 19908 29372
rect 19740 29204 19796 29214
rect 19068 29202 19796 29204
rect 19068 29150 19742 29202
rect 19794 29150 19796 29202
rect 19068 29148 19796 29150
rect 18956 28418 19012 28430
rect 18956 28366 18958 28418
rect 19010 28366 19012 28418
rect 18956 27074 19012 28366
rect 18956 27022 18958 27074
rect 19010 27022 19012 27074
rect 18956 27010 19012 27022
rect 18844 23986 18900 23996
rect 18284 23538 18340 23548
rect 18620 23940 18676 23950
rect 18172 22530 18228 22540
rect 18396 23156 18452 23166
rect 18060 22484 18116 22494
rect 18060 22390 18116 22428
rect 18396 22370 18452 23100
rect 18396 22318 18398 22370
rect 18450 22318 18452 22370
rect 18396 22306 18452 22318
rect 16884 21308 17220 21364
rect 17276 21700 17332 21710
rect 18172 21700 18228 21710
rect 16828 21298 16884 21308
rect 16940 20914 16996 20926
rect 16940 20862 16942 20914
rect 16994 20862 16996 20914
rect 16828 20804 16884 20814
rect 16828 20710 16884 20748
rect 16940 19460 16996 20862
rect 17052 19906 17108 21308
rect 17276 20914 17332 21644
rect 17724 21698 18228 21700
rect 17724 21646 18174 21698
rect 18226 21646 18228 21698
rect 17724 21644 18228 21646
rect 17276 20862 17278 20914
rect 17330 20862 17332 20914
rect 17276 20850 17332 20862
rect 17388 21588 17444 21598
rect 17052 19854 17054 19906
rect 17106 19854 17108 19906
rect 17052 19842 17108 19854
rect 17164 20802 17220 20814
rect 17164 20750 17166 20802
rect 17218 20750 17220 20802
rect 16828 19404 16996 19460
rect 16716 19348 16772 19358
rect 16716 18676 16772 19292
rect 16716 18610 16772 18620
rect 16604 18498 16660 18508
rect 16716 18452 16772 18462
rect 16828 18452 16884 19404
rect 16940 19236 16996 19246
rect 17164 19236 17220 20750
rect 17388 19458 17444 21532
rect 17612 21586 17668 21598
rect 17612 21534 17614 21586
rect 17666 21534 17668 21586
rect 17612 21364 17668 21534
rect 17612 21298 17668 21308
rect 17612 20578 17668 20590
rect 17612 20526 17614 20578
rect 17666 20526 17668 20578
rect 17612 19908 17668 20526
rect 17612 19842 17668 19852
rect 17388 19406 17390 19458
rect 17442 19406 17444 19458
rect 17388 19394 17444 19406
rect 16940 19234 17220 19236
rect 16940 19182 16942 19234
rect 16994 19182 17220 19234
rect 16940 19180 17220 19182
rect 17276 19234 17332 19246
rect 17276 19182 17278 19234
rect 17330 19182 17332 19234
rect 16940 19170 16996 19180
rect 16772 18396 16884 18452
rect 17276 19124 17332 19182
rect 17388 19236 17444 19246
rect 17388 19142 17444 19180
rect 17724 19234 17780 21644
rect 18172 21634 18228 21644
rect 18508 21700 18564 21710
rect 18508 21606 18564 21644
rect 18284 21364 18340 21374
rect 17948 21028 18004 21038
rect 17948 20934 18004 20972
rect 18284 20020 18340 21308
rect 18620 20244 18676 23884
rect 18956 23938 19012 23950
rect 18956 23886 18958 23938
rect 19010 23886 19012 23938
rect 18956 23828 19012 23886
rect 18956 23762 19012 23772
rect 19068 23548 19124 29148
rect 19740 29138 19796 29148
rect 19852 28642 19908 28654
rect 19852 28590 19854 28642
rect 19906 28590 19908 28642
rect 19180 28532 19236 28542
rect 19180 25618 19236 28476
rect 19404 28530 19460 28542
rect 19404 28478 19406 28530
rect 19458 28478 19460 28530
rect 19404 27076 19460 28478
rect 19180 25566 19182 25618
rect 19234 25566 19236 25618
rect 19180 25554 19236 25566
rect 19292 27074 19460 27076
rect 19292 27022 19406 27074
rect 19458 27022 19460 27074
rect 19292 27020 19460 27022
rect 19292 23828 19348 27020
rect 19404 27010 19460 27020
rect 19740 27634 19796 27646
rect 19740 27582 19742 27634
rect 19794 27582 19796 27634
rect 19740 26908 19796 27582
rect 19292 23762 19348 23772
rect 19628 26852 19796 26908
rect 19068 23492 19460 23548
rect 19292 22260 19348 22270
rect 19292 22166 19348 22204
rect 19068 22148 19124 22158
rect 18956 21700 19012 21710
rect 18844 21474 18900 21486
rect 18844 21422 18846 21474
rect 18898 21422 18900 21474
rect 18844 21028 18900 21422
rect 18844 20962 18900 20972
rect 18956 20804 19012 21644
rect 19068 21586 19124 22092
rect 19068 21534 19070 21586
rect 19122 21534 19124 21586
rect 19068 21028 19124 21534
rect 19292 21588 19348 21598
rect 19292 21494 19348 21532
rect 19068 20962 19124 20972
rect 19292 21028 19348 21038
rect 19068 20804 19124 20814
rect 18956 20802 19124 20804
rect 18956 20750 19070 20802
rect 19122 20750 19124 20802
rect 18956 20748 19124 20750
rect 19068 20738 19124 20748
rect 19292 20804 19348 20972
rect 18732 20692 18788 20702
rect 18732 20690 19012 20692
rect 18732 20638 18734 20690
rect 18786 20638 19012 20690
rect 18732 20636 19012 20638
rect 18732 20626 18788 20636
rect 18620 20178 18676 20188
rect 18060 19964 18340 20020
rect 17724 19182 17726 19234
rect 17778 19182 17780 19234
rect 17724 19170 17780 19182
rect 17836 19908 17892 19918
rect 16716 18358 16772 18396
rect 16828 17892 16884 17902
rect 16828 17798 16884 17836
rect 16716 17780 16772 17790
rect 16716 17668 16772 17724
rect 17164 17668 17220 17678
rect 16716 17666 17220 17668
rect 16716 17614 16718 17666
rect 16770 17614 17166 17666
rect 17218 17614 17220 17666
rect 16716 17612 17220 17614
rect 16716 17602 16772 17612
rect 16940 17332 16996 17342
rect 16940 16884 16996 17276
rect 17164 17220 17220 17612
rect 17164 17154 17220 17164
rect 16828 16882 16996 16884
rect 16828 16830 16942 16882
rect 16994 16830 16996 16882
rect 16828 16828 16996 16830
rect 16716 16100 16772 16110
rect 16380 16034 16436 16044
rect 16604 16098 16772 16100
rect 16604 16046 16718 16098
rect 16770 16046 16772 16098
rect 16604 16044 16772 16046
rect 16604 13972 16660 16044
rect 16716 16034 16772 16044
rect 16828 15314 16884 16828
rect 16940 16818 16996 16828
rect 17276 16772 17332 19068
rect 17388 18340 17444 18350
rect 17388 18246 17444 18284
rect 17836 18338 17892 19852
rect 17948 19796 18004 19806
rect 17948 18452 18004 19740
rect 17948 18358 18004 18396
rect 17836 18286 17838 18338
rect 17890 18286 17892 18338
rect 17836 18274 17892 18286
rect 17836 18116 17892 18126
rect 17500 17780 17556 17790
rect 17500 17686 17556 17724
rect 17836 17778 17892 18060
rect 17836 17726 17838 17778
rect 17890 17726 17892 17778
rect 17836 17714 17892 17726
rect 17388 17556 17444 17566
rect 17388 17462 17444 17500
rect 17948 17556 18004 17566
rect 17948 17220 18004 17500
rect 18060 17444 18116 19964
rect 18620 19908 18676 19918
rect 18620 19814 18676 19852
rect 18172 19794 18228 19806
rect 18172 19742 18174 19794
rect 18226 19742 18228 19794
rect 18172 18340 18228 19742
rect 18732 19794 18788 19806
rect 18732 19742 18734 19794
rect 18786 19742 18788 19794
rect 18172 17666 18228 18284
rect 18172 17614 18174 17666
rect 18226 17614 18228 17666
rect 18172 17556 18228 17614
rect 18172 17490 18228 17500
rect 18284 19234 18340 19246
rect 18284 19182 18286 19234
rect 18338 19182 18340 19234
rect 18060 17378 18116 17388
rect 18284 17332 18340 19182
rect 18732 18676 18788 19742
rect 18396 18620 18788 18676
rect 18844 19794 18900 19806
rect 18844 19742 18846 19794
rect 18898 19742 18900 19794
rect 18396 17444 18452 18620
rect 18844 18564 18900 19742
rect 18844 18498 18900 18508
rect 18508 18450 18564 18462
rect 18508 18398 18510 18450
rect 18562 18398 18564 18450
rect 18508 17668 18564 18398
rect 18620 18340 18676 18350
rect 18844 18338 18900 18350
rect 18844 18298 18846 18338
rect 18676 18286 18846 18298
rect 18898 18286 18900 18338
rect 18676 18284 18900 18286
rect 18620 18242 18900 18284
rect 18508 17602 18564 17612
rect 18620 18116 18676 18126
rect 18620 17666 18676 18060
rect 18844 17780 18900 17790
rect 18844 17686 18900 17724
rect 18620 17614 18622 17666
rect 18674 17614 18676 17666
rect 18620 17602 18676 17614
rect 18396 17388 18564 17444
rect 18284 17276 18452 17332
rect 17948 17164 18340 17220
rect 18284 17106 18340 17164
rect 18284 17054 18286 17106
rect 18338 17054 18340 17106
rect 18284 17042 18340 17054
rect 17276 16706 17332 16716
rect 17612 16877 17668 16889
rect 18396 16884 18452 17276
rect 18508 17106 18564 17388
rect 18508 17054 18510 17106
rect 18562 17054 18564 17106
rect 18508 17042 18564 17054
rect 17612 16825 17614 16877
rect 17666 16825 17668 16877
rect 17612 16436 17668 16825
rect 18172 16828 18452 16884
rect 18732 16882 18788 16894
rect 18732 16830 18734 16882
rect 18786 16830 18788 16882
rect 18956 16879 19012 20636
rect 19292 20020 19348 20748
rect 19404 20188 19460 23492
rect 19628 23044 19684 26852
rect 19852 26516 19908 28590
rect 19964 26516 20020 26526
rect 19852 26514 20020 26516
rect 19852 26462 19966 26514
rect 20018 26462 20020 26514
rect 19852 26460 20020 26462
rect 19964 26450 20020 26460
rect 20076 25732 20132 33966
rect 20300 31780 20356 34862
rect 20300 31714 20356 31724
rect 20188 31666 20244 31678
rect 20188 31614 20190 31666
rect 20242 31614 20244 31666
rect 20188 31444 20244 31614
rect 20188 31378 20244 31388
rect 20412 30996 20468 36430
rect 20300 30940 20468 30996
rect 20300 30100 20356 30940
rect 20300 30034 20356 30044
rect 20524 29764 20580 54124
rect 20636 53844 20692 54238
rect 21532 54068 21588 54350
rect 21532 54002 21588 54012
rect 20636 53778 20692 53788
rect 21420 52500 21476 52510
rect 21420 52386 21476 52444
rect 21420 52334 21422 52386
rect 21474 52334 21476 52386
rect 21420 52322 21476 52334
rect 21644 52276 21700 52286
rect 21756 52276 21812 56030
rect 22540 55860 22596 55870
rect 21868 55748 21924 55758
rect 21868 53842 21924 55692
rect 22428 55300 22484 55310
rect 22428 55206 22484 55244
rect 22540 54738 22596 55804
rect 22988 55522 23044 57372
rect 23520 57344 23632 57456
rect 24864 57344 24976 57456
rect 25564 57372 25956 57428
rect 23548 56308 23604 57344
rect 24332 57204 24388 57214
rect 24220 56756 24276 56766
rect 23804 56476 24068 56486
rect 23860 56420 23908 56476
rect 23964 56420 24012 56476
rect 23804 56410 24068 56420
rect 23548 56242 23604 56252
rect 22988 55470 22990 55522
rect 23042 55470 23044 55522
rect 22988 55458 23044 55470
rect 23548 55972 23604 55982
rect 22540 54686 22542 54738
rect 22594 54686 22596 54738
rect 22540 54674 22596 54686
rect 23324 55300 23380 55310
rect 21868 53790 21870 53842
rect 21922 53790 21924 53842
rect 21868 53778 21924 53790
rect 22316 53732 22372 53742
rect 22316 53638 22372 53676
rect 22764 53730 22820 53742
rect 22764 53678 22766 53730
rect 22818 53678 22820 53730
rect 22764 52388 22820 53678
rect 23100 52834 23156 52846
rect 23100 52782 23102 52834
rect 23154 52782 23156 52834
rect 23100 52612 23156 52782
rect 23100 52546 23156 52556
rect 22764 52322 22820 52332
rect 21980 52276 22036 52286
rect 21756 52274 22036 52276
rect 21756 52222 21982 52274
rect 22034 52222 22036 52274
rect 21756 52220 22036 52222
rect 20972 40964 21028 40974
rect 20972 38668 21028 40908
rect 20972 38612 21140 38668
rect 20748 38052 20804 38062
rect 20748 32674 20804 37996
rect 20748 32622 20750 32674
rect 20802 32622 20804 32674
rect 20748 32610 20804 32622
rect 20636 31780 20692 31790
rect 20636 31778 20916 31780
rect 20636 31726 20638 31778
rect 20690 31726 20916 31778
rect 20636 31724 20916 31726
rect 20636 31714 20692 31724
rect 20636 31444 20692 31454
rect 20636 30884 20692 31388
rect 20636 30882 20804 30884
rect 20636 30830 20638 30882
rect 20690 30830 20804 30882
rect 20636 30828 20804 30830
rect 20636 30818 20692 30828
rect 20300 29708 20580 29764
rect 20188 28642 20244 28654
rect 20188 28590 20190 28642
rect 20242 28590 20244 28642
rect 20188 26852 20244 28590
rect 20188 26786 20244 26796
rect 19852 25676 20132 25732
rect 19740 25396 19796 25406
rect 19740 25302 19796 25340
rect 19740 23940 19796 23950
rect 19740 23846 19796 23884
rect 19852 23380 19908 25676
rect 20188 25620 20244 25630
rect 19964 25618 20244 25620
rect 19964 25566 20190 25618
rect 20242 25566 20244 25618
rect 19964 25564 20244 25566
rect 19964 23492 20020 25564
rect 20188 25554 20244 25564
rect 19964 23426 20020 23436
rect 19852 23314 19908 23324
rect 19964 23156 20020 23166
rect 19516 23042 19684 23044
rect 19516 22990 19630 23042
rect 19682 22990 19684 23042
rect 19516 22988 19684 22990
rect 19516 21588 19572 22988
rect 19628 22978 19684 22988
rect 19740 23154 20020 23156
rect 19740 23102 19966 23154
rect 20018 23102 20020 23154
rect 19740 23100 20020 23102
rect 19628 22370 19684 22382
rect 19628 22318 19630 22370
rect 19682 22318 19684 22370
rect 19628 22148 19684 22318
rect 19628 22082 19684 22092
rect 19740 22036 19796 23100
rect 19964 23090 20020 23100
rect 19740 21970 19796 21980
rect 19852 22930 19908 22942
rect 19852 22878 19854 22930
rect 19906 22878 19908 22930
rect 19852 21812 19908 22878
rect 20076 22932 20132 22942
rect 20076 22930 20244 22932
rect 20076 22878 20078 22930
rect 20130 22878 20244 22930
rect 20076 22876 20244 22878
rect 20076 22866 20132 22876
rect 20076 22372 20132 22382
rect 20076 22278 20132 22316
rect 19516 21522 19572 21532
rect 19628 21756 19908 21812
rect 19628 21586 19684 21756
rect 19852 21700 19908 21756
rect 19852 21644 20020 21700
rect 19628 21534 19630 21586
rect 19682 21534 19684 21586
rect 19628 21522 19684 21534
rect 19628 21364 19684 21374
rect 19628 21270 19684 21308
rect 19964 21362 20020 21644
rect 19964 21310 19966 21362
rect 20018 21310 20020 21362
rect 19964 21298 20020 21310
rect 20076 21474 20132 21486
rect 20076 21422 20078 21474
rect 20130 21422 20132 21474
rect 19964 21140 20020 21150
rect 19740 21084 19964 21140
rect 19740 21026 19796 21084
rect 19964 21074 20020 21084
rect 19740 20974 19742 21026
rect 19794 20974 19796 21026
rect 19740 20962 19796 20974
rect 19516 20916 19572 20926
rect 19516 20802 19572 20860
rect 19516 20750 19518 20802
rect 19570 20750 19572 20802
rect 19516 20356 19572 20750
rect 19516 20290 19572 20300
rect 20076 20188 20132 21422
rect 20188 21140 20244 22876
rect 20300 22708 20356 29708
rect 20412 28756 20468 28766
rect 20412 28754 20692 28756
rect 20412 28702 20414 28754
rect 20466 28702 20692 28754
rect 20412 28700 20692 28702
rect 20412 28690 20468 28700
rect 20636 27858 20692 28700
rect 20636 27806 20638 27858
rect 20690 27806 20692 27858
rect 20636 27794 20692 27806
rect 20412 27074 20468 27086
rect 20412 27022 20414 27074
rect 20466 27022 20468 27074
rect 20412 26628 20468 27022
rect 20748 26908 20804 30828
rect 20860 30434 20916 31724
rect 20972 31778 21028 31790
rect 20972 31726 20974 31778
rect 21026 31726 21028 31778
rect 20972 31444 21028 31726
rect 20972 31378 21028 31388
rect 20972 31220 21028 31230
rect 20972 30994 21028 31164
rect 20972 30942 20974 30994
rect 21026 30942 21028 30994
rect 20972 30930 21028 30942
rect 21084 30772 21140 38612
rect 21308 34914 21364 34926
rect 21308 34862 21310 34914
rect 21362 34862 21364 34914
rect 21308 34132 21364 34862
rect 21308 34066 21364 34076
rect 21644 33684 21700 52220
rect 21980 52210 22036 52220
rect 22764 52164 22820 52174
rect 22764 52070 22820 52108
rect 21644 33618 21700 33628
rect 21756 40404 21812 40414
rect 21196 32338 21252 32350
rect 21532 32340 21588 32350
rect 21196 32286 21198 32338
rect 21250 32286 21252 32338
rect 21196 32228 21252 32286
rect 21196 32162 21252 32172
rect 21308 32338 21588 32340
rect 21308 32286 21534 32338
rect 21586 32286 21588 32338
rect 21308 32284 21588 32286
rect 21196 32004 21252 32014
rect 21308 32004 21364 32284
rect 21532 32274 21588 32284
rect 21756 32116 21812 40348
rect 22764 37716 22820 37726
rect 22316 35476 22372 35486
rect 22092 32676 22148 32686
rect 22092 32582 22148 32620
rect 21196 32002 21364 32004
rect 21196 31950 21198 32002
rect 21250 31950 21364 32002
rect 21196 31948 21364 31950
rect 21420 32060 21812 32116
rect 21868 32340 21924 32350
rect 21196 31938 21252 31948
rect 21420 31668 21476 32060
rect 21644 31892 21700 31902
rect 20860 30382 20862 30434
rect 20914 30382 20916 30434
rect 20860 30370 20916 30382
rect 20972 30716 21140 30772
rect 21196 31612 21476 31668
rect 21532 31780 21588 31790
rect 20748 26852 20916 26908
rect 20412 26562 20468 26572
rect 20748 26290 20804 26302
rect 20748 26238 20750 26290
rect 20802 26238 20804 26290
rect 20748 25732 20804 26238
rect 20524 25676 20804 25732
rect 20412 25396 20468 25406
rect 20524 25396 20580 25676
rect 20468 25340 20580 25396
rect 20412 23938 20468 25340
rect 20636 24836 20692 24846
rect 20636 24742 20692 24780
rect 20412 23886 20414 23938
rect 20466 23886 20468 23938
rect 20412 23874 20468 23886
rect 20860 23828 20916 26852
rect 20972 24948 21028 30716
rect 21084 28642 21140 28654
rect 21084 28590 21086 28642
rect 21138 28590 21140 28642
rect 21084 26908 21140 28590
rect 21196 27970 21252 31612
rect 21196 27918 21198 27970
rect 21250 27918 21252 27970
rect 21196 27906 21252 27918
rect 21308 31444 21364 31454
rect 21308 30996 21364 31388
rect 21420 30996 21476 31006
rect 21308 30994 21476 30996
rect 21308 30942 21422 30994
rect 21474 30942 21476 30994
rect 21308 30940 21476 30942
rect 21308 27412 21364 30940
rect 21420 30930 21476 30940
rect 21532 30660 21588 31724
rect 21644 30882 21700 31836
rect 21644 30830 21646 30882
rect 21698 30830 21700 30882
rect 21644 30818 21700 30830
rect 21756 31778 21812 31790
rect 21756 31726 21758 31778
rect 21810 31726 21812 31778
rect 21532 30604 21700 30660
rect 21308 27346 21364 27356
rect 21420 30212 21476 30222
rect 21420 28642 21476 30156
rect 21532 30100 21588 30110
rect 21532 30006 21588 30044
rect 21420 28590 21422 28642
rect 21474 28590 21476 28642
rect 21420 26908 21476 28590
rect 21644 27860 21700 30604
rect 21756 30212 21812 31726
rect 21756 30146 21812 30156
rect 21868 30322 21924 32284
rect 22092 30996 22148 31006
rect 22092 30902 22148 30940
rect 21868 30270 21870 30322
rect 21922 30270 21924 30322
rect 21644 27794 21700 27804
rect 21084 26852 21252 26908
rect 21420 26852 21700 26908
rect 21084 26628 21140 26638
rect 21084 25060 21140 26572
rect 21196 25732 21252 26852
rect 21532 26740 21588 26750
rect 21420 26516 21476 26526
rect 21308 26068 21364 26078
rect 21308 25974 21364 26012
rect 21308 25732 21364 25742
rect 21196 25730 21364 25732
rect 21196 25678 21310 25730
rect 21362 25678 21364 25730
rect 21196 25676 21364 25678
rect 21308 25666 21364 25676
rect 21084 25004 21364 25060
rect 20972 24892 21252 24948
rect 21084 24722 21140 24734
rect 21084 24670 21086 24722
rect 21138 24670 21140 24722
rect 21084 24164 21140 24670
rect 21084 24098 21140 24108
rect 20972 24052 21028 24062
rect 20972 23958 21028 23996
rect 20860 23772 21028 23828
rect 20300 22652 20468 22708
rect 20188 21074 20244 21084
rect 20300 22482 20356 22494
rect 20300 22430 20302 22482
rect 20354 22430 20356 22482
rect 20188 20804 20244 20814
rect 20188 20710 20244 20748
rect 20300 20356 20356 22430
rect 20300 20290 20356 20300
rect 19404 20132 20132 20188
rect 19292 19964 19684 20020
rect 19292 19234 19348 19246
rect 19292 19182 19294 19234
rect 19346 19182 19348 19234
rect 19068 18450 19124 18462
rect 19068 18398 19070 18450
rect 19122 18398 19124 18450
rect 19068 17780 19124 18398
rect 19292 18452 19348 19182
rect 19628 19236 19684 19964
rect 19740 20018 19796 20132
rect 19740 19966 19742 20018
rect 19794 19966 19796 20018
rect 19740 19796 19796 19966
rect 19964 20020 20020 20030
rect 20412 20020 20468 22652
rect 20748 22370 20804 22382
rect 20748 22318 20750 22370
rect 20802 22318 20804 22370
rect 20748 21700 20804 22318
rect 20636 21586 20692 21598
rect 20636 21534 20638 21586
rect 20690 21534 20692 21586
rect 20636 21364 20692 21534
rect 20636 21298 20692 21308
rect 20748 21028 20804 21644
rect 20636 20972 20804 21028
rect 20860 21586 20916 21598
rect 20860 21534 20862 21586
rect 20914 21534 20916 21586
rect 20524 20356 20580 20366
rect 20636 20356 20692 20972
rect 20748 20802 20804 20814
rect 20748 20750 20750 20802
rect 20802 20750 20804 20802
rect 20748 20580 20804 20750
rect 20748 20514 20804 20524
rect 20636 20300 20804 20356
rect 20524 20132 20580 20300
rect 20636 20132 20692 20142
rect 20524 20130 20692 20132
rect 20524 20078 20638 20130
rect 20690 20078 20692 20130
rect 20524 20076 20692 20078
rect 20636 20066 20692 20076
rect 20412 19964 20580 20020
rect 19964 19926 20020 19964
rect 20076 19908 20132 19918
rect 20076 19906 20356 19908
rect 20076 19854 20078 19906
rect 20130 19854 20356 19906
rect 20076 19852 20356 19854
rect 20076 19842 20132 19852
rect 19740 19730 19796 19740
rect 20300 19458 20356 19852
rect 20300 19406 20302 19458
rect 20354 19406 20356 19458
rect 20300 19394 20356 19406
rect 19628 19142 19684 19180
rect 20412 19234 20468 19246
rect 20412 19182 20414 19234
rect 20466 19182 20468 19234
rect 20412 18676 20468 19182
rect 20412 18610 20468 18620
rect 19292 18396 19908 18452
rect 19516 18226 19572 18238
rect 19516 18174 19518 18226
rect 19570 18174 19572 18226
rect 19516 18116 19572 18174
rect 19516 17892 19572 18060
rect 19516 17826 19572 17836
rect 19628 18226 19684 18238
rect 19628 18174 19630 18226
rect 19682 18174 19684 18226
rect 19068 17714 19124 17724
rect 19292 17668 19348 17678
rect 19292 17574 19348 17612
rect 19628 17444 19684 18174
rect 19180 17388 19684 17444
rect 19740 18226 19796 18238
rect 19740 18174 19742 18226
rect 19794 18174 19796 18226
rect 19068 16996 19124 17006
rect 19068 16902 19124 16940
rect 17052 16322 17108 16334
rect 17052 16270 17054 16322
rect 17106 16270 17108 16322
rect 16940 16100 16996 16110
rect 16940 15540 16996 16044
rect 17052 15652 17108 16270
rect 17500 16098 17556 16110
rect 17500 16046 17502 16098
rect 17554 16046 17556 16098
rect 17276 15874 17332 15886
rect 17276 15822 17278 15874
rect 17330 15822 17332 15874
rect 17276 15652 17332 15822
rect 17500 15764 17556 16046
rect 17500 15698 17556 15708
rect 17052 15596 17220 15652
rect 16940 15484 17108 15540
rect 16828 15262 16830 15314
rect 16882 15262 16884 15314
rect 16828 15148 16884 15262
rect 16828 15092 16996 15148
rect 16828 14756 16884 14766
rect 16828 14662 16884 14700
rect 16940 14642 16996 15092
rect 17052 15092 17108 15484
rect 17052 15026 17108 15036
rect 16940 14590 16942 14642
rect 16994 14590 16996 14642
rect 16716 14532 16772 14542
rect 16716 14438 16772 14476
rect 16604 13906 16660 13916
rect 16828 14420 16884 14430
rect 16716 13748 16772 13758
rect 16828 13748 16884 14364
rect 16716 13746 16884 13748
rect 16716 13694 16718 13746
rect 16770 13694 16884 13746
rect 16716 13692 16884 13694
rect 16716 13682 16772 13692
rect 16940 12964 16996 14590
rect 17164 14084 17220 15596
rect 17276 15586 17332 15596
rect 17612 15316 17668 16380
rect 18060 16772 18116 16782
rect 17836 16100 17892 16110
rect 17836 16098 18004 16100
rect 17836 16046 17838 16098
rect 17890 16046 18004 16098
rect 17836 16044 18004 16046
rect 17836 16034 17892 16044
rect 17948 15652 18004 16044
rect 18060 16098 18116 16716
rect 18060 16046 18062 16098
rect 18114 16046 18116 16098
rect 18060 15876 18116 16046
rect 18060 15810 18116 15820
rect 17948 15596 18116 15652
rect 17724 15316 17780 15326
rect 17612 15314 17780 15316
rect 17612 15262 17726 15314
rect 17778 15262 17780 15314
rect 17612 15260 17780 15262
rect 17500 15204 17556 15214
rect 17164 14018 17220 14028
rect 17276 14644 17332 14654
rect 16716 12908 16996 12964
rect 17164 13300 17220 13310
rect 17164 12962 17220 13244
rect 17164 12910 17166 12962
rect 17218 12910 17220 12962
rect 16492 12180 16548 12190
rect 16492 12086 16548 12124
rect 16716 12068 16772 12908
rect 16828 12738 16884 12750
rect 16828 12686 16830 12738
rect 16882 12686 16884 12738
rect 16828 12180 16884 12686
rect 16940 12180 16996 12190
rect 16828 12178 16996 12180
rect 16828 12126 16942 12178
rect 16994 12126 16996 12178
rect 16828 12124 16996 12126
rect 16940 12114 16996 12124
rect 16716 12012 16884 12068
rect 16268 11106 16324 11116
rect 16716 11506 16772 11518
rect 16716 11454 16718 11506
rect 16770 11454 16772 11506
rect 16604 10612 16660 10622
rect 15820 9090 15876 9100
rect 15932 10610 16660 10612
rect 15932 10558 16606 10610
rect 16658 10558 16660 10610
rect 15932 10556 16660 10558
rect 15708 8318 15710 8370
rect 15762 8318 15764 8370
rect 15484 8194 15540 8204
rect 15596 8258 15652 8270
rect 15596 8206 15598 8258
rect 15650 8206 15652 8258
rect 15596 8036 15652 8206
rect 15596 7970 15652 7980
rect 15708 7812 15764 8318
rect 15484 7756 15764 7812
rect 15484 7476 15540 7756
rect 15484 7410 15540 7420
rect 15596 7588 15652 7598
rect 15596 7474 15652 7532
rect 15596 7422 15598 7474
rect 15650 7422 15652 7474
rect 14924 7298 14980 7308
rect 15596 7364 15652 7422
rect 15932 7474 15988 10556
rect 16604 10546 16660 10556
rect 16268 10386 16324 10398
rect 16268 10334 16270 10386
rect 16322 10334 16324 10386
rect 16044 10164 16100 10174
rect 16044 10050 16100 10108
rect 16268 10164 16324 10334
rect 16268 10098 16324 10108
rect 16044 9998 16046 10050
rect 16098 9998 16100 10050
rect 16044 9986 16100 9998
rect 16492 10052 16548 10062
rect 16156 9940 16212 9950
rect 16156 9846 16212 9884
rect 16492 9266 16548 9996
rect 16604 9826 16660 9838
rect 16604 9774 16606 9826
rect 16658 9774 16660 9826
rect 16604 9492 16660 9774
rect 16604 9426 16660 9436
rect 16492 9214 16494 9266
rect 16546 9214 16548 9266
rect 16492 9202 16548 9214
rect 15932 7422 15934 7474
rect 15986 7422 15988 7474
rect 15932 7410 15988 7422
rect 16044 9156 16100 9166
rect 15596 7298 15652 7308
rect 15708 7252 15764 7262
rect 15708 7158 15764 7196
rect 14700 5854 14702 5906
rect 14754 5854 14756 5906
rect 14252 5842 14308 5852
rect 14700 5842 14756 5854
rect 15932 6468 15988 6478
rect 15260 5796 15316 5806
rect 14924 5794 15316 5796
rect 14924 5742 15262 5794
rect 15314 5742 15316 5794
rect 14924 5740 15316 5742
rect 14812 5684 14868 5694
rect 14812 5590 14868 5628
rect 14924 5346 14980 5740
rect 15260 5730 15316 5740
rect 14924 5294 14926 5346
rect 14978 5294 14980 5346
rect 14924 5282 14980 5294
rect 15372 5684 15428 5694
rect 15372 5346 15428 5628
rect 15372 5294 15374 5346
rect 15426 5294 15428 5346
rect 15372 5282 15428 5294
rect 13692 5182 13694 5234
rect 13746 5182 13748 5234
rect 13692 5170 13748 5182
rect 15932 5234 15988 6412
rect 16044 5906 16100 9100
rect 16716 8372 16772 11454
rect 16716 8306 16772 8316
rect 16156 8036 16212 8046
rect 16716 8036 16772 8046
rect 16156 8034 16772 8036
rect 16156 7982 16158 8034
rect 16210 7982 16718 8034
rect 16770 7982 16772 8034
rect 16156 7980 16772 7982
rect 16156 7970 16212 7980
rect 16716 7970 16772 7980
rect 16604 7812 16660 7822
rect 16604 7698 16660 7756
rect 16604 7646 16606 7698
rect 16658 7646 16660 7698
rect 16604 7634 16660 7646
rect 16716 7700 16772 7710
rect 16716 7606 16772 7644
rect 16380 7588 16436 7598
rect 16380 7494 16436 7532
rect 16156 7476 16212 7486
rect 16156 7382 16212 7420
rect 16268 7364 16324 7374
rect 16268 6020 16324 7308
rect 16268 5954 16324 5964
rect 16044 5854 16046 5906
rect 16098 5854 16100 5906
rect 16044 5842 16100 5854
rect 16828 5684 16884 12012
rect 17164 11788 17220 12910
rect 16940 11732 17220 11788
rect 17276 12178 17332 14588
rect 17388 13972 17444 13982
rect 17388 13878 17444 13916
rect 17276 12126 17278 12178
rect 17330 12126 17332 12178
rect 16940 11666 16996 11676
rect 17052 11394 17108 11406
rect 17052 11342 17054 11394
rect 17106 11342 17108 11394
rect 17052 11060 17108 11342
rect 17276 11396 17332 12126
rect 17276 11330 17332 11340
rect 17388 12964 17444 12974
rect 17052 10994 17108 11004
rect 17388 10612 17444 12908
rect 17500 12402 17556 15148
rect 17724 14642 17780 15260
rect 17724 14590 17726 14642
rect 17778 14590 17780 14642
rect 17724 14578 17780 14590
rect 17948 15316 18004 15326
rect 17948 14532 18004 15260
rect 18060 14756 18116 15596
rect 18172 15148 18228 16828
rect 18620 16660 18676 16670
rect 18284 16324 18340 16334
rect 18284 16322 18452 16324
rect 18284 16270 18286 16322
rect 18338 16270 18452 16322
rect 18284 16268 18452 16270
rect 18284 16258 18340 16268
rect 18284 16100 18340 16110
rect 18284 16006 18340 16044
rect 18396 15652 18452 16268
rect 18620 16098 18676 16604
rect 18732 16548 18788 16830
rect 18732 16482 18788 16492
rect 18844 16823 19012 16879
rect 19180 16882 19236 17388
rect 19740 17332 19796 18174
rect 19852 17666 19908 18396
rect 20300 18340 20356 18350
rect 19852 17614 19854 17666
rect 19906 17614 19908 17666
rect 19852 17602 19908 17614
rect 20076 17666 20132 17678
rect 20076 17614 20078 17666
rect 20130 17614 20132 17666
rect 19740 17276 19908 17332
rect 19628 16996 19684 17006
rect 19180 16830 19182 16882
rect 19234 16830 19236 16882
rect 18844 16212 18900 16823
rect 19180 16818 19236 16830
rect 19292 16994 19684 16996
rect 19292 16942 19630 16994
rect 19682 16942 19684 16994
rect 19292 16940 19684 16942
rect 18956 16658 19012 16670
rect 19292 16660 19348 16940
rect 19628 16930 19684 16940
rect 18956 16606 18958 16658
rect 19010 16606 19012 16658
rect 18956 16548 19012 16606
rect 19180 16604 19348 16660
rect 19740 16658 19796 16670
rect 19740 16606 19742 16658
rect 19794 16606 19796 16658
rect 19180 16548 19236 16604
rect 18956 16492 19236 16548
rect 19404 16548 19460 16558
rect 18956 16212 19012 16222
rect 18844 16210 19124 16212
rect 18844 16158 18958 16210
rect 19010 16158 19124 16210
rect 18844 16156 19124 16158
rect 18956 16146 19012 16156
rect 18620 16046 18622 16098
rect 18674 16046 18676 16098
rect 18620 16034 18676 16046
rect 18396 15586 18452 15596
rect 18844 15876 18900 15886
rect 18620 15538 18676 15550
rect 18620 15486 18622 15538
rect 18674 15486 18676 15538
rect 18508 15314 18564 15326
rect 18508 15262 18510 15314
rect 18562 15262 18564 15314
rect 18396 15204 18452 15214
rect 18172 15092 18340 15148
rect 18060 14700 18228 14756
rect 18060 14532 18116 14542
rect 18004 14530 18116 14532
rect 18004 14478 18062 14530
rect 18114 14478 18116 14530
rect 18004 14476 18116 14478
rect 17948 14438 18004 14476
rect 17724 13972 17780 13982
rect 17724 13878 17780 13916
rect 17836 13636 17892 13646
rect 17836 13074 17892 13580
rect 17836 13022 17838 13074
rect 17890 13022 17892 13074
rect 17836 12740 17892 13022
rect 17948 12964 18004 12974
rect 18060 12964 18116 14476
rect 18172 13746 18228 14700
rect 18284 14420 18340 15092
rect 18396 15090 18452 15148
rect 18396 15038 18398 15090
rect 18450 15038 18452 15090
rect 18396 15026 18452 15038
rect 18508 14756 18564 15262
rect 18508 14690 18564 14700
rect 18620 14644 18676 15486
rect 18844 15314 18900 15820
rect 18844 15262 18846 15314
rect 18898 15262 18900 15314
rect 18844 15250 18900 15262
rect 18956 15652 19012 15662
rect 18956 15148 19012 15596
rect 18844 15092 19012 15148
rect 18620 14578 18676 14588
rect 18732 14642 18788 14654
rect 18732 14590 18734 14642
rect 18786 14590 18788 14642
rect 18508 14532 18564 14542
rect 18508 14438 18564 14476
rect 18284 14354 18340 14364
rect 18172 13694 18174 13746
rect 18226 13694 18228 13746
rect 18172 13682 18228 13694
rect 18396 13748 18452 13758
rect 18396 13654 18452 13692
rect 18284 13636 18340 13646
rect 18284 13542 18340 13580
rect 18732 13074 18788 14590
rect 18732 13022 18734 13074
rect 18786 13022 18788 13074
rect 18732 13010 18788 13022
rect 18844 14532 18900 15092
rect 18396 12964 18452 12974
rect 17948 12962 18228 12964
rect 17948 12910 17950 12962
rect 18002 12910 18228 12962
rect 17948 12908 18228 12910
rect 17948 12898 18004 12908
rect 17836 12684 18004 12740
rect 17500 12350 17502 12402
rect 17554 12350 17556 12402
rect 17500 12338 17556 12350
rect 17612 12292 17668 12302
rect 17612 12178 17668 12236
rect 17612 12126 17614 12178
rect 17666 12126 17668 12178
rect 17612 12114 17668 12126
rect 17724 12068 17780 12078
rect 17724 11954 17780 12012
rect 17724 11902 17726 11954
rect 17778 11902 17780 11954
rect 17724 11890 17780 11902
rect 17948 11844 18004 12684
rect 18060 12178 18116 12190
rect 18060 12126 18062 12178
rect 18114 12126 18116 12178
rect 18060 12068 18116 12126
rect 18060 12002 18116 12012
rect 17948 11788 18116 11844
rect 17612 11732 17668 11742
rect 17612 10722 17668 11676
rect 17612 10670 17614 10722
rect 17666 10670 17668 10722
rect 17612 10658 17668 10670
rect 17724 11282 17780 11294
rect 17724 11230 17726 11282
rect 17778 11230 17780 11282
rect 17500 10612 17556 10622
rect 17388 10610 17556 10612
rect 17388 10558 17502 10610
rect 17554 10558 17556 10610
rect 17388 10556 17556 10558
rect 17500 10546 17556 10556
rect 17276 10500 17332 10510
rect 17276 10498 17444 10500
rect 17276 10446 17278 10498
rect 17330 10446 17444 10498
rect 17276 10444 17444 10446
rect 17276 10434 17332 10444
rect 16940 10388 16996 10398
rect 16940 10386 17108 10388
rect 16940 10334 16942 10386
rect 16994 10334 17108 10386
rect 16940 10332 17108 10334
rect 16940 10322 16996 10332
rect 17052 10052 17108 10332
rect 17164 10386 17220 10398
rect 17164 10334 17166 10386
rect 17218 10334 17220 10386
rect 17164 10276 17220 10334
rect 17164 10220 17332 10276
rect 17276 10052 17332 10220
rect 17388 10164 17444 10444
rect 17612 10388 17668 10398
rect 17388 10108 17556 10164
rect 17052 9996 17220 10052
rect 17164 9938 17220 9996
rect 17332 9996 17444 10052
rect 17276 9986 17332 9996
rect 17164 9886 17166 9938
rect 17218 9886 17220 9938
rect 17164 9874 17220 9886
rect 17052 9828 17108 9838
rect 17052 9734 17108 9772
rect 17276 9828 17332 9838
rect 16940 9716 16996 9726
rect 16940 9268 16996 9660
rect 17052 9268 17108 9278
rect 16940 9266 17108 9268
rect 16940 9214 17054 9266
rect 17106 9214 17108 9266
rect 16940 9212 17108 9214
rect 17052 9202 17108 9212
rect 17164 9268 17220 9278
rect 17276 9268 17332 9772
rect 17220 9212 17332 9268
rect 17164 9202 17220 9212
rect 17388 9156 17444 9996
rect 17276 9100 17444 9156
rect 16940 8260 16996 8270
rect 16940 8166 16996 8204
rect 17276 8258 17332 9100
rect 17500 8372 17556 10108
rect 17612 8708 17668 10332
rect 17724 8932 17780 11230
rect 17836 10498 17892 10510
rect 17836 10446 17838 10498
rect 17890 10446 17892 10498
rect 17836 10052 17892 10446
rect 17836 9986 17892 9996
rect 17948 9940 18004 9950
rect 17948 9716 18004 9884
rect 17948 9622 18004 9660
rect 17724 8866 17780 8876
rect 17612 8652 17780 8708
rect 17612 8372 17668 8382
rect 17500 8370 17668 8372
rect 17500 8318 17614 8370
rect 17666 8318 17668 8370
rect 17500 8316 17668 8318
rect 17612 8306 17668 8316
rect 17276 8206 17278 8258
rect 17330 8206 17332 8258
rect 17276 8194 17332 8206
rect 17388 8258 17444 8270
rect 17388 8206 17390 8258
rect 17442 8206 17444 8258
rect 17052 7812 17108 7822
rect 17052 7586 17108 7756
rect 17388 7700 17444 8206
rect 17388 7634 17444 7644
rect 17500 8146 17556 8158
rect 17500 8094 17502 8146
rect 17554 8094 17556 8146
rect 17052 7534 17054 7586
rect 17106 7534 17108 7586
rect 17052 7522 17108 7534
rect 16940 7476 16996 7486
rect 16940 5906 16996 7420
rect 17388 7476 17444 7486
rect 17388 7382 17444 7420
rect 16940 5854 16942 5906
rect 16994 5854 16996 5906
rect 16940 5842 16996 5854
rect 16828 5628 16996 5684
rect 15932 5182 15934 5234
rect 15986 5182 15988 5234
rect 15932 5170 15988 5182
rect 13244 5124 13300 5134
rect 13132 5122 13300 5124
rect 13132 5070 13246 5122
rect 13298 5070 13300 5122
rect 13132 5068 13300 5070
rect 13244 5058 13300 5068
rect 16828 4564 16884 4574
rect 15484 4452 15540 4462
rect 12012 3332 12180 3388
rect 12572 3332 12852 3388
rect 11452 2212 11508 2222
rect 11452 2098 11508 2156
rect 11452 2046 11454 2098
rect 11506 2046 11508 2098
rect 11452 2034 11508 2046
rect 12012 1986 12068 1998
rect 12012 1934 12014 1986
rect 12066 1934 12068 1986
rect 12012 1764 12068 1934
rect 12012 1698 12068 1708
rect 12124 1092 12180 3332
rect 12124 1026 12180 1036
rect 11452 196 11508 206
rect 11452 112 11508 140
rect 12796 112 12852 3332
rect 13244 2100 13300 2110
rect 13244 2006 13300 2044
rect 13804 1988 13860 1998
rect 13804 1894 13860 1932
rect 14140 980 14196 990
rect 14140 112 14196 924
rect 15484 112 15540 4396
rect 16828 112 16884 4508
rect 16940 4116 16996 5628
rect 17500 4228 17556 8094
rect 17724 5236 17780 8652
rect 17724 5170 17780 5180
rect 18060 4900 18116 11788
rect 18172 11394 18228 12908
rect 18396 12870 18452 12908
rect 18396 12738 18452 12750
rect 18396 12686 18398 12738
rect 18450 12686 18452 12738
rect 18284 12404 18340 12414
rect 18396 12404 18452 12686
rect 18284 12402 18452 12404
rect 18284 12350 18286 12402
rect 18338 12350 18452 12402
rect 18284 12348 18452 12350
rect 18284 12338 18340 12348
rect 18732 12292 18788 12302
rect 18620 12290 18788 12292
rect 18620 12238 18734 12290
rect 18786 12238 18788 12290
rect 18620 12236 18788 12238
rect 18508 12180 18564 12190
rect 18508 12086 18564 12124
rect 18508 11956 18564 11966
rect 18508 11788 18564 11900
rect 18284 11732 18564 11788
rect 18620 11788 18676 12236
rect 18732 12226 18788 12236
rect 18732 11956 18788 11966
rect 18844 11956 18900 14476
rect 19068 14420 19124 16156
rect 19404 16098 19460 16492
rect 19740 16548 19796 16606
rect 19740 16482 19796 16492
rect 19852 16324 19908 17276
rect 19964 17108 20020 17118
rect 19964 17014 20020 17052
rect 19964 16324 20020 16334
rect 19852 16322 20020 16324
rect 19852 16270 19966 16322
rect 20018 16270 20020 16322
rect 19852 16268 20020 16270
rect 19964 16258 20020 16268
rect 19404 16046 19406 16098
rect 19458 16046 19460 16098
rect 19404 16034 19460 16046
rect 19740 16212 19796 16222
rect 19740 16098 19796 16156
rect 19740 16046 19742 16098
rect 19794 16046 19796 16098
rect 19740 15652 19796 16046
rect 19740 15586 19796 15596
rect 19740 15426 19796 15438
rect 19740 15374 19742 15426
rect 19794 15374 19796 15426
rect 19180 15316 19236 15326
rect 19180 15222 19236 15260
rect 19740 15148 19796 15374
rect 20076 15428 20132 17614
rect 20076 15362 20132 15372
rect 20188 15652 20244 15662
rect 19292 15092 19796 15148
rect 20076 15204 20132 15242
rect 20076 15138 20132 15148
rect 19852 15092 19908 15102
rect 19180 14644 19236 14654
rect 19180 14550 19236 14588
rect 19068 14364 19236 14420
rect 19068 14084 19124 14094
rect 19068 13970 19124 14028
rect 19068 13918 19070 13970
rect 19122 13918 19124 13970
rect 19068 13906 19124 13918
rect 19180 13074 19236 14364
rect 19292 13970 19348 15092
rect 19852 15090 20020 15092
rect 19852 15038 19854 15090
rect 19906 15038 20020 15090
rect 19852 15036 20020 15038
rect 19852 15026 19908 15036
rect 19964 14756 20020 15036
rect 20188 14980 20244 15596
rect 19964 14690 20020 14700
rect 20076 14924 20244 14980
rect 19964 14532 20020 14542
rect 19964 14308 20020 14476
rect 19964 14242 20020 14252
rect 19292 13918 19294 13970
rect 19346 13918 19348 13970
rect 19292 13906 19348 13918
rect 19516 14084 19572 14094
rect 19180 13022 19182 13074
rect 19234 13022 19236 13074
rect 18956 12628 19012 12638
rect 18956 12178 19012 12572
rect 18956 12126 18958 12178
rect 19010 12126 19012 12178
rect 18956 12114 19012 12126
rect 19180 11956 19236 13022
rect 19516 13748 19572 14028
rect 19516 12962 19572 13692
rect 19516 12910 19518 12962
rect 19570 12910 19572 12962
rect 19292 12628 19348 12638
rect 19292 12292 19348 12572
rect 19516 12628 19572 12910
rect 19628 13746 19684 13758
rect 19628 13694 19630 13746
rect 19682 13694 19684 13746
rect 19628 12852 19684 13694
rect 19964 13636 20020 13646
rect 19964 13542 20020 13580
rect 19740 13524 19796 13534
rect 19740 13430 19796 13468
rect 19852 13522 19908 13534
rect 19852 13470 19854 13522
rect 19906 13470 19908 13522
rect 19684 12796 19796 12852
rect 19628 12786 19684 12796
rect 19516 12562 19572 12572
rect 19516 12292 19572 12302
rect 19292 12290 19572 12292
rect 19292 12238 19518 12290
rect 19570 12238 19572 12290
rect 19292 12236 19572 12238
rect 19516 12226 19572 12236
rect 19628 12292 19684 12302
rect 19628 12178 19684 12236
rect 19628 12126 19630 12178
rect 19682 12126 19684 12178
rect 19628 12114 19684 12126
rect 18844 11900 19124 11956
rect 19180 11900 19348 11956
rect 18732 11862 18788 11900
rect 19068 11844 19124 11900
rect 19068 11788 19236 11844
rect 18620 11732 19012 11788
rect 18284 11508 18340 11732
rect 18732 11618 18788 11630
rect 18732 11566 18734 11618
rect 18786 11566 18788 11618
rect 18732 11508 18788 11566
rect 18844 11508 18900 11518
rect 18732 11452 18844 11508
rect 18284 11442 18340 11452
rect 18844 11442 18900 11452
rect 18172 11342 18174 11394
rect 18226 11342 18228 11394
rect 18172 10164 18228 11342
rect 18396 11396 18452 11406
rect 18284 10836 18340 10846
rect 18284 10742 18340 10780
rect 18172 10098 18228 10108
rect 18396 9826 18452 11340
rect 18620 11396 18676 11406
rect 18620 11394 18788 11396
rect 18620 11342 18622 11394
rect 18674 11342 18788 11394
rect 18620 11340 18788 11342
rect 18620 11330 18676 11340
rect 18732 10948 18788 11340
rect 18956 11060 19012 11732
rect 19180 11620 19236 11788
rect 18956 10994 19012 11004
rect 19068 11564 19236 11620
rect 18732 10882 18788 10892
rect 18396 9774 18398 9826
rect 18450 9774 18452 9826
rect 18396 9762 18452 9774
rect 18620 10612 18676 10622
rect 18172 9380 18228 9390
rect 18172 8930 18228 9324
rect 18620 9154 18676 10556
rect 18956 10052 19012 10062
rect 18956 9958 19012 9996
rect 18620 9102 18622 9154
rect 18674 9102 18676 9154
rect 18620 9090 18676 9102
rect 18844 9826 18900 9838
rect 18844 9774 18846 9826
rect 18898 9774 18900 9826
rect 18172 8878 18174 8930
rect 18226 8878 18228 8930
rect 18172 8866 18228 8878
rect 18060 4834 18116 4844
rect 18508 8372 18564 8382
rect 17500 4162 17556 4172
rect 16940 4050 16996 4060
rect 18172 644 18228 654
rect 18172 112 18228 588
rect 18508 308 18564 8316
rect 18844 8260 18900 9774
rect 18844 8036 18900 8204
rect 18844 7970 18900 7980
rect 19068 3444 19124 11564
rect 19180 11396 19236 11406
rect 19180 11302 19236 11340
rect 19292 8932 19348 11900
rect 19404 11954 19460 11966
rect 19404 11902 19406 11954
rect 19458 11902 19460 11954
rect 19404 11508 19460 11902
rect 19740 11956 19796 12796
rect 19740 11890 19796 11900
rect 19404 11442 19460 11452
rect 19516 11844 19572 11854
rect 19404 10500 19460 10510
rect 19404 10406 19460 10444
rect 19404 10164 19460 10174
rect 19404 9938 19460 10108
rect 19404 9886 19406 9938
rect 19458 9886 19460 9938
rect 19404 9874 19460 9886
rect 19292 8866 19348 8876
rect 19516 9716 19572 11788
rect 19628 10836 19684 10846
rect 19852 10836 19908 13470
rect 20076 12962 20132 14924
rect 20188 13076 20244 13086
rect 20188 12982 20244 13020
rect 20076 12910 20078 12962
rect 20130 12910 20132 12962
rect 19964 12180 20020 12190
rect 19964 12086 20020 12124
rect 19964 11396 20020 11406
rect 19964 11302 20020 11340
rect 19628 10164 19684 10780
rect 19628 10098 19684 10108
rect 19740 10780 19908 10836
rect 20076 10948 20132 12910
rect 19516 8146 19572 9660
rect 19628 8932 19684 8942
rect 19628 8260 19684 8876
rect 19628 8194 19684 8204
rect 19516 8094 19518 8146
rect 19570 8094 19572 8146
rect 19516 6020 19572 8094
rect 19740 7924 19796 10780
rect 19964 10724 20020 10734
rect 19964 10610 20020 10668
rect 19964 10558 19966 10610
rect 20018 10558 20020 10610
rect 19964 10546 20020 10558
rect 19852 10164 19908 10174
rect 19852 8258 19908 10108
rect 19852 8206 19854 8258
rect 19906 8206 19908 8258
rect 19852 8194 19908 8206
rect 19964 9826 20020 9838
rect 19964 9774 19966 9826
rect 20018 9774 20020 9826
rect 19740 7858 19796 7868
rect 19964 7924 20020 9774
rect 20076 8820 20132 10892
rect 20076 8754 20132 8764
rect 20188 12628 20244 12638
rect 20188 8372 20244 12572
rect 20188 8306 20244 8316
rect 19964 7252 20020 7868
rect 19964 7186 20020 7196
rect 20300 8258 20356 18284
rect 20412 17668 20468 17678
rect 20412 16210 20468 17612
rect 20524 16772 20580 19964
rect 20748 19236 20804 20300
rect 20860 20020 20916 21534
rect 20972 21364 21028 23772
rect 21196 21700 21252 24892
rect 21308 22370 21364 25004
rect 21420 23548 21476 26460
rect 21532 24722 21588 26684
rect 21644 24836 21700 26852
rect 21868 26068 21924 30270
rect 21644 24770 21700 24780
rect 21756 25506 21812 25518
rect 21756 25454 21758 25506
rect 21810 25454 21812 25506
rect 21532 24670 21534 24722
rect 21586 24670 21588 24722
rect 21532 24658 21588 24670
rect 21644 24612 21700 24622
rect 21756 24612 21812 25454
rect 21644 24610 21812 24612
rect 21644 24558 21646 24610
rect 21698 24558 21812 24610
rect 21644 24556 21812 24558
rect 21644 24546 21700 24556
rect 21420 23492 21812 23548
rect 21308 22318 21310 22370
rect 21362 22318 21364 22370
rect 21308 22306 21364 22318
rect 21420 22372 21476 22382
rect 21196 21634 21252 21644
rect 21084 21588 21140 21598
rect 21084 21494 21140 21532
rect 20972 21298 21028 21308
rect 21196 20580 21252 20590
rect 20972 20132 21028 20142
rect 20972 20038 21028 20076
rect 20860 19954 20916 19964
rect 20860 19796 20916 19806
rect 20860 19702 20916 19740
rect 20860 19236 20916 19246
rect 20748 19234 20916 19236
rect 20748 19182 20862 19234
rect 20914 19182 20916 19234
rect 20748 19180 20916 19182
rect 20860 19170 20916 19180
rect 20972 18452 21028 18462
rect 20860 18450 21028 18452
rect 20860 18398 20974 18450
rect 21026 18398 21028 18450
rect 20860 18396 21028 18398
rect 20636 18338 20692 18350
rect 20636 18286 20638 18338
rect 20690 18286 20692 18338
rect 20636 18116 20692 18286
rect 20636 18050 20692 18060
rect 20860 17668 20916 18396
rect 20972 18386 21028 18396
rect 20860 17602 20916 17612
rect 20972 17668 21028 17678
rect 20972 17666 21140 17668
rect 20972 17614 20974 17666
rect 21026 17614 21140 17666
rect 20972 17612 21140 17614
rect 20972 17602 21028 17612
rect 20972 17332 21028 17342
rect 20972 17106 21028 17276
rect 20972 17054 20974 17106
rect 21026 17054 21028 17106
rect 20972 17042 21028 17054
rect 20524 16706 20580 16716
rect 20748 16658 20804 16670
rect 20748 16606 20750 16658
rect 20802 16606 20804 16658
rect 20412 16158 20414 16210
rect 20466 16158 20468 16210
rect 20412 16146 20468 16158
rect 20636 16436 20692 16446
rect 20636 15428 20692 16380
rect 20748 15652 20804 16606
rect 20860 16660 20916 16670
rect 20860 16566 20916 16604
rect 20748 15596 21028 15652
rect 20300 8206 20302 8258
rect 20354 8206 20356 8258
rect 20300 8036 20356 8206
rect 20412 15426 20692 15428
rect 20412 15374 20638 15426
rect 20690 15374 20692 15426
rect 20412 15372 20692 15374
rect 20412 8148 20468 15372
rect 20636 15362 20692 15372
rect 20972 15314 21028 15596
rect 20972 15262 20974 15314
rect 21026 15262 21028 15314
rect 20860 14756 20916 14766
rect 20748 14530 20804 14542
rect 20748 14478 20750 14530
rect 20802 14478 20804 14530
rect 20748 14420 20804 14478
rect 20748 14354 20804 14364
rect 20860 13748 20916 14700
rect 20972 14084 21028 15262
rect 21084 14420 21140 17612
rect 21084 14354 21140 14364
rect 21196 16098 21252 20524
rect 21308 19122 21364 19134
rect 21308 19070 21310 19122
rect 21362 19070 21364 19122
rect 21308 16436 21364 19070
rect 21420 18450 21476 22316
rect 21420 18398 21422 18450
rect 21474 18398 21476 18450
rect 21420 18340 21476 18398
rect 21532 22370 21588 22382
rect 21532 22318 21534 22370
rect 21586 22318 21588 22370
rect 21532 18452 21588 22318
rect 21756 20804 21812 23492
rect 21868 22484 21924 26012
rect 22316 25618 22372 35420
rect 22428 31778 22484 31790
rect 22428 31726 22430 31778
rect 22482 31726 22484 31778
rect 22428 30996 22484 31726
rect 22652 30996 22708 31006
rect 22428 30994 22708 30996
rect 22428 30942 22654 30994
rect 22706 30942 22708 30994
rect 22428 30940 22708 30942
rect 22652 30930 22708 30940
rect 22428 30772 22484 30782
rect 22428 28642 22484 30716
rect 22428 28590 22430 28642
rect 22482 28590 22484 28642
rect 22428 26908 22484 28590
rect 22428 26852 22596 26908
rect 22316 25566 22318 25618
rect 22370 25566 22372 25618
rect 22316 25554 22372 25566
rect 22428 26066 22484 26078
rect 22428 26014 22430 26066
rect 22482 26014 22484 26066
rect 22316 24724 22372 24734
rect 22428 24724 22484 26014
rect 22316 24722 22484 24724
rect 22316 24670 22318 24722
rect 22370 24670 22484 24722
rect 22316 24668 22484 24670
rect 22316 24658 22372 24668
rect 22092 24164 22148 24174
rect 22540 24164 22596 26852
rect 22092 24070 22148 24108
rect 22428 24108 22596 24164
rect 21868 22418 21924 22428
rect 22316 22370 22372 22382
rect 22316 22318 22318 22370
rect 22370 22318 22372 22370
rect 21980 21812 22036 21822
rect 21980 21586 22036 21756
rect 21980 21534 21982 21586
rect 22034 21534 22036 21586
rect 21980 21522 22036 21534
rect 22092 21810 22148 21822
rect 22092 21758 22094 21810
rect 22146 21758 22148 21810
rect 21756 20710 21812 20748
rect 22092 18564 22148 21758
rect 22204 21586 22260 21598
rect 22204 21534 22206 21586
rect 22258 21534 22260 21586
rect 22204 20132 22260 21534
rect 22204 20066 22260 20076
rect 22092 18498 22148 18508
rect 21532 18386 21588 18396
rect 21756 18452 21812 18462
rect 21420 18274 21476 18284
rect 21644 18226 21700 18238
rect 21644 18174 21646 18226
rect 21698 18174 21700 18226
rect 21532 17668 21588 17678
rect 21532 17574 21588 17612
rect 21644 17108 21700 18174
rect 21644 17042 21700 17052
rect 21308 16370 21364 16380
rect 21196 16046 21198 16098
rect 21250 16046 21252 16098
rect 20972 14018 21028 14028
rect 20636 13636 20692 13646
rect 20524 13634 20692 13636
rect 20524 13582 20638 13634
rect 20690 13582 20692 13634
rect 20524 13580 20692 13582
rect 20524 8370 20580 13580
rect 20636 13570 20692 13580
rect 20860 13634 20916 13692
rect 20860 13582 20862 13634
rect 20914 13582 20916 13634
rect 20860 13570 20916 13582
rect 20972 13636 21028 13646
rect 20748 13524 20804 13534
rect 20748 13430 20804 13468
rect 20860 13412 20916 13422
rect 20636 13076 20692 13086
rect 20636 12178 20692 13020
rect 20860 12962 20916 13356
rect 20860 12910 20862 12962
rect 20914 12910 20916 12962
rect 20860 12898 20916 12910
rect 20972 12740 21028 13580
rect 20748 12684 21028 12740
rect 21196 12962 21252 16046
rect 21532 15764 21588 15774
rect 21420 15540 21476 15550
rect 21420 15314 21476 15484
rect 21420 15262 21422 15314
rect 21474 15262 21476 15314
rect 21420 15250 21476 15262
rect 21196 12910 21198 12962
rect 21250 12910 21252 12962
rect 20748 12290 20804 12684
rect 20748 12238 20750 12290
rect 20802 12238 20804 12290
rect 20748 12226 20804 12238
rect 20636 12126 20638 12178
rect 20690 12126 20692 12178
rect 20636 12114 20692 12126
rect 20860 12180 20916 12218
rect 20860 12114 20916 12124
rect 21084 11956 21140 11966
rect 21084 11862 21140 11900
rect 20860 11394 20916 11406
rect 20860 11342 20862 11394
rect 20914 11342 20916 11394
rect 20860 10052 20916 11342
rect 20860 9986 20916 9996
rect 21196 11396 21252 12910
rect 21084 9826 21140 9838
rect 21084 9774 21086 9826
rect 21138 9774 21140 9826
rect 21084 8484 21140 9774
rect 21084 8418 21140 8428
rect 20524 8318 20526 8370
rect 20578 8318 20580 8370
rect 20524 8306 20580 8318
rect 20972 8372 21028 8382
rect 20972 8278 21028 8316
rect 20412 8092 21140 8148
rect 20300 7252 20356 7980
rect 20300 7186 20356 7196
rect 19516 5954 19572 5964
rect 20860 6804 20916 6814
rect 19068 3378 19124 3388
rect 18508 242 18564 252
rect 19516 420 19572 430
rect 19516 112 19572 364
rect 20860 112 20916 6748
rect 20972 6580 21028 6590
rect 20972 2100 21028 6524
rect 21084 2996 21140 8092
rect 21196 8036 21252 11340
rect 21308 15092 21364 15102
rect 21308 13524 21364 15036
rect 21420 14306 21476 14318
rect 21420 14254 21422 14306
rect 21474 14254 21476 14306
rect 21420 14084 21476 14254
rect 21420 14018 21476 14028
rect 21420 13748 21476 13758
rect 21420 13654 21476 13692
rect 21308 10836 21364 13468
rect 21532 12402 21588 15708
rect 21644 15204 21700 15242
rect 21644 15138 21700 15148
rect 21532 12350 21534 12402
rect 21586 12350 21588 12402
rect 21532 12180 21588 12350
rect 21532 12114 21588 12124
rect 21644 13748 21700 13758
rect 21644 12178 21700 13692
rect 21644 12126 21646 12178
rect 21698 12126 21700 12178
rect 21644 12114 21700 12126
rect 21308 10770 21364 10780
rect 21196 7970 21252 7980
rect 21308 8372 21364 8382
rect 21308 7476 21364 8316
rect 21308 7410 21364 7420
rect 21756 8258 21812 18396
rect 22316 18452 22372 22318
rect 22092 18338 22148 18350
rect 22092 18286 22094 18338
rect 22146 18286 22148 18338
rect 22092 17556 22148 18286
rect 22092 17490 22148 17500
rect 22204 16658 22260 16670
rect 22204 16606 22206 16658
rect 22258 16606 22260 16658
rect 22204 16324 22260 16606
rect 21868 16268 22260 16324
rect 21868 9044 21924 16268
rect 21980 16100 22036 16110
rect 21980 12964 22036 16044
rect 22092 15202 22148 15214
rect 22092 15150 22094 15202
rect 22146 15150 22148 15202
rect 22092 15092 22148 15150
rect 22092 15026 22148 15036
rect 22204 12964 22260 12974
rect 21980 12962 22260 12964
rect 21980 12910 22206 12962
rect 22258 12910 22260 12962
rect 21980 12908 22260 12910
rect 22092 10052 22148 12908
rect 22204 12898 22260 12908
rect 21868 8978 21924 8988
rect 21980 9268 22036 9278
rect 21756 8206 21758 8258
rect 21810 8206 21812 8258
rect 21756 7924 21812 8206
rect 21756 6132 21812 7868
rect 21868 7700 21924 7710
rect 21868 6244 21924 7644
rect 21868 6178 21924 6188
rect 21756 6066 21812 6076
rect 21084 2930 21140 2940
rect 20972 2034 21028 2044
rect 21980 196 22036 9212
rect 22092 7476 22148 9996
rect 22316 8372 22372 18396
rect 22316 8306 22372 8316
rect 22092 7410 22148 7420
rect 22428 3388 22484 24108
rect 22652 24052 22708 24062
rect 22652 23938 22708 23996
rect 22652 23886 22654 23938
rect 22706 23886 22708 23938
rect 22652 23874 22708 23886
rect 22652 18450 22708 18462
rect 22652 18398 22654 18450
rect 22706 18398 22708 18450
rect 22652 18340 22708 18398
rect 22652 18274 22708 18284
rect 22652 17778 22708 17790
rect 22652 17726 22654 17778
rect 22706 17726 22708 17778
rect 22652 17556 22708 17726
rect 22764 17780 22820 37660
rect 23212 31778 23268 31790
rect 23212 31726 23214 31778
rect 23266 31726 23268 31778
rect 23212 31332 23268 31726
rect 23212 31266 23268 31276
rect 22876 30994 22932 31006
rect 22876 30942 22878 30994
rect 22930 30942 22932 30994
rect 22876 29876 22932 30942
rect 23100 30212 23156 30222
rect 23100 30118 23156 30156
rect 22876 29820 23268 29876
rect 23100 29428 23156 29438
rect 22876 24724 22932 24734
rect 22876 24722 23044 24724
rect 22876 24670 22878 24722
rect 22930 24670 23044 24722
rect 22876 24668 23044 24670
rect 22876 24658 22932 24668
rect 22764 17714 22820 17724
rect 22876 22484 22932 22494
rect 22876 22370 22932 22428
rect 22876 22318 22878 22370
rect 22930 22318 22932 22370
rect 22876 17556 22932 22318
rect 22652 17500 22932 17556
rect 22540 16884 22596 16894
rect 22540 15540 22596 16828
rect 22988 16884 23044 24668
rect 23100 24050 23156 29372
rect 23100 23998 23102 24050
rect 23154 23998 23156 24050
rect 23100 23986 23156 23998
rect 23212 20580 23268 29820
rect 23212 20514 23268 20524
rect 23324 20132 23380 55244
rect 23548 50482 23604 55916
rect 23884 55970 23940 55982
rect 23884 55918 23886 55970
rect 23938 55918 23940 55970
rect 23884 55748 23940 55918
rect 23884 55682 23940 55692
rect 23804 54908 24068 54918
rect 23860 54852 23908 54908
rect 23964 54852 24012 54908
rect 23804 54842 24068 54852
rect 23772 54740 23828 54750
rect 23772 54646 23828 54684
rect 23660 54628 23716 54638
rect 23660 52050 23716 54572
rect 24108 54514 24164 54526
rect 24108 54462 24110 54514
rect 24162 54462 24164 54514
rect 23772 54404 23828 54414
rect 23772 53618 23828 54348
rect 24108 54180 24164 54462
rect 24108 54114 24164 54124
rect 23772 53566 23774 53618
rect 23826 53566 23828 53618
rect 23772 53554 23828 53566
rect 23804 53340 24068 53350
rect 23860 53284 23908 53340
rect 23964 53284 24012 53340
rect 23804 53274 24068 53284
rect 24108 53172 24164 53182
rect 24220 53172 24276 56700
rect 24332 54628 24388 57148
rect 24444 56308 24500 56318
rect 24444 56214 24500 56252
rect 24892 56308 24948 57344
rect 24892 56242 24948 56252
rect 25452 55972 25508 55982
rect 25452 55878 25508 55916
rect 24464 55692 24728 55702
rect 24520 55636 24568 55692
rect 24624 55636 24672 55692
rect 24464 55626 24728 55636
rect 25004 55412 25060 55422
rect 24668 55300 24724 55310
rect 24668 55206 24724 55244
rect 24332 54562 24388 54572
rect 24668 54402 24724 54414
rect 24668 54350 24670 54402
rect 24722 54350 24724 54402
rect 24668 54292 24724 54350
rect 25004 54404 25060 55356
rect 25564 54626 25620 57372
rect 25900 57316 25956 57372
rect 26208 57344 26320 57456
rect 27552 57344 27664 57456
rect 25900 57250 25956 57260
rect 26236 57316 26292 57344
rect 26236 57250 26292 57260
rect 27580 56644 27636 57344
rect 27580 56578 27636 56588
rect 26012 56308 26068 56318
rect 26012 56214 26068 56252
rect 25788 56196 25844 56206
rect 25564 54574 25566 54626
rect 25618 54574 25620 54626
rect 25564 54562 25620 54574
rect 25676 55074 25732 55086
rect 25676 55022 25678 55074
rect 25730 55022 25732 55074
rect 25676 54516 25732 55022
rect 25676 54450 25732 54460
rect 25004 54338 25060 54348
rect 24668 54226 24724 54236
rect 24464 54124 24728 54134
rect 24520 54068 24568 54124
rect 24624 54068 24672 54124
rect 24464 54058 24728 54068
rect 24668 53730 24724 53742
rect 24668 53678 24670 53730
rect 24722 53678 24724 53730
rect 24668 53620 24724 53678
rect 24668 53554 24724 53564
rect 25676 53620 25732 53630
rect 25676 53526 25732 53564
rect 24108 53170 24276 53172
rect 24108 53118 24110 53170
rect 24162 53118 24276 53170
rect 24108 53116 24276 53118
rect 24108 53106 24164 53116
rect 24668 52834 24724 52846
rect 24668 52782 24670 52834
rect 24722 52782 24724 52834
rect 24668 52724 24724 52782
rect 24668 52658 24724 52668
rect 25452 52834 25508 52846
rect 25452 52782 25454 52834
rect 25506 52782 25508 52834
rect 25452 52724 25508 52782
rect 25452 52658 25508 52668
rect 24464 52556 24728 52566
rect 24520 52500 24568 52556
rect 24624 52500 24672 52556
rect 24464 52490 24728 52500
rect 24668 52276 24724 52286
rect 24668 52182 24724 52220
rect 23660 51998 23662 52050
rect 23714 51998 23716 52050
rect 23660 51986 23716 51998
rect 25676 51938 25732 51950
rect 25676 51886 25678 51938
rect 25730 51886 25732 51938
rect 25676 51828 25732 51886
rect 23804 51772 24068 51782
rect 23860 51716 23908 51772
rect 23964 51716 24012 51772
rect 25676 51762 25732 51772
rect 23804 51706 24068 51716
rect 25676 51604 25732 51614
rect 25788 51604 25844 56140
rect 26460 55298 26516 55310
rect 26460 55246 26462 55298
rect 26514 55246 26516 55298
rect 26236 54402 26292 54414
rect 26236 54350 26238 54402
rect 26290 54350 26292 54402
rect 26236 53956 26292 54350
rect 26236 53890 26292 53900
rect 26236 53730 26292 53742
rect 26236 53678 26238 53730
rect 26290 53678 26292 53730
rect 26236 53508 26292 53678
rect 26236 53442 26292 53452
rect 26236 52836 26292 52846
rect 26236 52742 26292 52780
rect 26236 52164 26292 52174
rect 25676 51602 25844 51604
rect 25676 51550 25678 51602
rect 25730 51550 25844 51602
rect 25676 51548 25844 51550
rect 25900 52162 26292 52164
rect 25900 52110 26238 52162
rect 26290 52110 26292 52162
rect 25900 52108 26292 52110
rect 25676 51538 25732 51548
rect 24668 51268 24724 51278
rect 24668 51174 24724 51212
rect 24464 50988 24728 50998
rect 24520 50932 24568 50988
rect 24624 50932 24672 50988
rect 24464 50922 24728 50932
rect 23996 50596 24052 50606
rect 23996 50502 24052 50540
rect 24668 50594 24724 50606
rect 24668 50542 24670 50594
rect 24722 50542 24724 50594
rect 23548 50430 23550 50482
rect 23602 50430 23604 50482
rect 23548 50418 23604 50430
rect 24668 50484 24724 50542
rect 24668 50418 24724 50428
rect 25676 50484 25732 50494
rect 25676 50390 25732 50428
rect 23804 50204 24068 50214
rect 23860 50148 23908 50204
rect 23964 50148 24012 50204
rect 23804 50138 24068 50148
rect 25676 49922 25732 49934
rect 25676 49870 25678 49922
rect 25730 49870 25732 49922
rect 24668 49700 24724 49710
rect 24668 49606 24724 49644
rect 25676 49588 25732 49870
rect 25676 49522 25732 49532
rect 24464 49420 24728 49430
rect 24520 49364 24568 49420
rect 24624 49364 24672 49420
rect 24464 49354 24728 49364
rect 24668 49028 24724 49038
rect 24668 48934 24724 48972
rect 25676 48802 25732 48814
rect 25676 48750 25678 48802
rect 25730 48750 25732 48802
rect 25676 48692 25732 48750
rect 23804 48636 24068 48646
rect 23860 48580 23908 48636
rect 23964 48580 24012 48636
rect 25676 48626 25732 48636
rect 23804 48570 24068 48580
rect 24464 47852 24728 47862
rect 24520 47796 24568 47852
rect 24624 47796 24672 47852
rect 24464 47786 24728 47796
rect 24668 47458 24724 47470
rect 24668 47406 24670 47458
rect 24722 47406 24724 47458
rect 24668 47348 24724 47406
rect 24668 47282 24724 47292
rect 25676 47348 25732 47358
rect 25676 47254 25732 47292
rect 23804 47068 24068 47078
rect 23860 47012 23908 47068
rect 23964 47012 24012 47068
rect 23804 47002 24068 47012
rect 25676 46786 25732 46798
rect 25676 46734 25678 46786
rect 25730 46734 25732 46786
rect 24668 46564 24724 46574
rect 24332 46562 24724 46564
rect 24332 46510 24670 46562
rect 24722 46510 24724 46562
rect 24332 46508 24724 46510
rect 23804 45500 24068 45510
rect 23860 45444 23908 45500
rect 23964 45444 24012 45500
rect 23804 45434 24068 45444
rect 23804 43932 24068 43942
rect 23860 43876 23908 43932
rect 23964 43876 24012 43932
rect 23804 43866 24068 43876
rect 23804 42364 24068 42374
rect 23860 42308 23908 42364
rect 23964 42308 24012 42364
rect 23804 42298 24068 42308
rect 24332 41972 24388 46508
rect 24668 46498 24724 46508
rect 25676 46452 25732 46734
rect 25900 46788 25956 52108
rect 26236 52098 26292 52108
rect 26460 51492 26516 55246
rect 27244 55074 27300 55086
rect 27244 55022 27246 55074
rect 27298 55022 27300 55074
rect 27020 54402 27076 54414
rect 27020 54350 27022 54402
rect 27074 54350 27076 54402
rect 27020 53172 27076 54350
rect 27244 54068 27300 55022
rect 27244 54002 27300 54012
rect 27020 53106 27076 53116
rect 27244 53506 27300 53518
rect 27244 53454 27246 53506
rect 27298 53454 27300 53506
rect 26460 51426 26516 51436
rect 27132 53058 27188 53070
rect 27132 53006 27134 53058
rect 27186 53006 27188 53058
rect 26348 51378 26404 51390
rect 26348 51326 26350 51378
rect 26402 51326 26404 51378
rect 26236 50594 26292 50606
rect 26236 50542 26238 50594
rect 26290 50542 26292 50594
rect 26236 49924 26292 50542
rect 26236 49858 26292 49868
rect 26236 49028 26292 49038
rect 25900 46722 25956 46732
rect 26012 49026 26292 49028
rect 26012 48974 26238 49026
rect 26290 48974 26292 49026
rect 26012 48972 26292 48974
rect 25676 46386 25732 46396
rect 24464 46284 24728 46294
rect 24520 46228 24568 46284
rect 24624 46228 24672 46284
rect 24464 46218 24728 46228
rect 24892 45890 24948 45902
rect 24892 45838 24894 45890
rect 24946 45838 24948 45890
rect 24464 44716 24728 44726
rect 24520 44660 24568 44716
rect 24624 44660 24672 44716
rect 24464 44650 24728 44660
rect 24892 44548 24948 45838
rect 25676 45666 25732 45678
rect 25676 45614 25678 45666
rect 25730 45614 25732 45666
rect 25676 45556 25732 45614
rect 25676 45490 25732 45500
rect 24892 44482 24948 44492
rect 24892 44322 24948 44334
rect 24892 44270 24894 44322
rect 24946 44270 24948 44322
rect 24892 43708 24948 44270
rect 25676 44212 25732 44222
rect 25676 44118 25732 44156
rect 24892 43652 25060 43708
rect 24892 43538 24948 43550
rect 24892 43486 24894 43538
rect 24946 43486 24948 43538
rect 24464 43148 24728 43158
rect 24520 43092 24568 43148
rect 24624 43092 24672 43148
rect 24464 43082 24728 43092
rect 24332 41906 24388 41916
rect 24668 42754 24724 42766
rect 24668 42702 24670 42754
rect 24722 42702 24724 42754
rect 24668 41748 24724 42702
rect 24668 41682 24724 41692
rect 24464 41580 24728 41590
rect 24520 41524 24568 41580
rect 24624 41524 24672 41580
rect 24464 41514 24728 41524
rect 24780 41186 24836 41198
rect 24780 41134 24782 41186
rect 24834 41134 24836 41186
rect 23804 40796 24068 40806
rect 23860 40740 23908 40796
rect 23964 40740 24012 40796
rect 23804 40730 24068 40740
rect 24668 40404 24724 40414
rect 24668 40310 24724 40348
rect 24780 40180 24836 41134
rect 24780 40114 24836 40124
rect 24464 40012 24728 40022
rect 24520 39956 24568 40012
rect 24624 39956 24672 40012
rect 24464 39946 24728 39956
rect 24892 39844 24948 43486
rect 24892 39778 24948 39788
rect 24892 39618 24948 39630
rect 24892 39566 24894 39618
rect 24946 39566 24948 39618
rect 23804 39228 24068 39238
rect 23860 39172 23908 39228
rect 23964 39172 24012 39228
rect 23804 39162 24068 39172
rect 24464 38444 24728 38454
rect 24520 38388 24568 38444
rect 24624 38388 24672 38444
rect 24464 38378 24728 38388
rect 24668 38050 24724 38062
rect 24668 37998 24670 38050
rect 24722 37998 24724 38050
rect 23804 37660 24068 37670
rect 23860 37604 23908 37660
rect 23964 37604 24012 37660
rect 23804 37594 24068 37604
rect 24668 37492 24724 37998
rect 24668 37426 24724 37436
rect 24668 37154 24724 37166
rect 24668 37102 24670 37154
rect 24722 37102 24724 37154
rect 24668 37044 24724 37102
rect 24668 36978 24724 36988
rect 24464 36876 24728 36886
rect 24520 36820 24568 36876
rect 24624 36820 24672 36876
rect 24464 36810 24728 36820
rect 24668 36708 24724 36718
rect 24668 36594 24724 36652
rect 24668 36542 24670 36594
rect 24722 36542 24724 36594
rect 24668 36530 24724 36542
rect 23804 36092 24068 36102
rect 23860 36036 23908 36092
rect 23964 36036 24012 36092
rect 23804 36026 24068 36036
rect 24892 35476 24948 39566
rect 25004 35812 25060 43652
rect 25676 43650 25732 43662
rect 25676 43598 25678 43650
rect 25730 43598 25732 43650
rect 25676 43316 25732 43598
rect 25676 43250 25732 43260
rect 25676 42530 25732 42542
rect 25676 42478 25678 42530
rect 25730 42478 25732 42530
rect 25676 42420 25732 42478
rect 25676 42354 25732 42364
rect 25676 41076 25732 41086
rect 25676 40982 25732 41020
rect 25788 40964 25844 40974
rect 25676 40514 25732 40526
rect 25676 40462 25678 40514
rect 25730 40462 25732 40514
rect 25676 40180 25732 40462
rect 25676 40114 25732 40124
rect 25676 39394 25732 39406
rect 25676 39342 25678 39394
rect 25730 39342 25732 39394
rect 25676 39284 25732 39342
rect 25676 39218 25732 39228
rect 25004 35746 25060 35756
rect 25340 38724 25396 38734
rect 24892 35410 24948 35420
rect 24464 35308 24728 35318
rect 24520 35252 24568 35308
rect 24624 35252 24672 35308
rect 24464 35242 24728 35252
rect 24668 34916 24724 34926
rect 24332 34914 24724 34916
rect 24332 34862 24670 34914
rect 24722 34862 24724 34914
rect 24332 34860 24724 34862
rect 23804 34524 24068 34534
rect 23860 34468 23908 34524
rect 23964 34468 24012 34524
rect 23804 34458 24068 34468
rect 23436 33684 23492 33694
rect 23436 22482 23492 33628
rect 23804 32956 24068 32966
rect 23860 32900 23908 32956
rect 23964 32900 24012 32956
rect 23804 32890 24068 32900
rect 24332 31556 24388 34860
rect 24668 34850 24724 34860
rect 24668 34018 24724 34030
rect 24668 33966 24670 34018
rect 24722 33966 24724 34018
rect 24668 33908 24724 33966
rect 24668 33842 24724 33852
rect 25228 34020 25284 34030
rect 24464 33740 24728 33750
rect 24520 33684 24568 33740
rect 24624 33684 24672 33740
rect 24464 33674 24728 33684
rect 24892 33572 24948 33582
rect 24668 33346 24724 33358
rect 24668 33294 24670 33346
rect 24722 33294 24724 33346
rect 24668 33236 24724 33294
rect 24668 33170 24724 33180
rect 24464 32172 24728 32182
rect 24520 32116 24568 32172
rect 24624 32116 24672 32172
rect 24464 32106 24728 32116
rect 24892 31778 24948 33516
rect 24892 31726 24894 31778
rect 24946 31726 24948 31778
rect 24892 31714 24948 31726
rect 24332 31490 24388 31500
rect 23804 31388 24068 31398
rect 23660 31332 23716 31342
rect 23860 31332 23908 31388
rect 23964 31332 24012 31388
rect 23804 31322 24068 31332
rect 23660 30996 23716 31276
rect 23660 30902 23716 30940
rect 24892 30994 24948 31006
rect 24892 30942 24894 30994
rect 24946 30942 24948 30994
rect 24464 30604 24728 30614
rect 24520 30548 24568 30604
rect 24624 30548 24672 30604
rect 24464 30538 24728 30548
rect 23804 29820 24068 29830
rect 23860 29764 23908 29820
rect 23964 29764 24012 29820
rect 23804 29754 24068 29764
rect 24464 29036 24728 29046
rect 24520 28980 24568 29036
rect 24624 28980 24672 29036
rect 24464 28970 24728 28980
rect 23436 22430 23438 22482
rect 23490 22430 23492 22482
rect 23436 22418 23492 22430
rect 23548 28420 23604 28430
rect 23436 22036 23492 22046
rect 23436 21700 23492 21980
rect 23548 21812 23604 28364
rect 23804 28252 24068 28262
rect 23860 28196 23908 28252
rect 23964 28196 24012 28252
rect 23804 28186 24068 28196
rect 24668 27748 24724 27758
rect 24332 27746 24724 27748
rect 24332 27694 24670 27746
rect 24722 27694 24724 27746
rect 24332 27692 24724 27694
rect 24332 27300 24388 27692
rect 24668 27682 24724 27692
rect 24464 27468 24728 27478
rect 24520 27412 24568 27468
rect 24624 27412 24672 27468
rect 24464 27402 24728 27412
rect 24332 27234 24388 27244
rect 24668 27074 24724 27086
rect 24668 27022 24670 27074
rect 24722 27022 24724 27074
rect 24668 26908 24724 27022
rect 24220 26852 24724 26908
rect 24892 26908 24948 30942
rect 25116 30996 25172 31006
rect 24892 26852 25060 26908
rect 23804 26684 24068 26694
rect 23860 26628 23908 26684
rect 23964 26628 24012 26684
rect 23804 26618 24068 26628
rect 23804 25116 24068 25126
rect 23860 25060 23908 25116
rect 23964 25060 24012 25116
rect 23804 25050 24068 25060
rect 23772 24722 23828 24734
rect 23772 24670 23774 24722
rect 23826 24670 23828 24722
rect 23772 23940 23828 24670
rect 23772 23874 23828 23884
rect 23804 23548 24068 23558
rect 23660 23492 23716 23502
rect 23860 23492 23908 23548
rect 23964 23492 24012 23548
rect 23804 23482 24068 23492
rect 23660 22036 23716 23436
rect 23660 21970 23716 21980
rect 23804 21980 24068 21990
rect 23860 21924 23908 21980
rect 23964 21924 24012 21980
rect 23804 21914 24068 21924
rect 23548 21756 23940 21812
rect 23436 21644 23604 21700
rect 23212 20076 23380 20132
rect 23548 21586 23604 21644
rect 23884 21698 23940 21756
rect 23884 21646 23886 21698
rect 23938 21646 23940 21698
rect 23884 21634 23940 21646
rect 23548 21534 23550 21586
rect 23602 21534 23604 21586
rect 22988 16818 23044 16828
rect 23100 17554 23156 17566
rect 23100 17502 23102 17554
rect 23154 17502 23156 17554
rect 22540 15474 22596 15484
rect 22876 15314 22932 15326
rect 22876 15262 22878 15314
rect 22930 15262 22932 15314
rect 22652 15092 22708 15102
rect 22540 14868 22596 14878
rect 22540 14754 22596 14812
rect 22540 14702 22542 14754
rect 22594 14702 22596 14754
rect 22540 14690 22596 14702
rect 22652 13634 22708 15036
rect 22652 13582 22654 13634
rect 22706 13582 22708 13634
rect 22652 13570 22708 13582
rect 22876 14532 22932 15262
rect 23100 15148 23156 17502
rect 22540 11956 22596 11966
rect 22540 11954 22708 11956
rect 22540 11902 22542 11954
rect 22594 11902 22708 11954
rect 22540 11900 22708 11902
rect 22540 11890 22596 11900
rect 22540 8372 22596 8382
rect 22540 8258 22596 8316
rect 22540 8206 22542 8258
rect 22594 8206 22596 8258
rect 22540 5684 22596 8206
rect 22652 6916 22708 11900
rect 22652 6850 22708 6860
rect 22540 5618 22596 5628
rect 22876 3388 22932 14476
rect 22988 15092 23156 15148
rect 22988 14418 23044 15092
rect 22988 14366 22990 14418
rect 23042 14366 23044 14418
rect 22988 13746 23044 14366
rect 22988 13694 22990 13746
rect 23042 13694 23044 13746
rect 22988 10724 23044 13694
rect 22988 10658 23044 10668
rect 23100 12292 23156 12302
rect 23100 3556 23156 12236
rect 23212 11620 23268 20076
rect 23324 18788 23380 18798
rect 23324 16770 23380 18732
rect 23324 16718 23326 16770
rect 23378 16718 23380 16770
rect 23324 15092 23380 16718
rect 23324 15026 23380 15036
rect 23436 18564 23492 18574
rect 23212 11554 23268 11564
rect 23324 14868 23380 14878
rect 23324 11956 23380 14812
rect 23436 12292 23492 18508
rect 23548 14532 23604 21534
rect 23804 20412 24068 20422
rect 23860 20356 23908 20412
rect 23964 20356 24012 20412
rect 23804 20346 24068 20356
rect 24220 19796 24276 26852
rect 25004 26292 25060 26852
rect 25004 26226 25060 26236
rect 24332 26180 24388 26190
rect 24332 24164 24388 26124
rect 24464 25900 24728 25910
rect 24520 25844 24568 25900
rect 24624 25844 24672 25900
rect 24464 25834 24728 25844
rect 24668 25506 24724 25518
rect 24668 25454 24670 25506
rect 24722 25454 24724 25506
rect 24668 24612 24724 25454
rect 25004 24948 25060 24958
rect 24668 24546 24724 24556
rect 24892 24722 24948 24734
rect 24892 24670 24894 24722
rect 24946 24670 24948 24722
rect 24464 24332 24728 24342
rect 24520 24276 24568 24332
rect 24624 24276 24672 24332
rect 24464 24266 24728 24276
rect 24332 24108 24724 24164
rect 24668 24050 24724 24108
rect 24668 23998 24670 24050
rect 24722 23998 24724 24050
rect 24668 23986 24724 23998
rect 24332 23940 24388 23950
rect 24332 19908 24388 23884
rect 24892 23268 24948 24670
rect 24892 23202 24948 23212
rect 24464 22764 24728 22774
rect 24520 22708 24568 22764
rect 24624 22708 24672 22764
rect 24464 22698 24728 22708
rect 24892 22372 24948 22382
rect 25004 22372 25060 24892
rect 24892 22370 25060 22372
rect 24892 22318 24894 22370
rect 24946 22318 25060 22370
rect 24892 22316 25060 22318
rect 24892 22306 24948 22316
rect 24464 21196 24728 21206
rect 24520 21140 24568 21196
rect 24624 21140 24672 21196
rect 24464 21130 24728 21140
rect 24332 19852 25060 19908
rect 24220 19740 24388 19796
rect 24220 19572 24276 19582
rect 23804 18844 24068 18854
rect 23860 18788 23908 18844
rect 23964 18788 24012 18844
rect 23804 18778 24068 18788
rect 23660 18452 23716 18462
rect 23660 18358 23716 18396
rect 23804 17276 24068 17286
rect 23860 17220 23908 17276
rect 23964 17220 24012 17276
rect 23804 17210 24068 17220
rect 23772 16884 23828 16894
rect 23660 16882 23828 16884
rect 23660 16830 23774 16882
rect 23826 16830 23828 16882
rect 23660 16828 23828 16830
rect 23660 15540 23716 16828
rect 23772 16818 23828 16828
rect 23804 15708 24068 15718
rect 23860 15652 23908 15708
rect 23964 15652 24012 15708
rect 23804 15642 24068 15652
rect 23660 15484 23828 15540
rect 23548 14466 23604 14476
rect 23660 15314 23716 15326
rect 23660 15262 23662 15314
rect 23714 15262 23716 15314
rect 23660 14420 23716 15262
rect 23772 14644 23828 15484
rect 24220 15092 24276 19516
rect 24332 16548 24388 19740
rect 24464 19628 24728 19638
rect 24520 19572 24568 19628
rect 24624 19572 24672 19628
rect 24464 19562 24728 19572
rect 25004 19236 25060 19852
rect 25116 19572 25172 30940
rect 25228 24724 25284 33964
rect 25228 24658 25284 24668
rect 25340 21588 25396 38668
rect 25676 37940 25732 37950
rect 25676 37846 25732 37884
rect 25452 37154 25508 37166
rect 25452 37102 25454 37154
rect 25506 37102 25508 37154
rect 25452 37044 25508 37102
rect 25452 36978 25508 36988
rect 25676 36258 25732 36270
rect 25676 36206 25678 36258
rect 25730 36206 25732 36258
rect 25676 36148 25732 36206
rect 25676 36082 25732 36092
rect 25564 34916 25620 34926
rect 25452 30882 25508 30894
rect 25452 30830 25454 30882
rect 25506 30830 25508 30882
rect 25452 30772 25508 30830
rect 25452 30706 25508 30716
rect 25564 26908 25620 34860
rect 25676 34804 25732 34814
rect 25676 34710 25732 34748
rect 25676 34242 25732 34254
rect 25676 34190 25678 34242
rect 25730 34190 25732 34242
rect 25676 33908 25732 34190
rect 25676 33842 25732 33852
rect 25676 33122 25732 33134
rect 25676 33070 25678 33122
rect 25730 33070 25732 33122
rect 25676 33012 25732 33070
rect 25676 32946 25732 32956
rect 25676 31668 25732 31678
rect 25676 31574 25732 31612
rect 25676 27970 25732 27982
rect 25676 27918 25678 27970
rect 25730 27918 25732 27970
rect 25676 27188 25732 27918
rect 25676 27122 25732 27132
rect 25228 21532 25396 21588
rect 25452 26852 25620 26908
rect 25676 26962 25732 26974
rect 25676 26910 25678 26962
rect 25730 26910 25732 26962
rect 25228 21028 25284 21532
rect 25228 20962 25284 20972
rect 25340 21362 25396 21374
rect 25340 21310 25342 21362
rect 25394 21310 25396 21362
rect 25116 19506 25172 19516
rect 25004 19180 25172 19236
rect 24464 18060 24728 18070
rect 24520 18004 24568 18060
rect 24624 18004 24672 18060
rect 24464 17994 24728 18004
rect 24556 17780 24612 17790
rect 24556 17686 24612 17724
rect 25004 17666 25060 17678
rect 25004 17614 25006 17666
rect 25058 17614 25060 17666
rect 24892 16772 24948 16782
rect 24332 16482 24388 16492
rect 24464 16492 24728 16502
rect 24520 16436 24568 16492
rect 24624 16436 24672 16492
rect 24464 16426 24728 16436
rect 24220 15026 24276 15036
rect 24464 14924 24728 14934
rect 24520 14868 24568 14924
rect 24624 14868 24672 14924
rect 24464 14858 24728 14868
rect 23772 14578 23828 14588
rect 24780 14644 24836 14654
rect 24668 14532 24724 14542
rect 23660 14354 23716 14364
rect 24332 14420 24388 14430
rect 23804 14140 24068 14150
rect 23860 14084 23908 14140
rect 23964 14084 24012 14140
rect 23804 14074 24068 14084
rect 23660 13972 23716 13982
rect 23660 13878 23716 13916
rect 24220 13748 24276 13758
rect 23804 12572 24068 12582
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 23804 12506 24068 12516
rect 23436 12226 23492 12236
rect 24108 12180 24164 12190
rect 24220 12180 24276 13692
rect 24108 12178 24276 12180
rect 24108 12126 24110 12178
rect 24162 12126 24276 12178
rect 24108 12124 24276 12126
rect 24108 12068 24164 12124
rect 24108 12002 24164 12012
rect 23660 11956 23716 11966
rect 23324 11954 23716 11956
rect 23324 11902 23662 11954
rect 23714 11902 23716 11954
rect 23324 11900 23716 11902
rect 23324 11394 23380 11900
rect 23660 11890 23716 11900
rect 23772 11620 23828 11630
rect 23772 11506 23828 11564
rect 23772 11454 23774 11506
rect 23826 11454 23828 11506
rect 23772 11442 23828 11454
rect 23324 11342 23326 11394
rect 23378 11342 23380 11394
rect 23324 11330 23380 11342
rect 23804 11004 24068 11014
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 23804 10938 24068 10948
rect 23804 9436 24068 9446
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 23804 9370 24068 9380
rect 23804 7868 24068 7878
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 23804 7802 24068 7812
rect 23804 6300 24068 6310
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 23804 6234 24068 6244
rect 23804 4732 24068 4742
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 23804 4666 24068 4676
rect 23100 3490 23156 3500
rect 22428 3332 22596 3388
rect 21980 130 22036 140
rect 22204 1988 22260 1998
rect 22204 112 22260 1932
rect 22540 1428 22596 3332
rect 22652 3332 22932 3388
rect 22652 2548 22708 3332
rect 23804 3164 24068 3174
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 23804 3098 24068 3108
rect 22652 2482 22708 2492
rect 24332 2100 24388 14364
rect 24668 13636 24724 14476
rect 24780 14418 24836 14588
rect 24780 14366 24782 14418
rect 24834 14366 24836 14418
rect 24780 13860 24836 14366
rect 24780 13794 24836 13804
rect 24780 13636 24836 13646
rect 24668 13634 24836 13636
rect 24668 13582 24782 13634
rect 24834 13582 24836 13634
rect 24668 13580 24836 13582
rect 24780 13570 24836 13580
rect 24464 13356 24728 13366
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24464 13290 24728 13300
rect 24668 12852 24724 12862
rect 24892 12852 24948 16716
rect 25004 14644 25060 17614
rect 25004 14578 25060 14588
rect 25116 17668 25172 19180
rect 25116 13524 25172 17612
rect 25340 15148 25396 21310
rect 25452 15876 25508 26852
rect 25676 26292 25732 26910
rect 25676 26226 25732 26236
rect 25676 25284 25732 25294
rect 25676 25190 25732 25228
rect 25676 24834 25732 24846
rect 25676 24782 25678 24834
rect 25730 24782 25732 24834
rect 25676 24052 25732 24782
rect 25676 23986 25732 23996
rect 25676 23714 25732 23726
rect 25676 23662 25678 23714
rect 25730 23662 25732 23714
rect 25676 23156 25732 23662
rect 25676 23090 25732 23100
rect 25788 22372 25844 40908
rect 26012 36036 26068 48972
rect 26236 48962 26292 48972
rect 26236 48132 26292 48142
rect 26236 48038 26292 48076
rect 26348 47684 26404 51326
rect 27132 51380 27188 53006
rect 27244 52276 27300 53454
rect 27244 52210 27300 52220
rect 27132 51314 27188 51324
rect 27244 51938 27300 51950
rect 27244 51886 27246 51938
rect 27298 51886 27300 51938
rect 27020 51266 27076 51278
rect 27020 51214 27022 51266
rect 27074 51214 27076 51266
rect 27020 50036 27076 51214
rect 27244 50932 27300 51886
rect 27244 50866 27300 50876
rect 27020 49970 27076 49980
rect 27244 50370 27300 50382
rect 27244 50318 27246 50370
rect 27298 50318 27300 50370
rect 27132 49922 27188 49934
rect 27132 49870 27134 49922
rect 27186 49870 27188 49922
rect 26460 49812 26516 49822
rect 26460 49810 26740 49812
rect 26460 49758 26462 49810
rect 26514 49758 26740 49810
rect 26460 49756 26740 49758
rect 26460 49746 26516 49756
rect 26124 47628 26404 47684
rect 26124 40964 26180 47628
rect 26236 47460 26292 47470
rect 26236 47366 26292 47404
rect 26236 46564 26292 46574
rect 26236 46470 26292 46508
rect 26236 45892 26292 45902
rect 26236 45798 26292 45836
rect 26460 45106 26516 45118
rect 26460 45054 26462 45106
rect 26514 45054 26516 45106
rect 26348 44322 26404 44334
rect 26348 44270 26350 44322
rect 26402 44270 26404 44322
rect 26236 43428 26292 43438
rect 26236 43334 26292 43372
rect 26348 42980 26404 44270
rect 26348 42914 26404 42924
rect 26236 42756 26292 42766
rect 26236 42662 26292 42700
rect 26236 41860 26292 41870
rect 26236 41766 26292 41804
rect 26236 41188 26292 41198
rect 26236 41094 26292 41132
rect 26124 40898 26180 40908
rect 26236 40516 26292 40526
rect 26236 40402 26292 40460
rect 26236 40350 26238 40402
rect 26290 40350 26292 40402
rect 26236 40338 26292 40350
rect 26236 39620 26292 39630
rect 26236 39526 26292 39564
rect 26236 38724 26292 38734
rect 26236 38630 26292 38668
rect 26236 38052 26292 38062
rect 26236 37958 26292 37996
rect 26236 37156 26292 37166
rect 26236 37062 26292 37100
rect 26012 35970 26068 35980
rect 26348 36482 26404 36494
rect 26348 36430 26350 36482
rect 26402 36430 26404 36482
rect 26012 35588 26068 35598
rect 26236 35588 26292 35598
rect 26012 28196 26068 35532
rect 26124 35586 26292 35588
rect 26124 35534 26238 35586
rect 26290 35534 26292 35586
rect 26124 35532 26292 35534
rect 26124 32452 26180 35532
rect 26236 35522 26292 35532
rect 26236 34916 26292 34926
rect 26236 34822 26292 34860
rect 26348 34692 26404 36430
rect 26460 36372 26516 45054
rect 26460 36306 26516 36316
rect 26572 41412 26628 41422
rect 26348 34626 26404 34636
rect 26348 34356 26404 34366
rect 26236 34020 26292 34030
rect 26236 33926 26292 33964
rect 26236 33346 26292 33358
rect 26236 33294 26238 33346
rect 26290 33294 26292 33346
rect 26236 32676 26292 33294
rect 26236 32610 26292 32620
rect 26348 32562 26404 34300
rect 26348 32510 26350 32562
rect 26402 32510 26404 32562
rect 26348 32498 26404 32510
rect 26124 32386 26180 32396
rect 26460 31778 26516 31790
rect 26460 31726 26462 31778
rect 26514 31726 26516 31778
rect 26348 30994 26404 31006
rect 26348 30942 26350 30994
rect 26402 30942 26404 30994
rect 26236 30212 26292 30222
rect 26124 30210 26292 30212
rect 26124 30158 26238 30210
rect 26290 30158 26292 30210
rect 26124 30156 26292 30158
rect 26124 28532 26180 30156
rect 26236 30146 26292 30156
rect 26236 29540 26292 29550
rect 26236 29426 26292 29484
rect 26236 29374 26238 29426
rect 26290 29374 26292 29426
rect 26236 29362 26292 29374
rect 26236 28644 26292 28654
rect 26236 28550 26292 28588
rect 26124 28466 26180 28476
rect 26012 28140 26180 28196
rect 25900 27748 25956 27758
rect 25900 22932 25956 27692
rect 26124 27636 26180 28140
rect 26236 27748 26292 27758
rect 26236 27654 26292 27692
rect 25900 22866 25956 22876
rect 26012 27580 26180 27636
rect 25564 22316 25844 22372
rect 25564 20916 25620 22316
rect 25676 22146 25732 22158
rect 25676 22094 25678 22146
rect 25730 22094 25732 22146
rect 25676 21812 25732 22094
rect 25676 21746 25732 21756
rect 25788 21700 25844 21710
rect 25788 21606 25844 21644
rect 25564 20850 25620 20860
rect 25900 20804 25956 20814
rect 25452 15810 25508 15820
rect 25676 20802 25956 20804
rect 25676 20750 25902 20802
rect 25954 20750 25956 20802
rect 25676 20748 25956 20750
rect 25340 15092 25620 15148
rect 24668 12850 24948 12852
rect 24668 12798 24670 12850
rect 24722 12798 24948 12850
rect 24668 12796 24948 12798
rect 25004 13468 25172 13524
rect 25228 14642 25284 14654
rect 25228 14590 25230 14642
rect 25282 14590 25284 14642
rect 24668 12786 24724 12796
rect 25004 11956 25060 13468
rect 25228 13412 25284 14590
rect 25340 13748 25396 13758
rect 25340 13654 25396 13692
rect 25004 11890 25060 11900
rect 25116 13356 25284 13412
rect 25116 12962 25172 13356
rect 25116 12910 25118 12962
rect 25170 12910 25172 12962
rect 24464 11788 24728 11798
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24464 11722 24728 11732
rect 25116 10500 25172 12910
rect 25116 10434 25172 10444
rect 24464 10220 24728 10230
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24464 10154 24728 10164
rect 25564 9268 25620 15092
rect 25564 9202 25620 9212
rect 24464 8652 24728 8662
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24464 8586 24728 8596
rect 24464 7084 24728 7094
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 24464 7018 24728 7028
rect 24464 5516 24728 5526
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24464 5450 24728 5460
rect 24464 3948 24728 3958
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24464 3882 24728 3892
rect 24464 2380 24728 2390
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24464 2314 24728 2324
rect 24332 2034 24388 2044
rect 24892 1652 24948 1662
rect 23804 1596 24068 1606
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 23804 1530 24068 1540
rect 22540 1362 22596 1372
rect 24464 812 24728 822
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24464 746 24728 756
rect 23548 532 23604 542
rect 23548 112 23604 476
rect 24892 112 24948 1596
rect 25676 980 25732 20748
rect 25900 20738 25956 20748
rect 25788 20580 25844 20590
rect 25788 6468 25844 20524
rect 25900 19460 25956 19470
rect 25900 19366 25956 19404
rect 25788 6402 25844 6412
rect 26012 5908 26068 27580
rect 26348 27524 26404 30942
rect 26124 27468 26404 27524
rect 26124 7700 26180 27468
rect 26460 27412 26516 31726
rect 26348 27356 26516 27412
rect 26236 27076 26292 27086
rect 26236 26982 26292 27020
rect 26236 26178 26292 26190
rect 26236 26126 26238 26178
rect 26290 26126 26292 26178
rect 26236 25732 26292 26126
rect 26236 25666 26292 25676
rect 26236 25508 26292 25518
rect 26236 25414 26292 25452
rect 26236 24610 26292 24622
rect 26236 24558 26238 24610
rect 26290 24558 26292 24610
rect 26236 24500 26292 24558
rect 26236 24434 26292 24444
rect 26236 23938 26292 23950
rect 26236 23886 26238 23938
rect 26290 23886 26292 23938
rect 26236 23716 26292 23886
rect 26236 23650 26292 23660
rect 26236 23044 26292 23054
rect 26236 22950 26292 22988
rect 26236 22596 26292 22606
rect 26236 22482 26292 22540
rect 26236 22430 26238 22482
rect 26290 22430 26292 22482
rect 26236 22418 26292 22430
rect 26236 21476 26292 21486
rect 26236 21382 26292 21420
rect 26348 20580 26404 27356
rect 26572 26908 26628 41356
rect 26460 26852 26628 26908
rect 26460 20914 26516 26852
rect 26460 20862 26462 20914
rect 26514 20862 26516 20914
rect 26460 20850 26516 20862
rect 26348 20514 26404 20524
rect 26460 19348 26516 19358
rect 26460 19254 26516 19292
rect 26348 14306 26404 14318
rect 26348 14254 26350 14306
rect 26402 14254 26404 14306
rect 26348 11508 26404 14254
rect 26348 11442 26404 11452
rect 26124 7634 26180 7644
rect 26012 5842 26068 5852
rect 26572 6692 26628 6702
rect 26572 2098 26628 6636
rect 26684 5796 26740 49756
rect 27132 48244 27188 49870
rect 27244 49140 27300 50318
rect 27244 49074 27300 49084
rect 27132 48178 27188 48188
rect 27244 48802 27300 48814
rect 27244 48750 27246 48802
rect 27298 48750 27300 48802
rect 27020 48130 27076 48142
rect 27020 48078 27022 48130
rect 27074 48078 27076 48130
rect 27020 46900 27076 48078
rect 27244 47796 27300 48750
rect 27244 47730 27300 47740
rect 27020 46834 27076 46844
rect 27244 47234 27300 47246
rect 27244 47182 27246 47234
rect 27298 47182 27300 47234
rect 27132 46786 27188 46798
rect 27132 46734 27134 46786
rect 27186 46734 27188 46786
rect 27132 45108 27188 46734
rect 27244 46004 27300 47182
rect 27244 45938 27300 45948
rect 27132 45042 27188 45052
rect 27244 45666 27300 45678
rect 27244 45614 27246 45666
rect 27298 45614 27300 45666
rect 27020 44994 27076 45006
rect 27020 44942 27022 44994
rect 27074 44942 27076 44994
rect 27020 43764 27076 44942
rect 27244 44660 27300 45614
rect 27244 44594 27300 44604
rect 27020 43698 27076 43708
rect 27244 44098 27300 44110
rect 27244 44046 27246 44098
rect 27298 44046 27300 44098
rect 27132 43650 27188 43662
rect 27132 43598 27134 43650
rect 27186 43598 27188 43650
rect 27132 41972 27188 43598
rect 27244 42868 27300 44046
rect 27244 42802 27300 42812
rect 27132 41906 27188 41916
rect 27244 42530 27300 42542
rect 27244 42478 27246 42530
rect 27298 42478 27300 42530
rect 27020 41858 27076 41870
rect 27020 41806 27022 41858
rect 27074 41806 27076 41858
rect 27020 40628 27076 41806
rect 27244 41524 27300 42478
rect 27244 41458 27300 41468
rect 27020 40562 27076 40572
rect 27244 40962 27300 40974
rect 27244 40910 27246 40962
rect 27298 40910 27300 40962
rect 27132 40514 27188 40526
rect 27132 40462 27134 40514
rect 27186 40462 27188 40514
rect 27132 38836 27188 40462
rect 27244 39732 27300 40910
rect 27244 39666 27300 39676
rect 27132 38770 27188 38780
rect 27244 39394 27300 39406
rect 27244 39342 27246 39394
rect 27298 39342 27300 39394
rect 27020 38722 27076 38734
rect 27020 38670 27022 38722
rect 27074 38670 27076 38722
rect 27020 37492 27076 38670
rect 27244 38388 27300 39342
rect 27244 38322 27300 38332
rect 27020 37426 27076 37436
rect 27244 37826 27300 37838
rect 27244 37774 27246 37826
rect 27298 37774 27300 37826
rect 27132 37378 27188 37390
rect 27132 37326 27134 37378
rect 27186 37326 27188 37378
rect 27132 35700 27188 37326
rect 27244 36596 27300 37774
rect 27244 36530 27300 36540
rect 27132 35634 27188 35644
rect 27244 36258 27300 36270
rect 27244 36206 27246 36258
rect 27298 36206 27300 36258
rect 27020 35586 27076 35598
rect 27020 35534 27022 35586
rect 27074 35534 27076 35586
rect 27020 34356 27076 35534
rect 27244 35252 27300 36206
rect 27244 35186 27300 35196
rect 27020 34290 27076 34300
rect 27244 34690 27300 34702
rect 27244 34638 27246 34690
rect 27298 34638 27300 34690
rect 27132 34242 27188 34254
rect 27132 34190 27134 34242
rect 27186 34190 27188 34242
rect 27132 32564 27188 34190
rect 27244 33460 27300 34638
rect 27244 33394 27300 33404
rect 27132 32498 27188 32508
rect 27244 33122 27300 33134
rect 27244 33070 27246 33122
rect 27298 33070 27300 33122
rect 27020 32450 27076 32462
rect 27020 32398 27022 32450
rect 27074 32398 27076 32450
rect 27020 31220 27076 32398
rect 27244 32116 27300 33070
rect 27244 32050 27300 32060
rect 28364 32340 28420 32350
rect 27020 31154 27076 31164
rect 27244 31554 27300 31566
rect 27244 31502 27246 31554
rect 27298 31502 27300 31554
rect 27020 30882 27076 30894
rect 27020 30830 27022 30882
rect 27074 30830 27076 30882
rect 27020 29876 27076 30830
rect 27244 30324 27300 31502
rect 27244 30258 27300 30268
rect 27020 29810 27076 29820
rect 27132 30098 27188 30110
rect 27132 30046 27134 30098
rect 27186 30046 27188 30098
rect 27132 29428 27188 30046
rect 28140 29652 28196 29662
rect 27132 29362 27188 29372
rect 27244 29538 27300 29550
rect 27244 29486 27246 29538
rect 27298 29486 27300 29538
rect 27244 28980 27300 29486
rect 27244 28914 27300 28924
rect 27244 28532 27300 28542
rect 27244 28438 27300 28476
rect 27244 28084 27300 28094
rect 27244 27990 27300 28028
rect 27020 27636 27076 27646
rect 27020 27186 27076 27580
rect 27020 27134 27022 27186
rect 27074 27134 27076 27186
rect 27020 27122 27076 27134
rect 27244 26740 27300 26750
rect 27244 26514 27300 26684
rect 27244 26462 27246 26514
rect 27298 26462 27300 26514
rect 27244 26450 27300 26462
rect 27244 25844 27300 25854
rect 27132 25396 27188 25406
rect 27132 24834 27188 25340
rect 27244 25394 27300 25788
rect 27244 25342 27246 25394
rect 27298 25342 27300 25394
rect 27244 25330 27300 25342
rect 27132 24782 27134 24834
rect 27186 24782 27188 24834
rect 27132 24770 27188 24782
rect 27244 24500 27300 24510
rect 27244 23826 27300 24444
rect 27244 23774 27246 23826
rect 27298 23774 27300 23826
rect 27244 23762 27300 23774
rect 27244 23604 27300 23614
rect 27244 23378 27300 23548
rect 27244 23326 27246 23378
rect 27298 23326 27300 23378
rect 27244 23314 27300 23326
rect 27244 22708 27300 22718
rect 27132 22260 27188 22270
rect 27132 21698 27188 22204
rect 27244 22258 27300 22652
rect 27244 22206 27246 22258
rect 27298 22206 27300 22258
rect 27244 22194 27300 22206
rect 27132 21646 27134 21698
rect 27186 21646 27188 21698
rect 27132 21634 27188 21646
rect 27356 20916 27412 20926
rect 27356 20822 27412 20860
rect 28140 20916 28196 29596
rect 28140 20850 28196 20860
rect 26908 20802 26964 20814
rect 26908 20750 26910 20802
rect 26962 20750 26964 20802
rect 26908 20188 26964 20750
rect 26908 20132 27076 20188
rect 26684 5730 26740 5740
rect 27020 4452 27076 20132
rect 28364 20020 28420 32284
rect 28364 19954 28420 19964
rect 27020 4386 27076 4396
rect 27580 5124 27636 5134
rect 26572 2046 26574 2098
rect 26626 2046 26628 2098
rect 26572 2034 26628 2046
rect 27468 2212 27524 2222
rect 27468 2098 27524 2156
rect 27468 2046 27470 2098
rect 27522 2046 27524 2098
rect 27468 2034 27524 2046
rect 25676 914 25732 924
rect 26012 1986 26068 1998
rect 26012 1934 26014 1986
rect 26066 1934 26068 1986
rect 26012 644 26068 1934
rect 26908 1986 26964 1998
rect 26908 1934 26910 1986
rect 26962 1934 26964 1986
rect 26012 578 26068 588
rect 26236 1764 26292 1774
rect 26236 112 26292 1708
rect 26908 420 26964 1934
rect 26908 354 26964 364
rect 27580 112 27636 5068
rect 5292 28 5908 84
rect 6048 0 6160 112
rect 7392 0 7504 112
rect 8736 0 8848 112
rect 10080 0 10192 112
rect 11424 0 11536 112
rect 12768 0 12880 112
rect 14112 0 14224 112
rect 15456 0 15568 112
rect 16800 0 16912 112
rect 18144 0 18256 112
rect 19488 0 19600 112
rect 20832 0 20944 112
rect 22176 0 22288 112
rect 23520 0 23632 112
rect 24864 0 24976 112
rect 26208 0 26320 112
rect 27552 0 27664 112
<< via2 >>
rect 3804 56474 3860 56476
rect 3804 56422 3806 56474
rect 3806 56422 3858 56474
rect 3858 56422 3860 56474
rect 3804 56420 3860 56422
rect 3908 56474 3964 56476
rect 3908 56422 3910 56474
rect 3910 56422 3962 56474
rect 3962 56422 3964 56474
rect 3908 56420 3964 56422
rect 4012 56474 4068 56476
rect 4012 56422 4014 56474
rect 4014 56422 4066 56474
rect 4066 56422 4068 56474
rect 4012 56420 4068 56422
rect 4464 55690 4520 55692
rect 4464 55638 4466 55690
rect 4466 55638 4518 55690
rect 4518 55638 4520 55690
rect 4464 55636 4520 55638
rect 4568 55690 4624 55692
rect 4568 55638 4570 55690
rect 4570 55638 4622 55690
rect 4622 55638 4624 55690
rect 4568 55636 4624 55638
rect 4672 55690 4728 55692
rect 4672 55638 4674 55690
rect 4674 55638 4726 55690
rect 4726 55638 4728 55690
rect 4672 55636 4728 55638
rect 1372 53788 1428 53844
rect 2044 53340 2100 53396
rect 1484 52444 1540 52500
rect 588 41692 644 41748
rect 252 39564 308 39620
rect 588 38556 644 38612
rect 364 37324 420 37380
rect 364 23212 420 23268
rect 476 29372 532 29428
rect 924 40908 980 40964
rect 812 38108 868 38164
rect 812 28476 868 28532
rect 588 21756 644 21812
rect 700 18396 756 18452
rect 700 9212 756 9268
rect 812 12124 868 12180
rect 1596 45164 1652 45220
rect 1932 42588 1988 42644
rect 1820 40796 1876 40852
rect 1708 39004 1764 39060
rect 1148 38556 1204 38612
rect 1148 38220 1204 38276
rect 1372 35756 1428 35812
rect 1148 34018 1204 34020
rect 1148 33966 1150 34018
rect 1150 33966 1202 34018
rect 1202 33966 1204 34018
rect 1148 33964 1204 33966
rect 1036 32620 1092 32676
rect 1484 32620 1540 32676
rect 1484 31724 1540 31780
rect 1932 40124 1988 40180
rect 1820 37660 1876 37716
rect 1708 36876 1764 36932
rect 1708 36428 1764 36484
rect 1708 36204 1764 36260
rect 1708 31948 1764 32004
rect 1596 30268 1652 30324
rect 1708 31778 1764 31780
rect 1708 31726 1710 31778
rect 1710 31726 1762 31778
rect 1762 31726 1764 31778
rect 1708 31724 1764 31726
rect 1036 29932 1092 29988
rect 1148 29538 1204 29540
rect 1148 29486 1150 29538
rect 1150 29486 1202 29538
rect 1202 29486 1204 29538
rect 1148 29484 1204 29486
rect 1484 29426 1540 29428
rect 1484 29374 1486 29426
rect 1486 29374 1538 29426
rect 1538 29374 1540 29426
rect 1484 29372 1540 29374
rect 1484 28476 1540 28532
rect 1484 27244 1540 27300
rect 1596 28364 1652 28420
rect 1596 27916 1652 27972
rect 1260 27074 1316 27076
rect 1260 27022 1262 27074
rect 1262 27022 1314 27074
rect 1314 27022 1316 27074
rect 1260 27020 1316 27022
rect 1932 37100 1988 37156
rect 2828 55244 2884 55300
rect 2156 39900 2212 39956
rect 2604 40124 2660 40180
rect 2604 38780 2660 38836
rect 2716 39788 2772 39844
rect 2156 37436 2212 37492
rect 1932 34860 1988 34916
rect 2492 36876 2548 36932
rect 2940 48860 2996 48916
rect 2940 40236 2996 40292
rect 3052 46732 3108 46788
rect 3164 40460 3220 40516
rect 2828 37436 2884 37492
rect 2716 36988 2772 37044
rect 2828 36540 2884 36596
rect 2716 35810 2772 35812
rect 2716 35758 2718 35810
rect 2718 35758 2770 35810
rect 2770 35758 2772 35810
rect 2716 35756 2772 35758
rect 2604 35196 2660 35252
rect 2268 34412 2324 34468
rect 2380 34748 2436 34804
rect 1820 28700 1876 28756
rect 1932 33852 1988 33908
rect 1708 27298 1764 27300
rect 1708 27246 1710 27298
rect 1710 27246 1762 27298
rect 1762 27246 1764 27298
rect 1708 27244 1764 27246
rect 1260 26460 1316 26516
rect 1372 23772 1428 23828
rect 1148 23266 1204 23268
rect 1148 23214 1150 23266
rect 1150 23214 1202 23266
rect 1202 23214 1204 23266
rect 1148 23212 1204 23214
rect 1260 23100 1316 23156
rect 1148 19292 1204 19348
rect 1036 17500 1092 17556
rect 1820 27020 1876 27076
rect 2492 34300 2548 34356
rect 2380 33964 2436 34020
rect 2492 34076 2548 34132
rect 2268 32284 2324 32340
rect 2044 28364 2100 28420
rect 2380 31948 2436 32004
rect 2828 34802 2884 34804
rect 2828 34750 2830 34802
rect 2830 34750 2882 34802
rect 2882 34750 2884 34802
rect 2828 34748 2884 34750
rect 2716 34076 2772 34132
rect 6188 55970 6244 55972
rect 6188 55918 6190 55970
rect 6190 55918 6242 55970
rect 6242 55918 6244 55970
rect 6188 55916 6244 55918
rect 6300 55298 6356 55300
rect 6300 55246 6302 55298
rect 6302 55246 6354 55298
rect 6354 55246 6356 55298
rect 6300 55244 6356 55246
rect 6076 55132 6132 55188
rect 6860 55186 6916 55188
rect 6860 55134 6862 55186
rect 6862 55134 6914 55186
rect 6914 55134 6916 55186
rect 6860 55132 6916 55134
rect 3804 54906 3860 54908
rect 3804 54854 3806 54906
rect 3806 54854 3858 54906
rect 3858 54854 3860 54906
rect 3804 54852 3860 54854
rect 3908 54906 3964 54908
rect 3908 54854 3910 54906
rect 3910 54854 3962 54906
rect 3962 54854 3964 54906
rect 3908 54852 3964 54854
rect 4012 54906 4068 54908
rect 4012 54854 4014 54906
rect 4014 54854 4066 54906
rect 4066 54854 4068 54906
rect 4012 54852 4068 54854
rect 5964 54236 6020 54292
rect 4464 54122 4520 54124
rect 4464 54070 4466 54122
rect 4466 54070 4518 54122
rect 4518 54070 4520 54122
rect 4464 54068 4520 54070
rect 4568 54122 4624 54124
rect 4568 54070 4570 54122
rect 4570 54070 4622 54122
rect 4622 54070 4624 54122
rect 4568 54068 4624 54070
rect 4672 54122 4728 54124
rect 4672 54070 4674 54122
rect 4674 54070 4726 54122
rect 4726 54070 4728 54122
rect 4672 54068 4728 54070
rect 3804 53338 3860 53340
rect 3804 53286 3806 53338
rect 3806 53286 3858 53338
rect 3858 53286 3860 53338
rect 3804 53284 3860 53286
rect 3908 53338 3964 53340
rect 3908 53286 3910 53338
rect 3910 53286 3962 53338
rect 3962 53286 3964 53338
rect 3908 53284 3964 53286
rect 4012 53338 4068 53340
rect 4012 53286 4014 53338
rect 4014 53286 4066 53338
rect 4066 53286 4068 53338
rect 4012 53284 4068 53286
rect 4464 52554 4520 52556
rect 4464 52502 4466 52554
rect 4466 52502 4518 52554
rect 4518 52502 4520 52554
rect 4464 52500 4520 52502
rect 4568 52554 4624 52556
rect 4568 52502 4570 52554
rect 4570 52502 4622 52554
rect 4622 52502 4624 52554
rect 4568 52500 4624 52502
rect 4672 52554 4728 52556
rect 4672 52502 4674 52554
rect 4674 52502 4726 52554
rect 4726 52502 4728 52554
rect 4672 52500 4728 52502
rect 3804 51770 3860 51772
rect 3804 51718 3806 51770
rect 3806 51718 3858 51770
rect 3858 51718 3860 51770
rect 3804 51716 3860 51718
rect 3908 51770 3964 51772
rect 3908 51718 3910 51770
rect 3910 51718 3962 51770
rect 3962 51718 3964 51770
rect 3908 51716 3964 51718
rect 4012 51770 4068 51772
rect 4012 51718 4014 51770
rect 4014 51718 4066 51770
rect 4066 51718 4068 51770
rect 4012 51716 4068 51718
rect 4464 50986 4520 50988
rect 4464 50934 4466 50986
rect 4466 50934 4518 50986
rect 4518 50934 4520 50986
rect 4464 50932 4520 50934
rect 4568 50986 4624 50988
rect 4568 50934 4570 50986
rect 4570 50934 4622 50986
rect 4622 50934 4624 50986
rect 4568 50932 4624 50934
rect 4672 50986 4728 50988
rect 4672 50934 4674 50986
rect 4674 50934 4726 50986
rect 4726 50934 4728 50986
rect 4672 50932 4728 50934
rect 6748 54012 6804 54068
rect 3804 50202 3860 50204
rect 3804 50150 3806 50202
rect 3806 50150 3858 50202
rect 3858 50150 3860 50202
rect 3804 50148 3860 50150
rect 3908 50202 3964 50204
rect 3908 50150 3910 50202
rect 3910 50150 3962 50202
rect 3962 50150 3964 50202
rect 3908 50148 3964 50150
rect 4012 50202 4068 50204
rect 4012 50150 4014 50202
rect 4014 50150 4066 50202
rect 4066 50150 4068 50202
rect 4012 50148 4068 50150
rect 5292 49756 5348 49812
rect 4464 49418 4520 49420
rect 4464 49366 4466 49418
rect 4466 49366 4518 49418
rect 4518 49366 4520 49418
rect 4464 49364 4520 49366
rect 4568 49418 4624 49420
rect 4568 49366 4570 49418
rect 4570 49366 4622 49418
rect 4622 49366 4624 49418
rect 4568 49364 4624 49366
rect 4672 49418 4728 49420
rect 4672 49366 4674 49418
rect 4674 49366 4726 49418
rect 4726 49366 4728 49418
rect 4672 49364 4728 49366
rect 3804 48634 3860 48636
rect 3804 48582 3806 48634
rect 3806 48582 3858 48634
rect 3858 48582 3860 48634
rect 3804 48580 3860 48582
rect 3908 48634 3964 48636
rect 3908 48582 3910 48634
rect 3910 48582 3962 48634
rect 3962 48582 3964 48634
rect 3908 48580 3964 48582
rect 4012 48634 4068 48636
rect 4012 48582 4014 48634
rect 4014 48582 4066 48634
rect 4066 48582 4068 48634
rect 4012 48580 4068 48582
rect 4464 47850 4520 47852
rect 4464 47798 4466 47850
rect 4466 47798 4518 47850
rect 4518 47798 4520 47850
rect 4464 47796 4520 47798
rect 4568 47850 4624 47852
rect 4568 47798 4570 47850
rect 4570 47798 4622 47850
rect 4622 47798 4624 47850
rect 4568 47796 4624 47798
rect 4672 47850 4728 47852
rect 4672 47798 4674 47850
rect 4674 47798 4726 47850
rect 4726 47798 4728 47850
rect 4672 47796 4728 47798
rect 3804 47066 3860 47068
rect 3804 47014 3806 47066
rect 3806 47014 3858 47066
rect 3858 47014 3860 47066
rect 3804 47012 3860 47014
rect 3908 47066 3964 47068
rect 3908 47014 3910 47066
rect 3910 47014 3962 47066
rect 3962 47014 3964 47066
rect 3908 47012 3964 47014
rect 4012 47066 4068 47068
rect 4012 47014 4014 47066
rect 4014 47014 4066 47066
rect 4066 47014 4068 47066
rect 4012 47012 4068 47014
rect 4464 46282 4520 46284
rect 4464 46230 4466 46282
rect 4466 46230 4518 46282
rect 4518 46230 4520 46282
rect 4464 46228 4520 46230
rect 4568 46282 4624 46284
rect 4568 46230 4570 46282
rect 4570 46230 4622 46282
rect 4622 46230 4624 46282
rect 4568 46228 4624 46230
rect 4672 46282 4728 46284
rect 4672 46230 4674 46282
rect 4674 46230 4726 46282
rect 4726 46230 4728 46282
rect 4672 46228 4728 46230
rect 3804 45498 3860 45500
rect 3804 45446 3806 45498
rect 3806 45446 3858 45498
rect 3858 45446 3860 45498
rect 3804 45444 3860 45446
rect 3908 45498 3964 45500
rect 3908 45446 3910 45498
rect 3910 45446 3962 45498
rect 3962 45446 3964 45498
rect 3908 45444 3964 45446
rect 4012 45498 4068 45500
rect 4012 45446 4014 45498
rect 4014 45446 4066 45498
rect 4066 45446 4068 45498
rect 4012 45444 4068 45446
rect 4464 44714 4520 44716
rect 4464 44662 4466 44714
rect 4466 44662 4518 44714
rect 4518 44662 4520 44714
rect 4464 44660 4520 44662
rect 4568 44714 4624 44716
rect 4568 44662 4570 44714
rect 4570 44662 4622 44714
rect 4622 44662 4624 44714
rect 4568 44660 4624 44662
rect 4672 44714 4728 44716
rect 4672 44662 4674 44714
rect 4674 44662 4726 44714
rect 4726 44662 4728 44714
rect 4672 44660 4728 44662
rect 3804 43930 3860 43932
rect 3804 43878 3806 43930
rect 3806 43878 3858 43930
rect 3858 43878 3860 43930
rect 3804 43876 3860 43878
rect 3908 43930 3964 43932
rect 3908 43878 3910 43930
rect 3910 43878 3962 43930
rect 3962 43878 3964 43930
rect 3908 43876 3964 43878
rect 4012 43930 4068 43932
rect 4012 43878 4014 43930
rect 4014 43878 4066 43930
rect 4066 43878 4068 43930
rect 4012 43876 4068 43878
rect 4464 43146 4520 43148
rect 4464 43094 4466 43146
rect 4466 43094 4518 43146
rect 4518 43094 4520 43146
rect 4464 43092 4520 43094
rect 4568 43146 4624 43148
rect 4568 43094 4570 43146
rect 4570 43094 4622 43146
rect 4622 43094 4624 43146
rect 4568 43092 4624 43094
rect 4672 43146 4728 43148
rect 4672 43094 4674 43146
rect 4674 43094 4726 43146
rect 4726 43094 4728 43146
rect 4672 43092 4728 43094
rect 3804 42362 3860 42364
rect 3804 42310 3806 42362
rect 3806 42310 3858 42362
rect 3858 42310 3860 42362
rect 3804 42308 3860 42310
rect 3908 42362 3964 42364
rect 3908 42310 3910 42362
rect 3910 42310 3962 42362
rect 3962 42310 3964 42362
rect 3908 42308 3964 42310
rect 4012 42362 4068 42364
rect 4012 42310 4014 42362
rect 4014 42310 4066 42362
rect 4066 42310 4068 42362
rect 4012 42308 4068 42310
rect 4464 41578 4520 41580
rect 4464 41526 4466 41578
rect 4466 41526 4518 41578
rect 4518 41526 4520 41578
rect 4464 41524 4520 41526
rect 4568 41578 4624 41580
rect 4568 41526 4570 41578
rect 4570 41526 4622 41578
rect 4622 41526 4624 41578
rect 4568 41524 4624 41526
rect 4672 41578 4728 41580
rect 4672 41526 4674 41578
rect 4674 41526 4726 41578
rect 4726 41526 4728 41578
rect 4672 41524 4728 41526
rect 3804 40794 3860 40796
rect 3804 40742 3806 40794
rect 3806 40742 3858 40794
rect 3858 40742 3860 40794
rect 3804 40740 3860 40742
rect 3908 40794 3964 40796
rect 3908 40742 3910 40794
rect 3910 40742 3962 40794
rect 3962 40742 3964 40794
rect 3908 40740 3964 40742
rect 4012 40794 4068 40796
rect 4012 40742 4014 40794
rect 4014 40742 4066 40794
rect 4066 40742 4068 40794
rect 4012 40740 4068 40742
rect 5180 40124 5236 40180
rect 4464 40010 4520 40012
rect 4464 39958 4466 40010
rect 4466 39958 4518 40010
rect 4518 39958 4520 40010
rect 4464 39956 4520 39958
rect 4568 40010 4624 40012
rect 4568 39958 4570 40010
rect 4570 39958 4622 40010
rect 4622 39958 4624 40010
rect 4568 39956 4624 39958
rect 4672 40010 4728 40012
rect 4672 39958 4674 40010
rect 4674 39958 4726 40010
rect 4726 39958 4728 40010
rect 4672 39956 4728 39958
rect 3500 39676 3556 39732
rect 4172 39788 4228 39844
rect 3836 39618 3892 39620
rect 3836 39566 3838 39618
rect 3838 39566 3890 39618
rect 3890 39566 3892 39618
rect 3836 39564 3892 39566
rect 4172 39564 4228 39620
rect 3804 39226 3860 39228
rect 3804 39174 3806 39226
rect 3806 39174 3858 39226
rect 3858 39174 3860 39226
rect 3804 39172 3860 39174
rect 3908 39226 3964 39228
rect 3908 39174 3910 39226
rect 3910 39174 3962 39226
rect 3962 39174 3964 39226
rect 3908 39172 3964 39174
rect 4012 39226 4068 39228
rect 4012 39174 4014 39226
rect 4014 39174 4066 39226
rect 4066 39174 4068 39226
rect 4012 39172 4068 39174
rect 3500 38892 3556 38948
rect 5068 38892 5124 38948
rect 3804 37658 3860 37660
rect 3804 37606 3806 37658
rect 3806 37606 3858 37658
rect 3858 37606 3860 37658
rect 3804 37604 3860 37606
rect 3908 37658 3964 37660
rect 3908 37606 3910 37658
rect 3910 37606 3962 37658
rect 3962 37606 3964 37658
rect 3908 37604 3964 37606
rect 4012 37658 4068 37660
rect 4012 37606 4014 37658
rect 4014 37606 4066 37658
rect 4066 37606 4068 37658
rect 4012 37604 4068 37606
rect 3164 37324 3220 37380
rect 3164 36540 3220 36596
rect 3388 36988 3444 37044
rect 3052 34412 3108 34468
rect 2716 30828 2772 30884
rect 3612 36540 3668 36596
rect 4464 38442 4520 38444
rect 4464 38390 4466 38442
rect 4466 38390 4518 38442
rect 4518 38390 4520 38442
rect 4464 38388 4520 38390
rect 4568 38442 4624 38444
rect 4568 38390 4570 38442
rect 4570 38390 4622 38442
rect 4622 38390 4624 38442
rect 4568 38388 4624 38390
rect 4672 38442 4728 38444
rect 4672 38390 4674 38442
rect 4674 38390 4726 38442
rect 4726 38390 4728 38442
rect 4672 38388 4728 38390
rect 4844 38274 4900 38276
rect 4844 38222 4846 38274
rect 4846 38222 4898 38274
rect 4898 38222 4900 38274
rect 4844 38220 4900 38222
rect 4396 37938 4452 37940
rect 4396 37886 4398 37938
rect 4398 37886 4450 37938
rect 4450 37886 4452 37938
rect 4396 37884 4452 37886
rect 4844 37324 4900 37380
rect 4172 36594 4228 36596
rect 4172 36542 4174 36594
rect 4174 36542 4226 36594
rect 4226 36542 4228 36594
rect 4172 36540 4228 36542
rect 3804 36090 3860 36092
rect 3804 36038 3806 36090
rect 3806 36038 3858 36090
rect 3858 36038 3860 36090
rect 3804 36036 3860 36038
rect 3908 36090 3964 36092
rect 3908 36038 3910 36090
rect 3910 36038 3962 36090
rect 3962 36038 3964 36090
rect 3908 36036 3964 36038
rect 4012 36090 4068 36092
rect 4012 36038 4014 36090
rect 4014 36038 4066 36090
rect 4066 36038 4068 36090
rect 4012 36036 4068 36038
rect 3388 33740 3444 33796
rect 3836 35196 3892 35252
rect 3164 33516 3220 33572
rect 3276 33180 3332 33236
rect 3724 34972 3780 35028
rect 4844 36988 4900 37044
rect 4464 36874 4520 36876
rect 4464 36822 4466 36874
rect 4466 36822 4518 36874
rect 4518 36822 4520 36874
rect 4464 36820 4520 36822
rect 4568 36874 4624 36876
rect 4568 36822 4570 36874
rect 4570 36822 4622 36874
rect 4622 36822 4624 36874
rect 4568 36820 4624 36822
rect 4672 36874 4728 36876
rect 4672 36822 4674 36874
rect 4674 36822 4726 36874
rect 4726 36822 4728 36874
rect 4672 36820 4728 36822
rect 4396 35810 4452 35812
rect 4396 35758 4398 35810
rect 4398 35758 4450 35810
rect 4450 35758 4452 35810
rect 4396 35756 4452 35758
rect 4464 35306 4520 35308
rect 4464 35254 4466 35306
rect 4466 35254 4518 35306
rect 4518 35254 4520 35306
rect 4464 35252 4520 35254
rect 4568 35306 4624 35308
rect 4568 35254 4570 35306
rect 4570 35254 4622 35306
rect 4622 35254 4624 35306
rect 4568 35252 4624 35254
rect 4672 35306 4728 35308
rect 4672 35254 4674 35306
rect 4674 35254 4726 35306
rect 4726 35254 4728 35306
rect 4672 35252 4728 35254
rect 3804 34522 3860 34524
rect 3804 34470 3806 34522
rect 3806 34470 3858 34522
rect 3858 34470 3860 34522
rect 3804 34468 3860 34470
rect 3908 34522 3964 34524
rect 3908 34470 3910 34522
rect 3910 34470 3962 34522
rect 3962 34470 3964 34522
rect 3908 34468 3964 34470
rect 4012 34522 4068 34524
rect 4012 34470 4014 34522
rect 4014 34470 4066 34522
rect 4066 34470 4068 34522
rect 4012 34468 4068 34470
rect 4172 34130 4228 34132
rect 4172 34078 4174 34130
rect 4174 34078 4226 34130
rect 4226 34078 4228 34130
rect 4172 34076 4228 34078
rect 3612 33740 3668 33796
rect 2604 30492 2660 30548
rect 3164 30770 3220 30772
rect 3164 30718 3166 30770
rect 3166 30718 3218 30770
rect 3218 30718 3220 30770
rect 3164 30716 3220 30718
rect 2940 30380 2996 30436
rect 2828 30268 2884 30324
rect 2492 30044 2548 30100
rect 2268 29484 2324 29540
rect 2716 29538 2772 29540
rect 2716 29486 2718 29538
rect 2718 29486 2770 29538
rect 2770 29486 2772 29538
rect 2716 29484 2772 29486
rect 2492 28812 2548 28868
rect 2380 28754 2436 28756
rect 2380 28702 2382 28754
rect 2382 28702 2434 28754
rect 2434 28702 2436 28754
rect 2380 28700 2436 28702
rect 2156 26124 2212 26180
rect 3052 30492 3108 30548
rect 3276 30156 3332 30212
rect 2940 29036 2996 29092
rect 2380 26178 2436 26180
rect 2380 26126 2382 26178
rect 2382 26126 2434 26178
rect 2434 26126 2436 26178
rect 2380 26124 2436 26126
rect 2044 25228 2100 25284
rect 1484 23212 1540 23268
rect 1596 23996 1652 24052
rect 1708 23212 1764 23268
rect 1484 21980 1540 22036
rect 1372 18620 1428 18676
rect 1260 17388 1316 17444
rect 1372 14476 1428 14532
rect 1372 13916 1428 13972
rect 1260 9266 1316 9268
rect 1260 9214 1262 9266
rect 1262 9214 1314 9266
rect 1314 9214 1316 9266
rect 1260 9212 1316 9214
rect 1596 21756 1652 21812
rect 1820 20914 1876 20916
rect 1820 20862 1822 20914
rect 1822 20862 1874 20914
rect 1874 20862 1876 20914
rect 1820 20860 1876 20862
rect 1932 20412 1988 20468
rect 1708 18172 1764 18228
rect 1708 17388 1764 17444
rect 1820 17052 1876 17108
rect 1596 16770 1652 16772
rect 1596 16718 1598 16770
rect 1598 16718 1650 16770
rect 1650 16718 1652 16770
rect 1596 16716 1652 16718
rect 1820 16322 1876 16324
rect 1820 16270 1822 16322
rect 1822 16270 1874 16322
rect 1874 16270 1876 16322
rect 1820 16268 1876 16270
rect 1708 15314 1764 15316
rect 1708 15262 1710 15314
rect 1710 15262 1762 15314
rect 1762 15262 1764 15314
rect 1708 15260 1764 15262
rect 1596 14530 1652 14532
rect 1596 14478 1598 14530
rect 1598 14478 1650 14530
rect 1650 14478 1652 14530
rect 1596 14476 1652 14478
rect 2940 28812 2996 28868
rect 3724 33180 3780 33236
rect 3804 32954 3860 32956
rect 3804 32902 3806 32954
rect 3806 32902 3858 32954
rect 3858 32902 3860 32954
rect 3804 32900 3860 32902
rect 3908 32954 3964 32956
rect 3908 32902 3910 32954
rect 3910 32902 3962 32954
rect 3962 32902 3964 32954
rect 3908 32900 3964 32902
rect 4012 32954 4068 32956
rect 4012 32902 4014 32954
rect 4014 32902 4066 32954
rect 4066 32902 4068 32954
rect 4012 32900 4068 32902
rect 3836 32450 3892 32452
rect 3836 32398 3838 32450
rect 3838 32398 3890 32450
rect 3890 32398 3892 32450
rect 3836 32396 3892 32398
rect 3804 31386 3860 31388
rect 3804 31334 3806 31386
rect 3806 31334 3858 31386
rect 3858 31334 3860 31386
rect 3804 31332 3860 31334
rect 3908 31386 3964 31388
rect 3908 31334 3910 31386
rect 3910 31334 3962 31386
rect 3962 31334 3964 31386
rect 3908 31332 3964 31334
rect 4012 31386 4068 31388
rect 4012 31334 4014 31386
rect 4014 31334 4066 31386
rect 4066 31334 4068 31386
rect 4012 31332 4068 31334
rect 3500 29372 3556 29428
rect 3388 29260 3444 29316
rect 3276 29036 3332 29092
rect 3164 28476 3220 28532
rect 3276 26962 3332 26964
rect 3276 26910 3278 26962
rect 3278 26910 3330 26962
rect 3330 26910 3332 26962
rect 3276 26908 3332 26910
rect 3164 26236 3220 26292
rect 2716 25228 2772 25284
rect 2604 24556 2660 24612
rect 2380 23826 2436 23828
rect 2380 23774 2382 23826
rect 2382 23774 2434 23826
rect 2434 23774 2436 23826
rect 2380 23772 2436 23774
rect 2268 23266 2324 23268
rect 2268 23214 2270 23266
rect 2270 23214 2322 23266
rect 2322 23214 2324 23266
rect 2268 23212 2324 23214
rect 2156 19794 2212 19796
rect 2156 19742 2158 19794
rect 2158 19742 2210 19794
rect 2210 19742 2212 19794
rect 2156 19740 2212 19742
rect 2268 19346 2324 19348
rect 2268 19294 2270 19346
rect 2270 19294 2322 19346
rect 2322 19294 2324 19346
rect 2268 19292 2324 19294
rect 2156 18450 2212 18452
rect 2156 18398 2158 18450
rect 2158 18398 2210 18450
rect 2210 18398 2212 18450
rect 2156 18396 2212 18398
rect 2044 16716 2100 16772
rect 2156 16940 2212 16996
rect 2268 16716 2324 16772
rect 1596 11618 1652 11620
rect 1596 11566 1598 11618
rect 1598 11566 1650 11618
rect 1650 11566 1652 11618
rect 1596 11564 1652 11566
rect 1596 8540 1652 8596
rect 924 6860 980 6916
rect 1484 6748 1540 6804
rect 2156 15484 2212 15540
rect 1820 11676 1876 11732
rect 1708 7644 1764 7700
rect 1820 8372 1876 8428
rect 1484 4060 1540 4116
rect 1260 3164 1316 3220
rect 2268 13132 2324 13188
rect 2156 12124 2212 12180
rect 2044 11676 2100 11732
rect 2268 11564 2324 11620
rect 2268 11340 2324 11396
rect 2044 10610 2100 10612
rect 2044 10558 2046 10610
rect 2046 10558 2098 10610
rect 2098 10558 2100 10610
rect 2044 10556 2100 10558
rect 2044 8988 2100 9044
rect 2716 23100 2772 23156
rect 2604 22316 2660 22372
rect 2828 22204 2884 22260
rect 2492 19740 2548 19796
rect 2940 21644 2996 21700
rect 2828 20412 2884 20468
rect 2940 20188 2996 20244
rect 2716 17500 2772 17556
rect 4464 33738 4520 33740
rect 4464 33686 4466 33738
rect 4466 33686 4518 33738
rect 4518 33686 4520 33738
rect 4464 33684 4520 33686
rect 4568 33738 4624 33740
rect 4568 33686 4570 33738
rect 4570 33686 4622 33738
rect 4622 33686 4624 33738
rect 4568 33684 4624 33686
rect 4672 33738 4728 33740
rect 4672 33686 4674 33738
rect 4674 33686 4726 33738
rect 4726 33686 4728 33738
rect 4672 33684 4728 33686
rect 4844 33628 4900 33684
rect 4508 33516 4564 33572
rect 4508 32508 4564 32564
rect 4464 32170 4520 32172
rect 4464 32118 4466 32170
rect 4466 32118 4518 32170
rect 4518 32118 4520 32170
rect 4464 32116 4520 32118
rect 4568 32170 4624 32172
rect 4568 32118 4570 32170
rect 4570 32118 4622 32170
rect 4622 32118 4624 32170
rect 4568 32116 4624 32118
rect 4672 32170 4728 32172
rect 4672 32118 4674 32170
rect 4674 32118 4726 32170
rect 4726 32118 4728 32170
rect 4672 32116 4728 32118
rect 4284 31218 4340 31220
rect 4284 31166 4286 31218
rect 4286 31166 4338 31218
rect 4338 31166 4340 31218
rect 4284 31164 4340 31166
rect 5068 33964 5124 34020
rect 4956 33516 5012 33572
rect 5292 38668 5348 38724
rect 5404 42028 5460 42084
rect 6076 40124 6132 40180
rect 5852 38780 5908 38836
rect 5404 37884 5460 37940
rect 5628 37436 5684 37492
rect 5516 35196 5572 35252
rect 5292 33852 5348 33908
rect 5404 34636 5460 34692
rect 5404 34076 5460 34132
rect 5292 33516 5348 33572
rect 5516 33516 5572 33572
rect 4464 30602 4520 30604
rect 4464 30550 4466 30602
rect 4466 30550 4518 30602
rect 4518 30550 4520 30602
rect 4464 30548 4520 30550
rect 4568 30602 4624 30604
rect 4568 30550 4570 30602
rect 4570 30550 4622 30602
rect 4622 30550 4624 30602
rect 4568 30548 4624 30550
rect 4672 30602 4728 30604
rect 4672 30550 4674 30602
rect 4674 30550 4726 30602
rect 4726 30550 4728 30602
rect 4672 30548 4728 30550
rect 4172 30268 4228 30324
rect 4284 30210 4340 30212
rect 4284 30158 4286 30210
rect 4286 30158 4338 30210
rect 4338 30158 4340 30210
rect 4284 30156 4340 30158
rect 3804 29818 3860 29820
rect 3804 29766 3806 29818
rect 3806 29766 3858 29818
rect 3858 29766 3860 29818
rect 3804 29764 3860 29766
rect 3908 29818 3964 29820
rect 3908 29766 3910 29818
rect 3910 29766 3962 29818
rect 3962 29766 3964 29818
rect 3908 29764 3964 29766
rect 4012 29818 4068 29820
rect 4012 29766 4014 29818
rect 4014 29766 4066 29818
rect 4066 29766 4068 29818
rect 4012 29764 4068 29766
rect 4284 29650 4340 29652
rect 4284 29598 4286 29650
rect 4286 29598 4338 29650
rect 4338 29598 4340 29650
rect 4284 29596 4340 29598
rect 4060 28700 4116 28756
rect 4844 30156 4900 30212
rect 3804 28250 3860 28252
rect 3804 28198 3806 28250
rect 3806 28198 3858 28250
rect 3858 28198 3860 28250
rect 3804 28196 3860 28198
rect 3908 28250 3964 28252
rect 3908 28198 3910 28250
rect 3910 28198 3962 28250
rect 3962 28198 3964 28250
rect 3908 28196 3964 28198
rect 4012 28250 4068 28252
rect 4012 28198 4014 28250
rect 4014 28198 4066 28250
rect 4066 28198 4068 28250
rect 4012 28196 4068 28198
rect 4464 29034 4520 29036
rect 4464 28982 4466 29034
rect 4466 28982 4518 29034
rect 4518 28982 4520 29034
rect 4464 28980 4520 28982
rect 4568 29034 4624 29036
rect 4568 28982 4570 29034
rect 4570 28982 4622 29034
rect 4622 28982 4624 29034
rect 4568 28980 4624 28982
rect 4672 29034 4728 29036
rect 4672 28982 4674 29034
rect 4674 28982 4726 29034
rect 4726 28982 4728 29034
rect 4672 28980 4728 28982
rect 4508 28754 4564 28756
rect 4508 28702 4510 28754
rect 4510 28702 4562 28754
rect 4562 28702 4564 28754
rect 4508 28700 4564 28702
rect 3948 27020 4004 27076
rect 4060 27356 4116 27412
rect 4464 27466 4520 27468
rect 4464 27414 4466 27466
rect 4466 27414 4518 27466
rect 4518 27414 4520 27466
rect 4464 27412 4520 27414
rect 4568 27466 4624 27468
rect 4568 27414 4570 27466
rect 4570 27414 4622 27466
rect 4622 27414 4624 27466
rect 4568 27412 4624 27414
rect 4672 27466 4728 27468
rect 4672 27414 4674 27466
rect 4674 27414 4726 27466
rect 4726 27414 4728 27466
rect 4672 27412 4728 27414
rect 4284 27298 4340 27300
rect 4284 27246 4286 27298
rect 4286 27246 4338 27298
rect 4338 27246 4340 27298
rect 4284 27244 4340 27246
rect 3804 26682 3860 26684
rect 3804 26630 3806 26682
rect 3806 26630 3858 26682
rect 3858 26630 3860 26682
rect 3804 26628 3860 26630
rect 3908 26682 3964 26684
rect 3908 26630 3910 26682
rect 3910 26630 3962 26682
rect 3962 26630 3964 26682
rect 3908 26628 3964 26630
rect 4012 26682 4068 26684
rect 4012 26630 4014 26682
rect 4014 26630 4066 26682
rect 4066 26630 4068 26682
rect 4012 26628 4068 26630
rect 3612 25730 3668 25732
rect 3612 25678 3614 25730
rect 3614 25678 3666 25730
rect 3666 25678 3668 25730
rect 3612 25676 3668 25678
rect 3804 25114 3860 25116
rect 3804 25062 3806 25114
rect 3806 25062 3858 25114
rect 3858 25062 3860 25114
rect 3804 25060 3860 25062
rect 3908 25114 3964 25116
rect 3908 25062 3910 25114
rect 3910 25062 3962 25114
rect 3962 25062 3964 25114
rect 3908 25060 3964 25062
rect 4012 25114 4068 25116
rect 4012 25062 4014 25114
rect 4014 25062 4066 25114
rect 4066 25062 4068 25114
rect 4012 25060 4068 25062
rect 3388 24892 3444 24948
rect 3500 24834 3556 24836
rect 3500 24782 3502 24834
rect 3502 24782 3554 24834
rect 3554 24782 3556 24834
rect 3500 24780 3556 24782
rect 3500 24332 3556 24388
rect 3388 24050 3444 24052
rect 3388 23998 3390 24050
rect 3390 23998 3442 24050
rect 3442 23998 3444 24050
rect 3388 23996 3444 23998
rect 3276 23772 3332 23828
rect 3164 22204 3220 22260
rect 3164 21756 3220 21812
rect 4172 24780 4228 24836
rect 3804 23546 3860 23548
rect 3804 23494 3806 23546
rect 3806 23494 3858 23546
rect 3858 23494 3860 23546
rect 3804 23492 3860 23494
rect 3908 23546 3964 23548
rect 3908 23494 3910 23546
rect 3910 23494 3962 23546
rect 3962 23494 3964 23546
rect 3908 23492 3964 23494
rect 4012 23546 4068 23548
rect 4012 23494 4014 23546
rect 4014 23494 4066 23546
rect 4066 23494 4068 23546
rect 4012 23492 4068 23494
rect 4732 27074 4788 27076
rect 4732 27022 4734 27074
rect 4734 27022 4786 27074
rect 4786 27022 4788 27074
rect 4732 27020 4788 27022
rect 4396 26012 4452 26068
rect 4464 25898 4520 25900
rect 4464 25846 4466 25898
rect 4466 25846 4518 25898
rect 4518 25846 4520 25898
rect 4464 25844 4520 25846
rect 4568 25898 4624 25900
rect 4568 25846 4570 25898
rect 4570 25846 4622 25898
rect 4622 25846 4624 25898
rect 4568 25844 4624 25846
rect 4672 25898 4728 25900
rect 4672 25846 4674 25898
rect 4674 25846 4726 25898
rect 4726 25846 4728 25898
rect 4672 25844 4728 25846
rect 4732 24780 4788 24836
rect 4956 29596 5012 29652
rect 5068 29484 5124 29540
rect 5516 31500 5572 31556
rect 5404 31164 5460 31220
rect 5292 30828 5348 30884
rect 5628 30044 5684 30100
rect 5292 29372 5348 29428
rect 5628 29426 5684 29428
rect 5628 29374 5630 29426
rect 5630 29374 5682 29426
rect 5682 29374 5684 29426
rect 5628 29372 5684 29374
rect 5180 28364 5236 28420
rect 5516 27356 5572 27412
rect 4956 27244 5012 27300
rect 5292 27074 5348 27076
rect 5292 27022 5294 27074
rect 5294 27022 5346 27074
rect 5346 27022 5348 27074
rect 5292 27020 5348 27022
rect 5404 26908 5460 26964
rect 4956 25676 5012 25732
rect 5292 26012 5348 26068
rect 4464 24330 4520 24332
rect 4464 24278 4466 24330
rect 4466 24278 4518 24330
rect 4518 24278 4520 24330
rect 4464 24276 4520 24278
rect 4568 24330 4624 24332
rect 4568 24278 4570 24330
rect 4570 24278 4622 24330
rect 4622 24278 4624 24330
rect 4568 24276 4624 24278
rect 4672 24330 4728 24332
rect 4672 24278 4674 24330
rect 4674 24278 4726 24330
rect 4726 24278 4728 24330
rect 4672 24276 4728 24278
rect 4620 23938 4676 23940
rect 4620 23886 4622 23938
rect 4622 23886 4674 23938
rect 4674 23886 4676 23938
rect 4620 23884 4676 23886
rect 5068 23884 5124 23940
rect 4844 23548 4900 23604
rect 4464 22762 4520 22764
rect 4464 22710 4466 22762
rect 4466 22710 4518 22762
rect 4518 22710 4520 22762
rect 4464 22708 4520 22710
rect 4568 22762 4624 22764
rect 4568 22710 4570 22762
rect 4570 22710 4622 22762
rect 4622 22710 4624 22762
rect 4568 22708 4624 22710
rect 4672 22762 4728 22764
rect 4672 22710 4674 22762
rect 4674 22710 4726 22762
rect 4726 22710 4728 22762
rect 4672 22708 4728 22710
rect 3804 21978 3860 21980
rect 3804 21926 3806 21978
rect 3806 21926 3858 21978
rect 3858 21926 3860 21978
rect 3804 21924 3860 21926
rect 3908 21978 3964 21980
rect 3908 21926 3910 21978
rect 3910 21926 3962 21978
rect 3962 21926 3964 21978
rect 3908 21924 3964 21926
rect 4012 21978 4068 21980
rect 4012 21926 4014 21978
rect 4014 21926 4066 21978
rect 4066 21926 4068 21978
rect 4012 21924 4068 21926
rect 3612 21084 3668 21140
rect 4172 21756 4228 21812
rect 3164 20914 3220 20916
rect 3164 20862 3166 20914
rect 3166 20862 3218 20914
rect 3218 20862 3220 20914
rect 3164 20860 3220 20862
rect 3804 20410 3860 20412
rect 3804 20358 3806 20410
rect 3806 20358 3858 20410
rect 3858 20358 3860 20410
rect 3804 20356 3860 20358
rect 3908 20410 3964 20412
rect 3908 20358 3910 20410
rect 3910 20358 3962 20410
rect 3962 20358 3964 20410
rect 3908 20356 3964 20358
rect 4012 20410 4068 20412
rect 4012 20358 4014 20410
rect 4014 20358 4066 20410
rect 4066 20358 4068 20410
rect 4012 20356 4068 20358
rect 3052 19122 3108 19124
rect 3052 19070 3054 19122
rect 3054 19070 3106 19122
rect 3106 19070 3108 19122
rect 3052 19068 3108 19070
rect 2940 17612 2996 17668
rect 2716 16156 2772 16212
rect 2604 15202 2660 15204
rect 2604 15150 2606 15202
rect 2606 15150 2658 15202
rect 2658 15150 2660 15202
rect 2604 15148 2660 15150
rect 2492 12066 2548 12068
rect 2492 12014 2494 12066
rect 2494 12014 2546 12066
rect 2546 12014 2548 12066
rect 2492 12012 2548 12014
rect 2604 12124 2660 12180
rect 2380 8764 2436 8820
rect 2492 11788 2548 11844
rect 2716 11900 2772 11956
rect 2828 15708 2884 15764
rect 2492 9996 2548 10052
rect 2156 8372 2212 8428
rect 2604 10668 2660 10724
rect 2940 13020 2996 13076
rect 2604 8652 2660 8708
rect 2716 9436 2772 9492
rect 1932 4956 1988 5012
rect 2044 6860 2100 6916
rect 1820 2268 1876 2324
rect 476 1596 532 1652
rect 252 476 308 532
rect 700 588 756 644
rect 2268 7980 2324 8036
rect 2380 6860 2436 6916
rect 2268 6076 2324 6132
rect 3804 18842 3860 18844
rect 3804 18790 3806 18842
rect 3806 18790 3858 18842
rect 3858 18790 3860 18842
rect 3804 18788 3860 18790
rect 3908 18842 3964 18844
rect 3908 18790 3910 18842
rect 3910 18790 3962 18842
rect 3962 18790 3964 18842
rect 3908 18788 3964 18790
rect 4012 18842 4068 18844
rect 4012 18790 4014 18842
rect 4014 18790 4066 18842
rect 4066 18790 4068 18842
rect 4012 18788 4068 18790
rect 3500 18172 3556 18228
rect 3948 18396 4004 18452
rect 3724 17890 3780 17892
rect 3724 17838 3726 17890
rect 3726 17838 3778 17890
rect 3778 17838 3780 17890
rect 3724 17836 3780 17838
rect 3836 17724 3892 17780
rect 3164 15260 3220 15316
rect 3804 17274 3860 17276
rect 3804 17222 3806 17274
rect 3806 17222 3858 17274
rect 3858 17222 3860 17274
rect 3804 17220 3860 17222
rect 3908 17274 3964 17276
rect 3908 17222 3910 17274
rect 3910 17222 3962 17274
rect 3962 17222 3964 17274
rect 3908 17220 3964 17222
rect 4012 17274 4068 17276
rect 4012 17222 4014 17274
rect 4014 17222 4066 17274
rect 4066 17222 4068 17274
rect 4012 17220 4068 17222
rect 3388 16882 3444 16884
rect 3388 16830 3390 16882
rect 3390 16830 3442 16882
rect 3442 16830 3444 16882
rect 3388 16828 3444 16830
rect 3836 16828 3892 16884
rect 3612 16156 3668 16212
rect 4060 16210 4116 16212
rect 4060 16158 4062 16210
rect 4062 16158 4114 16210
rect 4114 16158 4116 16210
rect 4060 16156 4116 16158
rect 3388 15820 3444 15876
rect 3388 15148 3444 15204
rect 3804 15706 3860 15708
rect 3804 15654 3806 15706
rect 3806 15654 3858 15706
rect 3858 15654 3860 15706
rect 3804 15652 3860 15654
rect 3908 15706 3964 15708
rect 3908 15654 3910 15706
rect 3910 15654 3962 15706
rect 3962 15654 3964 15706
rect 3908 15652 3964 15654
rect 4012 15706 4068 15708
rect 4012 15654 4014 15706
rect 4014 15654 4066 15706
rect 4066 15654 4068 15706
rect 4012 15652 4068 15654
rect 4284 21362 4340 21364
rect 4284 21310 4286 21362
rect 4286 21310 4338 21362
rect 4338 21310 4340 21362
rect 4284 21308 4340 21310
rect 4464 21194 4520 21196
rect 4464 21142 4466 21194
rect 4466 21142 4518 21194
rect 4518 21142 4520 21194
rect 4464 21140 4520 21142
rect 4568 21194 4624 21196
rect 4568 21142 4570 21194
rect 4570 21142 4622 21194
rect 4622 21142 4624 21194
rect 4568 21140 4624 21142
rect 4672 21194 4728 21196
rect 4672 21142 4674 21194
rect 4674 21142 4726 21194
rect 4726 21142 4728 21194
rect 4672 21140 4728 21142
rect 4396 20802 4452 20804
rect 4396 20750 4398 20802
rect 4398 20750 4450 20802
rect 4450 20750 4452 20802
rect 4396 20748 4452 20750
rect 4464 19626 4520 19628
rect 4464 19574 4466 19626
rect 4466 19574 4518 19626
rect 4518 19574 4520 19626
rect 4464 19572 4520 19574
rect 4568 19626 4624 19628
rect 4568 19574 4570 19626
rect 4570 19574 4622 19626
rect 4622 19574 4624 19626
rect 4568 19572 4624 19574
rect 4672 19626 4728 19628
rect 4672 19574 4674 19626
rect 4674 19574 4726 19626
rect 4726 19574 4728 19626
rect 4672 19572 4728 19574
rect 4620 19234 4676 19236
rect 4620 19182 4622 19234
rect 4622 19182 4674 19234
rect 4674 19182 4676 19234
rect 4620 19180 4676 19182
rect 4844 18396 4900 18452
rect 4956 21644 5012 21700
rect 4464 18058 4520 18060
rect 4464 18006 4466 18058
rect 4466 18006 4518 18058
rect 4518 18006 4520 18058
rect 4464 18004 4520 18006
rect 4568 18058 4624 18060
rect 4568 18006 4570 18058
rect 4570 18006 4622 18058
rect 4622 18006 4624 18058
rect 4568 18004 4624 18006
rect 4672 18058 4728 18060
rect 4672 18006 4674 18058
rect 4674 18006 4726 18058
rect 4726 18006 4728 18058
rect 4672 18004 4728 18006
rect 5516 26178 5572 26180
rect 5516 26126 5518 26178
rect 5518 26126 5570 26178
rect 5570 26126 5572 26178
rect 5516 26124 5572 26126
rect 5516 25564 5572 25620
rect 5516 23938 5572 23940
rect 5516 23886 5518 23938
rect 5518 23886 5570 23938
rect 5570 23886 5572 23938
rect 5516 23884 5572 23886
rect 5292 23100 5348 23156
rect 5180 23042 5236 23044
rect 5180 22990 5182 23042
rect 5182 22990 5234 23042
rect 5234 22990 5236 23042
rect 5180 22988 5236 22990
rect 5628 23324 5684 23380
rect 5964 38274 6020 38276
rect 5964 38222 5966 38274
rect 5966 38222 6018 38274
rect 6018 38222 6020 38274
rect 5964 38220 6020 38222
rect 5964 36316 6020 36372
rect 5852 34636 5908 34692
rect 5852 32844 5908 32900
rect 5852 32674 5908 32676
rect 5852 32622 5854 32674
rect 5854 32622 5906 32674
rect 5906 32622 5908 32674
rect 5852 32620 5908 32622
rect 5852 31778 5908 31780
rect 5852 31726 5854 31778
rect 5854 31726 5906 31778
rect 5906 31726 5908 31778
rect 5852 31724 5908 31726
rect 5740 23100 5796 23156
rect 5852 31500 5908 31556
rect 5180 22092 5236 22148
rect 5516 22876 5572 22932
rect 5180 21420 5236 21476
rect 5404 21586 5460 21588
rect 5404 21534 5406 21586
rect 5406 21534 5458 21586
rect 5458 21534 5460 21586
rect 5404 21532 5460 21534
rect 5292 20972 5348 21028
rect 5068 18732 5124 18788
rect 5068 18562 5124 18564
rect 5068 18510 5070 18562
rect 5070 18510 5122 18562
rect 5122 18510 5124 18562
rect 5068 18508 5124 18510
rect 4284 17836 4340 17892
rect 4284 17666 4340 17668
rect 4284 17614 4286 17666
rect 4286 17614 4338 17666
rect 4338 17614 4340 17666
rect 4284 17612 4340 17614
rect 5628 22540 5684 22596
rect 5628 22370 5684 22372
rect 5628 22318 5630 22370
rect 5630 22318 5682 22370
rect 5682 22318 5684 22370
rect 5628 22316 5684 22318
rect 5628 22092 5684 22148
rect 5404 19234 5460 19236
rect 5404 19182 5406 19234
rect 5406 19182 5458 19234
rect 5458 19182 5460 19234
rect 5404 19180 5460 19182
rect 5404 18396 5460 18452
rect 5516 18732 5572 18788
rect 4732 17666 4788 17668
rect 4732 17614 4734 17666
rect 4734 17614 4786 17666
rect 4786 17614 4788 17666
rect 4732 17612 4788 17614
rect 5068 17554 5124 17556
rect 5068 17502 5070 17554
rect 5070 17502 5122 17554
rect 5122 17502 5124 17554
rect 5068 17500 5124 17502
rect 4956 16882 5012 16884
rect 4956 16830 4958 16882
rect 4958 16830 5010 16882
rect 5010 16830 5012 16882
rect 4956 16828 5012 16830
rect 4464 16490 4520 16492
rect 4464 16438 4466 16490
rect 4466 16438 4518 16490
rect 4518 16438 4520 16490
rect 4464 16436 4520 16438
rect 4568 16490 4624 16492
rect 4568 16438 4570 16490
rect 4570 16438 4622 16490
rect 4622 16438 4624 16490
rect 4568 16436 4624 16438
rect 4672 16490 4728 16492
rect 4672 16438 4674 16490
rect 4674 16438 4726 16490
rect 4726 16438 4728 16490
rect 4672 16436 4728 16438
rect 4284 15372 4340 15428
rect 3500 14252 3556 14308
rect 3388 13634 3444 13636
rect 3388 13582 3390 13634
rect 3390 13582 3442 13634
rect 3442 13582 3444 13634
rect 3388 13580 3444 13582
rect 3164 13074 3220 13076
rect 3164 13022 3166 13074
rect 3166 13022 3218 13074
rect 3218 13022 3220 13074
rect 3164 13020 3220 13022
rect 4284 15036 4340 15092
rect 4464 14922 4520 14924
rect 4464 14870 4466 14922
rect 4466 14870 4518 14922
rect 4518 14870 4520 14922
rect 4464 14868 4520 14870
rect 4568 14922 4624 14924
rect 4568 14870 4570 14922
rect 4570 14870 4622 14922
rect 4622 14870 4624 14922
rect 4568 14868 4624 14870
rect 4672 14922 4728 14924
rect 4672 14870 4674 14922
rect 4674 14870 4726 14922
rect 4726 14870 4728 14922
rect 4672 14868 4728 14870
rect 4172 14530 4228 14532
rect 4172 14478 4174 14530
rect 4174 14478 4226 14530
rect 4226 14478 4228 14530
rect 4172 14476 4228 14478
rect 3804 14138 3860 14140
rect 3804 14086 3806 14138
rect 3806 14086 3858 14138
rect 3858 14086 3860 14138
rect 3804 14084 3860 14086
rect 3908 14138 3964 14140
rect 3908 14086 3910 14138
rect 3910 14086 3962 14138
rect 3962 14086 3964 14138
rect 3908 14084 3964 14086
rect 4012 14138 4068 14140
rect 4012 14086 4014 14138
rect 4014 14086 4066 14138
rect 4066 14086 4068 14138
rect 4012 14084 4068 14086
rect 3724 13916 3780 13972
rect 3948 13916 4004 13972
rect 4732 14306 4788 14308
rect 4732 14254 4734 14306
rect 4734 14254 4786 14306
rect 4786 14254 4788 14306
rect 4732 14252 4788 14254
rect 4396 13916 4452 13972
rect 4464 13354 4520 13356
rect 4464 13302 4466 13354
rect 4466 13302 4518 13354
rect 4518 13302 4520 13354
rect 4464 13300 4520 13302
rect 4568 13354 4624 13356
rect 4568 13302 4570 13354
rect 4570 13302 4622 13354
rect 4622 13302 4624 13354
rect 4568 13300 4624 13302
rect 4672 13354 4728 13356
rect 4672 13302 4674 13354
rect 4674 13302 4726 13354
rect 4726 13302 4728 13354
rect 4672 13300 4728 13302
rect 4620 13132 4676 13188
rect 4956 13634 5012 13636
rect 4956 13582 4958 13634
rect 4958 13582 5010 13634
rect 5010 13582 5012 13634
rect 4956 13580 5012 13582
rect 4956 13132 5012 13188
rect 3804 12570 3860 12572
rect 3804 12518 3806 12570
rect 3806 12518 3858 12570
rect 3858 12518 3860 12570
rect 3804 12516 3860 12518
rect 3908 12570 3964 12572
rect 3908 12518 3910 12570
rect 3910 12518 3962 12570
rect 3962 12518 3964 12570
rect 3908 12516 3964 12518
rect 4012 12570 4068 12572
rect 4012 12518 4014 12570
rect 4014 12518 4066 12570
rect 4066 12518 4068 12570
rect 4012 12516 4068 12518
rect 3724 12236 3780 12292
rect 3276 11676 3332 11732
rect 3052 11228 3108 11284
rect 4172 11900 4228 11956
rect 3276 11228 3332 11284
rect 3612 11452 3668 11508
rect 3164 10332 3220 10388
rect 3276 11004 3332 11060
rect 3804 11002 3860 11004
rect 3804 10950 3806 11002
rect 3806 10950 3858 11002
rect 3858 10950 3860 11002
rect 3804 10948 3860 10950
rect 3908 11002 3964 11004
rect 3908 10950 3910 11002
rect 3910 10950 3962 11002
rect 3962 10950 3964 11002
rect 3908 10948 3964 10950
rect 4012 11002 4068 11004
rect 4012 10950 4014 11002
rect 4014 10950 4066 11002
rect 4066 10950 4068 11002
rect 4012 10948 4068 10950
rect 3836 9660 3892 9716
rect 3804 9434 3860 9436
rect 3804 9382 3806 9434
rect 3806 9382 3858 9434
rect 3858 9382 3860 9434
rect 3804 9380 3860 9382
rect 3908 9434 3964 9436
rect 3908 9382 3910 9434
rect 3910 9382 3962 9434
rect 3962 9382 3964 9434
rect 3908 9380 3964 9382
rect 4012 9434 4068 9436
rect 4012 9382 4014 9434
rect 4014 9382 4066 9434
rect 4066 9382 4068 9434
rect 4012 9380 4068 9382
rect 4464 11786 4520 11788
rect 4464 11734 4466 11786
rect 4466 11734 4518 11786
rect 4518 11734 4520 11786
rect 4464 11732 4520 11734
rect 4568 11786 4624 11788
rect 4568 11734 4570 11786
rect 4570 11734 4622 11786
rect 4622 11734 4624 11786
rect 4568 11732 4624 11734
rect 4672 11786 4728 11788
rect 4672 11734 4674 11786
rect 4674 11734 4726 11786
rect 4726 11734 4728 11786
rect 4672 11732 4728 11734
rect 4284 11394 4340 11396
rect 4284 11342 4286 11394
rect 4286 11342 4338 11394
rect 4338 11342 4340 11394
rect 4284 11340 4340 11342
rect 4464 10218 4520 10220
rect 4464 10166 4466 10218
rect 4466 10166 4518 10218
rect 4518 10166 4520 10218
rect 4464 10164 4520 10166
rect 4568 10218 4624 10220
rect 4568 10166 4570 10218
rect 4570 10166 4622 10218
rect 4622 10166 4624 10218
rect 4568 10164 4624 10166
rect 4672 10218 4728 10220
rect 4672 10166 4674 10218
rect 4674 10166 4726 10218
rect 4726 10166 4728 10218
rect 4672 10164 4728 10166
rect 4956 12236 5012 12292
rect 5404 17388 5460 17444
rect 5292 16604 5348 16660
rect 5180 15426 5236 15428
rect 5180 15374 5182 15426
rect 5182 15374 5234 15426
rect 5234 15374 5236 15426
rect 5180 15372 5236 15374
rect 5068 11452 5124 11508
rect 5180 10780 5236 10836
rect 5516 16268 5572 16324
rect 5740 21980 5796 22036
rect 6188 33964 6244 34020
rect 5964 31164 6020 31220
rect 5964 30492 6020 30548
rect 5964 27580 6020 27636
rect 5852 20578 5908 20580
rect 5852 20526 5854 20578
rect 5854 20526 5906 20578
rect 5906 20526 5908 20578
rect 5852 20524 5908 20526
rect 6076 30268 6132 30324
rect 6524 38220 6580 38276
rect 6636 39452 6692 39508
rect 6636 38892 6692 38948
rect 6524 37378 6580 37380
rect 6524 37326 6526 37378
rect 6526 37326 6578 37378
rect 6578 37326 6580 37378
rect 6524 37324 6580 37326
rect 6412 36706 6468 36708
rect 6412 36654 6414 36706
rect 6414 36654 6466 36706
rect 6466 36654 6468 36706
rect 6412 36652 6468 36654
rect 6524 36428 6580 36484
rect 6636 33628 6692 33684
rect 6300 33516 6356 33572
rect 6524 31612 6580 31668
rect 6412 31500 6468 31556
rect 6300 31164 6356 31220
rect 6300 30268 6356 30324
rect 6524 30828 6580 30884
rect 6524 29820 6580 29876
rect 6188 23436 6244 23492
rect 6076 22764 6132 22820
rect 6076 22092 6132 22148
rect 6412 27074 6468 27076
rect 6412 27022 6414 27074
rect 6414 27022 6466 27074
rect 6466 27022 6468 27074
rect 6412 27020 6468 27022
rect 6636 29596 6692 29652
rect 6636 28588 6692 28644
rect 6860 50428 6916 50484
rect 6860 45164 6916 45220
rect 7644 47180 7700 47236
rect 7756 40796 7812 40852
rect 7308 39730 7364 39732
rect 7308 39678 7310 39730
rect 7310 39678 7362 39730
rect 7362 39678 7364 39730
rect 7308 39676 7364 39678
rect 6860 39004 6916 39060
rect 6860 38668 6916 38724
rect 6972 37660 7028 37716
rect 6860 36204 6916 36260
rect 7084 35196 7140 35252
rect 7084 35026 7140 35028
rect 7084 34974 7086 35026
rect 7086 34974 7138 35026
rect 7138 34974 7140 35026
rect 7084 34972 7140 34974
rect 6972 33404 7028 33460
rect 7084 31276 7140 31332
rect 7756 39116 7812 39172
rect 9212 55916 9268 55972
rect 8540 46060 8596 46116
rect 8316 42700 8372 42756
rect 7980 40124 8036 40180
rect 8316 39116 8372 39172
rect 7868 37772 7924 37828
rect 8204 38556 8260 38612
rect 7868 36482 7924 36484
rect 7868 36430 7870 36482
rect 7870 36430 7922 36482
rect 7922 36430 7924 36482
rect 7868 36428 7924 36430
rect 7868 36204 7924 36260
rect 7756 34972 7812 35028
rect 7868 33964 7924 34020
rect 7644 33458 7700 33460
rect 7644 33406 7646 33458
rect 7646 33406 7698 33458
rect 7698 33406 7700 33458
rect 7644 33404 7700 33406
rect 7532 32620 7588 32676
rect 7644 31948 7700 32004
rect 7420 31276 7476 31332
rect 7308 31164 7364 31220
rect 7420 30492 7476 30548
rect 6972 29820 7028 29876
rect 7308 30156 7364 30212
rect 7196 29650 7252 29652
rect 7196 29598 7198 29650
rect 7198 29598 7250 29650
rect 7250 29598 7252 29650
rect 7196 29596 7252 29598
rect 7084 29484 7140 29540
rect 7644 29820 7700 29876
rect 7532 29708 7588 29764
rect 7308 28642 7364 28644
rect 7308 28590 7310 28642
rect 7310 28590 7362 28642
rect 7362 28590 7364 28642
rect 7308 28588 7364 28590
rect 7420 28476 7476 28532
rect 7084 28028 7140 28084
rect 6748 26348 6804 26404
rect 6748 23884 6804 23940
rect 6412 23436 6468 23492
rect 6412 22764 6468 22820
rect 6188 20076 6244 20132
rect 5740 18956 5796 19012
rect 5964 18732 6020 18788
rect 6076 18620 6132 18676
rect 6188 18396 6244 18452
rect 5964 18060 6020 18116
rect 5852 17724 5908 17780
rect 6076 17778 6132 17780
rect 6076 17726 6078 17778
rect 6078 17726 6130 17778
rect 6130 17726 6132 17778
rect 6076 17724 6132 17726
rect 5852 17500 5908 17556
rect 5852 17164 5908 17220
rect 6188 16492 6244 16548
rect 5852 15820 5908 15876
rect 5740 15260 5796 15316
rect 5852 13468 5908 13524
rect 5740 12850 5796 12852
rect 5740 12798 5742 12850
rect 5742 12798 5794 12850
rect 5794 12798 5796 12850
rect 5740 12796 5796 12798
rect 5516 12124 5572 12180
rect 5516 11788 5572 11844
rect 5628 12012 5684 12068
rect 6188 14812 6244 14868
rect 5964 11788 6020 11844
rect 4464 8650 4520 8652
rect 4464 8598 4466 8650
rect 4466 8598 4518 8650
rect 4518 8598 4520 8650
rect 4464 8596 4520 8598
rect 4568 8650 4624 8652
rect 4568 8598 4570 8650
rect 4570 8598 4622 8650
rect 4622 8598 4624 8650
rect 4568 8596 4624 8598
rect 4672 8650 4728 8652
rect 4672 8598 4674 8650
rect 4674 8598 4726 8650
rect 4726 8598 4728 8650
rect 4672 8596 4728 8598
rect 3612 8204 3668 8260
rect 2828 5852 2884 5908
rect 3836 8092 3892 8148
rect 5068 8034 5124 8036
rect 5068 7982 5070 8034
rect 5070 7982 5122 8034
rect 5122 7982 5124 8034
rect 5068 7980 5124 7982
rect 3804 7866 3860 7868
rect 3804 7814 3806 7866
rect 3806 7814 3858 7866
rect 3858 7814 3860 7866
rect 3804 7812 3860 7814
rect 3908 7866 3964 7868
rect 3908 7814 3910 7866
rect 3910 7814 3962 7866
rect 3962 7814 3964 7866
rect 3908 7812 3964 7814
rect 4012 7866 4068 7868
rect 4012 7814 4014 7866
rect 4014 7814 4066 7866
rect 4066 7814 4068 7866
rect 4012 7812 4068 7814
rect 3836 7474 3892 7476
rect 3836 7422 3838 7474
rect 3838 7422 3890 7474
rect 3890 7422 3892 7474
rect 3836 7420 3892 7422
rect 4464 7082 4520 7084
rect 4464 7030 4466 7082
rect 4466 7030 4518 7082
rect 4518 7030 4520 7082
rect 4464 7028 4520 7030
rect 4568 7082 4624 7084
rect 4568 7030 4570 7082
rect 4570 7030 4622 7082
rect 4622 7030 4624 7082
rect 4568 7028 4624 7030
rect 4672 7082 4728 7084
rect 4672 7030 4674 7082
rect 4674 7030 4726 7082
rect 4726 7030 4728 7082
rect 4672 7028 4728 7030
rect 3052 6412 3108 6468
rect 3804 6298 3860 6300
rect 3804 6246 3806 6298
rect 3806 6246 3858 6298
rect 3858 6246 3860 6298
rect 3804 6244 3860 6246
rect 3908 6298 3964 6300
rect 3908 6246 3910 6298
rect 3910 6246 3962 6298
rect 3962 6246 3964 6298
rect 3908 6244 3964 6246
rect 4012 6298 4068 6300
rect 4012 6246 4014 6298
rect 4014 6246 4066 6298
rect 4066 6246 4068 6298
rect 4012 6244 4068 6246
rect 3164 6018 3220 6020
rect 3164 5966 3166 6018
rect 3166 5966 3218 6018
rect 3218 5966 3220 6018
rect 3164 5964 3220 5966
rect 4464 5514 4520 5516
rect 4464 5462 4466 5514
rect 4466 5462 4518 5514
rect 4518 5462 4520 5514
rect 4464 5460 4520 5462
rect 4568 5514 4624 5516
rect 4568 5462 4570 5514
rect 4570 5462 4622 5514
rect 4622 5462 4624 5514
rect 4568 5460 4624 5462
rect 4672 5514 4728 5516
rect 4672 5462 4674 5514
rect 4674 5462 4726 5514
rect 4726 5462 4728 5514
rect 4672 5460 4728 5462
rect 3612 5346 3668 5348
rect 3612 5294 3614 5346
rect 3614 5294 3666 5346
rect 3666 5294 3668 5346
rect 3612 5292 3668 5294
rect 3804 4730 3860 4732
rect 3804 4678 3806 4730
rect 3806 4678 3858 4730
rect 3858 4678 3860 4730
rect 3804 4676 3860 4678
rect 3908 4730 3964 4732
rect 3908 4678 3910 4730
rect 3910 4678 3962 4730
rect 3962 4678 3964 4730
rect 3908 4676 3964 4678
rect 4012 4730 4068 4732
rect 4012 4678 4014 4730
rect 4014 4678 4066 4730
rect 4066 4678 4068 4730
rect 4012 4676 4068 4678
rect 2268 4226 2324 4228
rect 2268 4174 2270 4226
rect 2270 4174 2322 4226
rect 2322 4174 2324 4226
rect 2268 4172 2324 4174
rect 4464 3946 4520 3948
rect 4464 3894 4466 3946
rect 4466 3894 4518 3946
rect 4518 3894 4520 3946
rect 4464 3892 4520 3894
rect 4568 3946 4624 3948
rect 4568 3894 4570 3946
rect 4570 3894 4622 3946
rect 4622 3894 4624 3946
rect 4568 3892 4624 3894
rect 4672 3946 4728 3948
rect 4672 3894 4674 3946
rect 4674 3894 4726 3946
rect 4726 3894 4728 3946
rect 4672 3892 4728 3894
rect 2268 3554 2324 3556
rect 2268 3502 2270 3554
rect 2270 3502 2322 3554
rect 2322 3502 2324 3554
rect 2268 3500 2324 3502
rect 3804 3162 3860 3164
rect 3804 3110 3806 3162
rect 3806 3110 3858 3162
rect 3858 3110 3860 3162
rect 3804 3108 3860 3110
rect 3908 3162 3964 3164
rect 3908 3110 3910 3162
rect 3910 3110 3962 3162
rect 3962 3110 3964 3162
rect 3908 3108 3964 3110
rect 4012 3162 4068 3164
rect 4012 3110 4014 3162
rect 4014 3110 4066 3162
rect 4066 3110 4068 3162
rect 4012 3108 4068 3110
rect 4464 2378 4520 2380
rect 4464 2326 4466 2378
rect 4466 2326 4518 2378
rect 4518 2326 4520 2378
rect 4464 2324 4520 2326
rect 4568 2378 4624 2380
rect 4568 2326 4570 2378
rect 4570 2326 4622 2378
rect 4622 2326 4624 2378
rect 4568 2324 4624 2326
rect 4672 2378 4728 2380
rect 4672 2326 4674 2378
rect 4674 2326 4726 2378
rect 4726 2326 4728 2378
rect 4672 2324 4728 2326
rect 3388 1596 3444 1652
rect 3804 1594 3860 1596
rect 3804 1542 3806 1594
rect 3806 1542 3858 1594
rect 3858 1542 3860 1594
rect 3804 1540 3860 1542
rect 3908 1594 3964 1596
rect 3908 1542 3910 1594
rect 3910 1542 3962 1594
rect 3962 1542 3964 1594
rect 3908 1540 3964 1542
rect 4012 1594 4068 1596
rect 4012 1542 4014 1594
rect 4014 1542 4066 1594
rect 4066 1542 4068 1594
rect 4012 1540 4068 1542
rect 4464 810 4520 812
rect 4464 758 4466 810
rect 4466 758 4518 810
rect 4518 758 4520 810
rect 4464 756 4520 758
rect 4568 810 4624 812
rect 4568 758 4570 810
rect 4570 758 4622 810
rect 4622 758 4624 810
rect 4568 756 4624 758
rect 4672 810 4728 812
rect 4672 758 4674 810
rect 4674 758 4726 810
rect 4726 758 4728 810
rect 4672 756 4728 758
rect 4732 476 4788 532
rect 5404 10050 5460 10052
rect 5404 9998 5406 10050
rect 5406 9998 5458 10050
rect 5458 9998 5460 10050
rect 5404 9996 5460 9998
rect 6748 21196 6804 21252
rect 6524 20748 6580 20804
rect 6524 20524 6580 20580
rect 6748 19628 6804 19684
rect 6524 18338 6580 18340
rect 6524 18286 6526 18338
rect 6526 18286 6578 18338
rect 6578 18286 6580 18338
rect 6524 18284 6580 18286
rect 6524 17836 6580 17892
rect 6412 17388 6468 17444
rect 6412 16716 6468 16772
rect 7084 25730 7140 25732
rect 7084 25678 7086 25730
rect 7086 25678 7138 25730
rect 7138 25678 7140 25730
rect 7084 25676 7140 25678
rect 6972 24610 7028 24612
rect 6972 24558 6974 24610
rect 6974 24558 7026 24610
rect 7026 24558 7028 24610
rect 6972 24556 7028 24558
rect 6972 24220 7028 24276
rect 7196 24108 7252 24164
rect 7084 23660 7140 23716
rect 6972 23266 7028 23268
rect 6972 23214 6974 23266
rect 6974 23214 7026 23266
rect 7026 23214 7028 23266
rect 6972 23212 7028 23214
rect 6972 21644 7028 21700
rect 7196 23436 7252 23492
rect 7084 21196 7140 21252
rect 6972 19628 7028 19684
rect 7532 28364 7588 28420
rect 7420 27804 7476 27860
rect 7420 27132 7476 27188
rect 7420 26348 7476 26404
rect 7420 26012 7476 26068
rect 8204 34690 8260 34692
rect 8204 34638 8206 34690
rect 8206 34638 8258 34690
rect 8258 34638 8260 34690
rect 8204 34636 8260 34638
rect 8092 34076 8148 34132
rect 8204 33964 8260 34020
rect 7980 33404 8036 33460
rect 7756 28028 7812 28084
rect 7868 31052 7924 31108
rect 7868 30044 7924 30100
rect 7980 27804 8036 27860
rect 8092 33234 8148 33236
rect 8092 33182 8094 33234
rect 8094 33182 8146 33234
rect 8146 33182 8148 33234
rect 8092 33180 8148 33182
rect 8092 32172 8148 32228
rect 7868 27132 7924 27188
rect 8316 29932 8372 29988
rect 8428 34860 8484 34916
rect 8204 28252 8260 28308
rect 8316 29596 8372 29652
rect 8204 27970 8260 27972
rect 8204 27918 8206 27970
rect 8206 27918 8258 27970
rect 8258 27918 8260 27970
rect 8204 27916 8260 27918
rect 8092 27132 8148 27188
rect 7980 26066 8036 26068
rect 7980 26014 7982 26066
rect 7982 26014 8034 26066
rect 8034 26014 8036 26066
rect 7980 26012 8036 26014
rect 7644 24892 7700 24948
rect 7980 24610 8036 24612
rect 7980 24558 7982 24610
rect 7982 24558 8034 24610
rect 8034 24558 8036 24610
rect 7980 24556 8036 24558
rect 7756 23714 7812 23716
rect 7756 23662 7758 23714
rect 7758 23662 7810 23714
rect 7810 23662 7812 23714
rect 7756 23660 7812 23662
rect 8764 45276 8820 45332
rect 9212 41132 9268 41188
rect 9884 41692 9940 41748
rect 9772 41020 9828 41076
rect 9100 40236 9156 40292
rect 8876 39004 8932 39060
rect 8652 37266 8708 37268
rect 8652 37214 8654 37266
rect 8654 37214 8706 37266
rect 8706 37214 8708 37266
rect 8652 37212 8708 37214
rect 8652 33404 8708 33460
rect 8652 32844 8708 32900
rect 8540 30044 8596 30100
rect 8540 29538 8596 29540
rect 8540 29486 8542 29538
rect 8542 29486 8594 29538
rect 8594 29486 8596 29538
rect 8540 29484 8596 29486
rect 8204 23884 8260 23940
rect 7532 21980 7588 22036
rect 7196 20636 7252 20692
rect 7308 21308 7364 21364
rect 7756 22930 7812 22932
rect 7756 22878 7758 22930
rect 7758 22878 7810 22930
rect 7810 22878 7812 22930
rect 7756 22876 7812 22878
rect 7308 19234 7364 19236
rect 7308 19182 7310 19234
rect 7310 19182 7362 19234
rect 7362 19182 7364 19234
rect 7308 19180 7364 19182
rect 7420 19068 7476 19124
rect 8092 22876 8148 22932
rect 7980 20076 8036 20132
rect 7868 20018 7924 20020
rect 7868 19966 7870 20018
rect 7870 19966 7922 20018
rect 7922 19966 7924 20018
rect 7868 19964 7924 19966
rect 7980 19906 8036 19908
rect 7980 19854 7982 19906
rect 7982 19854 8034 19906
rect 8034 19854 8036 19906
rect 7980 19852 8036 19854
rect 8652 25676 8708 25732
rect 8540 21474 8596 21476
rect 8540 21422 8542 21474
rect 8542 21422 8594 21474
rect 8594 21422 8596 21474
rect 8540 21420 8596 21422
rect 8316 21084 8372 21140
rect 8204 19516 8260 19572
rect 7868 19180 7924 19236
rect 6636 16716 6692 16772
rect 6636 16492 6692 16548
rect 6636 15986 6692 15988
rect 6636 15934 6638 15986
rect 6638 15934 6690 15986
rect 6690 15934 6692 15986
rect 6636 15932 6692 15934
rect 6412 15596 6468 15652
rect 6412 14700 6468 14756
rect 6748 15314 6804 15316
rect 6748 15262 6750 15314
rect 6750 15262 6802 15314
rect 6802 15262 6804 15314
rect 6748 15260 6804 15262
rect 7308 17948 7364 18004
rect 7308 17666 7364 17668
rect 7308 17614 7310 17666
rect 7310 17614 7362 17666
rect 7362 17614 7364 17666
rect 7308 17612 7364 17614
rect 7532 17388 7588 17444
rect 7532 16940 7588 16996
rect 7756 16940 7812 16996
rect 7084 16322 7140 16324
rect 7084 16270 7086 16322
rect 7086 16270 7138 16322
rect 7138 16270 7140 16322
rect 7084 16268 7140 16270
rect 7532 15820 7588 15876
rect 7084 15314 7140 15316
rect 7084 15262 7086 15314
rect 7086 15262 7138 15314
rect 7138 15262 7140 15314
rect 7084 15260 7140 15262
rect 6636 13468 6692 13524
rect 6300 11788 6356 11844
rect 6524 11676 6580 11732
rect 7084 14924 7140 14980
rect 6860 14642 6916 14644
rect 6860 14590 6862 14642
rect 6862 14590 6914 14642
rect 6914 14590 6916 14642
rect 6860 14588 6916 14590
rect 6972 13746 7028 13748
rect 6972 13694 6974 13746
rect 6974 13694 7026 13746
rect 7026 13694 7028 13746
rect 6972 13692 7028 13694
rect 6972 12348 7028 12404
rect 7756 15148 7812 15204
rect 8428 20636 8484 20692
rect 7980 18284 8036 18340
rect 8204 17666 8260 17668
rect 8204 17614 8206 17666
rect 8206 17614 8258 17666
rect 8258 17614 8260 17666
rect 8204 17612 8260 17614
rect 8204 16828 8260 16884
rect 8092 15484 8148 15540
rect 8204 15932 8260 15988
rect 9212 39228 9268 39284
rect 9324 39676 9380 39732
rect 9100 34860 9156 34916
rect 9100 34636 9156 34692
rect 8876 33740 8932 33796
rect 8876 33346 8932 33348
rect 8876 33294 8878 33346
rect 8878 33294 8930 33346
rect 8930 33294 8932 33346
rect 8876 33292 8932 33294
rect 9660 37212 9716 37268
rect 9548 36764 9604 36820
rect 9436 35308 9492 35364
rect 15484 56252 15540 56308
rect 16492 56306 16548 56308
rect 16492 56254 16494 56306
rect 16494 56254 16546 56306
rect 16546 56254 16548 56306
rect 16492 56252 16548 56254
rect 11452 55132 11508 55188
rect 14028 55692 14084 55748
rect 11900 55186 11956 55188
rect 11900 55134 11902 55186
rect 11902 55134 11954 55186
rect 11954 55134 11956 55186
rect 11900 55132 11956 55134
rect 11564 54460 11620 54516
rect 10220 53788 10276 53844
rect 9996 41244 10052 41300
rect 10108 40236 10164 40292
rect 9884 39228 9940 39284
rect 9884 38780 9940 38836
rect 9324 34412 9380 34468
rect 9548 34412 9604 34468
rect 9436 33404 9492 33460
rect 9324 32620 9380 32676
rect 8876 30940 8932 30996
rect 9100 30828 9156 30884
rect 8876 30210 8932 30212
rect 8876 30158 8878 30210
rect 8878 30158 8930 30210
rect 8930 30158 8932 30210
rect 8876 30156 8932 30158
rect 8988 28924 9044 28980
rect 10108 39116 10164 39172
rect 10892 52556 10948 52612
rect 10780 50652 10836 50708
rect 10444 39452 10500 39508
rect 10332 37324 10388 37380
rect 10444 37996 10500 38052
rect 10220 34130 10276 34132
rect 10220 34078 10222 34130
rect 10222 34078 10274 34130
rect 10274 34078 10276 34130
rect 10220 34076 10276 34078
rect 10668 37660 10724 37716
rect 9660 30604 9716 30660
rect 9436 30210 9492 30212
rect 9436 30158 9438 30210
rect 9438 30158 9490 30210
rect 9490 30158 9492 30210
rect 9436 30156 9492 30158
rect 9548 28530 9604 28532
rect 9548 28478 9550 28530
rect 9550 28478 9602 28530
rect 9602 28478 9604 28530
rect 9548 28476 9604 28478
rect 9436 27468 9492 27524
rect 9772 29708 9828 29764
rect 9324 26908 9380 26964
rect 9436 27244 9492 27300
rect 9100 25506 9156 25508
rect 9100 25454 9102 25506
rect 9102 25454 9154 25506
rect 9154 25454 9156 25506
rect 9100 25452 9156 25454
rect 9212 24780 9268 24836
rect 8988 23996 9044 24052
rect 8988 23772 9044 23828
rect 8876 23436 8932 23492
rect 8764 20076 8820 20132
rect 8876 19852 8932 19908
rect 8764 18338 8820 18340
rect 8764 18286 8766 18338
rect 8766 18286 8818 18338
rect 8818 18286 8820 18338
rect 8764 18284 8820 18286
rect 8316 15484 8372 15540
rect 7644 14700 7700 14756
rect 7868 14588 7924 14644
rect 7308 14306 7364 14308
rect 7308 14254 7310 14306
rect 7310 14254 7362 14306
rect 7362 14254 7364 14306
rect 7308 14252 7364 14254
rect 7308 13804 7364 13860
rect 6748 11900 6804 11956
rect 7196 12908 7252 12964
rect 6636 11394 6692 11396
rect 6636 11342 6638 11394
rect 6638 11342 6690 11394
rect 6690 11342 6692 11394
rect 6636 11340 6692 11342
rect 6748 11228 6804 11284
rect 6524 10556 6580 10612
rect 6188 10220 6244 10276
rect 6524 9938 6580 9940
rect 6524 9886 6526 9938
rect 6526 9886 6578 9938
rect 6578 9886 6580 9938
rect 6524 9884 6580 9886
rect 6412 9154 6468 9156
rect 6412 9102 6414 9154
rect 6414 9102 6466 9154
rect 6466 9102 6468 9154
rect 6412 9100 6468 9102
rect 6300 8370 6356 8372
rect 6300 8318 6302 8370
rect 6302 8318 6354 8370
rect 6354 8318 6356 8370
rect 6300 8316 6356 8318
rect 6748 10498 6804 10500
rect 6748 10446 6750 10498
rect 6750 10446 6802 10498
rect 6802 10446 6804 10498
rect 6748 10444 6804 10446
rect 6748 9996 6804 10052
rect 6748 8876 6804 8932
rect 6748 8316 6804 8372
rect 6076 6748 6132 6804
rect 7420 13522 7476 13524
rect 7420 13470 7422 13522
rect 7422 13470 7474 13522
rect 7474 13470 7476 13522
rect 7420 13468 7476 13470
rect 7420 12684 7476 12740
rect 7308 11788 7364 11844
rect 6972 10108 7028 10164
rect 7084 11228 7140 11284
rect 7196 10892 7252 10948
rect 7084 10332 7140 10388
rect 6972 9884 7028 9940
rect 8204 14530 8260 14532
rect 8204 14478 8206 14530
rect 8206 14478 8258 14530
rect 8258 14478 8260 14530
rect 8204 14476 8260 14478
rect 7756 12908 7812 12964
rect 7868 12738 7924 12740
rect 7868 12686 7870 12738
rect 7870 12686 7922 12738
rect 7922 12686 7924 12738
rect 7868 12684 7924 12686
rect 8204 14252 8260 14308
rect 8204 13468 8260 13524
rect 8204 12738 8260 12740
rect 8204 12686 8206 12738
rect 8206 12686 8258 12738
rect 8258 12686 8260 12738
rect 8204 12684 8260 12686
rect 8428 14364 8484 14420
rect 8540 15932 8596 15988
rect 8876 17778 8932 17780
rect 8876 17726 8878 17778
rect 8878 17726 8930 17778
rect 8930 17726 8932 17778
rect 8876 17724 8932 17726
rect 9100 23660 9156 23716
rect 9324 23266 9380 23268
rect 9324 23214 9326 23266
rect 9326 23214 9378 23266
rect 9378 23214 9380 23266
rect 9324 23212 9380 23214
rect 9100 20188 9156 20244
rect 9212 21420 9268 21476
rect 9548 26236 9604 26292
rect 9660 27468 9716 27524
rect 9548 25730 9604 25732
rect 9548 25678 9550 25730
rect 9550 25678 9602 25730
rect 9602 25678 9604 25730
rect 9548 25676 9604 25678
rect 9772 26290 9828 26292
rect 9772 26238 9774 26290
rect 9774 26238 9826 26290
rect 9826 26238 9828 26290
rect 9772 26236 9828 26238
rect 9660 25452 9716 25508
rect 9772 26012 9828 26068
rect 9660 23660 9716 23716
rect 9548 23212 9604 23268
rect 9548 21868 9604 21924
rect 8988 16940 9044 16996
rect 9100 17612 9156 17668
rect 9772 23436 9828 23492
rect 9772 23212 9828 23268
rect 9324 18284 9380 18340
rect 9772 20188 9828 20244
rect 9996 32172 10052 32228
rect 10892 41580 10948 41636
rect 11228 47964 11284 48020
rect 10892 40290 10948 40292
rect 10892 40238 10894 40290
rect 10894 40238 10946 40290
rect 10946 40238 10948 40290
rect 10892 40236 10948 40238
rect 11004 38834 11060 38836
rect 11004 38782 11006 38834
rect 11006 38782 11058 38834
rect 11058 38782 11060 38834
rect 11004 38780 11060 38782
rect 11900 47292 11956 47348
rect 11788 40908 11844 40964
rect 11788 38892 11844 38948
rect 10892 37996 10948 38052
rect 10892 34914 10948 34916
rect 10892 34862 10894 34914
rect 10894 34862 10946 34914
rect 10946 34862 10948 34914
rect 10892 34860 10948 34862
rect 11228 35196 11284 35252
rect 10892 34130 10948 34132
rect 10892 34078 10894 34130
rect 10894 34078 10946 34130
rect 10946 34078 10948 34130
rect 10892 34076 10948 34078
rect 10332 31836 10388 31892
rect 10108 31724 10164 31780
rect 10220 31612 10276 31668
rect 10108 31388 10164 31444
rect 9996 31052 10052 31108
rect 10444 32956 10500 33012
rect 10108 29932 10164 29988
rect 9996 28924 10052 28980
rect 10108 27916 10164 27972
rect 10220 27692 10276 27748
rect 9996 27244 10052 27300
rect 10220 27020 10276 27076
rect 9996 26066 10052 26068
rect 9996 26014 9998 26066
rect 9998 26014 10050 26066
rect 10050 26014 10052 26066
rect 9996 26012 10052 26014
rect 9996 23436 10052 23492
rect 10108 23324 10164 23380
rect 9996 23100 10052 23156
rect 10556 29932 10612 29988
rect 10444 29820 10500 29876
rect 10444 28476 10500 28532
rect 10332 22764 10388 22820
rect 10220 20972 10276 21028
rect 10556 28364 10612 28420
rect 10556 27468 10612 27524
rect 10892 31724 10948 31780
rect 10892 30716 10948 30772
rect 10780 30156 10836 30212
rect 10892 28700 10948 28756
rect 10892 28028 10948 28084
rect 11228 34076 11284 34132
rect 11116 31890 11172 31892
rect 11116 31838 11118 31890
rect 11118 31838 11170 31890
rect 11170 31838 11172 31890
rect 11116 31836 11172 31838
rect 11788 36652 11844 36708
rect 11676 35420 11732 35476
rect 11788 34130 11844 34132
rect 11788 34078 11790 34130
rect 11790 34078 11842 34130
rect 11842 34078 11844 34130
rect 11788 34076 11844 34078
rect 11676 32172 11732 32228
rect 11452 31666 11508 31668
rect 11452 31614 11454 31666
rect 11454 31614 11506 31666
rect 11506 31614 11508 31666
rect 11452 31612 11508 31614
rect 11340 31388 11396 31444
rect 11676 31388 11732 31444
rect 11228 31052 11284 31108
rect 11116 28642 11172 28644
rect 11116 28590 11118 28642
rect 11118 28590 11170 28642
rect 11170 28590 11172 28642
rect 11116 28588 11172 28590
rect 11004 27804 11060 27860
rect 11116 28364 11172 28420
rect 10556 26012 10612 26068
rect 10668 25452 10724 25508
rect 10444 22540 10500 22596
rect 9996 20018 10052 20020
rect 9996 19966 9998 20018
rect 9998 19966 10050 20018
rect 10050 19966 10052 20018
rect 9996 19964 10052 19966
rect 9884 19346 9940 19348
rect 9884 19294 9886 19346
rect 9886 19294 9938 19346
rect 9938 19294 9940 19346
rect 9884 19292 9940 19294
rect 9884 17724 9940 17780
rect 9100 17052 9156 17108
rect 9324 16882 9380 16884
rect 9324 16830 9326 16882
rect 9326 16830 9378 16882
rect 9378 16830 9380 16882
rect 9324 16828 9380 16830
rect 8988 16156 9044 16212
rect 9100 15986 9156 15988
rect 9100 15934 9102 15986
rect 9102 15934 9154 15986
rect 9154 15934 9156 15986
rect 9100 15932 9156 15934
rect 8876 15874 8932 15876
rect 8876 15822 8878 15874
rect 8878 15822 8930 15874
rect 8930 15822 8932 15874
rect 8876 15820 8932 15822
rect 9324 14812 9380 14868
rect 9100 14754 9156 14756
rect 9100 14702 9102 14754
rect 9102 14702 9154 14754
rect 9154 14702 9156 14754
rect 9100 14700 9156 14702
rect 8876 14642 8932 14644
rect 8876 14590 8878 14642
rect 8878 14590 8930 14642
rect 8930 14590 8932 14642
rect 8876 14588 8932 14590
rect 8764 14530 8820 14532
rect 8764 14478 8766 14530
rect 8766 14478 8818 14530
rect 8818 14478 8820 14530
rect 8764 14476 8820 14478
rect 8652 14252 8708 14308
rect 8316 12572 8372 12628
rect 8540 13746 8596 13748
rect 8540 13694 8542 13746
rect 8542 13694 8594 13746
rect 8594 13694 8596 13746
rect 8540 13692 8596 13694
rect 9324 13746 9380 13748
rect 9324 13694 9326 13746
rect 9326 13694 9378 13746
rect 9378 13694 9380 13746
rect 9324 13692 9380 13694
rect 8764 13580 8820 13636
rect 7644 11116 7700 11172
rect 8988 13634 9044 13636
rect 8988 13582 8990 13634
rect 8990 13582 9042 13634
rect 9042 13582 9044 13634
rect 8988 13580 9044 13582
rect 8540 12066 8596 12068
rect 8540 12014 8542 12066
rect 8542 12014 8594 12066
rect 8594 12014 8596 12066
rect 8540 12012 8596 12014
rect 8764 11788 8820 11844
rect 8204 11506 8260 11508
rect 8204 11454 8206 11506
rect 8206 11454 8258 11506
rect 8258 11454 8260 11506
rect 8204 11452 8260 11454
rect 7756 10892 7812 10948
rect 8652 11116 8708 11172
rect 7980 10722 8036 10724
rect 7980 10670 7982 10722
rect 7982 10670 8034 10722
rect 8034 10670 8036 10722
rect 7980 10668 8036 10670
rect 7868 10610 7924 10612
rect 7868 10558 7870 10610
rect 7870 10558 7922 10610
rect 7922 10558 7924 10610
rect 7868 10556 7924 10558
rect 7756 10444 7812 10500
rect 7644 10332 7700 10388
rect 7532 9884 7588 9940
rect 7420 9154 7476 9156
rect 7420 9102 7422 9154
rect 7422 9102 7474 9154
rect 7474 9102 7476 9154
rect 7420 9100 7476 9102
rect 8092 10386 8148 10388
rect 8092 10334 8094 10386
rect 8094 10334 8146 10386
rect 8146 10334 8148 10386
rect 8092 10332 8148 10334
rect 8204 10220 8260 10276
rect 7868 9826 7924 9828
rect 7868 9774 7870 9826
rect 7870 9774 7922 9826
rect 7922 9774 7924 9826
rect 7868 9772 7924 9774
rect 7308 8930 7364 8932
rect 7308 8878 7310 8930
rect 7310 8878 7362 8930
rect 7362 8878 7364 8930
rect 7308 8876 7364 8878
rect 7196 8652 7252 8708
rect 8092 8540 8148 8596
rect 8540 8652 8596 8708
rect 8428 8482 8484 8484
rect 8428 8430 8430 8482
rect 8430 8430 8482 8482
rect 8482 8430 8484 8482
rect 8428 8428 8484 8430
rect 7756 8146 7812 8148
rect 7756 8094 7758 8146
rect 7758 8094 7810 8146
rect 7810 8094 7812 8146
rect 7756 8092 7812 8094
rect 7084 7756 7140 7812
rect 7308 7586 7364 7588
rect 7308 7534 7310 7586
rect 7310 7534 7362 7586
rect 7362 7534 7364 7586
rect 7308 7532 7364 7534
rect 7756 6748 7812 6804
rect 7756 5628 7812 5684
rect 8316 5234 8372 5236
rect 8316 5182 8318 5234
rect 8318 5182 8370 5234
rect 8370 5182 8372 5234
rect 8316 5180 8372 5182
rect 8764 10892 8820 10948
rect 8764 10668 8820 10724
rect 8988 12012 9044 12068
rect 9212 11452 9268 11508
rect 9324 12684 9380 12740
rect 9436 12348 9492 12404
rect 9324 11900 9380 11956
rect 9660 16940 9716 16996
rect 9996 17276 10052 17332
rect 10108 17500 10164 17556
rect 10108 16940 10164 16996
rect 9884 16828 9940 16884
rect 9660 16268 9716 16324
rect 9660 15148 9716 15204
rect 10108 16716 10164 16772
rect 10108 16380 10164 16436
rect 9996 15484 10052 15540
rect 9996 14700 10052 14756
rect 9884 14252 9940 14308
rect 10108 13692 10164 13748
rect 10108 13468 10164 13524
rect 10556 21586 10612 21588
rect 10556 21534 10558 21586
rect 10558 21534 10610 21586
rect 10610 21534 10612 21586
rect 10556 21532 10612 21534
rect 10556 18620 10612 18676
rect 11004 26684 11060 26740
rect 11004 26012 11060 26068
rect 11340 30604 11396 30660
rect 11564 29484 11620 29540
rect 11564 29036 11620 29092
rect 12348 45836 12404 45892
rect 12124 40796 12180 40852
rect 15036 53452 15092 53508
rect 14140 52332 14196 52388
rect 12908 40796 12964 40852
rect 13692 51548 13748 51604
rect 12124 38780 12180 38836
rect 12012 37378 12068 37380
rect 12012 37326 12014 37378
rect 12014 37326 12066 37378
rect 12066 37326 12068 37378
rect 12012 37324 12068 37326
rect 12124 37212 12180 37268
rect 12012 31948 12068 32004
rect 12124 31724 12180 31780
rect 12236 36092 12292 36148
rect 12796 37324 12852 37380
rect 12460 32844 12516 32900
rect 12572 32620 12628 32676
rect 12460 32060 12516 32116
rect 12908 31948 12964 32004
rect 12348 31388 12404 31444
rect 11788 29708 11844 29764
rect 11676 28364 11732 28420
rect 11228 26684 11284 26740
rect 11340 28028 11396 28084
rect 11228 26460 11284 26516
rect 10780 24892 10836 24948
rect 11004 25676 11060 25732
rect 11116 25788 11172 25844
rect 11116 25228 11172 25284
rect 11228 26012 11284 26068
rect 11116 24722 11172 24724
rect 11116 24670 11118 24722
rect 11118 24670 11170 24722
rect 11170 24670 11172 24722
rect 11116 24668 11172 24670
rect 10892 22988 10948 23044
rect 11004 22764 11060 22820
rect 11564 27692 11620 27748
rect 11452 27132 11508 27188
rect 11228 23826 11284 23828
rect 11228 23774 11230 23826
rect 11230 23774 11282 23826
rect 11282 23774 11284 23826
rect 11228 23772 11284 23774
rect 11340 25228 11396 25284
rect 11340 22988 11396 23044
rect 11116 22652 11172 22708
rect 11340 22764 11396 22820
rect 10892 22316 10948 22372
rect 11228 21980 11284 22036
rect 10892 21868 10948 21924
rect 11116 21756 11172 21812
rect 11004 21362 11060 21364
rect 11004 21310 11006 21362
rect 11006 21310 11058 21362
rect 11058 21310 11060 21362
rect 11004 21308 11060 21310
rect 11116 20188 11172 20244
rect 11228 21532 11284 21588
rect 11900 28642 11956 28644
rect 11900 28590 11902 28642
rect 11902 28590 11954 28642
rect 11954 28590 11956 28642
rect 11900 28588 11956 28590
rect 12348 30604 12404 30660
rect 12236 30492 12292 30548
rect 12124 29986 12180 29988
rect 12124 29934 12126 29986
rect 12126 29934 12178 29986
rect 12178 29934 12180 29986
rect 12124 29932 12180 29934
rect 12796 30604 12852 30660
rect 11788 25618 11844 25620
rect 11788 25566 11790 25618
rect 11790 25566 11842 25618
rect 11842 25566 11844 25618
rect 11788 25564 11844 25566
rect 11788 23996 11844 24052
rect 11564 23938 11620 23940
rect 11564 23886 11566 23938
rect 11566 23886 11618 23938
rect 11618 23886 11620 23938
rect 11564 23884 11620 23886
rect 11676 23772 11732 23828
rect 11452 22428 11508 22484
rect 11340 20076 11396 20132
rect 10892 19740 10948 19796
rect 11116 19068 11172 19124
rect 10780 18620 10836 18676
rect 11004 18338 11060 18340
rect 11004 18286 11006 18338
rect 11006 18286 11058 18338
rect 11058 18286 11060 18338
rect 11004 18284 11060 18286
rect 11004 18060 11060 18116
rect 10332 17276 10388 17332
rect 10444 16882 10500 16884
rect 10444 16830 10446 16882
rect 10446 16830 10498 16882
rect 10498 16830 10500 16882
rect 10444 16828 10500 16830
rect 10332 16268 10388 16324
rect 10444 16210 10500 16212
rect 10444 16158 10446 16210
rect 10446 16158 10498 16210
rect 10498 16158 10500 16210
rect 10444 16156 10500 16158
rect 11004 17388 11060 17444
rect 11116 17276 11172 17332
rect 11228 16716 11284 16772
rect 9884 11900 9940 11956
rect 9884 11506 9940 11508
rect 9884 11454 9886 11506
rect 9886 11454 9938 11506
rect 9938 11454 9940 11506
rect 9884 11452 9940 11454
rect 9548 11228 9604 11284
rect 8988 9884 9044 9940
rect 9100 11004 9156 11060
rect 9212 10892 9268 10948
rect 8876 9772 8932 9828
rect 9436 10556 9492 10612
rect 9660 10498 9716 10500
rect 9660 10446 9662 10498
rect 9662 10446 9714 10498
rect 9714 10446 9716 10498
rect 9660 10444 9716 10446
rect 9548 10386 9604 10388
rect 9548 10334 9550 10386
rect 9550 10334 9602 10386
rect 9602 10334 9604 10386
rect 9548 10332 9604 10334
rect 9772 9996 9828 10052
rect 9324 9212 9380 9268
rect 10108 12460 10164 12516
rect 10108 10108 10164 10164
rect 9884 9100 9940 9156
rect 9772 8652 9828 8708
rect 9324 8540 9380 8596
rect 9772 7362 9828 7364
rect 9772 7310 9774 7362
rect 9774 7310 9826 7362
rect 9826 7310 9828 7362
rect 9772 7308 9828 7310
rect 10220 8428 10276 8484
rect 10332 8316 10388 8372
rect 10556 15484 10612 15540
rect 11004 15260 11060 15316
rect 10668 13244 10724 13300
rect 10556 12908 10612 12964
rect 11116 11900 11172 11956
rect 11452 18284 11508 18340
rect 11116 11676 11172 11732
rect 10668 10668 10724 10724
rect 10892 10892 10948 10948
rect 10556 9436 10612 9492
rect 10556 9212 10612 9268
rect 10892 9436 10948 9492
rect 11116 11340 11172 11396
rect 11116 10780 11172 10836
rect 11340 13468 11396 13524
rect 11788 22540 11844 22596
rect 11564 18060 11620 18116
rect 11676 22316 11732 22372
rect 11564 17442 11620 17444
rect 11564 17390 11566 17442
rect 11566 17390 11618 17442
rect 11618 17390 11620 17442
rect 11564 17388 11620 17390
rect 12236 28812 12292 28868
rect 12572 28866 12628 28868
rect 12572 28814 12574 28866
rect 12574 28814 12626 28866
rect 12626 28814 12628 28866
rect 12572 28812 12628 28814
rect 12348 28252 12404 28308
rect 12684 28252 12740 28308
rect 12124 28082 12180 28084
rect 12124 28030 12126 28082
rect 12126 28030 12178 28082
rect 12178 28030 12180 28082
rect 12124 28028 12180 28030
rect 12908 30044 12964 30100
rect 13132 38668 13188 38724
rect 13356 38668 13412 38724
rect 13468 40124 13524 40180
rect 13468 39564 13524 39620
rect 13580 39116 13636 39172
rect 13244 33404 13300 33460
rect 13356 33852 13412 33908
rect 13244 33068 13300 33124
rect 13244 31724 13300 31780
rect 13244 30716 13300 30772
rect 13468 33068 13524 33124
rect 13580 31388 13636 31444
rect 13468 31164 13524 31220
rect 13468 30716 13524 30772
rect 13356 30604 13412 30660
rect 13468 30492 13524 30548
rect 13020 29484 13076 29540
rect 13020 28028 13076 28084
rect 13580 28252 13636 28308
rect 13468 27916 13524 27972
rect 12796 27692 12852 27748
rect 12908 27804 12964 27860
rect 12124 26796 12180 26852
rect 12236 26236 12292 26292
rect 12572 26908 12628 26964
rect 12572 26236 12628 26292
rect 12572 25340 12628 25396
rect 12012 23772 12068 23828
rect 11452 13020 11508 13076
rect 11676 16380 11732 16436
rect 11564 12908 11620 12964
rect 11340 10780 11396 10836
rect 11452 11394 11508 11396
rect 11452 11342 11454 11394
rect 11454 11342 11506 11394
rect 11506 11342 11508 11394
rect 11452 11340 11508 11342
rect 11564 10892 11620 10948
rect 11228 10386 11284 10388
rect 11228 10334 11230 10386
rect 11230 10334 11282 10386
rect 11282 10334 11284 10386
rect 11228 10332 11284 10334
rect 11452 10610 11508 10612
rect 11452 10558 11454 10610
rect 11454 10558 11506 10610
rect 11506 10558 11508 10610
rect 11452 10556 11508 10558
rect 11564 10444 11620 10500
rect 11340 9548 11396 9604
rect 11452 9996 11508 10052
rect 11116 8370 11172 8372
rect 11116 8318 11118 8370
rect 11118 8318 11170 8370
rect 11170 8318 11172 8370
rect 11116 8316 11172 8318
rect 10444 7308 10500 7364
rect 11004 7308 11060 7364
rect 11004 6748 11060 6804
rect 9772 6188 9828 6244
rect 8876 5682 8932 5684
rect 8876 5630 8878 5682
rect 8878 5630 8930 5682
rect 8930 5630 8932 5682
rect 8876 5628 8932 5630
rect 11676 10108 11732 10164
rect 11564 9100 11620 9156
rect 11452 8540 11508 8596
rect 11228 7196 11284 7252
rect 12236 24444 12292 24500
rect 12460 23884 12516 23940
rect 12348 23772 12404 23828
rect 12236 22316 12292 22372
rect 12124 21586 12180 21588
rect 12124 21534 12126 21586
rect 12126 21534 12178 21586
rect 12178 21534 12180 21586
rect 12124 21532 12180 21534
rect 12348 21756 12404 21812
rect 12348 20802 12404 20804
rect 12348 20750 12350 20802
rect 12350 20750 12402 20802
rect 12402 20750 12404 20802
rect 12348 20748 12404 20750
rect 12572 20524 12628 20580
rect 13020 27692 13076 27748
rect 13132 27298 13188 27300
rect 13132 27246 13134 27298
rect 13134 27246 13186 27298
rect 13186 27246 13188 27298
rect 13132 27244 13188 27246
rect 13580 27468 13636 27524
rect 12908 25452 12964 25508
rect 13020 26684 13076 26740
rect 12796 24498 12852 24500
rect 12796 24446 12798 24498
rect 12798 24446 12850 24498
rect 12850 24446 12852 24498
rect 12796 24444 12852 24446
rect 13244 25900 13300 25956
rect 12796 19964 12852 20020
rect 12796 19404 12852 19460
rect 12012 19346 12068 19348
rect 12012 19294 12014 19346
rect 12014 19294 12066 19346
rect 12066 19294 12068 19346
rect 12012 19292 12068 19294
rect 12572 19292 12628 19348
rect 11900 12460 11956 12516
rect 12460 19122 12516 19124
rect 12460 19070 12462 19122
rect 12462 19070 12514 19122
rect 12514 19070 12516 19122
rect 12460 19068 12516 19070
rect 12124 18844 12180 18900
rect 13468 23938 13524 23940
rect 13468 23886 13470 23938
rect 13470 23886 13522 23938
rect 13522 23886 13524 23938
rect 13468 23884 13524 23886
rect 13356 22764 13412 22820
rect 13356 22594 13412 22596
rect 13356 22542 13358 22594
rect 13358 22542 13410 22594
rect 13410 22542 13412 22594
rect 13356 22540 13412 22542
rect 13356 21868 13412 21924
rect 13020 18844 13076 18900
rect 13356 20524 13412 20580
rect 12684 17890 12740 17892
rect 12684 17838 12686 17890
rect 12686 17838 12738 17890
rect 12738 17838 12740 17890
rect 12684 17836 12740 17838
rect 13020 18620 13076 18676
rect 12124 17276 12180 17332
rect 11900 12290 11956 12292
rect 11900 12238 11902 12290
rect 11902 12238 11954 12290
rect 11954 12238 11956 12290
rect 11900 12236 11956 12238
rect 12796 16828 12852 16884
rect 12124 16492 12180 16548
rect 13020 16716 13076 16772
rect 13244 19234 13300 19236
rect 13244 19182 13246 19234
rect 13246 19182 13298 19234
rect 13298 19182 13300 19234
rect 13244 19180 13300 19182
rect 14028 43372 14084 43428
rect 13804 40908 13860 40964
rect 13804 38722 13860 38724
rect 13804 38670 13806 38722
rect 13806 38670 13858 38722
rect 13858 38670 13860 38722
rect 13804 38668 13860 38670
rect 13916 32284 13972 32340
rect 13804 30380 13860 30436
rect 13804 29932 13860 29988
rect 13916 29596 13972 29652
rect 13804 28700 13860 28756
rect 13916 27244 13972 27300
rect 13916 27020 13972 27076
rect 14252 42082 14308 42084
rect 14252 42030 14254 42082
rect 14254 42030 14306 42082
rect 14306 42030 14308 42082
rect 14252 42028 14308 42030
rect 14476 40908 14532 40964
rect 14924 40178 14980 40180
rect 14924 40126 14926 40178
rect 14926 40126 14978 40178
rect 14978 40126 14980 40178
rect 14924 40124 14980 40126
rect 14364 38892 14420 38948
rect 14252 38834 14308 38836
rect 14252 38782 14254 38834
rect 14254 38782 14306 38834
rect 14306 38782 14308 38834
rect 14252 38780 14308 38782
rect 19516 57260 19572 57316
rect 19852 57260 19908 57316
rect 20860 56252 20916 56308
rect 21644 56588 21700 56644
rect 16828 53564 16884 53620
rect 15596 41356 15652 41412
rect 15708 44492 15764 44548
rect 14364 36988 14420 37044
rect 14252 30210 14308 30212
rect 14252 30158 14254 30210
rect 14254 30158 14306 30210
rect 14306 30158 14308 30210
rect 14252 30156 14308 30158
rect 14476 31778 14532 31780
rect 14476 31726 14478 31778
rect 14478 31726 14530 31778
rect 14530 31726 14532 31778
rect 14476 31724 14532 31726
rect 14476 30828 14532 30884
rect 14588 30492 14644 30548
rect 13692 25004 13748 25060
rect 14364 27858 14420 27860
rect 14364 27806 14366 27858
rect 14366 27806 14418 27858
rect 14418 27806 14420 27858
rect 14364 27804 14420 27806
rect 13580 20860 13636 20916
rect 13692 24556 13748 24612
rect 13580 20018 13636 20020
rect 13580 19966 13582 20018
rect 13582 19966 13634 20018
rect 13634 19966 13636 20018
rect 13580 19964 13636 19966
rect 13580 19180 13636 19236
rect 12460 15260 12516 15316
rect 13580 18172 13636 18228
rect 12796 15036 12852 15092
rect 13356 17836 13412 17892
rect 12124 14252 12180 14308
rect 13244 15484 13300 15540
rect 13132 14140 13188 14196
rect 12572 13074 12628 13076
rect 12572 13022 12574 13074
rect 12574 13022 12626 13074
rect 12626 13022 12628 13074
rect 12572 13020 12628 13022
rect 12572 12460 12628 12516
rect 12236 12348 12292 12404
rect 12012 11004 12068 11060
rect 12348 10556 12404 10612
rect 11900 9996 11956 10052
rect 12236 10444 12292 10500
rect 11676 5906 11732 5908
rect 11676 5854 11678 5906
rect 11678 5854 11730 5906
rect 11730 5854 11732 5906
rect 11676 5852 11732 5854
rect 11116 5628 11172 5684
rect 10108 3836 10164 3892
rect 6860 140 6916 196
rect 7420 140 7476 196
rect 12124 9996 12180 10052
rect 12236 9884 12292 9940
rect 12124 9324 12180 9380
rect 12348 9324 12404 9380
rect 12460 9212 12516 9268
rect 12236 7698 12292 7700
rect 12236 7646 12238 7698
rect 12238 7646 12290 7698
rect 12290 7646 12292 7698
rect 12236 7644 12292 7646
rect 12236 7308 12292 7364
rect 12124 5794 12180 5796
rect 12124 5742 12126 5794
rect 12126 5742 12178 5794
rect 12178 5742 12180 5794
rect 12124 5740 12180 5742
rect 12684 11340 12740 11396
rect 12908 13244 12964 13300
rect 13020 11676 13076 11732
rect 12908 11452 12964 11508
rect 12796 11004 12852 11060
rect 13020 11340 13076 11396
rect 13020 11004 13076 11060
rect 13244 10780 13300 10836
rect 13020 10444 13076 10500
rect 13132 9996 13188 10052
rect 13132 9772 13188 9828
rect 12796 9212 12852 9268
rect 12796 8428 12852 8484
rect 13132 8428 13188 8484
rect 12684 6802 12740 6804
rect 12684 6750 12686 6802
rect 12686 6750 12738 6802
rect 12738 6750 12740 6802
rect 12684 6748 12740 6750
rect 12796 5292 12852 5348
rect 13244 7644 13300 7700
rect 13468 16716 13524 16772
rect 13468 14140 13524 14196
rect 13468 12908 13524 12964
rect 13804 23548 13860 23604
rect 13916 26684 13972 26740
rect 14252 26684 14308 26740
rect 14028 25004 14084 25060
rect 14252 26348 14308 26404
rect 14252 24332 14308 24388
rect 14588 26236 14644 26292
rect 14476 25900 14532 25956
rect 14588 24610 14644 24612
rect 14588 24558 14590 24610
rect 14590 24558 14642 24610
rect 14642 24558 14644 24610
rect 14588 24556 14644 24558
rect 15148 38050 15204 38052
rect 15148 37998 15150 38050
rect 15150 37998 15202 38050
rect 15202 37998 15204 38050
rect 15148 37996 15204 37998
rect 15596 39004 15652 39060
rect 15036 30882 15092 30884
rect 15036 30830 15038 30882
rect 15038 30830 15090 30882
rect 15090 30830 15092 30882
rect 15036 30828 15092 30830
rect 14812 26348 14868 26404
rect 14924 25452 14980 25508
rect 14700 24332 14756 24388
rect 15036 24556 15092 24612
rect 14364 23938 14420 23940
rect 14364 23886 14366 23938
rect 14366 23886 14418 23938
rect 14418 23886 14420 23938
rect 14364 23884 14420 23886
rect 14140 22092 14196 22148
rect 14028 21644 14084 21700
rect 14028 21474 14084 21476
rect 14028 21422 14030 21474
rect 14030 21422 14082 21474
rect 14082 21422 14084 21474
rect 14028 21420 14084 21422
rect 14700 23154 14756 23156
rect 14700 23102 14702 23154
rect 14702 23102 14754 23154
rect 14754 23102 14756 23154
rect 14700 23100 14756 23102
rect 13916 19740 13972 19796
rect 14812 22482 14868 22484
rect 14812 22430 14814 22482
rect 14814 22430 14866 22482
rect 14866 22430 14868 22482
rect 14812 22428 14868 22430
rect 14700 21980 14756 22036
rect 14812 21586 14868 21588
rect 14812 21534 14814 21586
rect 14814 21534 14866 21586
rect 14866 21534 14868 21586
rect 14812 21532 14868 21534
rect 14812 20914 14868 20916
rect 14812 20862 14814 20914
rect 14814 20862 14866 20914
rect 14866 20862 14868 20914
rect 14812 20860 14868 20862
rect 14588 20188 14644 20244
rect 15596 34972 15652 35028
rect 15596 33628 15652 33684
rect 15596 32674 15652 32676
rect 15596 32622 15598 32674
rect 15598 32622 15650 32674
rect 15650 32622 15652 32674
rect 15596 32620 15652 32622
rect 15932 37266 15988 37268
rect 15932 37214 15934 37266
rect 15934 37214 15986 37266
rect 15986 37214 15988 37266
rect 15932 37212 15988 37214
rect 15484 29372 15540 29428
rect 15260 28924 15316 28980
rect 15932 31612 15988 31668
rect 15820 30994 15876 30996
rect 15820 30942 15822 30994
rect 15822 30942 15874 30994
rect 15874 30942 15876 30994
rect 15820 30940 15876 30942
rect 15708 30210 15764 30212
rect 15708 30158 15710 30210
rect 15710 30158 15762 30210
rect 15762 30158 15764 30210
rect 15708 30156 15764 30158
rect 15708 28924 15764 28980
rect 15260 26290 15316 26292
rect 15260 26238 15262 26290
rect 15262 26238 15314 26290
rect 15314 26238 15316 26290
rect 15260 26236 15316 26238
rect 15484 25228 15540 25284
rect 15372 24556 15428 24612
rect 15148 24220 15204 24276
rect 15148 23436 15204 23492
rect 15148 23042 15204 23044
rect 15148 22990 15150 23042
rect 15150 22990 15202 23042
rect 15202 22990 15204 23042
rect 15148 22988 15204 22990
rect 15148 21756 15204 21812
rect 14476 19516 14532 19572
rect 14364 16940 14420 16996
rect 13804 15148 13860 15204
rect 13804 14812 13860 14868
rect 13804 13580 13860 13636
rect 13692 12684 13748 12740
rect 14028 12908 14084 12964
rect 14028 12178 14084 12180
rect 14028 12126 14030 12178
rect 14030 12126 14082 12178
rect 14082 12126 14084 12178
rect 14028 12124 14084 12126
rect 13468 7980 13524 8036
rect 13692 10386 13748 10388
rect 13692 10334 13694 10386
rect 13694 10334 13746 10386
rect 13746 10334 13748 10386
rect 13692 10332 13748 10334
rect 13580 7420 13636 7476
rect 13692 9996 13748 10052
rect 13356 7362 13412 7364
rect 13356 7310 13358 7362
rect 13358 7310 13410 7362
rect 13410 7310 13412 7362
rect 13356 7308 13412 7310
rect 14364 14924 14420 14980
rect 14700 19964 14756 20020
rect 14812 19852 14868 19908
rect 14812 19516 14868 19572
rect 14924 19964 14980 20020
rect 14700 18396 14756 18452
rect 14700 17052 14756 17108
rect 15596 24610 15652 24612
rect 15596 24558 15598 24610
rect 15598 24558 15650 24610
rect 15650 24558 15652 24610
rect 15596 24556 15652 24558
rect 15372 22316 15428 22372
rect 15372 21868 15428 21924
rect 15260 20636 15316 20692
rect 15372 21420 15428 21476
rect 15036 16882 15092 16884
rect 15036 16830 15038 16882
rect 15038 16830 15090 16882
rect 15090 16830 15092 16882
rect 15036 16828 15092 16830
rect 15036 15874 15092 15876
rect 15036 15822 15038 15874
rect 15038 15822 15090 15874
rect 15090 15822 15092 15874
rect 15036 15820 15092 15822
rect 14924 15484 14980 15540
rect 15148 15314 15204 15316
rect 15148 15262 15150 15314
rect 15150 15262 15202 15314
rect 15202 15262 15204 15314
rect 15148 15260 15204 15262
rect 14700 14642 14756 14644
rect 14700 14590 14702 14642
rect 14702 14590 14754 14642
rect 14754 14590 14756 14642
rect 14700 14588 14756 14590
rect 14476 14140 14532 14196
rect 14700 14364 14756 14420
rect 14364 12962 14420 12964
rect 14364 12910 14366 12962
rect 14366 12910 14418 12962
rect 14418 12910 14420 12962
rect 14364 12908 14420 12910
rect 15484 19292 15540 19348
rect 16380 37660 16436 37716
rect 16156 36652 16212 36708
rect 16268 36988 16324 37044
rect 16716 36706 16772 36708
rect 16716 36654 16718 36706
rect 16718 36654 16770 36706
rect 16770 36654 16772 36706
rect 16716 36652 16772 36654
rect 16380 34860 16436 34916
rect 16044 28642 16100 28644
rect 16044 28590 16046 28642
rect 16046 28590 16098 28642
rect 16098 28590 16100 28642
rect 16044 28588 16100 28590
rect 15820 26178 15876 26180
rect 15820 26126 15822 26178
rect 15822 26126 15874 26178
rect 15874 26126 15876 26178
rect 15820 26124 15876 26126
rect 16044 24444 16100 24500
rect 15820 24332 15876 24388
rect 16044 22146 16100 22148
rect 16044 22094 16046 22146
rect 16046 22094 16098 22146
rect 16098 22094 16100 22146
rect 16044 22092 16100 22094
rect 16380 26796 16436 26852
rect 16268 25676 16324 25732
rect 16380 25228 16436 25284
rect 16492 30156 16548 30212
rect 16940 46508 16996 46564
rect 17276 42924 17332 42980
rect 17052 41804 17108 41860
rect 17052 39228 17108 39284
rect 17164 37324 17220 37380
rect 19516 55970 19572 55972
rect 19516 55918 19518 55970
rect 19518 55918 19570 55970
rect 19570 55918 19572 55970
rect 19516 55916 19572 55918
rect 21308 55970 21364 55972
rect 21308 55918 21310 55970
rect 21310 55918 21362 55970
rect 21362 55918 21364 55970
rect 21308 55916 21364 55918
rect 19516 55692 19572 55748
rect 18284 55298 18340 55300
rect 18284 55246 18286 55298
rect 18286 55246 18338 55298
rect 18338 55246 18340 55298
rect 18284 55244 18340 55246
rect 22204 56306 22260 56308
rect 22204 56254 22206 56306
rect 22206 56254 22258 56306
rect 22258 56254 22260 56306
rect 22204 56252 22260 56254
rect 20524 55298 20580 55300
rect 20524 55246 20526 55298
rect 20526 55246 20578 55298
rect 20578 55246 20580 55298
rect 20524 55244 20580 55246
rect 20860 55298 20916 55300
rect 20860 55246 20862 55298
rect 20862 55246 20914 55298
rect 20914 55246 20916 55298
rect 20860 55244 20916 55246
rect 20076 55132 20132 55188
rect 21196 54514 21252 54516
rect 21196 54462 21198 54514
rect 21198 54462 21250 54514
rect 21250 54462 21252 54514
rect 21196 54460 21252 54462
rect 19068 54290 19124 54292
rect 19068 54238 19070 54290
rect 19070 54238 19122 54290
rect 19122 54238 19124 54290
rect 19068 54236 19124 54238
rect 20524 54124 20580 54180
rect 20076 52780 20132 52836
rect 19740 47404 19796 47460
rect 17724 44380 17780 44436
rect 17500 37772 17556 37828
rect 17612 39564 17668 39620
rect 19180 43484 19236 43540
rect 18284 41916 18340 41972
rect 18396 40124 18452 40180
rect 17500 35196 17556 35252
rect 17500 34748 17556 34804
rect 18060 34748 18116 34804
rect 18060 34188 18116 34244
rect 16940 30882 16996 30884
rect 16940 30830 16942 30882
rect 16942 30830 16994 30882
rect 16994 30830 16996 30882
rect 16940 30828 16996 30830
rect 17052 30098 17108 30100
rect 17052 30046 17054 30098
rect 17054 30046 17106 30098
rect 17106 30046 17108 30098
rect 17052 30044 17108 30046
rect 17500 33628 17556 33684
rect 17388 32732 17444 32788
rect 17836 33404 17892 33460
rect 17836 32732 17892 32788
rect 17948 32284 18004 32340
rect 18060 32172 18116 32228
rect 18284 35196 18340 35252
rect 18284 35026 18340 35028
rect 18284 34974 18286 35026
rect 18286 34974 18338 35026
rect 18338 34974 18340 35026
rect 18284 34972 18340 34974
rect 17500 30156 17556 30212
rect 17276 29932 17332 29988
rect 16268 23378 16324 23380
rect 16268 23326 16270 23378
rect 16270 23326 16322 23378
rect 16322 23326 16324 23378
rect 16268 23324 16324 23326
rect 16156 21756 16212 21812
rect 16156 21586 16212 21588
rect 16156 21534 16158 21586
rect 16158 21534 16210 21586
rect 16210 21534 16212 21586
rect 16156 21532 16212 21534
rect 16044 20802 16100 20804
rect 16044 20750 16046 20802
rect 16046 20750 16098 20802
rect 16098 20750 16100 20802
rect 16044 20748 16100 20750
rect 15596 17276 15652 17332
rect 15036 14364 15092 14420
rect 14812 13692 14868 13748
rect 15260 14028 15316 14084
rect 15148 13634 15204 13636
rect 15148 13582 15150 13634
rect 15150 13582 15202 13634
rect 15202 13582 15204 13634
rect 15148 13580 15204 13582
rect 15036 13468 15092 13524
rect 14924 13186 14980 13188
rect 14924 13134 14926 13186
rect 14926 13134 14978 13186
rect 14978 13134 14980 13186
rect 14924 13132 14980 13134
rect 14812 12178 14868 12180
rect 14812 12126 14814 12178
rect 14814 12126 14866 12178
rect 14866 12126 14868 12178
rect 14812 12124 14868 12126
rect 14812 10668 14868 10724
rect 13804 9826 13860 9828
rect 13804 9774 13806 9826
rect 13806 9774 13858 9826
rect 13858 9774 13860 9826
rect 13804 9772 13860 9774
rect 13804 9266 13860 9268
rect 13804 9214 13806 9266
rect 13806 9214 13858 9266
rect 13858 9214 13860 9266
rect 13804 9212 13860 9214
rect 14028 9324 14084 9380
rect 13916 8428 13972 8484
rect 14252 7756 14308 7812
rect 14140 6076 14196 6132
rect 13692 5852 13748 5908
rect 14588 7474 14644 7476
rect 14588 7422 14590 7474
rect 14590 7422 14642 7474
rect 14642 7422 14644 7474
rect 14588 7420 14644 7422
rect 15036 9996 15092 10052
rect 15148 10108 15204 10164
rect 15932 19292 15988 19348
rect 16268 19404 16324 19460
rect 15932 19068 15988 19124
rect 16156 19122 16212 19124
rect 16156 19070 16158 19122
rect 16158 19070 16210 19122
rect 16210 19070 16212 19122
rect 16156 19068 16212 19070
rect 16044 18844 16100 18900
rect 16156 17388 16212 17444
rect 15932 16604 15988 16660
rect 15932 16268 15988 16324
rect 16044 16210 16100 16212
rect 16044 16158 16046 16210
rect 16046 16158 16098 16210
rect 16098 16158 16100 16210
rect 16044 16156 16100 16158
rect 15932 16044 15988 16100
rect 16156 15820 16212 15876
rect 15484 11004 15540 11060
rect 15596 11676 15652 11732
rect 15596 10332 15652 10388
rect 14812 9212 14868 9268
rect 15260 9772 15316 9828
rect 15372 9436 15428 9492
rect 15372 8818 15428 8820
rect 15372 8766 15374 8818
rect 15374 8766 15426 8818
rect 15426 8766 15428 8818
rect 15372 8764 15428 8766
rect 14924 8428 14980 8484
rect 15708 9436 15764 9492
rect 16044 12908 16100 12964
rect 16156 12236 16212 12292
rect 16716 29372 16772 29428
rect 16604 27858 16660 27860
rect 16604 27806 16606 27858
rect 16606 27806 16658 27858
rect 16658 27806 16660 27858
rect 16604 27804 16660 27806
rect 16604 27356 16660 27412
rect 16716 27132 16772 27188
rect 16940 27804 16996 27860
rect 16828 24556 16884 24612
rect 16716 24220 16772 24276
rect 17388 28530 17444 28532
rect 17388 28478 17390 28530
rect 17390 28478 17442 28530
rect 17442 28478 17444 28530
rect 17388 28476 17444 28478
rect 17388 27186 17444 27188
rect 17388 27134 17390 27186
rect 17390 27134 17442 27186
rect 17442 27134 17444 27186
rect 17388 27132 17444 27134
rect 17612 27804 17668 27860
rect 17724 29932 17780 29988
rect 17836 28754 17892 28756
rect 17836 28702 17838 28754
rect 17838 28702 17890 28754
rect 17890 28702 17892 28754
rect 17836 28700 17892 28702
rect 17836 26460 17892 26516
rect 19404 36258 19460 36260
rect 19404 36206 19406 36258
rect 19406 36206 19458 36258
rect 19458 36206 19460 36258
rect 19404 36204 19460 36206
rect 19068 34914 19124 34916
rect 19068 34862 19070 34914
rect 19070 34862 19122 34914
rect 19122 34862 19124 34914
rect 19068 34860 19124 34862
rect 18732 33458 18788 33460
rect 18732 33406 18734 33458
rect 18734 33406 18786 33458
rect 18786 33406 18788 33458
rect 18732 33404 18788 33406
rect 18620 32172 18676 32228
rect 17948 25900 18004 25956
rect 18508 31612 18564 31668
rect 17276 25788 17332 25844
rect 18508 30994 18564 30996
rect 18508 30942 18510 30994
rect 18510 30942 18562 30994
rect 18562 30942 18564 30994
rect 18508 30940 18564 30942
rect 18284 29820 18340 29876
rect 18172 29260 18228 29316
rect 18620 29986 18676 29988
rect 18620 29934 18622 29986
rect 18622 29934 18674 29986
rect 18674 29934 18676 29986
rect 18620 29932 18676 29934
rect 19180 33404 19236 33460
rect 19852 41132 19908 41188
rect 19852 36204 19908 36260
rect 19740 30940 19796 30996
rect 18508 28700 18564 28756
rect 18732 25788 18788 25844
rect 18396 25340 18452 25396
rect 18732 25452 18788 25508
rect 18172 24780 18228 24836
rect 17612 24444 17668 24500
rect 17164 23996 17220 24052
rect 16940 23884 16996 23940
rect 17052 23324 17108 23380
rect 16492 21420 16548 21476
rect 16604 22988 16660 23044
rect 16492 20018 16548 20020
rect 16492 19966 16494 20018
rect 16494 19966 16546 20018
rect 16546 19966 16548 20018
rect 16492 19964 16548 19966
rect 16828 21532 16884 21588
rect 17612 23548 17668 23604
rect 19292 30098 19348 30100
rect 19292 30046 19294 30098
rect 19294 30046 19346 30098
rect 19346 30046 19348 30098
rect 19292 30044 19348 30046
rect 19964 31164 20020 31220
rect 19852 29372 19908 29428
rect 18844 23996 18900 24052
rect 18284 23548 18340 23604
rect 18620 23884 18676 23940
rect 18172 22540 18228 22596
rect 18396 23100 18452 23156
rect 18060 22482 18116 22484
rect 18060 22430 18062 22482
rect 18062 22430 18114 22482
rect 18114 22430 18116 22482
rect 18060 22428 18116 22430
rect 16828 21308 16884 21364
rect 17276 21644 17332 21700
rect 16828 20802 16884 20804
rect 16828 20750 16830 20802
rect 16830 20750 16882 20802
rect 16882 20750 16884 20802
rect 16828 20748 16884 20750
rect 17388 21532 17444 21588
rect 16716 19292 16772 19348
rect 16716 18620 16772 18676
rect 16604 18508 16660 18564
rect 17612 21308 17668 21364
rect 17612 19852 17668 19908
rect 16716 18450 16772 18452
rect 16716 18398 16718 18450
rect 16718 18398 16770 18450
rect 16770 18398 16772 18450
rect 16716 18396 16772 18398
rect 17388 19234 17444 19236
rect 17388 19182 17390 19234
rect 17390 19182 17442 19234
rect 17442 19182 17444 19234
rect 17388 19180 17444 19182
rect 18508 21698 18564 21700
rect 18508 21646 18510 21698
rect 18510 21646 18562 21698
rect 18562 21646 18564 21698
rect 18508 21644 18564 21646
rect 18284 21362 18340 21364
rect 18284 21310 18286 21362
rect 18286 21310 18338 21362
rect 18338 21310 18340 21362
rect 18284 21308 18340 21310
rect 17948 21026 18004 21028
rect 17948 20974 17950 21026
rect 17950 20974 18002 21026
rect 18002 20974 18004 21026
rect 17948 20972 18004 20974
rect 18956 23772 19012 23828
rect 19180 28476 19236 28532
rect 19292 23772 19348 23828
rect 19292 22258 19348 22260
rect 19292 22206 19294 22258
rect 19294 22206 19346 22258
rect 19346 22206 19348 22258
rect 19292 22204 19348 22206
rect 19068 22092 19124 22148
rect 18956 21644 19012 21700
rect 18844 20972 18900 21028
rect 19292 21586 19348 21588
rect 19292 21534 19294 21586
rect 19294 21534 19346 21586
rect 19346 21534 19348 21586
rect 19292 21532 19348 21534
rect 19068 20972 19124 21028
rect 19292 20972 19348 21028
rect 19292 20748 19348 20804
rect 18620 20188 18676 20244
rect 17836 19852 17892 19908
rect 17276 19068 17332 19124
rect 16828 17890 16884 17892
rect 16828 17838 16830 17890
rect 16830 17838 16882 17890
rect 16882 17838 16884 17890
rect 16828 17836 16884 17838
rect 16716 17724 16772 17780
rect 16940 17276 16996 17332
rect 17164 17164 17220 17220
rect 16380 16044 16436 16100
rect 17388 18338 17444 18340
rect 17388 18286 17390 18338
rect 17390 18286 17442 18338
rect 17442 18286 17444 18338
rect 17388 18284 17444 18286
rect 17948 19740 18004 19796
rect 17948 18450 18004 18452
rect 17948 18398 17950 18450
rect 17950 18398 18002 18450
rect 18002 18398 18004 18450
rect 17948 18396 18004 18398
rect 17836 18060 17892 18116
rect 17500 17778 17556 17780
rect 17500 17726 17502 17778
rect 17502 17726 17554 17778
rect 17554 17726 17556 17778
rect 17500 17724 17556 17726
rect 17388 17554 17444 17556
rect 17388 17502 17390 17554
rect 17390 17502 17442 17554
rect 17442 17502 17444 17554
rect 17388 17500 17444 17502
rect 17948 17500 18004 17556
rect 18620 19906 18676 19908
rect 18620 19854 18622 19906
rect 18622 19854 18674 19906
rect 18674 19854 18676 19906
rect 18620 19852 18676 19854
rect 18172 18284 18228 18340
rect 18172 17500 18228 17556
rect 18060 17388 18116 17444
rect 18844 18508 18900 18564
rect 18620 18284 18676 18340
rect 18508 17612 18564 17668
rect 18620 18060 18676 18116
rect 18844 17778 18900 17780
rect 18844 17726 18846 17778
rect 18846 17726 18898 17778
rect 18898 17726 18900 17778
rect 18844 17724 18900 17726
rect 17276 16716 17332 16772
rect 20300 31724 20356 31780
rect 20188 31388 20244 31444
rect 20300 30044 20356 30100
rect 21532 54012 21588 54068
rect 20636 53788 20692 53844
rect 21420 52444 21476 52500
rect 21644 52220 21700 52276
rect 22540 55804 22596 55860
rect 21868 55692 21924 55748
rect 22428 55298 22484 55300
rect 22428 55246 22430 55298
rect 22430 55246 22482 55298
rect 22482 55246 22484 55298
rect 22428 55244 22484 55246
rect 24332 57148 24388 57204
rect 24220 56700 24276 56756
rect 23804 56474 23860 56476
rect 23804 56422 23806 56474
rect 23806 56422 23858 56474
rect 23858 56422 23860 56474
rect 23804 56420 23860 56422
rect 23908 56474 23964 56476
rect 23908 56422 23910 56474
rect 23910 56422 23962 56474
rect 23962 56422 23964 56474
rect 23908 56420 23964 56422
rect 24012 56474 24068 56476
rect 24012 56422 24014 56474
rect 24014 56422 24066 56474
rect 24066 56422 24068 56474
rect 24012 56420 24068 56422
rect 23548 56252 23604 56308
rect 23548 55916 23604 55972
rect 23324 55244 23380 55300
rect 22316 53730 22372 53732
rect 22316 53678 22318 53730
rect 22318 53678 22370 53730
rect 22370 53678 22372 53730
rect 22316 53676 22372 53678
rect 23100 52556 23156 52612
rect 22764 52332 22820 52388
rect 20972 40908 21028 40964
rect 20748 37996 20804 38052
rect 20636 31388 20692 31444
rect 20188 26796 20244 26852
rect 19740 25394 19796 25396
rect 19740 25342 19742 25394
rect 19742 25342 19794 25394
rect 19794 25342 19796 25394
rect 19740 25340 19796 25342
rect 19740 23938 19796 23940
rect 19740 23886 19742 23938
rect 19742 23886 19794 23938
rect 19794 23886 19796 23938
rect 19740 23884 19796 23886
rect 19964 23436 20020 23492
rect 19852 23324 19908 23380
rect 19628 22092 19684 22148
rect 19740 21980 19796 22036
rect 20076 22370 20132 22372
rect 20076 22318 20078 22370
rect 20078 22318 20130 22370
rect 20130 22318 20132 22370
rect 20076 22316 20132 22318
rect 19516 21532 19572 21588
rect 19628 21362 19684 21364
rect 19628 21310 19630 21362
rect 19630 21310 19682 21362
rect 19682 21310 19684 21362
rect 19628 21308 19684 21310
rect 19964 21084 20020 21140
rect 19516 20860 19572 20916
rect 19516 20300 19572 20356
rect 20972 31388 21028 31444
rect 20972 31164 21028 31220
rect 21308 34076 21364 34132
rect 22764 52162 22820 52164
rect 22764 52110 22766 52162
rect 22766 52110 22818 52162
rect 22818 52110 22820 52162
rect 22764 52108 22820 52110
rect 21644 33628 21700 33684
rect 21756 40348 21812 40404
rect 21196 32172 21252 32228
rect 22764 37660 22820 37716
rect 22316 35420 22372 35476
rect 22092 32674 22148 32676
rect 22092 32622 22094 32674
rect 22094 32622 22146 32674
rect 22146 32622 22148 32674
rect 22092 32620 22148 32622
rect 21868 32284 21924 32340
rect 21644 31836 21700 31892
rect 21532 31724 21588 31780
rect 20412 26572 20468 26628
rect 20412 25340 20468 25396
rect 20636 24834 20692 24836
rect 20636 24782 20638 24834
rect 20638 24782 20690 24834
rect 20690 24782 20692 24834
rect 20636 24780 20692 24782
rect 21308 31388 21364 31444
rect 21308 27356 21364 27412
rect 21420 30156 21476 30212
rect 21532 30098 21588 30100
rect 21532 30046 21534 30098
rect 21534 30046 21586 30098
rect 21586 30046 21588 30098
rect 21532 30044 21588 30046
rect 21756 30156 21812 30212
rect 22092 30994 22148 30996
rect 22092 30942 22094 30994
rect 22094 30942 22146 30994
rect 22146 30942 22148 30994
rect 22092 30940 22148 30942
rect 21644 27804 21700 27860
rect 21084 26572 21140 26628
rect 21532 26684 21588 26740
rect 21420 26460 21476 26516
rect 21308 26066 21364 26068
rect 21308 26014 21310 26066
rect 21310 26014 21362 26066
rect 21362 26014 21364 26066
rect 21308 26012 21364 26014
rect 21084 24108 21140 24164
rect 20972 24050 21028 24052
rect 20972 23998 20974 24050
rect 20974 23998 21026 24050
rect 21026 23998 21028 24050
rect 20972 23996 21028 23998
rect 20188 21084 20244 21140
rect 20188 20802 20244 20804
rect 20188 20750 20190 20802
rect 20190 20750 20242 20802
rect 20242 20750 20244 20802
rect 20188 20748 20244 20750
rect 20300 20300 20356 20356
rect 19964 20018 20020 20020
rect 19964 19966 19966 20018
rect 19966 19966 20018 20018
rect 20018 19966 20020 20018
rect 19964 19964 20020 19966
rect 20748 21644 20804 21700
rect 20636 21308 20692 21364
rect 20524 20300 20580 20356
rect 20748 20524 20804 20580
rect 19740 19740 19796 19796
rect 19628 19234 19684 19236
rect 19628 19182 19630 19234
rect 19630 19182 19682 19234
rect 19682 19182 19684 19234
rect 19628 19180 19684 19182
rect 20412 18620 20468 18676
rect 19516 18060 19572 18116
rect 19516 17836 19572 17892
rect 19068 17724 19124 17780
rect 19292 17666 19348 17668
rect 19292 17614 19294 17666
rect 19294 17614 19346 17666
rect 19346 17614 19348 17666
rect 19292 17612 19348 17614
rect 19068 16994 19124 16996
rect 19068 16942 19070 16994
rect 19070 16942 19122 16994
rect 19122 16942 19124 16994
rect 19068 16940 19124 16942
rect 17612 16380 17668 16436
rect 16940 16098 16996 16100
rect 16940 16046 16942 16098
rect 16942 16046 16994 16098
rect 16994 16046 16996 16098
rect 16940 16044 16996 16046
rect 17500 15708 17556 15764
rect 16828 14754 16884 14756
rect 16828 14702 16830 14754
rect 16830 14702 16882 14754
rect 16882 14702 16884 14754
rect 16828 14700 16884 14702
rect 17052 15036 17108 15092
rect 16716 14530 16772 14532
rect 16716 14478 16718 14530
rect 16718 14478 16770 14530
rect 16770 14478 16772 14530
rect 16716 14476 16772 14478
rect 16604 13916 16660 13972
rect 16828 14364 16884 14420
rect 17276 15596 17332 15652
rect 18060 16716 18116 16772
rect 18060 15820 18116 15876
rect 17500 15148 17556 15204
rect 17164 14028 17220 14084
rect 17276 14588 17332 14644
rect 17164 13244 17220 13300
rect 16492 12178 16548 12180
rect 16492 12126 16494 12178
rect 16494 12126 16546 12178
rect 16546 12126 16548 12178
rect 16492 12124 16548 12126
rect 16268 11116 16324 11172
rect 15820 9100 15876 9156
rect 15484 8204 15540 8260
rect 15596 7980 15652 8036
rect 15484 7420 15540 7476
rect 15596 7532 15652 7588
rect 14924 7308 14980 7364
rect 16044 10108 16100 10164
rect 16268 10108 16324 10164
rect 16492 9996 16548 10052
rect 16156 9938 16212 9940
rect 16156 9886 16158 9938
rect 16158 9886 16210 9938
rect 16210 9886 16212 9938
rect 16156 9884 16212 9886
rect 16604 9436 16660 9492
rect 16044 9100 16100 9156
rect 15596 7308 15652 7364
rect 15708 7250 15764 7252
rect 15708 7198 15710 7250
rect 15710 7198 15762 7250
rect 15762 7198 15764 7250
rect 15708 7196 15764 7198
rect 15932 6412 15988 6468
rect 14812 5682 14868 5684
rect 14812 5630 14814 5682
rect 14814 5630 14866 5682
rect 14866 5630 14868 5682
rect 14812 5628 14868 5630
rect 15372 5628 15428 5684
rect 16716 8316 16772 8372
rect 16604 7756 16660 7812
rect 16716 7698 16772 7700
rect 16716 7646 16718 7698
rect 16718 7646 16770 7698
rect 16770 7646 16772 7698
rect 16716 7644 16772 7646
rect 16380 7586 16436 7588
rect 16380 7534 16382 7586
rect 16382 7534 16434 7586
rect 16434 7534 16436 7586
rect 16380 7532 16436 7534
rect 16156 7474 16212 7476
rect 16156 7422 16158 7474
rect 16158 7422 16210 7474
rect 16210 7422 16212 7474
rect 16156 7420 16212 7422
rect 16268 7308 16324 7364
rect 16268 5964 16324 6020
rect 17388 13970 17444 13972
rect 17388 13918 17390 13970
rect 17390 13918 17442 13970
rect 17442 13918 17444 13970
rect 17388 13916 17444 13918
rect 16940 11676 16996 11732
rect 17276 11340 17332 11396
rect 17388 12908 17444 12964
rect 17052 11004 17108 11060
rect 17948 15260 18004 15316
rect 18620 16604 18676 16660
rect 18284 16098 18340 16100
rect 18284 16046 18286 16098
rect 18286 16046 18338 16098
rect 18338 16046 18340 16098
rect 18284 16044 18340 16046
rect 18732 16492 18788 16548
rect 20300 18284 20356 18340
rect 19404 16492 19460 16548
rect 18396 15596 18452 15652
rect 18844 15820 18900 15876
rect 18396 15148 18452 15204
rect 17948 14476 18004 14532
rect 17724 13970 17780 13972
rect 17724 13918 17726 13970
rect 17726 13918 17778 13970
rect 17778 13918 17780 13970
rect 17724 13916 17780 13918
rect 17836 13580 17892 13636
rect 18508 14700 18564 14756
rect 18956 15596 19012 15652
rect 18620 14588 18676 14644
rect 18508 14530 18564 14532
rect 18508 14478 18510 14530
rect 18510 14478 18562 14530
rect 18562 14478 18564 14530
rect 18508 14476 18564 14478
rect 18284 14364 18340 14420
rect 18396 13746 18452 13748
rect 18396 13694 18398 13746
rect 18398 13694 18450 13746
rect 18450 13694 18452 13746
rect 18396 13692 18452 13694
rect 18284 13634 18340 13636
rect 18284 13582 18286 13634
rect 18286 13582 18338 13634
rect 18338 13582 18340 13634
rect 18284 13580 18340 13582
rect 18844 14476 18900 14532
rect 17612 12236 17668 12292
rect 17724 12012 17780 12068
rect 18060 12012 18116 12068
rect 17612 11676 17668 11732
rect 17612 10332 17668 10388
rect 17276 9996 17332 10052
rect 17052 9826 17108 9828
rect 17052 9774 17054 9826
rect 17054 9774 17106 9826
rect 17106 9774 17108 9826
rect 17052 9772 17108 9774
rect 17276 9826 17332 9828
rect 17276 9774 17278 9826
rect 17278 9774 17330 9826
rect 17330 9774 17332 9826
rect 17276 9772 17332 9774
rect 16940 9660 16996 9716
rect 17164 9212 17220 9268
rect 16940 8258 16996 8260
rect 16940 8206 16942 8258
rect 16942 8206 16994 8258
rect 16994 8206 16996 8258
rect 16940 8204 16996 8206
rect 17836 9996 17892 10052
rect 17948 9884 18004 9940
rect 17948 9714 18004 9716
rect 17948 9662 17950 9714
rect 17950 9662 18002 9714
rect 18002 9662 18004 9714
rect 17948 9660 18004 9662
rect 17724 8876 17780 8932
rect 17052 7756 17108 7812
rect 17388 7644 17444 7700
rect 16940 7420 16996 7476
rect 17388 7474 17444 7476
rect 17388 7422 17390 7474
rect 17390 7422 17442 7474
rect 17442 7422 17444 7474
rect 17388 7420 17444 7422
rect 16828 4508 16884 4564
rect 15484 4396 15540 4452
rect 11452 2156 11508 2212
rect 12012 1708 12068 1764
rect 12124 1036 12180 1092
rect 11452 140 11508 196
rect 13244 2098 13300 2100
rect 13244 2046 13246 2098
rect 13246 2046 13298 2098
rect 13298 2046 13300 2098
rect 13244 2044 13300 2046
rect 13804 1986 13860 1988
rect 13804 1934 13806 1986
rect 13806 1934 13858 1986
rect 13858 1934 13860 1986
rect 13804 1932 13860 1934
rect 14140 924 14196 980
rect 17724 5180 17780 5236
rect 18396 12962 18452 12964
rect 18396 12910 18398 12962
rect 18398 12910 18450 12962
rect 18450 12910 18452 12962
rect 18396 12908 18452 12910
rect 18508 12178 18564 12180
rect 18508 12126 18510 12178
rect 18510 12126 18562 12178
rect 18562 12126 18564 12178
rect 18508 12124 18564 12126
rect 18508 11900 18564 11956
rect 18732 11954 18788 11956
rect 18732 11902 18734 11954
rect 18734 11902 18786 11954
rect 18786 11902 18788 11954
rect 18732 11900 18788 11902
rect 19740 16492 19796 16548
rect 19964 17106 20020 17108
rect 19964 17054 19966 17106
rect 19966 17054 20018 17106
rect 20018 17054 20020 17106
rect 19964 17052 20020 17054
rect 19740 16156 19796 16212
rect 19740 15596 19796 15652
rect 19180 15314 19236 15316
rect 19180 15262 19182 15314
rect 19182 15262 19234 15314
rect 19234 15262 19236 15314
rect 19180 15260 19236 15262
rect 20076 15372 20132 15428
rect 20188 15596 20244 15652
rect 20076 15202 20132 15204
rect 20076 15150 20078 15202
rect 20078 15150 20130 15202
rect 20130 15150 20132 15202
rect 20076 15148 20132 15150
rect 19180 14642 19236 14644
rect 19180 14590 19182 14642
rect 19182 14590 19234 14642
rect 19234 14590 19236 14642
rect 19180 14588 19236 14590
rect 19068 14028 19124 14084
rect 19964 14700 20020 14756
rect 19964 14530 20020 14532
rect 19964 14478 19966 14530
rect 19966 14478 20018 14530
rect 20018 14478 20020 14530
rect 19964 14476 20020 14478
rect 19964 14252 20020 14308
rect 19516 14028 19572 14084
rect 18956 12572 19012 12628
rect 19516 13692 19572 13748
rect 19292 12572 19348 12628
rect 19964 13634 20020 13636
rect 19964 13582 19966 13634
rect 19966 13582 20018 13634
rect 20018 13582 20020 13634
rect 19964 13580 20020 13582
rect 19740 13522 19796 13524
rect 19740 13470 19742 13522
rect 19742 13470 19794 13522
rect 19794 13470 19796 13522
rect 19740 13468 19796 13470
rect 19628 12796 19684 12852
rect 19516 12572 19572 12628
rect 19628 12236 19684 12292
rect 18284 11452 18340 11508
rect 18844 11452 18900 11508
rect 18396 11340 18452 11396
rect 18284 10834 18340 10836
rect 18284 10782 18286 10834
rect 18286 10782 18338 10834
rect 18338 10782 18340 10834
rect 18284 10780 18340 10782
rect 18172 10108 18228 10164
rect 18956 11004 19012 11060
rect 18732 10892 18788 10948
rect 18620 10556 18676 10612
rect 18172 9324 18228 9380
rect 18956 10050 19012 10052
rect 18956 9998 18958 10050
rect 18958 9998 19010 10050
rect 19010 9998 19012 10050
rect 18956 9996 19012 9998
rect 18060 4844 18116 4900
rect 18508 8316 18564 8372
rect 17500 4172 17556 4228
rect 16940 4060 16996 4116
rect 18172 588 18228 644
rect 18844 8204 18900 8260
rect 18844 7980 18900 8036
rect 19180 11394 19236 11396
rect 19180 11342 19182 11394
rect 19182 11342 19234 11394
rect 19234 11342 19236 11394
rect 19180 11340 19236 11342
rect 19740 11900 19796 11956
rect 19404 11452 19460 11508
rect 19516 11788 19572 11844
rect 19404 10498 19460 10500
rect 19404 10446 19406 10498
rect 19406 10446 19458 10498
rect 19458 10446 19460 10498
rect 19404 10444 19460 10446
rect 19404 10108 19460 10164
rect 19292 8876 19348 8932
rect 20188 13074 20244 13076
rect 20188 13022 20190 13074
rect 20190 13022 20242 13074
rect 20242 13022 20244 13074
rect 20188 13020 20244 13022
rect 19964 12178 20020 12180
rect 19964 12126 19966 12178
rect 19966 12126 20018 12178
rect 20018 12126 20020 12178
rect 19964 12124 20020 12126
rect 19964 11394 20020 11396
rect 19964 11342 19966 11394
rect 19966 11342 20018 11394
rect 20018 11342 20020 11394
rect 19964 11340 20020 11342
rect 19628 10780 19684 10836
rect 19628 10108 19684 10164
rect 20076 10892 20132 10948
rect 19516 9660 19572 9716
rect 19628 8876 19684 8932
rect 19628 8204 19684 8260
rect 19964 10668 20020 10724
rect 19852 10108 19908 10164
rect 19740 7868 19796 7924
rect 20076 8764 20132 8820
rect 20188 12572 20244 12628
rect 20188 8316 20244 8372
rect 19964 7868 20020 7924
rect 19964 7196 20020 7252
rect 20412 17612 20468 17668
rect 21868 26012 21924 26068
rect 21644 24780 21700 24836
rect 21420 22316 21476 22372
rect 21196 21644 21252 21700
rect 21084 21586 21140 21588
rect 21084 21534 21086 21586
rect 21086 21534 21138 21586
rect 21138 21534 21140 21586
rect 21084 21532 21140 21534
rect 20972 21308 21028 21364
rect 21196 20524 21252 20580
rect 20972 20130 21028 20132
rect 20972 20078 20974 20130
rect 20974 20078 21026 20130
rect 21026 20078 21028 20130
rect 20972 20076 21028 20078
rect 20860 19964 20916 20020
rect 20860 19794 20916 19796
rect 20860 19742 20862 19794
rect 20862 19742 20914 19794
rect 20914 19742 20916 19794
rect 20860 19740 20916 19742
rect 20636 18060 20692 18116
rect 20860 17612 20916 17668
rect 20972 17276 21028 17332
rect 20524 16716 20580 16772
rect 20636 16380 20692 16436
rect 20860 16658 20916 16660
rect 20860 16606 20862 16658
rect 20862 16606 20914 16658
rect 20914 16606 20916 16658
rect 20860 16604 20916 16606
rect 20860 14700 20916 14756
rect 20748 14364 20804 14420
rect 21084 14364 21140 14420
rect 22428 30716 22484 30772
rect 22092 24162 22148 24164
rect 22092 24110 22094 24162
rect 22094 24110 22146 24162
rect 22146 24110 22148 24162
rect 22092 24108 22148 24110
rect 21868 22428 21924 22484
rect 21980 21756 22036 21812
rect 21756 20802 21812 20804
rect 21756 20750 21758 20802
rect 21758 20750 21810 20802
rect 21810 20750 21812 20802
rect 21756 20748 21812 20750
rect 22204 20076 22260 20132
rect 22092 18508 22148 18564
rect 21532 18396 21588 18452
rect 21756 18396 21812 18452
rect 21420 18284 21476 18340
rect 21532 17666 21588 17668
rect 21532 17614 21534 17666
rect 21534 17614 21586 17666
rect 21586 17614 21588 17666
rect 21532 17612 21588 17614
rect 21644 17052 21700 17108
rect 21308 16380 21364 16436
rect 20972 14028 21028 14084
rect 20860 13692 20916 13748
rect 20972 13580 21028 13636
rect 20748 13522 20804 13524
rect 20748 13470 20750 13522
rect 20750 13470 20802 13522
rect 20802 13470 20804 13522
rect 20748 13468 20804 13470
rect 20860 13356 20916 13412
rect 20636 13020 20692 13076
rect 21532 15708 21588 15764
rect 21420 15484 21476 15540
rect 20860 12178 20916 12180
rect 20860 12126 20862 12178
rect 20862 12126 20914 12178
rect 20914 12126 20916 12178
rect 20860 12124 20916 12126
rect 21084 11954 21140 11956
rect 21084 11902 21086 11954
rect 21086 11902 21138 11954
rect 21138 11902 21140 11954
rect 21084 11900 21140 11902
rect 20860 9996 20916 10052
rect 21196 11340 21252 11396
rect 21084 8428 21140 8484
rect 20972 8370 21028 8372
rect 20972 8318 20974 8370
rect 20974 8318 21026 8370
rect 21026 8318 21028 8370
rect 20972 8316 21028 8318
rect 20300 7980 20356 8036
rect 20300 7196 20356 7252
rect 19516 5964 19572 6020
rect 20860 6748 20916 6804
rect 19068 3388 19124 3444
rect 18508 252 18564 308
rect 19516 364 19572 420
rect 20972 6524 21028 6580
rect 21308 15036 21364 15092
rect 21420 14028 21476 14084
rect 21420 13746 21476 13748
rect 21420 13694 21422 13746
rect 21422 13694 21474 13746
rect 21474 13694 21476 13746
rect 21420 13692 21476 13694
rect 21308 13468 21364 13524
rect 21644 15202 21700 15204
rect 21644 15150 21646 15202
rect 21646 15150 21698 15202
rect 21698 15150 21700 15202
rect 21644 15148 21700 15150
rect 21532 12124 21588 12180
rect 21644 13692 21700 13748
rect 21308 10780 21364 10836
rect 21196 7980 21252 8036
rect 21308 8316 21364 8372
rect 21308 7420 21364 7476
rect 22316 18396 22372 18452
rect 22092 17500 22148 17556
rect 21980 16098 22036 16100
rect 21980 16046 21982 16098
rect 21982 16046 22034 16098
rect 22034 16046 22036 16098
rect 21980 16044 22036 16046
rect 22092 15036 22148 15092
rect 22092 9996 22148 10052
rect 21868 8988 21924 9044
rect 21980 9212 22036 9268
rect 21756 7868 21812 7924
rect 21868 7644 21924 7700
rect 21868 6188 21924 6244
rect 21756 6076 21812 6132
rect 21084 2940 21140 2996
rect 20972 2044 21028 2100
rect 22316 8316 22372 8372
rect 22092 7420 22148 7476
rect 22652 23996 22708 24052
rect 22652 18284 22708 18340
rect 23212 31276 23268 31332
rect 23100 30210 23156 30212
rect 23100 30158 23102 30210
rect 23102 30158 23154 30210
rect 23154 30158 23156 30210
rect 23100 30156 23156 30158
rect 23100 29372 23156 29428
rect 22764 17724 22820 17780
rect 22876 22428 22932 22484
rect 22540 16828 22596 16884
rect 23212 20524 23268 20580
rect 23884 55692 23940 55748
rect 23804 54906 23860 54908
rect 23804 54854 23806 54906
rect 23806 54854 23858 54906
rect 23858 54854 23860 54906
rect 23804 54852 23860 54854
rect 23908 54906 23964 54908
rect 23908 54854 23910 54906
rect 23910 54854 23962 54906
rect 23962 54854 23964 54906
rect 23908 54852 23964 54854
rect 24012 54906 24068 54908
rect 24012 54854 24014 54906
rect 24014 54854 24066 54906
rect 24066 54854 24068 54906
rect 24012 54852 24068 54854
rect 23772 54738 23828 54740
rect 23772 54686 23774 54738
rect 23774 54686 23826 54738
rect 23826 54686 23828 54738
rect 23772 54684 23828 54686
rect 23660 54572 23716 54628
rect 23772 54348 23828 54404
rect 24108 54124 24164 54180
rect 23804 53338 23860 53340
rect 23804 53286 23806 53338
rect 23806 53286 23858 53338
rect 23858 53286 23860 53338
rect 23804 53284 23860 53286
rect 23908 53338 23964 53340
rect 23908 53286 23910 53338
rect 23910 53286 23962 53338
rect 23962 53286 23964 53338
rect 23908 53284 23964 53286
rect 24012 53338 24068 53340
rect 24012 53286 24014 53338
rect 24014 53286 24066 53338
rect 24066 53286 24068 53338
rect 24012 53284 24068 53286
rect 24444 56306 24500 56308
rect 24444 56254 24446 56306
rect 24446 56254 24498 56306
rect 24498 56254 24500 56306
rect 24444 56252 24500 56254
rect 24892 56252 24948 56308
rect 25452 55970 25508 55972
rect 25452 55918 25454 55970
rect 25454 55918 25506 55970
rect 25506 55918 25508 55970
rect 25452 55916 25508 55918
rect 24464 55690 24520 55692
rect 24464 55638 24466 55690
rect 24466 55638 24518 55690
rect 24518 55638 24520 55690
rect 24464 55636 24520 55638
rect 24568 55690 24624 55692
rect 24568 55638 24570 55690
rect 24570 55638 24622 55690
rect 24622 55638 24624 55690
rect 24568 55636 24624 55638
rect 24672 55690 24728 55692
rect 24672 55638 24674 55690
rect 24674 55638 24726 55690
rect 24726 55638 24728 55690
rect 24672 55636 24728 55638
rect 25004 55356 25060 55412
rect 24668 55298 24724 55300
rect 24668 55246 24670 55298
rect 24670 55246 24722 55298
rect 24722 55246 24724 55298
rect 24668 55244 24724 55246
rect 24332 54572 24388 54628
rect 25900 57260 25956 57316
rect 26236 57260 26292 57316
rect 27580 56588 27636 56644
rect 26012 56306 26068 56308
rect 26012 56254 26014 56306
rect 26014 56254 26066 56306
rect 26066 56254 26068 56306
rect 26012 56252 26068 56254
rect 25788 56140 25844 56196
rect 25676 54460 25732 54516
rect 25004 54348 25060 54404
rect 24668 54236 24724 54292
rect 24464 54122 24520 54124
rect 24464 54070 24466 54122
rect 24466 54070 24518 54122
rect 24518 54070 24520 54122
rect 24464 54068 24520 54070
rect 24568 54122 24624 54124
rect 24568 54070 24570 54122
rect 24570 54070 24622 54122
rect 24622 54070 24624 54122
rect 24568 54068 24624 54070
rect 24672 54122 24728 54124
rect 24672 54070 24674 54122
rect 24674 54070 24726 54122
rect 24726 54070 24728 54122
rect 24672 54068 24728 54070
rect 24668 53564 24724 53620
rect 25676 53618 25732 53620
rect 25676 53566 25678 53618
rect 25678 53566 25730 53618
rect 25730 53566 25732 53618
rect 25676 53564 25732 53566
rect 24668 52668 24724 52724
rect 25452 52668 25508 52724
rect 24464 52554 24520 52556
rect 24464 52502 24466 52554
rect 24466 52502 24518 52554
rect 24518 52502 24520 52554
rect 24464 52500 24520 52502
rect 24568 52554 24624 52556
rect 24568 52502 24570 52554
rect 24570 52502 24622 52554
rect 24622 52502 24624 52554
rect 24568 52500 24624 52502
rect 24672 52554 24728 52556
rect 24672 52502 24674 52554
rect 24674 52502 24726 52554
rect 24726 52502 24728 52554
rect 24672 52500 24728 52502
rect 24668 52274 24724 52276
rect 24668 52222 24670 52274
rect 24670 52222 24722 52274
rect 24722 52222 24724 52274
rect 24668 52220 24724 52222
rect 23804 51770 23860 51772
rect 23804 51718 23806 51770
rect 23806 51718 23858 51770
rect 23858 51718 23860 51770
rect 23804 51716 23860 51718
rect 23908 51770 23964 51772
rect 23908 51718 23910 51770
rect 23910 51718 23962 51770
rect 23962 51718 23964 51770
rect 23908 51716 23964 51718
rect 24012 51770 24068 51772
rect 24012 51718 24014 51770
rect 24014 51718 24066 51770
rect 24066 51718 24068 51770
rect 25676 51772 25732 51828
rect 24012 51716 24068 51718
rect 26236 53900 26292 53956
rect 26236 53452 26292 53508
rect 26236 52834 26292 52836
rect 26236 52782 26238 52834
rect 26238 52782 26290 52834
rect 26290 52782 26292 52834
rect 26236 52780 26292 52782
rect 24668 51266 24724 51268
rect 24668 51214 24670 51266
rect 24670 51214 24722 51266
rect 24722 51214 24724 51266
rect 24668 51212 24724 51214
rect 24464 50986 24520 50988
rect 24464 50934 24466 50986
rect 24466 50934 24518 50986
rect 24518 50934 24520 50986
rect 24464 50932 24520 50934
rect 24568 50986 24624 50988
rect 24568 50934 24570 50986
rect 24570 50934 24622 50986
rect 24622 50934 24624 50986
rect 24568 50932 24624 50934
rect 24672 50986 24728 50988
rect 24672 50934 24674 50986
rect 24674 50934 24726 50986
rect 24726 50934 24728 50986
rect 24672 50932 24728 50934
rect 23996 50594 24052 50596
rect 23996 50542 23998 50594
rect 23998 50542 24050 50594
rect 24050 50542 24052 50594
rect 23996 50540 24052 50542
rect 24668 50428 24724 50484
rect 25676 50482 25732 50484
rect 25676 50430 25678 50482
rect 25678 50430 25730 50482
rect 25730 50430 25732 50482
rect 25676 50428 25732 50430
rect 23804 50202 23860 50204
rect 23804 50150 23806 50202
rect 23806 50150 23858 50202
rect 23858 50150 23860 50202
rect 23804 50148 23860 50150
rect 23908 50202 23964 50204
rect 23908 50150 23910 50202
rect 23910 50150 23962 50202
rect 23962 50150 23964 50202
rect 23908 50148 23964 50150
rect 24012 50202 24068 50204
rect 24012 50150 24014 50202
rect 24014 50150 24066 50202
rect 24066 50150 24068 50202
rect 24012 50148 24068 50150
rect 24668 49698 24724 49700
rect 24668 49646 24670 49698
rect 24670 49646 24722 49698
rect 24722 49646 24724 49698
rect 24668 49644 24724 49646
rect 25676 49532 25732 49588
rect 24464 49418 24520 49420
rect 24464 49366 24466 49418
rect 24466 49366 24518 49418
rect 24518 49366 24520 49418
rect 24464 49364 24520 49366
rect 24568 49418 24624 49420
rect 24568 49366 24570 49418
rect 24570 49366 24622 49418
rect 24622 49366 24624 49418
rect 24568 49364 24624 49366
rect 24672 49418 24728 49420
rect 24672 49366 24674 49418
rect 24674 49366 24726 49418
rect 24726 49366 24728 49418
rect 24672 49364 24728 49366
rect 24668 49026 24724 49028
rect 24668 48974 24670 49026
rect 24670 48974 24722 49026
rect 24722 48974 24724 49026
rect 24668 48972 24724 48974
rect 23804 48634 23860 48636
rect 23804 48582 23806 48634
rect 23806 48582 23858 48634
rect 23858 48582 23860 48634
rect 23804 48580 23860 48582
rect 23908 48634 23964 48636
rect 23908 48582 23910 48634
rect 23910 48582 23962 48634
rect 23962 48582 23964 48634
rect 23908 48580 23964 48582
rect 24012 48634 24068 48636
rect 24012 48582 24014 48634
rect 24014 48582 24066 48634
rect 24066 48582 24068 48634
rect 25676 48636 25732 48692
rect 24012 48580 24068 48582
rect 24464 47850 24520 47852
rect 24464 47798 24466 47850
rect 24466 47798 24518 47850
rect 24518 47798 24520 47850
rect 24464 47796 24520 47798
rect 24568 47850 24624 47852
rect 24568 47798 24570 47850
rect 24570 47798 24622 47850
rect 24622 47798 24624 47850
rect 24568 47796 24624 47798
rect 24672 47850 24728 47852
rect 24672 47798 24674 47850
rect 24674 47798 24726 47850
rect 24726 47798 24728 47850
rect 24672 47796 24728 47798
rect 24668 47292 24724 47348
rect 25676 47346 25732 47348
rect 25676 47294 25678 47346
rect 25678 47294 25730 47346
rect 25730 47294 25732 47346
rect 25676 47292 25732 47294
rect 23804 47066 23860 47068
rect 23804 47014 23806 47066
rect 23806 47014 23858 47066
rect 23858 47014 23860 47066
rect 23804 47012 23860 47014
rect 23908 47066 23964 47068
rect 23908 47014 23910 47066
rect 23910 47014 23962 47066
rect 23962 47014 23964 47066
rect 23908 47012 23964 47014
rect 24012 47066 24068 47068
rect 24012 47014 24014 47066
rect 24014 47014 24066 47066
rect 24066 47014 24068 47066
rect 24012 47012 24068 47014
rect 23804 45498 23860 45500
rect 23804 45446 23806 45498
rect 23806 45446 23858 45498
rect 23858 45446 23860 45498
rect 23804 45444 23860 45446
rect 23908 45498 23964 45500
rect 23908 45446 23910 45498
rect 23910 45446 23962 45498
rect 23962 45446 23964 45498
rect 23908 45444 23964 45446
rect 24012 45498 24068 45500
rect 24012 45446 24014 45498
rect 24014 45446 24066 45498
rect 24066 45446 24068 45498
rect 24012 45444 24068 45446
rect 23804 43930 23860 43932
rect 23804 43878 23806 43930
rect 23806 43878 23858 43930
rect 23858 43878 23860 43930
rect 23804 43876 23860 43878
rect 23908 43930 23964 43932
rect 23908 43878 23910 43930
rect 23910 43878 23962 43930
rect 23962 43878 23964 43930
rect 23908 43876 23964 43878
rect 24012 43930 24068 43932
rect 24012 43878 24014 43930
rect 24014 43878 24066 43930
rect 24066 43878 24068 43930
rect 24012 43876 24068 43878
rect 23804 42362 23860 42364
rect 23804 42310 23806 42362
rect 23806 42310 23858 42362
rect 23858 42310 23860 42362
rect 23804 42308 23860 42310
rect 23908 42362 23964 42364
rect 23908 42310 23910 42362
rect 23910 42310 23962 42362
rect 23962 42310 23964 42362
rect 23908 42308 23964 42310
rect 24012 42362 24068 42364
rect 24012 42310 24014 42362
rect 24014 42310 24066 42362
rect 24066 42310 24068 42362
rect 24012 42308 24068 42310
rect 27244 54012 27300 54068
rect 27020 53116 27076 53172
rect 26460 51436 26516 51492
rect 26236 49868 26292 49924
rect 25900 46732 25956 46788
rect 25676 46396 25732 46452
rect 24464 46282 24520 46284
rect 24464 46230 24466 46282
rect 24466 46230 24518 46282
rect 24518 46230 24520 46282
rect 24464 46228 24520 46230
rect 24568 46282 24624 46284
rect 24568 46230 24570 46282
rect 24570 46230 24622 46282
rect 24622 46230 24624 46282
rect 24568 46228 24624 46230
rect 24672 46282 24728 46284
rect 24672 46230 24674 46282
rect 24674 46230 24726 46282
rect 24726 46230 24728 46282
rect 24672 46228 24728 46230
rect 24464 44714 24520 44716
rect 24464 44662 24466 44714
rect 24466 44662 24518 44714
rect 24518 44662 24520 44714
rect 24464 44660 24520 44662
rect 24568 44714 24624 44716
rect 24568 44662 24570 44714
rect 24570 44662 24622 44714
rect 24622 44662 24624 44714
rect 24568 44660 24624 44662
rect 24672 44714 24728 44716
rect 24672 44662 24674 44714
rect 24674 44662 24726 44714
rect 24726 44662 24728 44714
rect 24672 44660 24728 44662
rect 25676 45500 25732 45556
rect 24892 44492 24948 44548
rect 25676 44210 25732 44212
rect 25676 44158 25678 44210
rect 25678 44158 25730 44210
rect 25730 44158 25732 44210
rect 25676 44156 25732 44158
rect 24464 43146 24520 43148
rect 24464 43094 24466 43146
rect 24466 43094 24518 43146
rect 24518 43094 24520 43146
rect 24464 43092 24520 43094
rect 24568 43146 24624 43148
rect 24568 43094 24570 43146
rect 24570 43094 24622 43146
rect 24622 43094 24624 43146
rect 24568 43092 24624 43094
rect 24672 43146 24728 43148
rect 24672 43094 24674 43146
rect 24674 43094 24726 43146
rect 24726 43094 24728 43146
rect 24672 43092 24728 43094
rect 24332 41916 24388 41972
rect 24668 41692 24724 41748
rect 24464 41578 24520 41580
rect 24464 41526 24466 41578
rect 24466 41526 24518 41578
rect 24518 41526 24520 41578
rect 24464 41524 24520 41526
rect 24568 41578 24624 41580
rect 24568 41526 24570 41578
rect 24570 41526 24622 41578
rect 24622 41526 24624 41578
rect 24568 41524 24624 41526
rect 24672 41578 24728 41580
rect 24672 41526 24674 41578
rect 24674 41526 24726 41578
rect 24726 41526 24728 41578
rect 24672 41524 24728 41526
rect 23804 40794 23860 40796
rect 23804 40742 23806 40794
rect 23806 40742 23858 40794
rect 23858 40742 23860 40794
rect 23804 40740 23860 40742
rect 23908 40794 23964 40796
rect 23908 40742 23910 40794
rect 23910 40742 23962 40794
rect 23962 40742 23964 40794
rect 23908 40740 23964 40742
rect 24012 40794 24068 40796
rect 24012 40742 24014 40794
rect 24014 40742 24066 40794
rect 24066 40742 24068 40794
rect 24012 40740 24068 40742
rect 24668 40402 24724 40404
rect 24668 40350 24670 40402
rect 24670 40350 24722 40402
rect 24722 40350 24724 40402
rect 24668 40348 24724 40350
rect 24780 40124 24836 40180
rect 24464 40010 24520 40012
rect 24464 39958 24466 40010
rect 24466 39958 24518 40010
rect 24518 39958 24520 40010
rect 24464 39956 24520 39958
rect 24568 40010 24624 40012
rect 24568 39958 24570 40010
rect 24570 39958 24622 40010
rect 24622 39958 24624 40010
rect 24568 39956 24624 39958
rect 24672 40010 24728 40012
rect 24672 39958 24674 40010
rect 24674 39958 24726 40010
rect 24726 39958 24728 40010
rect 24672 39956 24728 39958
rect 24892 39788 24948 39844
rect 23804 39226 23860 39228
rect 23804 39174 23806 39226
rect 23806 39174 23858 39226
rect 23858 39174 23860 39226
rect 23804 39172 23860 39174
rect 23908 39226 23964 39228
rect 23908 39174 23910 39226
rect 23910 39174 23962 39226
rect 23962 39174 23964 39226
rect 23908 39172 23964 39174
rect 24012 39226 24068 39228
rect 24012 39174 24014 39226
rect 24014 39174 24066 39226
rect 24066 39174 24068 39226
rect 24012 39172 24068 39174
rect 24464 38442 24520 38444
rect 24464 38390 24466 38442
rect 24466 38390 24518 38442
rect 24518 38390 24520 38442
rect 24464 38388 24520 38390
rect 24568 38442 24624 38444
rect 24568 38390 24570 38442
rect 24570 38390 24622 38442
rect 24622 38390 24624 38442
rect 24568 38388 24624 38390
rect 24672 38442 24728 38444
rect 24672 38390 24674 38442
rect 24674 38390 24726 38442
rect 24726 38390 24728 38442
rect 24672 38388 24728 38390
rect 23804 37658 23860 37660
rect 23804 37606 23806 37658
rect 23806 37606 23858 37658
rect 23858 37606 23860 37658
rect 23804 37604 23860 37606
rect 23908 37658 23964 37660
rect 23908 37606 23910 37658
rect 23910 37606 23962 37658
rect 23962 37606 23964 37658
rect 23908 37604 23964 37606
rect 24012 37658 24068 37660
rect 24012 37606 24014 37658
rect 24014 37606 24066 37658
rect 24066 37606 24068 37658
rect 24012 37604 24068 37606
rect 24668 37436 24724 37492
rect 24668 36988 24724 37044
rect 24464 36874 24520 36876
rect 24464 36822 24466 36874
rect 24466 36822 24518 36874
rect 24518 36822 24520 36874
rect 24464 36820 24520 36822
rect 24568 36874 24624 36876
rect 24568 36822 24570 36874
rect 24570 36822 24622 36874
rect 24622 36822 24624 36874
rect 24568 36820 24624 36822
rect 24672 36874 24728 36876
rect 24672 36822 24674 36874
rect 24674 36822 24726 36874
rect 24726 36822 24728 36874
rect 24672 36820 24728 36822
rect 24668 36652 24724 36708
rect 23804 36090 23860 36092
rect 23804 36038 23806 36090
rect 23806 36038 23858 36090
rect 23858 36038 23860 36090
rect 23804 36036 23860 36038
rect 23908 36090 23964 36092
rect 23908 36038 23910 36090
rect 23910 36038 23962 36090
rect 23962 36038 23964 36090
rect 23908 36036 23964 36038
rect 24012 36090 24068 36092
rect 24012 36038 24014 36090
rect 24014 36038 24066 36090
rect 24066 36038 24068 36090
rect 24012 36036 24068 36038
rect 25676 43260 25732 43316
rect 25676 42364 25732 42420
rect 25676 41074 25732 41076
rect 25676 41022 25678 41074
rect 25678 41022 25730 41074
rect 25730 41022 25732 41074
rect 25676 41020 25732 41022
rect 25788 40908 25844 40964
rect 25676 40124 25732 40180
rect 25676 39228 25732 39284
rect 25004 35756 25060 35812
rect 25340 38668 25396 38724
rect 24892 35420 24948 35476
rect 24464 35306 24520 35308
rect 24464 35254 24466 35306
rect 24466 35254 24518 35306
rect 24518 35254 24520 35306
rect 24464 35252 24520 35254
rect 24568 35306 24624 35308
rect 24568 35254 24570 35306
rect 24570 35254 24622 35306
rect 24622 35254 24624 35306
rect 24568 35252 24624 35254
rect 24672 35306 24728 35308
rect 24672 35254 24674 35306
rect 24674 35254 24726 35306
rect 24726 35254 24728 35306
rect 24672 35252 24728 35254
rect 23804 34522 23860 34524
rect 23804 34470 23806 34522
rect 23806 34470 23858 34522
rect 23858 34470 23860 34522
rect 23804 34468 23860 34470
rect 23908 34522 23964 34524
rect 23908 34470 23910 34522
rect 23910 34470 23962 34522
rect 23962 34470 23964 34522
rect 23908 34468 23964 34470
rect 24012 34522 24068 34524
rect 24012 34470 24014 34522
rect 24014 34470 24066 34522
rect 24066 34470 24068 34522
rect 24012 34468 24068 34470
rect 23436 33628 23492 33684
rect 23804 32954 23860 32956
rect 23804 32902 23806 32954
rect 23806 32902 23858 32954
rect 23858 32902 23860 32954
rect 23804 32900 23860 32902
rect 23908 32954 23964 32956
rect 23908 32902 23910 32954
rect 23910 32902 23962 32954
rect 23962 32902 23964 32954
rect 23908 32900 23964 32902
rect 24012 32954 24068 32956
rect 24012 32902 24014 32954
rect 24014 32902 24066 32954
rect 24066 32902 24068 32954
rect 24012 32900 24068 32902
rect 24668 33852 24724 33908
rect 25228 33964 25284 34020
rect 24464 33738 24520 33740
rect 24464 33686 24466 33738
rect 24466 33686 24518 33738
rect 24518 33686 24520 33738
rect 24464 33684 24520 33686
rect 24568 33738 24624 33740
rect 24568 33686 24570 33738
rect 24570 33686 24622 33738
rect 24622 33686 24624 33738
rect 24568 33684 24624 33686
rect 24672 33738 24728 33740
rect 24672 33686 24674 33738
rect 24674 33686 24726 33738
rect 24726 33686 24728 33738
rect 24672 33684 24728 33686
rect 24892 33516 24948 33572
rect 24668 33180 24724 33236
rect 24464 32170 24520 32172
rect 24464 32118 24466 32170
rect 24466 32118 24518 32170
rect 24518 32118 24520 32170
rect 24464 32116 24520 32118
rect 24568 32170 24624 32172
rect 24568 32118 24570 32170
rect 24570 32118 24622 32170
rect 24622 32118 24624 32170
rect 24568 32116 24624 32118
rect 24672 32170 24728 32172
rect 24672 32118 24674 32170
rect 24674 32118 24726 32170
rect 24726 32118 24728 32170
rect 24672 32116 24728 32118
rect 24332 31500 24388 31556
rect 23804 31386 23860 31388
rect 23660 31276 23716 31332
rect 23804 31334 23806 31386
rect 23806 31334 23858 31386
rect 23858 31334 23860 31386
rect 23804 31332 23860 31334
rect 23908 31386 23964 31388
rect 23908 31334 23910 31386
rect 23910 31334 23962 31386
rect 23962 31334 23964 31386
rect 23908 31332 23964 31334
rect 24012 31386 24068 31388
rect 24012 31334 24014 31386
rect 24014 31334 24066 31386
rect 24066 31334 24068 31386
rect 24012 31332 24068 31334
rect 23660 30994 23716 30996
rect 23660 30942 23662 30994
rect 23662 30942 23714 30994
rect 23714 30942 23716 30994
rect 23660 30940 23716 30942
rect 24464 30602 24520 30604
rect 24464 30550 24466 30602
rect 24466 30550 24518 30602
rect 24518 30550 24520 30602
rect 24464 30548 24520 30550
rect 24568 30602 24624 30604
rect 24568 30550 24570 30602
rect 24570 30550 24622 30602
rect 24622 30550 24624 30602
rect 24568 30548 24624 30550
rect 24672 30602 24728 30604
rect 24672 30550 24674 30602
rect 24674 30550 24726 30602
rect 24726 30550 24728 30602
rect 24672 30548 24728 30550
rect 23804 29818 23860 29820
rect 23804 29766 23806 29818
rect 23806 29766 23858 29818
rect 23858 29766 23860 29818
rect 23804 29764 23860 29766
rect 23908 29818 23964 29820
rect 23908 29766 23910 29818
rect 23910 29766 23962 29818
rect 23962 29766 23964 29818
rect 23908 29764 23964 29766
rect 24012 29818 24068 29820
rect 24012 29766 24014 29818
rect 24014 29766 24066 29818
rect 24066 29766 24068 29818
rect 24012 29764 24068 29766
rect 24464 29034 24520 29036
rect 24464 28982 24466 29034
rect 24466 28982 24518 29034
rect 24518 28982 24520 29034
rect 24464 28980 24520 28982
rect 24568 29034 24624 29036
rect 24568 28982 24570 29034
rect 24570 28982 24622 29034
rect 24622 28982 24624 29034
rect 24568 28980 24624 28982
rect 24672 29034 24728 29036
rect 24672 28982 24674 29034
rect 24674 28982 24726 29034
rect 24726 28982 24728 29034
rect 24672 28980 24728 28982
rect 23548 28364 23604 28420
rect 23436 21980 23492 22036
rect 23804 28250 23860 28252
rect 23804 28198 23806 28250
rect 23806 28198 23858 28250
rect 23858 28198 23860 28250
rect 23804 28196 23860 28198
rect 23908 28250 23964 28252
rect 23908 28198 23910 28250
rect 23910 28198 23962 28250
rect 23962 28198 23964 28250
rect 23908 28196 23964 28198
rect 24012 28250 24068 28252
rect 24012 28198 24014 28250
rect 24014 28198 24066 28250
rect 24066 28198 24068 28250
rect 24012 28196 24068 28198
rect 24464 27466 24520 27468
rect 24464 27414 24466 27466
rect 24466 27414 24518 27466
rect 24518 27414 24520 27466
rect 24464 27412 24520 27414
rect 24568 27466 24624 27468
rect 24568 27414 24570 27466
rect 24570 27414 24622 27466
rect 24622 27414 24624 27466
rect 24568 27412 24624 27414
rect 24672 27466 24728 27468
rect 24672 27414 24674 27466
rect 24674 27414 24726 27466
rect 24726 27414 24728 27466
rect 24672 27412 24728 27414
rect 24332 27244 24388 27300
rect 25116 30940 25172 30996
rect 23804 26682 23860 26684
rect 23804 26630 23806 26682
rect 23806 26630 23858 26682
rect 23858 26630 23860 26682
rect 23804 26628 23860 26630
rect 23908 26682 23964 26684
rect 23908 26630 23910 26682
rect 23910 26630 23962 26682
rect 23962 26630 23964 26682
rect 23908 26628 23964 26630
rect 24012 26682 24068 26684
rect 24012 26630 24014 26682
rect 24014 26630 24066 26682
rect 24066 26630 24068 26682
rect 24012 26628 24068 26630
rect 23804 25114 23860 25116
rect 23804 25062 23806 25114
rect 23806 25062 23858 25114
rect 23858 25062 23860 25114
rect 23804 25060 23860 25062
rect 23908 25114 23964 25116
rect 23908 25062 23910 25114
rect 23910 25062 23962 25114
rect 23962 25062 23964 25114
rect 23908 25060 23964 25062
rect 24012 25114 24068 25116
rect 24012 25062 24014 25114
rect 24014 25062 24066 25114
rect 24066 25062 24068 25114
rect 24012 25060 24068 25062
rect 23772 23884 23828 23940
rect 23804 23546 23860 23548
rect 23660 23436 23716 23492
rect 23804 23494 23806 23546
rect 23806 23494 23858 23546
rect 23858 23494 23860 23546
rect 23804 23492 23860 23494
rect 23908 23546 23964 23548
rect 23908 23494 23910 23546
rect 23910 23494 23962 23546
rect 23962 23494 23964 23546
rect 23908 23492 23964 23494
rect 24012 23546 24068 23548
rect 24012 23494 24014 23546
rect 24014 23494 24066 23546
rect 24066 23494 24068 23546
rect 24012 23492 24068 23494
rect 23660 21980 23716 22036
rect 23804 21978 23860 21980
rect 23804 21926 23806 21978
rect 23806 21926 23858 21978
rect 23858 21926 23860 21978
rect 23804 21924 23860 21926
rect 23908 21978 23964 21980
rect 23908 21926 23910 21978
rect 23910 21926 23962 21978
rect 23962 21926 23964 21978
rect 23908 21924 23964 21926
rect 24012 21978 24068 21980
rect 24012 21926 24014 21978
rect 24014 21926 24066 21978
rect 24066 21926 24068 21978
rect 24012 21924 24068 21926
rect 22988 16828 23044 16884
rect 22540 15484 22596 15540
rect 22652 15036 22708 15092
rect 22540 14812 22596 14868
rect 22876 14476 22932 14532
rect 22540 8316 22596 8372
rect 22652 6860 22708 6916
rect 22540 5628 22596 5684
rect 22988 10668 23044 10724
rect 23100 12236 23156 12292
rect 23324 18732 23380 18788
rect 23324 15036 23380 15092
rect 23436 18508 23492 18564
rect 23212 11564 23268 11620
rect 23324 14812 23380 14868
rect 23804 20410 23860 20412
rect 23804 20358 23806 20410
rect 23806 20358 23858 20410
rect 23858 20358 23860 20410
rect 23804 20356 23860 20358
rect 23908 20410 23964 20412
rect 23908 20358 23910 20410
rect 23910 20358 23962 20410
rect 23962 20358 23964 20410
rect 23908 20356 23964 20358
rect 24012 20410 24068 20412
rect 24012 20358 24014 20410
rect 24014 20358 24066 20410
rect 24066 20358 24068 20410
rect 24012 20356 24068 20358
rect 25004 26236 25060 26292
rect 24332 26124 24388 26180
rect 24464 25898 24520 25900
rect 24464 25846 24466 25898
rect 24466 25846 24518 25898
rect 24518 25846 24520 25898
rect 24464 25844 24520 25846
rect 24568 25898 24624 25900
rect 24568 25846 24570 25898
rect 24570 25846 24622 25898
rect 24622 25846 24624 25898
rect 24568 25844 24624 25846
rect 24672 25898 24728 25900
rect 24672 25846 24674 25898
rect 24674 25846 24726 25898
rect 24726 25846 24728 25898
rect 24672 25844 24728 25846
rect 25004 24892 25060 24948
rect 24668 24556 24724 24612
rect 24464 24330 24520 24332
rect 24464 24278 24466 24330
rect 24466 24278 24518 24330
rect 24518 24278 24520 24330
rect 24464 24276 24520 24278
rect 24568 24330 24624 24332
rect 24568 24278 24570 24330
rect 24570 24278 24622 24330
rect 24622 24278 24624 24330
rect 24568 24276 24624 24278
rect 24672 24330 24728 24332
rect 24672 24278 24674 24330
rect 24674 24278 24726 24330
rect 24726 24278 24728 24330
rect 24672 24276 24728 24278
rect 24332 23884 24388 23940
rect 24892 23212 24948 23268
rect 24464 22762 24520 22764
rect 24464 22710 24466 22762
rect 24466 22710 24518 22762
rect 24518 22710 24520 22762
rect 24464 22708 24520 22710
rect 24568 22762 24624 22764
rect 24568 22710 24570 22762
rect 24570 22710 24622 22762
rect 24622 22710 24624 22762
rect 24568 22708 24624 22710
rect 24672 22762 24728 22764
rect 24672 22710 24674 22762
rect 24674 22710 24726 22762
rect 24726 22710 24728 22762
rect 24672 22708 24728 22710
rect 24464 21194 24520 21196
rect 24464 21142 24466 21194
rect 24466 21142 24518 21194
rect 24518 21142 24520 21194
rect 24464 21140 24520 21142
rect 24568 21194 24624 21196
rect 24568 21142 24570 21194
rect 24570 21142 24622 21194
rect 24622 21142 24624 21194
rect 24568 21140 24624 21142
rect 24672 21194 24728 21196
rect 24672 21142 24674 21194
rect 24674 21142 24726 21194
rect 24726 21142 24728 21194
rect 24672 21140 24728 21142
rect 24220 19516 24276 19572
rect 23804 18842 23860 18844
rect 23804 18790 23806 18842
rect 23806 18790 23858 18842
rect 23858 18790 23860 18842
rect 23804 18788 23860 18790
rect 23908 18842 23964 18844
rect 23908 18790 23910 18842
rect 23910 18790 23962 18842
rect 23962 18790 23964 18842
rect 23908 18788 23964 18790
rect 24012 18842 24068 18844
rect 24012 18790 24014 18842
rect 24014 18790 24066 18842
rect 24066 18790 24068 18842
rect 24012 18788 24068 18790
rect 23660 18450 23716 18452
rect 23660 18398 23662 18450
rect 23662 18398 23714 18450
rect 23714 18398 23716 18450
rect 23660 18396 23716 18398
rect 23804 17274 23860 17276
rect 23804 17222 23806 17274
rect 23806 17222 23858 17274
rect 23858 17222 23860 17274
rect 23804 17220 23860 17222
rect 23908 17274 23964 17276
rect 23908 17222 23910 17274
rect 23910 17222 23962 17274
rect 23962 17222 23964 17274
rect 23908 17220 23964 17222
rect 24012 17274 24068 17276
rect 24012 17222 24014 17274
rect 24014 17222 24066 17274
rect 24066 17222 24068 17274
rect 24012 17220 24068 17222
rect 23804 15706 23860 15708
rect 23804 15654 23806 15706
rect 23806 15654 23858 15706
rect 23858 15654 23860 15706
rect 23804 15652 23860 15654
rect 23908 15706 23964 15708
rect 23908 15654 23910 15706
rect 23910 15654 23962 15706
rect 23962 15654 23964 15706
rect 23908 15652 23964 15654
rect 24012 15706 24068 15708
rect 24012 15654 24014 15706
rect 24014 15654 24066 15706
rect 24066 15654 24068 15706
rect 24012 15652 24068 15654
rect 23548 14476 23604 14532
rect 24464 19626 24520 19628
rect 24464 19574 24466 19626
rect 24466 19574 24518 19626
rect 24518 19574 24520 19626
rect 24464 19572 24520 19574
rect 24568 19626 24624 19628
rect 24568 19574 24570 19626
rect 24570 19574 24622 19626
rect 24622 19574 24624 19626
rect 24568 19572 24624 19574
rect 24672 19626 24728 19628
rect 24672 19574 24674 19626
rect 24674 19574 24726 19626
rect 24726 19574 24728 19626
rect 24672 19572 24728 19574
rect 25228 24668 25284 24724
rect 25676 37938 25732 37940
rect 25676 37886 25678 37938
rect 25678 37886 25730 37938
rect 25730 37886 25732 37938
rect 25676 37884 25732 37886
rect 25452 36988 25508 37044
rect 25676 36092 25732 36148
rect 25564 34860 25620 34916
rect 25452 30716 25508 30772
rect 25676 34802 25732 34804
rect 25676 34750 25678 34802
rect 25678 34750 25730 34802
rect 25730 34750 25732 34802
rect 25676 34748 25732 34750
rect 25676 33852 25732 33908
rect 25676 32956 25732 33012
rect 25676 31666 25732 31668
rect 25676 31614 25678 31666
rect 25678 31614 25730 31666
rect 25730 31614 25732 31666
rect 25676 31612 25732 31614
rect 25676 27132 25732 27188
rect 25228 20972 25284 21028
rect 25116 19516 25172 19572
rect 24464 18058 24520 18060
rect 24464 18006 24466 18058
rect 24466 18006 24518 18058
rect 24518 18006 24520 18058
rect 24464 18004 24520 18006
rect 24568 18058 24624 18060
rect 24568 18006 24570 18058
rect 24570 18006 24622 18058
rect 24622 18006 24624 18058
rect 24568 18004 24624 18006
rect 24672 18058 24728 18060
rect 24672 18006 24674 18058
rect 24674 18006 24726 18058
rect 24726 18006 24728 18058
rect 24672 18004 24728 18006
rect 24556 17778 24612 17780
rect 24556 17726 24558 17778
rect 24558 17726 24610 17778
rect 24610 17726 24612 17778
rect 24556 17724 24612 17726
rect 24332 16492 24388 16548
rect 24892 16716 24948 16772
rect 24464 16490 24520 16492
rect 24464 16438 24466 16490
rect 24466 16438 24518 16490
rect 24518 16438 24520 16490
rect 24464 16436 24520 16438
rect 24568 16490 24624 16492
rect 24568 16438 24570 16490
rect 24570 16438 24622 16490
rect 24622 16438 24624 16490
rect 24568 16436 24624 16438
rect 24672 16490 24728 16492
rect 24672 16438 24674 16490
rect 24674 16438 24726 16490
rect 24726 16438 24728 16490
rect 24672 16436 24728 16438
rect 24220 15036 24276 15092
rect 24464 14922 24520 14924
rect 24464 14870 24466 14922
rect 24466 14870 24518 14922
rect 24518 14870 24520 14922
rect 24464 14868 24520 14870
rect 24568 14922 24624 14924
rect 24568 14870 24570 14922
rect 24570 14870 24622 14922
rect 24622 14870 24624 14922
rect 24568 14868 24624 14870
rect 24672 14922 24728 14924
rect 24672 14870 24674 14922
rect 24674 14870 24726 14922
rect 24726 14870 24728 14922
rect 24672 14868 24728 14870
rect 23772 14588 23828 14644
rect 24780 14588 24836 14644
rect 24668 14476 24724 14532
rect 23660 14364 23716 14420
rect 24332 14364 24388 14420
rect 23804 14138 23860 14140
rect 23804 14086 23806 14138
rect 23806 14086 23858 14138
rect 23858 14086 23860 14138
rect 23804 14084 23860 14086
rect 23908 14138 23964 14140
rect 23908 14086 23910 14138
rect 23910 14086 23962 14138
rect 23962 14086 23964 14138
rect 23908 14084 23964 14086
rect 24012 14138 24068 14140
rect 24012 14086 24014 14138
rect 24014 14086 24066 14138
rect 24066 14086 24068 14138
rect 24012 14084 24068 14086
rect 23660 13970 23716 13972
rect 23660 13918 23662 13970
rect 23662 13918 23714 13970
rect 23714 13918 23716 13970
rect 23660 13916 23716 13918
rect 24220 13692 24276 13748
rect 23804 12570 23860 12572
rect 23804 12518 23806 12570
rect 23806 12518 23858 12570
rect 23858 12518 23860 12570
rect 23804 12516 23860 12518
rect 23908 12570 23964 12572
rect 23908 12518 23910 12570
rect 23910 12518 23962 12570
rect 23962 12518 23964 12570
rect 23908 12516 23964 12518
rect 24012 12570 24068 12572
rect 24012 12518 24014 12570
rect 24014 12518 24066 12570
rect 24066 12518 24068 12570
rect 24012 12516 24068 12518
rect 23436 12236 23492 12292
rect 24108 12012 24164 12068
rect 23772 11564 23828 11620
rect 23804 11002 23860 11004
rect 23804 10950 23806 11002
rect 23806 10950 23858 11002
rect 23858 10950 23860 11002
rect 23804 10948 23860 10950
rect 23908 11002 23964 11004
rect 23908 10950 23910 11002
rect 23910 10950 23962 11002
rect 23962 10950 23964 11002
rect 23908 10948 23964 10950
rect 24012 11002 24068 11004
rect 24012 10950 24014 11002
rect 24014 10950 24066 11002
rect 24066 10950 24068 11002
rect 24012 10948 24068 10950
rect 23804 9434 23860 9436
rect 23804 9382 23806 9434
rect 23806 9382 23858 9434
rect 23858 9382 23860 9434
rect 23804 9380 23860 9382
rect 23908 9434 23964 9436
rect 23908 9382 23910 9434
rect 23910 9382 23962 9434
rect 23962 9382 23964 9434
rect 23908 9380 23964 9382
rect 24012 9434 24068 9436
rect 24012 9382 24014 9434
rect 24014 9382 24066 9434
rect 24066 9382 24068 9434
rect 24012 9380 24068 9382
rect 23804 7866 23860 7868
rect 23804 7814 23806 7866
rect 23806 7814 23858 7866
rect 23858 7814 23860 7866
rect 23804 7812 23860 7814
rect 23908 7866 23964 7868
rect 23908 7814 23910 7866
rect 23910 7814 23962 7866
rect 23962 7814 23964 7866
rect 23908 7812 23964 7814
rect 24012 7866 24068 7868
rect 24012 7814 24014 7866
rect 24014 7814 24066 7866
rect 24066 7814 24068 7866
rect 24012 7812 24068 7814
rect 23804 6298 23860 6300
rect 23804 6246 23806 6298
rect 23806 6246 23858 6298
rect 23858 6246 23860 6298
rect 23804 6244 23860 6246
rect 23908 6298 23964 6300
rect 23908 6246 23910 6298
rect 23910 6246 23962 6298
rect 23962 6246 23964 6298
rect 23908 6244 23964 6246
rect 24012 6298 24068 6300
rect 24012 6246 24014 6298
rect 24014 6246 24066 6298
rect 24066 6246 24068 6298
rect 24012 6244 24068 6246
rect 23804 4730 23860 4732
rect 23804 4678 23806 4730
rect 23806 4678 23858 4730
rect 23858 4678 23860 4730
rect 23804 4676 23860 4678
rect 23908 4730 23964 4732
rect 23908 4678 23910 4730
rect 23910 4678 23962 4730
rect 23962 4678 23964 4730
rect 23908 4676 23964 4678
rect 24012 4730 24068 4732
rect 24012 4678 24014 4730
rect 24014 4678 24066 4730
rect 24066 4678 24068 4730
rect 24012 4676 24068 4678
rect 23100 3500 23156 3556
rect 21980 140 22036 196
rect 22204 1932 22260 1988
rect 23804 3162 23860 3164
rect 23804 3110 23806 3162
rect 23806 3110 23858 3162
rect 23858 3110 23860 3162
rect 23804 3108 23860 3110
rect 23908 3162 23964 3164
rect 23908 3110 23910 3162
rect 23910 3110 23962 3162
rect 23962 3110 23964 3162
rect 23908 3108 23964 3110
rect 24012 3162 24068 3164
rect 24012 3110 24014 3162
rect 24014 3110 24066 3162
rect 24066 3110 24068 3162
rect 24012 3108 24068 3110
rect 22652 2492 22708 2548
rect 24780 13804 24836 13860
rect 24464 13354 24520 13356
rect 24464 13302 24466 13354
rect 24466 13302 24518 13354
rect 24518 13302 24520 13354
rect 24464 13300 24520 13302
rect 24568 13354 24624 13356
rect 24568 13302 24570 13354
rect 24570 13302 24622 13354
rect 24622 13302 24624 13354
rect 24568 13300 24624 13302
rect 24672 13354 24728 13356
rect 24672 13302 24674 13354
rect 24674 13302 24726 13354
rect 24726 13302 24728 13354
rect 24672 13300 24728 13302
rect 25004 14588 25060 14644
rect 25116 17612 25172 17668
rect 25676 26236 25732 26292
rect 25676 25282 25732 25284
rect 25676 25230 25678 25282
rect 25678 25230 25730 25282
rect 25730 25230 25732 25282
rect 25676 25228 25732 25230
rect 25676 23996 25732 24052
rect 25676 23100 25732 23156
rect 26236 48130 26292 48132
rect 26236 48078 26238 48130
rect 26238 48078 26290 48130
rect 26290 48078 26292 48130
rect 26236 48076 26292 48078
rect 27244 52220 27300 52276
rect 27132 51324 27188 51380
rect 27244 50876 27300 50932
rect 27020 49980 27076 50036
rect 26236 47458 26292 47460
rect 26236 47406 26238 47458
rect 26238 47406 26290 47458
rect 26290 47406 26292 47458
rect 26236 47404 26292 47406
rect 26236 46562 26292 46564
rect 26236 46510 26238 46562
rect 26238 46510 26290 46562
rect 26290 46510 26292 46562
rect 26236 46508 26292 46510
rect 26236 45890 26292 45892
rect 26236 45838 26238 45890
rect 26238 45838 26290 45890
rect 26290 45838 26292 45890
rect 26236 45836 26292 45838
rect 26236 43426 26292 43428
rect 26236 43374 26238 43426
rect 26238 43374 26290 43426
rect 26290 43374 26292 43426
rect 26236 43372 26292 43374
rect 26348 42924 26404 42980
rect 26236 42754 26292 42756
rect 26236 42702 26238 42754
rect 26238 42702 26290 42754
rect 26290 42702 26292 42754
rect 26236 42700 26292 42702
rect 26236 41858 26292 41860
rect 26236 41806 26238 41858
rect 26238 41806 26290 41858
rect 26290 41806 26292 41858
rect 26236 41804 26292 41806
rect 26236 41186 26292 41188
rect 26236 41134 26238 41186
rect 26238 41134 26290 41186
rect 26290 41134 26292 41186
rect 26236 41132 26292 41134
rect 26124 40908 26180 40964
rect 26236 40460 26292 40516
rect 26236 39618 26292 39620
rect 26236 39566 26238 39618
rect 26238 39566 26290 39618
rect 26290 39566 26292 39618
rect 26236 39564 26292 39566
rect 26236 38722 26292 38724
rect 26236 38670 26238 38722
rect 26238 38670 26290 38722
rect 26290 38670 26292 38722
rect 26236 38668 26292 38670
rect 26236 38050 26292 38052
rect 26236 37998 26238 38050
rect 26238 37998 26290 38050
rect 26290 37998 26292 38050
rect 26236 37996 26292 37998
rect 26236 37154 26292 37156
rect 26236 37102 26238 37154
rect 26238 37102 26290 37154
rect 26290 37102 26292 37154
rect 26236 37100 26292 37102
rect 26012 35980 26068 36036
rect 26012 35532 26068 35588
rect 26236 34914 26292 34916
rect 26236 34862 26238 34914
rect 26238 34862 26290 34914
rect 26290 34862 26292 34914
rect 26236 34860 26292 34862
rect 26460 36316 26516 36372
rect 26572 41356 26628 41412
rect 26348 34636 26404 34692
rect 26348 34300 26404 34356
rect 26236 34018 26292 34020
rect 26236 33966 26238 34018
rect 26238 33966 26290 34018
rect 26290 33966 26292 34018
rect 26236 33964 26292 33966
rect 26236 32620 26292 32676
rect 26124 32396 26180 32452
rect 26236 29484 26292 29540
rect 26236 28642 26292 28644
rect 26236 28590 26238 28642
rect 26238 28590 26290 28642
rect 26290 28590 26292 28642
rect 26236 28588 26292 28590
rect 26124 28476 26180 28532
rect 25900 27692 25956 27748
rect 26236 27746 26292 27748
rect 26236 27694 26238 27746
rect 26238 27694 26290 27746
rect 26290 27694 26292 27746
rect 26236 27692 26292 27694
rect 25900 22876 25956 22932
rect 25676 21756 25732 21812
rect 25788 21698 25844 21700
rect 25788 21646 25790 21698
rect 25790 21646 25842 21698
rect 25842 21646 25844 21698
rect 25788 21644 25844 21646
rect 25564 20860 25620 20916
rect 25452 15820 25508 15876
rect 25340 13746 25396 13748
rect 25340 13694 25342 13746
rect 25342 13694 25394 13746
rect 25394 13694 25396 13746
rect 25340 13692 25396 13694
rect 25004 11900 25060 11956
rect 24464 11786 24520 11788
rect 24464 11734 24466 11786
rect 24466 11734 24518 11786
rect 24518 11734 24520 11786
rect 24464 11732 24520 11734
rect 24568 11786 24624 11788
rect 24568 11734 24570 11786
rect 24570 11734 24622 11786
rect 24622 11734 24624 11786
rect 24568 11732 24624 11734
rect 24672 11786 24728 11788
rect 24672 11734 24674 11786
rect 24674 11734 24726 11786
rect 24726 11734 24728 11786
rect 24672 11732 24728 11734
rect 25116 10444 25172 10500
rect 24464 10218 24520 10220
rect 24464 10166 24466 10218
rect 24466 10166 24518 10218
rect 24518 10166 24520 10218
rect 24464 10164 24520 10166
rect 24568 10218 24624 10220
rect 24568 10166 24570 10218
rect 24570 10166 24622 10218
rect 24622 10166 24624 10218
rect 24568 10164 24624 10166
rect 24672 10218 24728 10220
rect 24672 10166 24674 10218
rect 24674 10166 24726 10218
rect 24726 10166 24728 10218
rect 24672 10164 24728 10166
rect 25564 9212 25620 9268
rect 24464 8650 24520 8652
rect 24464 8598 24466 8650
rect 24466 8598 24518 8650
rect 24518 8598 24520 8650
rect 24464 8596 24520 8598
rect 24568 8650 24624 8652
rect 24568 8598 24570 8650
rect 24570 8598 24622 8650
rect 24622 8598 24624 8650
rect 24568 8596 24624 8598
rect 24672 8650 24728 8652
rect 24672 8598 24674 8650
rect 24674 8598 24726 8650
rect 24726 8598 24728 8650
rect 24672 8596 24728 8598
rect 24464 7082 24520 7084
rect 24464 7030 24466 7082
rect 24466 7030 24518 7082
rect 24518 7030 24520 7082
rect 24464 7028 24520 7030
rect 24568 7082 24624 7084
rect 24568 7030 24570 7082
rect 24570 7030 24622 7082
rect 24622 7030 24624 7082
rect 24568 7028 24624 7030
rect 24672 7082 24728 7084
rect 24672 7030 24674 7082
rect 24674 7030 24726 7082
rect 24726 7030 24728 7082
rect 24672 7028 24728 7030
rect 24464 5514 24520 5516
rect 24464 5462 24466 5514
rect 24466 5462 24518 5514
rect 24518 5462 24520 5514
rect 24464 5460 24520 5462
rect 24568 5514 24624 5516
rect 24568 5462 24570 5514
rect 24570 5462 24622 5514
rect 24622 5462 24624 5514
rect 24568 5460 24624 5462
rect 24672 5514 24728 5516
rect 24672 5462 24674 5514
rect 24674 5462 24726 5514
rect 24726 5462 24728 5514
rect 24672 5460 24728 5462
rect 24464 3946 24520 3948
rect 24464 3894 24466 3946
rect 24466 3894 24518 3946
rect 24518 3894 24520 3946
rect 24464 3892 24520 3894
rect 24568 3946 24624 3948
rect 24568 3894 24570 3946
rect 24570 3894 24622 3946
rect 24622 3894 24624 3946
rect 24568 3892 24624 3894
rect 24672 3946 24728 3948
rect 24672 3894 24674 3946
rect 24674 3894 24726 3946
rect 24726 3894 24728 3946
rect 24672 3892 24728 3894
rect 24464 2378 24520 2380
rect 24464 2326 24466 2378
rect 24466 2326 24518 2378
rect 24518 2326 24520 2378
rect 24464 2324 24520 2326
rect 24568 2378 24624 2380
rect 24568 2326 24570 2378
rect 24570 2326 24622 2378
rect 24622 2326 24624 2378
rect 24568 2324 24624 2326
rect 24672 2378 24728 2380
rect 24672 2326 24674 2378
rect 24674 2326 24726 2378
rect 24726 2326 24728 2378
rect 24672 2324 24728 2326
rect 24332 2044 24388 2100
rect 23804 1594 23860 1596
rect 23804 1542 23806 1594
rect 23806 1542 23858 1594
rect 23858 1542 23860 1594
rect 23804 1540 23860 1542
rect 23908 1594 23964 1596
rect 23908 1542 23910 1594
rect 23910 1542 23962 1594
rect 23962 1542 23964 1594
rect 23908 1540 23964 1542
rect 24012 1594 24068 1596
rect 24012 1542 24014 1594
rect 24014 1542 24066 1594
rect 24066 1542 24068 1594
rect 24012 1540 24068 1542
rect 24892 1596 24948 1652
rect 22540 1372 22596 1428
rect 24464 810 24520 812
rect 24464 758 24466 810
rect 24466 758 24518 810
rect 24518 758 24520 810
rect 24464 756 24520 758
rect 24568 810 24624 812
rect 24568 758 24570 810
rect 24570 758 24622 810
rect 24622 758 24624 810
rect 24568 756 24624 758
rect 24672 810 24728 812
rect 24672 758 24674 810
rect 24674 758 24726 810
rect 24726 758 24728 810
rect 24672 756 24728 758
rect 23548 476 23604 532
rect 25788 20524 25844 20580
rect 25900 19458 25956 19460
rect 25900 19406 25902 19458
rect 25902 19406 25954 19458
rect 25954 19406 25956 19458
rect 25900 19404 25956 19406
rect 25788 6412 25844 6468
rect 26236 27074 26292 27076
rect 26236 27022 26238 27074
rect 26238 27022 26290 27074
rect 26290 27022 26292 27074
rect 26236 27020 26292 27022
rect 26236 25676 26292 25732
rect 26236 25506 26292 25508
rect 26236 25454 26238 25506
rect 26238 25454 26290 25506
rect 26290 25454 26292 25506
rect 26236 25452 26292 25454
rect 26236 24444 26292 24500
rect 26236 23660 26292 23716
rect 26236 23042 26292 23044
rect 26236 22990 26238 23042
rect 26238 22990 26290 23042
rect 26290 22990 26292 23042
rect 26236 22988 26292 22990
rect 26236 22540 26292 22596
rect 26236 21474 26292 21476
rect 26236 21422 26238 21474
rect 26238 21422 26290 21474
rect 26290 21422 26292 21474
rect 26236 21420 26292 21422
rect 26348 20524 26404 20580
rect 26460 19346 26516 19348
rect 26460 19294 26462 19346
rect 26462 19294 26514 19346
rect 26514 19294 26516 19346
rect 26460 19292 26516 19294
rect 26348 11452 26404 11508
rect 26124 7644 26180 7700
rect 26012 5852 26068 5908
rect 26572 6636 26628 6692
rect 27244 49084 27300 49140
rect 27132 48188 27188 48244
rect 27244 47740 27300 47796
rect 27020 46844 27076 46900
rect 27244 45948 27300 46004
rect 27132 45052 27188 45108
rect 27244 44604 27300 44660
rect 27020 43708 27076 43764
rect 27244 42812 27300 42868
rect 27132 41916 27188 41972
rect 27244 41468 27300 41524
rect 27020 40572 27076 40628
rect 27244 39676 27300 39732
rect 27132 38780 27188 38836
rect 27244 38332 27300 38388
rect 27020 37436 27076 37492
rect 27244 36540 27300 36596
rect 27132 35644 27188 35700
rect 27244 35196 27300 35252
rect 27020 34300 27076 34356
rect 27244 33404 27300 33460
rect 27132 32508 27188 32564
rect 27244 32060 27300 32116
rect 28364 32284 28420 32340
rect 27020 31164 27076 31220
rect 27244 30268 27300 30324
rect 27020 29820 27076 29876
rect 28140 29596 28196 29652
rect 27132 29372 27188 29428
rect 27244 28924 27300 28980
rect 27244 28530 27300 28532
rect 27244 28478 27246 28530
rect 27246 28478 27298 28530
rect 27298 28478 27300 28530
rect 27244 28476 27300 28478
rect 27244 28082 27300 28084
rect 27244 28030 27246 28082
rect 27246 28030 27298 28082
rect 27298 28030 27300 28082
rect 27244 28028 27300 28030
rect 27020 27580 27076 27636
rect 27244 26684 27300 26740
rect 27244 25788 27300 25844
rect 27132 25340 27188 25396
rect 27244 24444 27300 24500
rect 27244 23548 27300 23604
rect 27244 22652 27300 22708
rect 27132 22204 27188 22260
rect 27356 20914 27412 20916
rect 27356 20862 27358 20914
rect 27358 20862 27410 20914
rect 27410 20862 27412 20914
rect 27356 20860 27412 20862
rect 28140 20860 28196 20916
rect 26684 5740 26740 5796
rect 28364 19964 28420 20020
rect 27020 4396 27076 4452
rect 27580 5068 27636 5124
rect 27468 2156 27524 2212
rect 25676 924 25732 980
rect 26012 588 26068 644
rect 26236 1708 26292 1764
rect 26908 364 26964 420
<< metal3 >>
rect 19506 57260 19516 57316
rect 19572 57260 19852 57316
rect 19908 57260 19918 57316
rect 25890 57260 25900 57316
rect 25956 57260 26236 57316
rect 26292 57260 26302 57316
rect 28448 57204 28560 57232
rect 24322 57148 24332 57204
rect 24388 57148 28560 57204
rect 28448 57120 28560 57148
rect 28448 56756 28560 56784
rect 24210 56700 24220 56756
rect 24276 56700 28560 56756
rect 28448 56672 28560 56700
rect 21634 56588 21644 56644
rect 21700 56588 27580 56644
rect 27636 56588 27646 56644
rect 3794 56420 3804 56476
rect 3860 56420 3908 56476
rect 3964 56420 4012 56476
rect 4068 56420 4078 56476
rect 23794 56420 23804 56476
rect 23860 56420 23908 56476
rect 23964 56420 24012 56476
rect 24068 56420 24078 56476
rect 28448 56308 28560 56336
rect 15474 56252 15484 56308
rect 15540 56252 16492 56308
rect 16548 56252 16558 56308
rect 20850 56252 20860 56308
rect 20916 56252 22204 56308
rect 22260 56252 22270 56308
rect 23538 56252 23548 56308
rect 23604 56252 24444 56308
rect 24500 56252 24510 56308
rect 24882 56252 24892 56308
rect 24948 56252 26012 56308
rect 26068 56252 26078 56308
rect 27132 56252 28560 56308
rect 27132 56196 27188 56252
rect 28448 56224 28560 56252
rect 25778 56140 25788 56196
rect 25844 56140 27188 56196
rect 6178 55916 6188 55972
rect 6244 55916 9212 55972
rect 9268 55916 9278 55972
rect 19478 55916 19516 55972
rect 19572 55916 19582 55972
rect 21270 55916 21308 55972
rect 21364 55916 21374 55972
rect 23538 55916 23548 55972
rect 23604 55916 25452 55972
rect 25508 55916 25518 55972
rect 28448 55860 28560 55888
rect 22530 55804 22540 55860
rect 22596 55804 28560 55860
rect 28448 55776 28560 55804
rect 14018 55692 14028 55748
rect 14084 55692 19516 55748
rect 19572 55692 19582 55748
rect 21858 55692 21868 55748
rect 21924 55692 23884 55748
rect 23940 55692 23950 55748
rect 4454 55636 4464 55692
rect 4520 55636 4568 55692
rect 4624 55636 4672 55692
rect 4728 55636 4738 55692
rect 24454 55636 24464 55692
rect 24520 55636 24568 55692
rect 24624 55636 24672 55692
rect 24728 55636 24738 55692
rect 28448 55412 28560 55440
rect 24994 55356 25004 55412
rect 25060 55356 28560 55412
rect 28448 55328 28560 55356
rect 2818 55244 2828 55300
rect 2884 55244 6300 55300
rect 6356 55244 6366 55300
rect 18274 55244 18284 55300
rect 18340 55244 20524 55300
rect 20580 55244 20590 55300
rect 20822 55244 20860 55300
rect 20916 55244 20926 55300
rect 22390 55244 22428 55300
rect 22484 55244 22494 55300
rect 23314 55244 23324 55300
rect 23380 55244 24668 55300
rect 24724 55244 24734 55300
rect 0 55188 112 55216
rect 0 55132 3164 55188
rect 3220 55132 3230 55188
rect 6066 55132 6076 55188
rect 6132 55132 6860 55188
rect 6916 55132 6926 55188
rect 11442 55132 11452 55188
rect 11508 55132 11900 55188
rect 11956 55132 11966 55188
rect 20066 55132 20076 55188
rect 20132 55132 27020 55188
rect 27076 55132 27086 55188
rect 0 55104 112 55132
rect 28448 54964 28560 54992
rect 26124 54908 28560 54964
rect 3794 54852 3804 54908
rect 3860 54852 3908 54908
rect 3964 54852 4012 54908
rect 4068 54852 4078 54908
rect 23794 54852 23804 54908
rect 23860 54852 23908 54908
rect 23964 54852 24012 54908
rect 24068 54852 24078 54908
rect 26124 54740 26180 54908
rect 28448 54880 28560 54908
rect 23762 54684 23772 54740
rect 23828 54684 26180 54740
rect 23650 54572 23660 54628
rect 23716 54572 24332 54628
rect 24388 54572 24398 54628
rect 28448 54516 28560 54544
rect 11554 54460 11564 54516
rect 11620 54460 21196 54516
rect 21252 54460 21262 54516
rect 25666 54460 25676 54516
rect 25732 54460 28560 54516
rect 28448 54432 28560 54460
rect 23762 54348 23772 54404
rect 23828 54348 25004 54404
rect 25060 54348 25070 54404
rect 0 54292 112 54320
rect 0 54236 5964 54292
rect 6020 54236 6030 54292
rect 19030 54236 19068 54292
rect 19124 54236 19134 54292
rect 20132 54236 24668 54292
rect 24724 54236 24734 54292
rect 0 54208 112 54236
rect 20132 54180 20188 54236
rect 17714 54124 17724 54180
rect 17780 54124 20188 54180
rect 20514 54124 20524 54180
rect 20580 54124 24108 54180
rect 24164 54124 24174 54180
rect 4454 54068 4464 54124
rect 4520 54068 4568 54124
rect 4624 54068 4672 54124
rect 4728 54068 4738 54124
rect 24454 54068 24464 54124
rect 24520 54068 24568 54124
rect 24624 54068 24672 54124
rect 24728 54068 24738 54124
rect 28448 54068 28560 54096
rect 6738 54012 6748 54068
rect 6804 54012 21532 54068
rect 21588 54012 21598 54068
rect 27234 54012 27244 54068
rect 27300 54012 28560 54068
rect 28448 53984 28560 54012
rect 20066 53900 20076 53956
rect 20132 53900 26236 53956
rect 26292 53900 26302 53956
rect 1362 53788 1372 53844
rect 1428 53788 10220 53844
rect 10276 53788 10286 53844
rect 17938 53788 17948 53844
rect 18004 53788 20636 53844
rect 20692 53788 20702 53844
rect 16706 53676 16716 53732
rect 16772 53676 22316 53732
rect 22372 53676 22382 53732
rect 28448 53620 28560 53648
rect 16818 53564 16828 53620
rect 16884 53564 24668 53620
rect 24724 53564 24734 53620
rect 25666 53564 25676 53620
rect 25732 53564 28560 53620
rect 28448 53536 28560 53564
rect 15026 53452 15036 53508
rect 15092 53452 26236 53508
rect 26292 53452 26302 53508
rect 0 53396 112 53424
rect 0 53340 2044 53396
rect 2100 53340 2110 53396
rect 0 53312 112 53340
rect 3794 53284 3804 53340
rect 3860 53284 3908 53340
rect 3964 53284 4012 53340
rect 4068 53284 4078 53340
rect 23794 53284 23804 53340
rect 23860 53284 23908 53340
rect 23964 53284 24012 53340
rect 24068 53284 24078 53340
rect 28448 53172 28560 53200
rect 27010 53116 27020 53172
rect 27076 53116 28560 53172
rect 28448 53088 28560 53116
rect 20066 52780 20076 52836
rect 20132 52780 26236 52836
rect 26292 52780 26302 52836
rect 28448 52724 28560 52752
rect 12562 52668 12572 52724
rect 12628 52668 24668 52724
rect 24724 52668 24734 52724
rect 25442 52668 25452 52724
rect 25508 52668 28560 52724
rect 28448 52640 28560 52668
rect 10882 52556 10892 52612
rect 10948 52556 23100 52612
rect 23156 52556 23166 52612
rect 0 52500 112 52528
rect 4454 52500 4464 52556
rect 4520 52500 4568 52556
rect 4624 52500 4672 52556
rect 4728 52500 4738 52556
rect 24454 52500 24464 52556
rect 24520 52500 24568 52556
rect 24624 52500 24672 52556
rect 24728 52500 24738 52556
rect 0 52444 1484 52500
rect 1540 52444 1550 52500
rect 21410 52444 21420 52500
rect 21476 52444 24388 52500
rect 0 52416 112 52444
rect 24332 52388 24388 52444
rect 14130 52332 14140 52388
rect 14196 52332 22764 52388
rect 22820 52332 22830 52388
rect 24332 52332 27132 52388
rect 27188 52332 27198 52388
rect 28448 52276 28560 52304
rect 21634 52220 21644 52276
rect 21700 52220 24668 52276
rect 24724 52220 24734 52276
rect 27234 52220 27244 52276
rect 27300 52220 28560 52276
rect 28448 52192 28560 52220
rect 22726 52108 22764 52164
rect 22820 52108 22830 52164
rect 28448 51828 28560 51856
rect 25666 51772 25676 51828
rect 25732 51772 28560 51828
rect 3794 51716 3804 51772
rect 3860 51716 3908 51772
rect 3964 51716 4012 51772
rect 4068 51716 4078 51772
rect 23794 51716 23804 51772
rect 23860 51716 23908 51772
rect 23964 51716 24012 51772
rect 24068 51716 24078 51772
rect 28448 51744 28560 51772
rect 0 51604 112 51632
rect 0 51548 13692 51604
rect 13748 51548 13758 51604
rect 0 51520 112 51548
rect 9202 51436 9212 51492
rect 9268 51436 26460 51492
rect 26516 51436 26526 51492
rect 28448 51380 28560 51408
rect 27122 51324 27132 51380
rect 27188 51324 28560 51380
rect 28448 51296 28560 51324
rect 11330 51212 11340 51268
rect 11396 51212 24668 51268
rect 24724 51212 24734 51268
rect 4454 50932 4464 50988
rect 4520 50932 4568 50988
rect 4624 50932 4672 50988
rect 4728 50932 4738 50988
rect 24454 50932 24464 50988
rect 24520 50932 24568 50988
rect 24624 50932 24672 50988
rect 24728 50932 24738 50988
rect 28448 50932 28560 50960
rect 27234 50876 27244 50932
rect 27300 50876 28560 50932
rect 28448 50848 28560 50876
rect 0 50708 112 50736
rect 0 50652 10780 50708
rect 10836 50652 10846 50708
rect 0 50624 112 50652
rect 23986 50540 23996 50596
rect 24052 50540 26908 50596
rect 26964 50540 26974 50596
rect 28448 50484 28560 50512
rect 6850 50428 6860 50484
rect 6916 50428 24668 50484
rect 24724 50428 24734 50484
rect 25666 50428 25676 50484
rect 25732 50428 28560 50484
rect 28448 50400 28560 50428
rect 3794 50148 3804 50204
rect 3860 50148 3908 50204
rect 3964 50148 4012 50204
rect 4068 50148 4078 50204
rect 23794 50148 23804 50204
rect 23860 50148 23908 50204
rect 23964 50148 24012 50204
rect 24068 50148 24078 50204
rect 28448 50036 28560 50064
rect 27010 49980 27020 50036
rect 27076 49980 28560 50036
rect 28448 49952 28560 49980
rect 6178 49868 6188 49924
rect 6244 49868 26236 49924
rect 26292 49868 26302 49924
rect 0 49812 112 49840
rect 0 49756 5292 49812
rect 5348 49756 5358 49812
rect 0 49728 112 49756
rect 14242 49644 14252 49700
rect 14308 49644 24668 49700
rect 24724 49644 24734 49700
rect 28448 49588 28560 49616
rect 25666 49532 25676 49588
rect 25732 49532 28560 49588
rect 28448 49504 28560 49532
rect 4454 49364 4464 49420
rect 4520 49364 4568 49420
rect 4624 49364 4672 49420
rect 4728 49364 4738 49420
rect 24454 49364 24464 49420
rect 24520 49364 24568 49420
rect 24624 49364 24672 49420
rect 24728 49364 24738 49420
rect 28448 49140 28560 49168
rect 27234 49084 27244 49140
rect 27300 49084 28560 49140
rect 28448 49056 28560 49084
rect 2370 48972 2380 49028
rect 2436 48972 24668 49028
rect 24724 48972 24734 49028
rect 0 48916 112 48944
rect 0 48860 2940 48916
rect 2996 48860 3006 48916
rect 0 48832 112 48860
rect 28448 48692 28560 48720
rect 25666 48636 25676 48692
rect 25732 48636 28560 48692
rect 3794 48580 3804 48636
rect 3860 48580 3908 48636
rect 3964 48580 4012 48636
rect 4068 48580 4078 48636
rect 23794 48580 23804 48636
rect 23860 48580 23908 48636
rect 23964 48580 24012 48636
rect 24068 48580 24078 48636
rect 28448 48608 28560 48636
rect 28448 48244 28560 48272
rect 27122 48188 27132 48244
rect 27188 48188 28560 48244
rect 28448 48160 28560 48188
rect 15922 48076 15932 48132
rect 15988 48076 26236 48132
rect 26292 48076 26302 48132
rect 0 48020 112 48048
rect 0 47964 11228 48020
rect 11284 47964 11294 48020
rect 0 47936 112 47964
rect 4454 47796 4464 47852
rect 4520 47796 4568 47852
rect 4624 47796 4672 47852
rect 4728 47796 4738 47852
rect 24454 47796 24464 47852
rect 24520 47796 24568 47852
rect 24624 47796 24672 47852
rect 24728 47796 24738 47852
rect 28448 47796 28560 47824
rect 27234 47740 27244 47796
rect 27300 47740 28560 47796
rect 28448 47712 28560 47740
rect 19730 47404 19740 47460
rect 19796 47404 26236 47460
rect 26292 47404 26302 47460
rect 28448 47348 28560 47376
rect 11890 47292 11900 47348
rect 11956 47292 24668 47348
rect 24724 47292 24734 47348
rect 25666 47292 25676 47348
rect 25732 47292 28560 47348
rect 28448 47264 28560 47292
rect 1036 47180 7644 47236
rect 7700 47180 7710 47236
rect 0 47124 112 47152
rect 1036 47124 1092 47180
rect 0 47068 1092 47124
rect 0 47040 112 47068
rect 3794 47012 3804 47068
rect 3860 47012 3908 47068
rect 3964 47012 4012 47068
rect 4068 47012 4078 47068
rect 23794 47012 23804 47068
rect 23860 47012 23908 47068
rect 23964 47012 24012 47068
rect 24068 47012 24078 47068
rect 28448 46900 28560 46928
rect 27010 46844 27020 46900
rect 27076 46844 28560 46900
rect 28448 46816 28560 46844
rect 3042 46732 3052 46788
rect 3108 46732 25900 46788
rect 25956 46732 25966 46788
rect 16930 46508 16940 46564
rect 16996 46508 26236 46564
rect 26292 46508 26302 46564
rect 28448 46452 28560 46480
rect 25666 46396 25676 46452
rect 25732 46396 28560 46452
rect 28448 46368 28560 46396
rect 0 46228 112 46256
rect 4454 46228 4464 46284
rect 4520 46228 4568 46284
rect 4624 46228 4672 46284
rect 4728 46228 4738 46284
rect 24454 46228 24464 46284
rect 24520 46228 24568 46284
rect 24624 46228 24672 46284
rect 24728 46228 24738 46284
rect 0 46172 3388 46228
rect 0 46144 112 46172
rect 3332 46116 3388 46172
rect 3332 46060 8540 46116
rect 8596 46060 8606 46116
rect 28448 46004 28560 46032
rect 27234 45948 27244 46004
rect 27300 45948 28560 46004
rect 28448 45920 28560 45948
rect 12338 45836 12348 45892
rect 12404 45836 26236 45892
rect 26292 45836 26302 45892
rect 28448 45556 28560 45584
rect 25666 45500 25676 45556
rect 25732 45500 28560 45556
rect 3794 45444 3804 45500
rect 3860 45444 3908 45500
rect 3964 45444 4012 45500
rect 4068 45444 4078 45500
rect 23794 45444 23804 45500
rect 23860 45444 23908 45500
rect 23964 45444 24012 45500
rect 24068 45444 24078 45500
rect 28448 45472 28560 45500
rect 0 45332 112 45360
rect 0 45276 8764 45332
rect 8820 45276 8830 45332
rect 0 45248 112 45276
rect 1586 45164 1596 45220
rect 1652 45164 6860 45220
rect 6916 45164 6926 45220
rect 28448 45108 28560 45136
rect 27122 45052 27132 45108
rect 27188 45052 28560 45108
rect 28448 45024 28560 45052
rect 4454 44660 4464 44716
rect 4520 44660 4568 44716
rect 4624 44660 4672 44716
rect 4728 44660 4738 44716
rect 24454 44660 24464 44716
rect 24520 44660 24568 44716
rect 24624 44660 24672 44716
rect 24728 44660 24738 44716
rect 28448 44660 28560 44688
rect 27234 44604 27244 44660
rect 27300 44604 28560 44660
rect 28448 44576 28560 44604
rect 15698 44492 15708 44548
rect 15764 44492 24892 44548
rect 24948 44492 24958 44548
rect 0 44436 112 44464
rect 0 44380 17724 44436
rect 17780 44380 17790 44436
rect 0 44352 112 44380
rect 28448 44212 28560 44240
rect 25666 44156 25676 44212
rect 25732 44156 28560 44212
rect 28448 44128 28560 44156
rect 3794 43876 3804 43932
rect 3860 43876 3908 43932
rect 3964 43876 4012 43932
rect 4068 43876 4078 43932
rect 23794 43876 23804 43932
rect 23860 43876 23908 43932
rect 23964 43876 24012 43932
rect 24068 43876 24078 43932
rect 28448 43764 28560 43792
rect 27010 43708 27020 43764
rect 27076 43708 28560 43764
rect 28448 43680 28560 43708
rect 0 43540 112 43568
rect 0 43484 19180 43540
rect 19236 43484 19246 43540
rect 0 43456 112 43484
rect 14018 43372 14028 43428
rect 14084 43372 26236 43428
rect 26292 43372 26302 43428
rect 28448 43316 28560 43344
rect 25666 43260 25676 43316
rect 25732 43260 28560 43316
rect 28448 43232 28560 43260
rect 4454 43092 4464 43148
rect 4520 43092 4568 43148
rect 4624 43092 4672 43148
rect 4728 43092 4738 43148
rect 24454 43092 24464 43148
rect 24520 43092 24568 43148
rect 24624 43092 24672 43148
rect 24728 43092 24738 43148
rect 17266 42924 17276 42980
rect 17332 42924 26348 42980
rect 26404 42924 26414 42980
rect 28448 42868 28560 42896
rect 27234 42812 27244 42868
rect 27300 42812 28560 42868
rect 28448 42784 28560 42812
rect 8306 42700 8316 42756
rect 8372 42700 26236 42756
rect 26292 42700 26302 42756
rect 0 42644 112 42672
rect 0 42588 1932 42644
rect 1988 42588 1998 42644
rect 0 42560 112 42588
rect 28448 42420 28560 42448
rect 25666 42364 25676 42420
rect 25732 42364 28560 42420
rect 3794 42308 3804 42364
rect 3860 42308 3908 42364
rect 3964 42308 4012 42364
rect 4068 42308 4078 42364
rect 23794 42308 23804 42364
rect 23860 42308 23908 42364
rect 23964 42308 24012 42364
rect 24068 42308 24078 42364
rect 28448 42336 28560 42364
rect 5394 42028 5404 42084
rect 5460 42028 14252 42084
rect 14308 42028 14318 42084
rect 28448 41972 28560 42000
rect 18274 41916 18284 41972
rect 18340 41916 24332 41972
rect 24388 41916 24398 41972
rect 27122 41916 27132 41972
rect 27188 41916 28560 41972
rect 28448 41888 28560 41916
rect 17042 41804 17052 41860
rect 17108 41804 26236 41860
rect 26292 41804 26302 41860
rect 0 41748 112 41776
rect 0 41692 588 41748
rect 644 41692 654 41748
rect 9874 41692 9884 41748
rect 9940 41692 24668 41748
rect 24724 41692 24734 41748
rect 0 41664 112 41692
rect 6402 41580 6412 41636
rect 6468 41580 10892 41636
rect 10948 41580 10958 41636
rect 4454 41524 4464 41580
rect 4520 41524 4568 41580
rect 4624 41524 4672 41580
rect 4728 41524 4738 41580
rect 24454 41524 24464 41580
rect 24520 41524 24568 41580
rect 24624 41524 24672 41580
rect 24728 41524 24738 41580
rect 28448 41524 28560 41552
rect 27234 41468 27244 41524
rect 27300 41468 28560 41524
rect 28448 41440 28560 41468
rect 15586 41356 15596 41412
rect 15652 41356 26572 41412
rect 26628 41356 26638 41412
rect 9986 41244 9996 41300
rect 10052 41244 27244 41300
rect 27300 41244 27310 41300
rect 9202 41132 9212 41188
rect 9268 41132 19852 41188
rect 19908 41132 19918 41188
rect 20132 41132 26236 41188
rect 26292 41132 26302 41188
rect 20132 41076 20188 41132
rect 28448 41076 28560 41104
rect 9762 41020 9772 41076
rect 9828 41020 20188 41076
rect 25666 41020 25676 41076
rect 25732 41020 28560 41076
rect 28448 40992 28560 41020
rect 914 40908 924 40964
rect 980 40908 11788 40964
rect 11844 40908 11854 40964
rect 12124 40908 13804 40964
rect 13860 40908 14476 40964
rect 14532 40908 14542 40964
rect 20132 40908 20972 40964
rect 21028 40908 21038 40964
rect 25778 40908 25788 40964
rect 25844 40908 26124 40964
rect 26180 40908 26190 40964
rect 0 40852 112 40880
rect 12124 40852 12180 40908
rect 20132 40852 20188 40908
rect 0 40796 1820 40852
rect 1876 40796 1886 40852
rect 7746 40796 7756 40852
rect 7812 40796 12124 40852
rect 12180 40796 12190 40852
rect 12898 40796 12908 40852
rect 12964 40796 20188 40852
rect 0 40768 112 40796
rect 3794 40740 3804 40796
rect 3860 40740 3908 40796
rect 3964 40740 4012 40796
rect 4068 40740 4078 40796
rect 23794 40740 23804 40796
rect 23860 40740 23908 40796
rect 23964 40740 24012 40796
rect 24068 40740 24078 40796
rect 28448 40628 28560 40656
rect 27010 40572 27020 40628
rect 27076 40572 28560 40628
rect 28448 40544 28560 40572
rect 3154 40460 3164 40516
rect 3220 40460 26236 40516
rect 26292 40460 26302 40516
rect 21746 40348 21756 40404
rect 21812 40348 24668 40404
rect 24724 40348 24734 40404
rect 2930 40236 2940 40292
rect 2996 40236 9100 40292
rect 9156 40236 9166 40292
rect 10098 40236 10108 40292
rect 10164 40236 10892 40292
rect 10948 40236 10958 40292
rect 28448 40180 28560 40208
rect 1922 40124 1932 40180
rect 1988 40124 2604 40180
rect 2660 40124 2670 40180
rect 5170 40124 5180 40180
rect 5236 40124 6076 40180
rect 6132 40124 7980 40180
rect 8036 40124 8046 40180
rect 13458 40124 13468 40180
rect 13524 40124 14924 40180
rect 14980 40124 14990 40180
rect 18386 40124 18396 40180
rect 18452 40124 24780 40180
rect 24836 40124 24846 40180
rect 25666 40124 25676 40180
rect 25732 40124 28560 40180
rect 28448 40096 28560 40124
rect 0 39956 112 39984
rect 4454 39956 4464 40012
rect 4520 39956 4568 40012
rect 4624 39956 4672 40012
rect 4728 39956 4738 40012
rect 24454 39956 24464 40012
rect 24520 39956 24568 40012
rect 24624 39956 24672 40012
rect 24728 39956 24738 40012
rect 0 39900 2156 39956
rect 2212 39900 2222 39956
rect 0 39872 112 39900
rect 2706 39788 2716 39844
rect 2772 39788 4172 39844
rect 4228 39788 4238 39844
rect 20132 39788 24892 39844
rect 24948 39788 24958 39844
rect 20132 39732 20188 39788
rect 28448 39732 28560 39760
rect 3490 39676 3500 39732
rect 3556 39676 7308 39732
rect 7364 39676 7374 39732
rect 9314 39676 9324 39732
rect 9380 39676 20188 39732
rect 27234 39676 27244 39732
rect 27300 39676 28560 39732
rect 28448 39648 28560 39676
rect 242 39564 252 39620
rect 308 39564 3836 39620
rect 3892 39564 3902 39620
rect 4162 39564 4172 39620
rect 4228 39564 13468 39620
rect 13524 39564 13534 39620
rect 17602 39564 17612 39620
rect 17668 39564 26236 39620
rect 26292 39564 26302 39620
rect 6626 39452 6636 39508
rect 6692 39452 10444 39508
rect 10500 39452 10510 39508
rect 28448 39284 28560 39312
rect 9202 39228 9212 39284
rect 9268 39228 9884 39284
rect 9940 39228 9950 39284
rect 10434 39228 10444 39284
rect 10500 39228 17052 39284
rect 17108 39228 17118 39284
rect 25666 39228 25676 39284
rect 25732 39228 28560 39284
rect 3794 39172 3804 39228
rect 3860 39172 3908 39228
rect 3964 39172 4012 39228
rect 4068 39172 4078 39228
rect 23794 39172 23804 39228
rect 23860 39172 23908 39228
rect 23964 39172 24012 39228
rect 24068 39172 24078 39228
rect 28448 39200 28560 39228
rect 7746 39116 7756 39172
rect 7812 39116 8316 39172
rect 8372 39116 10108 39172
rect 10164 39116 13580 39172
rect 13636 39116 13646 39172
rect 0 39060 112 39088
rect 0 39004 1708 39060
rect 1764 39004 1774 39060
rect 6850 39004 6860 39060
rect 6916 39004 8876 39060
rect 8932 39004 15596 39060
rect 15652 39004 15662 39060
rect 0 38976 112 39004
rect 3490 38892 3500 38948
rect 3556 38892 5068 38948
rect 5124 38892 6636 38948
rect 6692 38892 6702 38948
rect 11778 38892 11788 38948
rect 11844 38892 14364 38948
rect 14420 38892 14430 38948
rect 28448 38836 28560 38864
rect 2594 38780 2604 38836
rect 2660 38780 5852 38836
rect 5908 38780 5918 38836
rect 9874 38780 9884 38836
rect 9940 38780 11004 38836
rect 11060 38780 11070 38836
rect 12114 38780 12124 38836
rect 12180 38780 14252 38836
rect 14308 38780 14318 38836
rect 27122 38780 27132 38836
rect 27188 38780 28560 38836
rect 28448 38752 28560 38780
rect 5282 38668 5292 38724
rect 5348 38668 6860 38724
rect 6916 38668 6926 38724
rect 8204 38668 13132 38724
rect 13188 38668 13198 38724
rect 13346 38668 13356 38724
rect 13412 38668 13804 38724
rect 13860 38668 13870 38724
rect 25330 38668 25340 38724
rect 25396 38668 26236 38724
rect 26292 38668 26302 38724
rect 8204 38612 8260 38668
rect 578 38556 588 38612
rect 644 38556 1148 38612
rect 1204 38556 1214 38612
rect 8194 38556 8204 38612
rect 8260 38556 8270 38612
rect 4454 38388 4464 38444
rect 4520 38388 4568 38444
rect 4624 38388 4672 38444
rect 4728 38388 4738 38444
rect 24454 38388 24464 38444
rect 24520 38388 24568 38444
rect 24624 38388 24672 38444
rect 24728 38388 24738 38444
rect 28448 38388 28560 38416
rect 27234 38332 27244 38388
rect 27300 38332 28560 38388
rect 28448 38304 28560 38332
rect 1138 38220 1148 38276
rect 1204 38220 4844 38276
rect 4900 38220 4910 38276
rect 5954 38220 5964 38276
rect 6020 38220 6524 38276
rect 6580 38220 6590 38276
rect 0 38164 112 38192
rect 0 38108 812 38164
rect 868 38108 878 38164
rect 0 38080 112 38108
rect 10434 37996 10444 38052
rect 10500 37996 10892 38052
rect 10948 37996 15148 38052
rect 15204 37996 15214 38052
rect 20738 37996 20748 38052
rect 20804 37996 26236 38052
rect 26292 37996 26302 38052
rect 28448 37940 28560 37968
rect 4386 37884 4396 37940
rect 4452 37884 5404 37940
rect 5460 37884 5470 37940
rect 25666 37884 25676 37940
rect 25732 37884 28560 37940
rect 28448 37856 28560 37884
rect 7858 37772 7868 37828
rect 7924 37772 17332 37828
rect 17490 37772 17500 37828
rect 17556 37772 27356 37828
rect 27412 37772 27422 37828
rect 17276 37716 17332 37772
rect 1782 37660 1820 37716
rect 1876 37660 1886 37716
rect 6962 37660 6972 37716
rect 7028 37660 10668 37716
rect 10724 37660 16380 37716
rect 16436 37660 16446 37716
rect 17276 37660 22764 37716
rect 22820 37660 22830 37716
rect 3794 37604 3804 37660
rect 3860 37604 3908 37660
rect 3964 37604 4012 37660
rect 4068 37604 4078 37660
rect 23794 37604 23804 37660
rect 23860 37604 23908 37660
rect 23964 37604 24012 37660
rect 24068 37604 24078 37660
rect 28448 37492 28560 37520
rect 2146 37436 2156 37492
rect 2212 37436 2828 37492
rect 2884 37436 2894 37492
rect 5618 37436 5628 37492
rect 5684 37436 24668 37492
rect 24724 37436 24734 37492
rect 27010 37436 27020 37492
rect 27076 37436 28560 37492
rect 28448 37408 28560 37436
rect 354 37324 364 37380
rect 420 37324 3164 37380
rect 3220 37324 3230 37380
rect 4834 37324 4844 37380
rect 4900 37324 6524 37380
rect 6580 37324 10332 37380
rect 10388 37324 10398 37380
rect 12002 37324 12012 37380
rect 12068 37324 12796 37380
rect 12852 37324 17164 37380
rect 17220 37324 17230 37380
rect 0 37268 112 37296
rect 0 37212 8372 37268
rect 8642 37212 8652 37268
rect 8708 37212 9660 37268
rect 9716 37212 9726 37268
rect 12114 37212 12124 37268
rect 12180 37212 15932 37268
rect 15988 37212 15998 37268
rect 0 37184 112 37212
rect 1922 37100 1932 37156
rect 1988 37100 8092 37156
rect 8148 37100 8158 37156
rect 8316 37044 8372 37212
rect 8530 37100 8540 37156
rect 8596 37100 26236 37156
rect 26292 37100 26302 37156
rect 28448 37044 28560 37072
rect 2706 36988 2716 37044
rect 2772 36988 3388 37044
rect 3444 36988 4844 37044
rect 4900 36988 4910 37044
rect 8316 36988 14364 37044
rect 14420 36988 14430 37044
rect 16258 36988 16268 37044
rect 16324 36988 24668 37044
rect 24724 36988 24734 37044
rect 25442 36988 25452 37044
rect 25508 36988 28560 37044
rect 28448 36960 28560 36988
rect 1698 36876 1708 36932
rect 1764 36876 2492 36932
rect 2548 36876 2558 36932
rect 4454 36820 4464 36876
rect 4520 36820 4568 36876
rect 4624 36820 4672 36876
rect 4728 36820 4738 36876
rect 24454 36820 24464 36876
rect 24520 36820 24568 36876
rect 24624 36820 24672 36876
rect 24728 36820 24738 36876
rect 9538 36764 9548 36820
rect 9604 36764 19908 36820
rect 19852 36708 19908 36764
rect 3332 36652 6412 36708
rect 6468 36652 11788 36708
rect 11844 36652 11854 36708
rect 16146 36652 16156 36708
rect 16212 36652 16716 36708
rect 16772 36652 16782 36708
rect 19852 36652 24668 36708
rect 24724 36652 24734 36708
rect 3332 36596 3388 36652
rect 28448 36596 28560 36624
rect 2818 36540 2828 36596
rect 2884 36540 3164 36596
rect 3220 36540 3388 36596
rect 3602 36540 3612 36596
rect 3668 36540 4172 36596
rect 4228 36540 4238 36596
rect 27234 36540 27244 36596
rect 27300 36540 28560 36596
rect 28448 36512 28560 36540
rect 1698 36428 1708 36484
rect 1764 36428 5796 36484
rect 6514 36428 6524 36484
rect 6580 36428 7868 36484
rect 7924 36428 7934 36484
rect 0 36372 112 36400
rect 0 36316 5684 36372
rect 0 36288 112 36316
rect 1698 36204 1708 36260
rect 1764 36204 1820 36260
rect 1876 36204 1886 36260
rect 5628 36148 5684 36316
rect 5740 36260 5796 36428
rect 5954 36316 5964 36372
rect 6020 36316 26460 36372
rect 26516 36316 26526 36372
rect 5740 36204 6860 36260
rect 6916 36204 7868 36260
rect 7924 36204 7934 36260
rect 19394 36204 19404 36260
rect 19460 36204 19852 36260
rect 19908 36204 19918 36260
rect 28448 36148 28560 36176
rect 5628 36092 12236 36148
rect 12292 36092 12302 36148
rect 25666 36092 25676 36148
rect 25732 36092 28560 36148
rect 3794 36036 3804 36092
rect 3860 36036 3908 36092
rect 3964 36036 4012 36092
rect 4068 36036 4078 36092
rect 23794 36036 23804 36092
rect 23860 36036 23908 36092
rect 23964 36036 24012 36092
rect 24068 36036 24078 36092
rect 28448 36064 28560 36092
rect 26002 35980 26012 36036
rect 26068 35980 26078 36036
rect 1362 35756 1372 35812
rect 1428 35756 2716 35812
rect 2772 35756 2782 35812
rect 4386 35756 4396 35812
rect 4452 35756 25004 35812
rect 25060 35756 25070 35812
rect 26012 35588 26068 35980
rect 28448 35700 28560 35728
rect 27122 35644 27132 35700
rect 27188 35644 28560 35700
rect 28448 35616 28560 35644
rect 26002 35532 26012 35588
rect 26068 35532 26078 35588
rect 0 35476 112 35504
rect 0 35420 11676 35476
rect 11732 35420 11742 35476
rect 22306 35420 22316 35476
rect 22372 35420 24892 35476
rect 24948 35420 24958 35476
rect 0 35392 112 35420
rect 9426 35308 9436 35364
rect 9492 35308 9502 35364
rect 4454 35252 4464 35308
rect 4520 35252 4568 35308
rect 4624 35252 4672 35308
rect 4728 35252 4738 35308
rect 9436 35252 9492 35308
rect 24454 35252 24464 35308
rect 24520 35252 24568 35308
rect 24624 35252 24672 35308
rect 24728 35252 24738 35308
rect 28448 35252 28560 35280
rect 2594 35196 2604 35252
rect 2660 35196 3836 35252
rect 3892 35196 3902 35252
rect 5506 35196 5516 35252
rect 5572 35196 7084 35252
rect 7140 35196 7150 35252
rect 9436 35196 11228 35252
rect 11284 35196 11294 35252
rect 17490 35196 17500 35252
rect 17556 35196 18284 35252
rect 18340 35196 18350 35252
rect 27234 35196 27244 35252
rect 27300 35196 28560 35252
rect 9436 35140 9492 35196
rect 28448 35168 28560 35196
rect 3724 35084 9492 35140
rect 3724 35028 3780 35084
rect 3332 34972 3724 35028
rect 3780 34972 3790 35028
rect 7074 34972 7084 35028
rect 7140 34972 7756 35028
rect 7812 34972 7822 35028
rect 15586 34972 15596 35028
rect 15652 34972 18284 35028
rect 18340 34972 18350 35028
rect 3332 34916 3388 34972
rect 1922 34860 1932 34916
rect 1988 34860 3388 34916
rect 8418 34860 8428 34916
rect 8484 34860 9100 34916
rect 9156 34860 9166 34916
rect 10854 34860 10892 34916
rect 10948 34860 10958 34916
rect 16370 34860 16380 34916
rect 16436 34860 19068 34916
rect 19124 34860 19134 34916
rect 25554 34860 25564 34916
rect 25620 34860 26236 34916
rect 26292 34860 26302 34916
rect 28448 34804 28560 34832
rect 2370 34748 2380 34804
rect 2436 34748 2828 34804
rect 2884 34748 2894 34804
rect 17490 34748 17500 34804
rect 17556 34748 18060 34804
rect 18116 34748 18126 34804
rect 25666 34748 25676 34804
rect 25732 34748 28560 34804
rect 28448 34720 28560 34748
rect 3332 34636 4844 34692
rect 4900 34636 4910 34692
rect 5394 34636 5404 34692
rect 5460 34636 5852 34692
rect 5908 34636 5918 34692
rect 8194 34636 8204 34692
rect 8260 34636 9100 34692
rect 9156 34636 9166 34692
rect 18386 34636 18396 34692
rect 18452 34636 26348 34692
rect 26404 34636 26414 34692
rect 0 34580 112 34608
rect 3332 34580 3388 34636
rect 0 34524 3388 34580
rect 0 34496 112 34524
rect 3794 34468 3804 34524
rect 3860 34468 3908 34524
rect 3964 34468 4012 34524
rect 4068 34468 4078 34524
rect 23794 34468 23804 34524
rect 23860 34468 23908 34524
rect 23964 34468 24012 34524
rect 24068 34468 24078 34524
rect 2258 34412 2268 34468
rect 2324 34412 3052 34468
rect 3108 34412 3118 34468
rect 9090 34412 9100 34468
rect 9156 34412 9324 34468
rect 9380 34412 9548 34468
rect 9604 34412 9614 34468
rect 28448 34356 28560 34384
rect 2482 34300 2492 34356
rect 2548 34300 26348 34356
rect 26404 34300 26414 34356
rect 27010 34300 27020 34356
rect 27076 34300 28560 34356
rect 28448 34272 28560 34300
rect 4274 34188 4284 34244
rect 4340 34188 18060 34244
rect 18116 34188 18126 34244
rect 2482 34076 2492 34132
rect 2548 34076 2716 34132
rect 2772 34076 2782 34132
rect 4162 34076 4172 34132
rect 4228 34076 5404 34132
rect 5460 34076 5470 34132
rect 8082 34076 8092 34132
rect 8148 34076 10220 34132
rect 10276 34076 10286 34132
rect 10882 34076 10892 34132
rect 10948 34076 11228 34132
rect 11284 34076 11294 34132
rect 11778 34076 11788 34132
rect 11844 34076 13580 34132
rect 13636 34076 21308 34132
rect 21364 34076 21374 34132
rect 1138 33964 1148 34020
rect 1204 33964 2380 34020
rect 2436 33964 2446 34020
rect 5058 33964 5068 34020
rect 5124 33964 6188 34020
rect 6244 33964 6254 34020
rect 7858 33964 7868 34020
rect 7924 33964 8204 34020
rect 8260 33964 8270 34020
rect 25218 33964 25228 34020
rect 25284 33964 26236 34020
rect 26292 33964 26302 34020
rect 28448 33908 28560 33936
rect 1922 33852 1932 33908
rect 1988 33852 5292 33908
rect 5348 33852 5358 33908
rect 13346 33852 13356 33908
rect 13412 33852 24668 33908
rect 24724 33852 24734 33908
rect 25666 33852 25676 33908
rect 25732 33852 28560 33908
rect 28448 33824 28560 33852
rect 3378 33740 3388 33796
rect 3444 33740 3612 33796
rect 3668 33740 3678 33796
rect 8866 33740 8876 33796
rect 8932 33740 8988 33796
rect 9044 33740 9054 33796
rect 0 33684 112 33712
rect 4454 33684 4464 33740
rect 4520 33684 4568 33740
rect 4624 33684 4672 33740
rect 4728 33684 4738 33740
rect 24454 33684 24464 33740
rect 24520 33684 24568 33740
rect 24624 33684 24672 33740
rect 24728 33684 24738 33740
rect 0 33628 4284 33684
rect 4340 33628 4350 33684
rect 4834 33628 4844 33684
rect 4900 33628 6636 33684
rect 6692 33628 6702 33684
rect 15586 33628 15596 33684
rect 15652 33628 17500 33684
rect 17556 33628 17566 33684
rect 21634 33628 21644 33684
rect 21700 33628 23436 33684
rect 23492 33628 23502 33684
rect 0 33600 112 33628
rect 3154 33516 3164 33572
rect 3220 33516 4508 33572
rect 4564 33516 4956 33572
rect 5012 33516 5022 33572
rect 5282 33516 5292 33572
rect 5348 33516 5516 33572
rect 5572 33516 5582 33572
rect 6290 33516 6300 33572
rect 6356 33516 24892 33572
rect 24948 33516 24958 33572
rect 28448 33460 28560 33488
rect 6962 33404 6972 33460
rect 7028 33404 7644 33460
rect 7700 33404 7980 33460
rect 8036 33404 8046 33460
rect 8642 33404 8652 33460
rect 8708 33404 9436 33460
rect 9492 33404 13244 33460
rect 13300 33404 13310 33460
rect 17826 33404 17836 33460
rect 17892 33404 18732 33460
rect 18788 33404 19180 33460
rect 19236 33404 19246 33460
rect 27234 33404 27244 33460
rect 27300 33404 28560 33460
rect 7980 33348 8036 33404
rect 28448 33376 28560 33404
rect 7980 33292 8876 33348
rect 8932 33292 8942 33348
rect 3266 33180 3276 33236
rect 3332 33180 3724 33236
rect 3780 33180 3790 33236
rect 8082 33180 8092 33236
rect 8148 33180 8204 33236
rect 8260 33180 8270 33236
rect 15092 33180 24668 33236
rect 24724 33180 24734 33236
rect 13234 33068 13244 33124
rect 13300 33068 13468 33124
rect 13524 33068 13534 33124
rect 15092 33012 15148 33180
rect 28448 33012 28560 33040
rect 10434 32956 10444 33012
rect 10500 32956 15148 33012
rect 25666 32956 25676 33012
rect 25732 32956 28560 33012
rect 3794 32900 3804 32956
rect 3860 32900 3908 32956
rect 3964 32900 4012 32956
rect 4068 32900 4078 32956
rect 23794 32900 23804 32956
rect 23860 32900 23908 32956
rect 23964 32900 24012 32956
rect 24068 32900 24078 32956
rect 28448 32928 28560 32956
rect 5842 32844 5852 32900
rect 5908 32844 8652 32900
rect 8708 32844 8718 32900
rect 12338 32844 12348 32900
rect 12404 32844 12460 32900
rect 12516 32844 12526 32900
rect 0 32788 112 32816
rect 0 32732 17388 32788
rect 17444 32732 17836 32788
rect 17892 32732 17902 32788
rect 0 32704 112 32732
rect 1026 32620 1036 32676
rect 1092 32620 1484 32676
rect 1540 32620 5852 32676
rect 5908 32620 5918 32676
rect 7522 32620 7532 32676
rect 7588 32620 9324 32676
rect 9380 32620 9390 32676
rect 12562 32620 12572 32676
rect 12628 32620 15596 32676
rect 15652 32620 15662 32676
rect 22082 32620 22092 32676
rect 22148 32620 26236 32676
rect 26292 32620 26302 32676
rect 28448 32564 28560 32592
rect 4498 32508 4508 32564
rect 4564 32508 26908 32564
rect 27122 32508 27132 32564
rect 27188 32508 28560 32564
rect 3826 32396 3836 32452
rect 3892 32396 26124 32452
rect 26180 32396 26190 32452
rect 26852 32340 26908 32508
rect 28448 32480 28560 32508
rect 2258 32284 2268 32340
rect 2324 32284 13916 32340
rect 13972 32284 13982 32340
rect 17938 32284 17948 32340
rect 18004 32284 21868 32340
rect 21924 32284 21934 32340
rect 26852 32284 28364 32340
rect 28420 32284 28430 32340
rect 8082 32172 8092 32228
rect 8148 32172 9996 32228
rect 10052 32172 10062 32228
rect 11638 32172 11676 32228
rect 11732 32172 11742 32228
rect 18050 32172 18060 32228
rect 18116 32172 18620 32228
rect 18676 32172 18686 32228
rect 21186 32172 21196 32228
rect 21252 32172 21700 32228
rect 4454 32116 4464 32172
rect 4520 32116 4568 32172
rect 4624 32116 4672 32172
rect 4728 32116 4738 32172
rect 11788 32060 12460 32116
rect 12516 32060 12526 32116
rect 1698 31948 1708 32004
rect 1764 31948 2380 32004
rect 2436 31948 7644 32004
rect 7700 31948 7710 32004
rect 0 31892 112 31920
rect 11788 31892 11844 32060
rect 12002 31948 12012 32004
rect 12068 31948 12908 32004
rect 12964 31948 12974 32004
rect 21644 31892 21700 32172
rect 24454 32116 24464 32172
rect 24520 32116 24568 32172
rect 24624 32116 24672 32172
rect 24728 32116 24738 32172
rect 28448 32116 28560 32144
rect 27234 32060 27244 32116
rect 27300 32060 28560 32116
rect 28448 32032 28560 32060
rect 0 31836 10332 31892
rect 10388 31836 10398 31892
rect 11106 31836 11116 31892
rect 11172 31836 11844 31892
rect 21634 31836 21644 31892
rect 21700 31836 21710 31892
rect 0 31808 112 31836
rect 1474 31724 1484 31780
rect 1540 31724 1708 31780
rect 1764 31724 1774 31780
rect 5842 31724 5852 31780
rect 5908 31724 9100 31780
rect 9156 31724 9166 31780
rect 10098 31724 10108 31780
rect 10164 31724 10892 31780
rect 10948 31724 10958 31780
rect 12114 31724 12124 31780
rect 12180 31724 13244 31780
rect 13300 31724 13310 31780
rect 14466 31724 14476 31780
rect 14532 31724 20300 31780
rect 20356 31724 21532 31780
rect 21588 31724 21598 31780
rect 28448 31668 28560 31696
rect 3332 31612 6524 31668
rect 6580 31612 6590 31668
rect 10182 31612 10220 31668
rect 10276 31612 10286 31668
rect 11442 31612 11452 31668
rect 11508 31612 15932 31668
rect 15988 31612 18508 31668
rect 18564 31612 18574 31668
rect 25666 31612 25676 31668
rect 25732 31612 28560 31668
rect 3332 31556 3388 31612
rect 28448 31584 28560 31612
rect 2258 31500 2268 31556
rect 2324 31500 3388 31556
rect 5506 31500 5516 31556
rect 5572 31500 5852 31556
rect 5908 31500 5918 31556
rect 6402 31500 6412 31556
rect 6468 31500 24332 31556
rect 24388 31500 24398 31556
rect 5740 31388 10108 31444
rect 10164 31388 10174 31444
rect 11330 31388 11340 31444
rect 11396 31388 11676 31444
rect 11732 31388 11742 31444
rect 12338 31388 12348 31444
rect 12404 31388 13580 31444
rect 13636 31388 13646 31444
rect 20178 31388 20188 31444
rect 20244 31388 20636 31444
rect 20692 31388 20702 31444
rect 20962 31388 20972 31444
rect 21028 31388 21308 31444
rect 21364 31388 21374 31444
rect 3794 31332 3804 31388
rect 3860 31332 3908 31388
rect 3964 31332 4012 31388
rect 4068 31332 4078 31388
rect 4274 31164 4284 31220
rect 4340 31164 5404 31220
rect 5460 31164 5470 31220
rect 0 30996 112 31024
rect 5740 30996 5796 31388
rect 23794 31332 23804 31388
rect 23860 31332 23908 31388
rect 23964 31332 24012 31388
rect 24068 31332 24078 31388
rect 7074 31276 7084 31332
rect 7140 31276 7420 31332
rect 7476 31276 23212 31332
rect 23268 31276 23660 31332
rect 23716 31276 23726 31332
rect 28448 31220 28560 31248
rect 5954 31164 5964 31220
rect 6020 31164 6300 31220
rect 6356 31164 7308 31220
rect 7364 31164 7374 31220
rect 9996 31164 13468 31220
rect 13524 31164 13534 31220
rect 19954 31164 19964 31220
rect 20020 31164 20972 31220
rect 21028 31164 21038 31220
rect 27010 31164 27020 31220
rect 27076 31164 28560 31220
rect 9996 31108 10052 31164
rect 28448 31136 28560 31164
rect 7858 31052 7868 31108
rect 7924 31052 9996 31108
rect 10052 31052 10062 31108
rect 10210 31052 10220 31108
rect 10276 31052 11228 31108
rect 11284 31052 11294 31108
rect 0 30940 5796 30996
rect 8866 30940 8876 30996
rect 8932 30940 15820 30996
rect 15876 30940 15886 30996
rect 18498 30940 18508 30996
rect 18564 30940 18574 30996
rect 19730 30940 19740 30996
rect 19796 30940 22092 30996
rect 22148 30940 22158 30996
rect 23650 30940 23660 30996
rect 23716 30940 25116 30996
rect 25172 30940 25182 30996
rect 0 30912 112 30940
rect 18508 30884 18564 30940
rect 2706 30828 2716 30884
rect 2772 30828 5292 30884
rect 5348 30828 5358 30884
rect 6514 30828 6524 30884
rect 6580 30828 9100 30884
rect 9156 30828 14476 30884
rect 14532 30828 14542 30884
rect 15026 30828 15036 30884
rect 15092 30828 16940 30884
rect 16996 30828 17006 30884
rect 18508 30828 22484 30884
rect 22428 30772 22484 30828
rect 28448 30772 28560 30800
rect 1810 30716 1820 30772
rect 1876 30716 3164 30772
rect 3220 30716 10892 30772
rect 10948 30716 10958 30772
rect 13206 30716 13244 30772
rect 13300 30716 13310 30772
rect 13430 30716 13468 30772
rect 13524 30716 13534 30772
rect 22418 30716 22428 30772
rect 22484 30716 22494 30772
rect 25442 30716 25452 30772
rect 25508 30716 28560 30772
rect 28448 30688 28560 30716
rect 9650 30604 9660 30660
rect 9716 30604 11340 30660
rect 11396 30604 12348 30660
rect 12404 30604 12414 30660
rect 12786 30604 12796 30660
rect 12852 30604 13356 30660
rect 13412 30604 13422 30660
rect 4454 30548 4464 30604
rect 4520 30548 4568 30604
rect 4624 30548 4672 30604
rect 4728 30548 4738 30604
rect 24454 30548 24464 30604
rect 24520 30548 24568 30604
rect 24624 30548 24672 30604
rect 24728 30548 24738 30604
rect 2594 30492 2604 30548
rect 2660 30492 3052 30548
rect 3108 30492 3118 30548
rect 5954 30492 5964 30548
rect 6020 30492 7420 30548
rect 7476 30492 7486 30548
rect 12226 30492 12236 30548
rect 12292 30492 13468 30548
rect 13524 30492 14588 30548
rect 14644 30492 22652 30548
rect 22708 30492 22718 30548
rect 2930 30380 2940 30436
rect 2996 30380 13804 30436
rect 13860 30380 13870 30436
rect 28448 30324 28560 30352
rect 1586 30268 1596 30324
rect 1652 30268 2828 30324
rect 2884 30268 2894 30324
rect 4162 30268 4172 30324
rect 4228 30268 4900 30324
rect 6066 30268 6076 30324
rect 6132 30268 6300 30324
rect 6356 30268 6366 30324
rect 27234 30268 27244 30324
rect 27300 30268 28560 30324
rect 4844 30212 4900 30268
rect 28448 30240 28560 30268
rect 3266 30156 3276 30212
rect 3332 30156 4284 30212
rect 4340 30156 4350 30212
rect 4834 30156 4844 30212
rect 4900 30156 4910 30212
rect 7298 30156 7308 30212
rect 7364 30156 8876 30212
rect 8932 30156 8942 30212
rect 9426 30156 9436 30212
rect 9492 30156 10780 30212
rect 10836 30156 10846 30212
rect 14242 30156 14252 30212
rect 14308 30156 14318 30212
rect 15698 30156 15708 30212
rect 15764 30156 16492 30212
rect 16548 30156 16558 30212
rect 17490 30156 17500 30212
rect 17556 30156 21420 30212
rect 21476 30156 21486 30212
rect 21746 30156 21756 30212
rect 21812 30156 23100 30212
rect 23156 30156 23166 30212
rect 0 30100 112 30128
rect 14252 30100 14308 30156
rect 0 30044 2492 30100
rect 2548 30044 2558 30100
rect 5618 30044 5628 30100
rect 5684 30044 7868 30100
rect 7924 30044 7934 30100
rect 8530 30044 8540 30100
rect 8596 30044 12908 30100
rect 12964 30044 12974 30100
rect 13580 30044 14308 30100
rect 15250 30044 15260 30100
rect 15316 30044 17052 30100
rect 17108 30044 19292 30100
rect 19348 30044 20300 30100
rect 20356 30044 21532 30100
rect 21588 30044 21598 30100
rect 0 30016 112 30044
rect 13580 29988 13636 30044
rect 1026 29932 1036 29988
rect 1092 29932 8316 29988
rect 8372 29932 8382 29988
rect 10098 29932 10108 29988
rect 10164 29932 10556 29988
rect 10612 29932 10622 29988
rect 12114 29932 12124 29988
rect 12180 29932 13636 29988
rect 13794 29932 13804 29988
rect 13860 29932 17276 29988
rect 17332 29932 17342 29988
rect 17714 29932 17724 29988
rect 17780 29932 18620 29988
rect 18676 29932 18686 29988
rect 28448 29876 28560 29904
rect 6514 29820 6524 29876
rect 6580 29820 6972 29876
rect 7028 29820 7644 29876
rect 7700 29820 10444 29876
rect 10500 29820 13468 29876
rect 13524 29820 18284 29876
rect 18340 29820 18350 29876
rect 27010 29820 27020 29876
rect 27076 29820 28560 29876
rect 3794 29764 3804 29820
rect 3860 29764 3908 29820
rect 3964 29764 4012 29820
rect 4068 29764 4078 29820
rect 23794 29764 23804 29820
rect 23860 29764 23908 29820
rect 23964 29764 24012 29820
rect 24068 29764 24078 29820
rect 28448 29792 28560 29820
rect 7522 29708 7532 29764
rect 7588 29708 8316 29764
rect 8372 29708 8382 29764
rect 9762 29708 9772 29764
rect 9828 29708 11788 29764
rect 11844 29708 11854 29764
rect 12012 29708 18396 29764
rect 18452 29708 18462 29764
rect 12012 29652 12068 29708
rect 4274 29596 4284 29652
rect 4340 29596 4956 29652
rect 5012 29596 5022 29652
rect 6626 29596 6636 29652
rect 6692 29596 7196 29652
rect 7252 29596 7262 29652
rect 8306 29596 8316 29652
rect 8372 29596 12068 29652
rect 13906 29596 13916 29652
rect 13972 29596 28140 29652
rect 28196 29596 28206 29652
rect 1138 29484 1148 29540
rect 1204 29484 2268 29540
rect 2324 29484 2716 29540
rect 2772 29484 5068 29540
rect 5124 29484 7084 29540
rect 7140 29484 8540 29540
rect 8596 29484 8606 29540
rect 11554 29484 11564 29540
rect 11620 29484 12348 29540
rect 12404 29484 12414 29540
rect 13010 29484 13020 29540
rect 13076 29484 26236 29540
rect 26292 29484 26302 29540
rect 28448 29428 28560 29456
rect 466 29372 476 29428
rect 532 29372 1484 29428
rect 1540 29372 1550 29428
rect 3490 29372 3500 29428
rect 3556 29372 5124 29428
rect 5282 29372 5292 29428
rect 5348 29372 5628 29428
rect 5684 29372 15260 29428
rect 15316 29372 15326 29428
rect 15474 29372 15484 29428
rect 15540 29372 16716 29428
rect 16772 29372 16782 29428
rect 19842 29372 19852 29428
rect 19908 29372 23100 29428
rect 23156 29372 23166 29428
rect 27122 29372 27132 29428
rect 27188 29372 28560 29428
rect 0 29204 112 29232
rect 3332 29204 3388 29316
rect 3444 29260 3454 29316
rect 0 29148 3388 29204
rect 0 29120 112 29148
rect 5068 29092 5124 29372
rect 28448 29344 28560 29372
rect 8306 29260 8316 29316
rect 8372 29260 18172 29316
rect 18228 29260 18238 29316
rect 2930 29036 2940 29092
rect 2996 29036 3276 29092
rect 3332 29036 3342 29092
rect 5068 29036 11564 29092
rect 11620 29036 11630 29092
rect 4454 28980 4464 29036
rect 4520 28980 4568 29036
rect 4624 28980 4672 29036
rect 4728 28980 4738 29036
rect 24454 28980 24464 29036
rect 24520 28980 24568 29036
rect 24624 28980 24672 29036
rect 24728 28980 24738 29036
rect 28448 28980 28560 29008
rect 8950 28924 8988 28980
rect 9044 28924 9996 28980
rect 10052 28924 10062 28980
rect 15250 28924 15260 28980
rect 15316 28924 15708 28980
rect 15764 28924 15774 28980
rect 27234 28924 27244 28980
rect 27300 28924 28560 28980
rect 28448 28896 28560 28924
rect 2482 28812 2492 28868
rect 2548 28812 2940 28868
rect 2996 28812 3006 28868
rect 12226 28812 12236 28868
rect 12292 28812 12572 28868
rect 12628 28812 12638 28868
rect 1810 28700 1820 28756
rect 1876 28700 2380 28756
rect 2436 28700 2446 28756
rect 4050 28700 4060 28756
rect 4116 28700 4508 28756
rect 4564 28700 4574 28756
rect 10882 28700 10892 28756
rect 10948 28700 13804 28756
rect 13860 28700 13870 28756
rect 17826 28700 17836 28756
rect 17892 28700 18508 28756
rect 18564 28700 18574 28756
rect 6626 28588 6636 28644
rect 6692 28588 7308 28644
rect 7364 28588 7374 28644
rect 11106 28588 11116 28644
rect 11172 28588 11900 28644
rect 11956 28588 11966 28644
rect 16034 28588 16044 28644
rect 16100 28588 26236 28644
rect 26292 28588 26302 28644
rect 28448 28532 28560 28560
rect 802 28476 812 28532
rect 868 28476 1484 28532
rect 1540 28476 3164 28532
rect 3220 28476 3230 28532
rect 7410 28476 7420 28532
rect 7476 28476 9548 28532
rect 9604 28476 10444 28532
rect 10500 28476 10510 28532
rect 10668 28476 17388 28532
rect 17444 28476 17454 28532
rect 19170 28476 19180 28532
rect 19236 28476 26124 28532
rect 26180 28476 26190 28532
rect 27234 28476 27244 28532
rect 27300 28476 28560 28532
rect 10668 28420 10724 28476
rect 28448 28448 28560 28476
rect 1586 28364 1596 28420
rect 1652 28364 2044 28420
rect 2100 28364 2110 28420
rect 5170 28364 5180 28420
rect 5236 28364 7532 28420
rect 7588 28364 7598 28420
rect 10546 28364 10556 28420
rect 10612 28364 10724 28420
rect 11106 28364 11116 28420
rect 11172 28364 11676 28420
rect 11732 28364 11742 28420
rect 20066 28364 20076 28420
rect 20132 28364 23548 28420
rect 23604 28364 23614 28420
rect 0 28308 112 28336
rect 0 28252 3668 28308
rect 8194 28252 8204 28308
rect 8260 28252 12348 28308
rect 12404 28252 12414 28308
rect 12674 28252 12684 28308
rect 12740 28252 13580 28308
rect 13636 28252 13646 28308
rect 15092 28252 22988 28308
rect 23044 28252 23054 28308
rect 0 28224 112 28252
rect 3612 28084 3668 28252
rect 3794 28196 3804 28252
rect 3860 28196 3908 28252
rect 3964 28196 4012 28252
rect 4068 28196 4078 28252
rect 12348 28196 12404 28252
rect 15092 28196 15148 28252
rect 23794 28196 23804 28252
rect 23860 28196 23908 28252
rect 23964 28196 24012 28252
rect 24068 28196 24078 28252
rect 12348 28140 15148 28196
rect 28448 28084 28560 28112
rect 3612 28028 7084 28084
rect 7140 28028 7756 28084
rect 7812 28028 7822 28084
rect 10882 28028 10892 28084
rect 10948 28028 11340 28084
rect 11396 28028 11406 28084
rect 12114 28028 12124 28084
rect 12180 28028 13020 28084
rect 13076 28028 13086 28084
rect 27234 28028 27244 28084
rect 27300 28028 28560 28084
rect 28448 28000 28560 28028
rect 1586 27916 1596 27972
rect 1652 27916 8204 27972
rect 8260 27916 8270 27972
rect 10098 27916 10108 27972
rect 10164 27916 13468 27972
rect 13524 27916 13534 27972
rect 7410 27804 7420 27860
rect 7476 27804 7980 27860
rect 8036 27804 8046 27860
rect 10994 27804 11004 27860
rect 11060 27804 12908 27860
rect 12964 27804 12974 27860
rect 13234 27804 13244 27860
rect 13300 27804 14364 27860
rect 14420 27804 15372 27860
rect 15428 27804 15438 27860
rect 16594 27804 16604 27860
rect 16660 27804 16940 27860
rect 16996 27804 17612 27860
rect 17668 27804 17678 27860
rect 21634 27804 21644 27860
rect 21700 27804 28364 27860
rect 28420 27804 28430 27860
rect 10210 27692 10220 27748
rect 10276 27692 11564 27748
rect 11620 27692 11630 27748
rect 12786 27692 12796 27748
rect 12852 27692 13020 27748
rect 13076 27692 13086 27748
rect 25890 27692 25900 27748
rect 25956 27692 26236 27748
rect 26292 27692 26302 27748
rect 28448 27636 28560 27664
rect 4284 27580 5964 27636
rect 6020 27580 6030 27636
rect 27010 27580 27020 27636
rect 27076 27580 28560 27636
rect 0 27412 112 27440
rect 4284 27412 4340 27580
rect 28448 27552 28560 27580
rect 9426 27468 9436 27524
rect 9492 27468 9660 27524
rect 9716 27468 10556 27524
rect 10612 27468 10622 27524
rect 13570 27468 13580 27524
rect 13636 27468 15148 27524
rect 4454 27412 4464 27468
rect 4520 27412 4568 27468
rect 4624 27412 4672 27468
rect 4728 27412 4738 27468
rect 15092 27412 15148 27468
rect 24454 27412 24464 27468
rect 24520 27412 24568 27468
rect 24624 27412 24672 27468
rect 24728 27412 24738 27468
rect 0 27356 3388 27412
rect 4050 27356 4060 27412
rect 4116 27356 4340 27412
rect 5506 27356 5516 27412
rect 5572 27356 14196 27412
rect 15092 27356 16604 27412
rect 16660 27356 21308 27412
rect 21364 27356 21374 27412
rect 0 27328 112 27356
rect 1474 27244 1484 27300
rect 1540 27244 1708 27300
rect 1764 27244 1774 27300
rect 3332 27188 3388 27356
rect 14140 27300 14196 27356
rect 4274 27244 4284 27300
rect 4340 27244 4956 27300
rect 5012 27244 5022 27300
rect 9426 27244 9436 27300
rect 9492 27244 9996 27300
rect 10052 27244 10062 27300
rect 13122 27244 13132 27300
rect 13188 27244 13916 27300
rect 13972 27244 13982 27300
rect 14140 27244 24332 27300
rect 24388 27244 24398 27300
rect 28448 27188 28560 27216
rect 3332 27132 7420 27188
rect 7476 27132 7486 27188
rect 7830 27132 7868 27188
rect 7924 27132 7934 27188
rect 8082 27132 8092 27188
rect 8148 27132 11452 27188
rect 11508 27132 11518 27188
rect 16706 27132 16716 27188
rect 16772 27132 17388 27188
rect 17444 27132 17454 27188
rect 25666 27132 25676 27188
rect 25732 27132 28560 27188
rect 28448 27104 28560 27132
rect 1250 27020 1260 27076
rect 1316 27020 1820 27076
rect 1876 27020 1886 27076
rect 3938 27020 3948 27076
rect 4004 27020 4732 27076
rect 4788 27020 4798 27076
rect 5254 27020 5292 27076
rect 5348 27020 5358 27076
rect 6402 27020 6412 27076
rect 6468 27020 10220 27076
rect 10276 27020 10286 27076
rect 13906 27020 13916 27076
rect 13972 27020 26236 27076
rect 26292 27020 26302 27076
rect 3266 26908 3276 26964
rect 3332 26908 5404 26964
rect 5460 26908 5470 26964
rect 9314 26908 9324 26964
rect 9380 26908 9436 26964
rect 9492 26908 9502 26964
rect 12562 26908 12572 26964
rect 12628 26908 19068 26964
rect 19124 26908 19134 26964
rect 12114 26796 12124 26852
rect 12180 26796 15988 26852
rect 16370 26796 16380 26852
rect 16436 26796 20188 26852
rect 20244 26796 21588 26852
rect 10994 26684 11004 26740
rect 11060 26684 11228 26740
rect 11284 26684 11294 26740
rect 12338 26684 12348 26740
rect 12404 26684 13020 26740
rect 13076 26684 13086 26740
rect 13906 26684 13916 26740
rect 13972 26684 14252 26740
rect 14308 26684 14318 26740
rect 3794 26628 3804 26684
rect 3860 26628 3908 26684
rect 3964 26628 4012 26684
rect 4068 26628 4078 26684
rect 15932 26628 15988 26796
rect 21532 26740 21588 26796
rect 28448 26740 28560 26768
rect 21522 26684 21532 26740
rect 21588 26684 21598 26740
rect 27234 26684 27244 26740
rect 27300 26684 28560 26740
rect 23794 26628 23804 26684
rect 23860 26628 23908 26684
rect 23964 26628 24012 26684
rect 24068 26628 24078 26684
rect 28448 26656 28560 26684
rect 15932 26572 20412 26628
rect 20468 26572 21084 26628
rect 21140 26572 21150 26628
rect 0 26516 112 26544
rect 0 26460 1260 26516
rect 1316 26460 1326 26516
rect 11218 26460 11228 26516
rect 11284 26460 17836 26516
rect 17892 26460 21420 26516
rect 21476 26460 21486 26516
rect 0 26432 112 26460
rect 6738 26348 6748 26404
rect 6804 26348 7420 26404
rect 7476 26348 7486 26404
rect 14242 26348 14252 26404
rect 14308 26348 14812 26404
rect 14868 26348 14878 26404
rect 28448 26292 28560 26320
rect 3154 26236 3164 26292
rect 3220 26236 9548 26292
rect 9604 26236 9772 26292
rect 9828 26236 9838 26292
rect 12226 26236 12236 26292
rect 12292 26236 12572 26292
rect 12628 26236 12638 26292
rect 14578 26236 14588 26292
rect 14644 26236 15260 26292
rect 15316 26236 15326 26292
rect 15596 26236 25004 26292
rect 25060 26236 25070 26292
rect 25666 26236 25676 26292
rect 25732 26236 28560 26292
rect 15596 26180 15652 26236
rect 28448 26208 28560 26236
rect 2118 26124 2156 26180
rect 2212 26124 2380 26180
rect 2436 26124 2446 26180
rect 5506 26124 5516 26180
rect 5572 26124 15652 26180
rect 15810 26124 15820 26180
rect 15876 26124 24332 26180
rect 24388 26124 24398 26180
rect 4386 26012 4396 26068
rect 4452 26012 5292 26068
rect 5348 26012 5358 26068
rect 7410 26012 7420 26068
rect 7476 26012 7980 26068
rect 8036 26012 8046 26068
rect 9426 26012 9436 26068
rect 9492 26012 9772 26068
rect 9828 26012 9838 26068
rect 9986 26012 9996 26068
rect 10052 26012 10556 26068
rect 10612 26012 10622 26068
rect 10994 26012 11004 26068
rect 11060 26012 11228 26068
rect 11284 26012 11294 26068
rect 21298 26012 21308 26068
rect 21364 26012 21868 26068
rect 21924 26012 21934 26068
rect 5292 25956 5348 26012
rect 5292 25900 13244 25956
rect 13300 25900 14476 25956
rect 14532 25900 17948 25956
rect 18004 25900 18014 25956
rect 4454 25844 4464 25900
rect 4520 25844 4568 25900
rect 4624 25844 4672 25900
rect 4728 25844 4738 25900
rect 24454 25844 24464 25900
rect 24520 25844 24568 25900
rect 24624 25844 24672 25900
rect 24728 25844 24738 25900
rect 28448 25844 28560 25872
rect 11106 25788 11116 25844
rect 11172 25788 17276 25844
rect 17332 25788 18732 25844
rect 18788 25788 18798 25844
rect 27234 25788 27244 25844
rect 27300 25788 28560 25844
rect 28448 25760 28560 25788
rect 3602 25676 3612 25732
rect 3668 25676 4956 25732
rect 5012 25676 5022 25732
rect 7074 25676 7084 25732
rect 7140 25676 7196 25732
rect 7252 25676 7262 25732
rect 8642 25676 8652 25732
rect 8708 25676 9548 25732
rect 9604 25676 11004 25732
rect 11060 25676 11070 25732
rect 16258 25676 16268 25732
rect 16324 25676 26236 25732
rect 26292 25676 26302 25732
rect 0 25620 112 25648
rect 0 25564 5516 25620
rect 5572 25564 5582 25620
rect 10668 25564 11676 25620
rect 11732 25564 11788 25620
rect 11844 25564 11854 25620
rect 0 25536 112 25564
rect 10668 25508 10724 25564
rect 9090 25452 9100 25508
rect 9156 25452 9660 25508
rect 9716 25452 9726 25508
rect 10658 25452 10668 25508
rect 10724 25452 10734 25508
rect 12572 25452 12908 25508
rect 12964 25452 14924 25508
rect 14980 25452 14990 25508
rect 18722 25452 18732 25508
rect 18788 25452 26236 25508
rect 26292 25452 26302 25508
rect 12572 25396 12628 25452
rect 28448 25396 28560 25424
rect 12562 25340 12572 25396
rect 12628 25340 12638 25396
rect 18386 25340 18396 25396
rect 18452 25340 19740 25396
rect 19796 25340 20412 25396
rect 20468 25340 20478 25396
rect 27122 25340 27132 25396
rect 27188 25340 28560 25396
rect 28448 25312 28560 25340
rect 2034 25228 2044 25284
rect 2100 25228 2716 25284
rect 2772 25228 2782 25284
rect 11106 25228 11116 25284
rect 11172 25228 11340 25284
rect 11396 25228 11406 25284
rect 15474 25228 15484 25284
rect 15540 25228 16380 25284
rect 16436 25228 16446 25284
rect 25666 25228 25676 25284
rect 25732 25228 26964 25284
rect 3794 25060 3804 25116
rect 3860 25060 3908 25116
rect 3964 25060 4012 25116
rect 4068 25060 4078 25116
rect 23794 25060 23804 25116
rect 23860 25060 23908 25116
rect 23964 25060 24012 25116
rect 24068 25060 24078 25116
rect 13682 25004 13692 25060
rect 13748 25004 14028 25060
rect 14084 25004 14094 25060
rect 26908 24948 26964 25228
rect 28448 24948 28560 24976
rect 3378 24892 3388 24948
rect 3444 24892 7644 24948
rect 7700 24892 7710 24948
rect 10770 24892 10780 24948
rect 10836 24892 25004 24948
rect 25060 24892 25070 24948
rect 26908 24892 28560 24948
rect 28448 24864 28560 24892
rect 3490 24780 3500 24836
rect 3556 24780 4172 24836
rect 4228 24780 4238 24836
rect 4722 24780 4732 24836
rect 4788 24780 9212 24836
rect 9268 24780 18172 24836
rect 18228 24780 18238 24836
rect 20626 24780 20636 24836
rect 20692 24780 21644 24836
rect 21700 24780 21710 24836
rect 0 24724 112 24752
rect 0 24668 3500 24724
rect 3556 24668 3566 24724
rect 11106 24668 11116 24724
rect 11172 24668 25228 24724
rect 25284 24668 25294 24724
rect 0 24640 112 24668
rect 2594 24556 2604 24612
rect 2660 24556 6972 24612
rect 7028 24556 7038 24612
rect 7858 24556 7868 24612
rect 7924 24556 7980 24612
rect 8036 24556 8046 24612
rect 13682 24556 13692 24612
rect 13748 24556 14588 24612
rect 14644 24556 14654 24612
rect 15026 24556 15036 24612
rect 15092 24556 15372 24612
rect 15428 24556 15438 24612
rect 15586 24556 15596 24612
rect 15652 24556 16828 24612
rect 16884 24556 16894 24612
rect 17052 24556 24668 24612
rect 24724 24556 24734 24612
rect 17052 24500 17108 24556
rect 28448 24500 28560 24528
rect 3154 24444 3164 24500
rect 3220 24444 11340 24500
rect 11396 24444 11406 24500
rect 12226 24444 12236 24500
rect 12292 24444 12796 24500
rect 12852 24444 12862 24500
rect 16034 24444 16044 24500
rect 16100 24444 17108 24500
rect 17602 24444 17612 24500
rect 17668 24444 17836 24500
rect 17892 24444 17902 24500
rect 18060 24444 26236 24500
rect 26292 24444 26302 24500
rect 27234 24444 27244 24500
rect 27300 24444 28560 24500
rect 18060 24388 18116 24444
rect 28448 24416 28560 24444
rect 3462 24332 3500 24388
rect 3556 24332 3566 24388
rect 9874 24332 9884 24388
rect 9940 24332 14252 24388
rect 14308 24332 14318 24388
rect 14690 24332 14700 24388
rect 14756 24332 15820 24388
rect 15876 24332 15886 24388
rect 16492 24332 18116 24388
rect 4454 24276 4464 24332
rect 4520 24276 4568 24332
rect 4624 24276 4672 24332
rect 4728 24276 4738 24332
rect 6962 24220 6972 24276
rect 7028 24220 15148 24276
rect 15204 24220 15214 24276
rect 16492 24164 16548 24332
rect 24454 24276 24464 24332
rect 24520 24276 24568 24332
rect 24624 24276 24672 24332
rect 24728 24276 24738 24332
rect 16706 24220 16716 24276
rect 16772 24220 22372 24276
rect 22316 24164 22372 24220
rect 7158 24108 7196 24164
rect 7252 24108 7262 24164
rect 15092 24108 16548 24164
rect 21074 24108 21084 24164
rect 21140 24108 22092 24164
rect 22148 24108 22158 24164
rect 22316 24108 26012 24164
rect 26068 24108 26078 24164
rect 15092 24052 15148 24108
rect 28448 24052 28560 24080
rect 1586 23996 1596 24052
rect 1652 23996 3388 24052
rect 3444 23996 3454 24052
rect 8950 23996 8988 24052
rect 9044 23996 9054 24052
rect 11778 23996 11788 24052
rect 11844 23996 15148 24052
rect 17154 23996 17164 24052
rect 17220 23996 18844 24052
rect 18900 23996 20972 24052
rect 21028 23996 22652 24052
rect 22708 23996 22718 24052
rect 25666 23996 25676 24052
rect 25732 23996 28560 24052
rect 28448 23968 28560 23996
rect 4610 23884 4620 23940
rect 4676 23884 5068 23940
rect 5124 23884 5292 23940
rect 5348 23884 5358 23940
rect 5506 23884 5516 23940
rect 5572 23884 6748 23940
rect 6804 23884 6814 23940
rect 8194 23884 8204 23940
rect 8260 23884 11564 23940
rect 11620 23884 11630 23940
rect 12450 23884 12460 23940
rect 12516 23884 13468 23940
rect 13524 23884 13580 23940
rect 13636 23884 13646 23940
rect 14354 23884 14364 23940
rect 14420 23884 16940 23940
rect 16996 23884 17836 23940
rect 17892 23884 17902 23940
rect 18610 23884 18620 23940
rect 18676 23884 19740 23940
rect 19796 23884 19806 23940
rect 23762 23884 23772 23940
rect 23828 23884 24332 23940
rect 24388 23884 24398 23940
rect 0 23828 112 23856
rect 0 23772 1372 23828
rect 1428 23772 1438 23828
rect 2370 23772 2380 23828
rect 2436 23772 3276 23828
rect 3332 23772 3342 23828
rect 8950 23772 8988 23828
rect 9044 23772 9054 23828
rect 11218 23772 11228 23828
rect 11284 23772 11676 23828
rect 11732 23772 11742 23828
rect 12002 23772 12012 23828
rect 12068 23772 12348 23828
rect 12404 23772 12414 23828
rect 18946 23772 18956 23828
rect 19012 23772 19292 23828
rect 19348 23772 24892 23828
rect 24948 23772 24958 23828
rect 0 23744 112 23772
rect 7074 23660 7084 23716
rect 7140 23660 7756 23716
rect 7812 23660 7822 23716
rect 9062 23660 9100 23716
rect 9156 23660 9166 23716
rect 9650 23660 9660 23716
rect 9716 23660 26236 23716
rect 26292 23660 26302 23716
rect 28448 23604 28560 23632
rect 4834 23548 4844 23604
rect 4900 23548 13804 23604
rect 13860 23548 13870 23604
rect 17602 23548 17612 23604
rect 17668 23548 18284 23604
rect 18340 23548 20188 23604
rect 20244 23548 20254 23604
rect 27234 23548 27244 23604
rect 27300 23548 28560 23604
rect 3794 23492 3804 23548
rect 3860 23492 3908 23548
rect 3964 23492 4012 23548
rect 4068 23492 4078 23548
rect 23794 23492 23804 23548
rect 23860 23492 23908 23548
rect 23964 23492 24012 23548
rect 24068 23492 24078 23548
rect 28448 23520 28560 23548
rect 6178 23436 6188 23492
rect 6244 23436 6412 23492
rect 6468 23436 6478 23492
rect 7186 23436 7196 23492
rect 7252 23436 8876 23492
rect 8932 23436 8942 23492
rect 9762 23436 9772 23492
rect 9828 23436 9996 23492
rect 10052 23436 10062 23492
rect 15138 23436 15148 23492
rect 15204 23436 19964 23492
rect 20020 23436 23660 23492
rect 23716 23436 23726 23492
rect 5618 23324 5628 23380
rect 5684 23324 10108 23380
rect 10164 23324 10174 23380
rect 16258 23324 16268 23380
rect 16324 23324 17052 23380
rect 17108 23324 17118 23380
rect 19814 23324 19852 23380
rect 19908 23324 19918 23380
rect 354 23212 364 23268
rect 420 23212 1148 23268
rect 1204 23212 1214 23268
rect 1474 23212 1484 23268
rect 1540 23212 1708 23268
rect 1764 23212 2268 23268
rect 2324 23212 2334 23268
rect 6962 23212 6972 23268
rect 7028 23212 9324 23268
rect 9380 23212 9548 23268
rect 9604 23212 9614 23268
rect 9762 23212 9772 23268
rect 9828 23212 24892 23268
rect 24948 23212 24958 23268
rect 1484 23156 1540 23212
rect 28448 23156 28560 23184
rect 1250 23100 1260 23156
rect 1316 23100 1540 23156
rect 2706 23100 2716 23156
rect 2772 23100 5292 23156
rect 5348 23100 5740 23156
rect 5796 23100 5806 23156
rect 9986 23100 9996 23156
rect 10052 23100 11620 23156
rect 14690 23100 14700 23156
rect 14756 23100 18396 23156
rect 18452 23100 18462 23156
rect 25666 23100 25676 23156
rect 25732 23100 28560 23156
rect 11564 23044 11620 23100
rect 28448 23072 28560 23100
rect 5170 22988 5180 23044
rect 5236 22988 10164 23044
rect 10882 22988 10892 23044
rect 10948 22988 11340 23044
rect 11396 22988 11406 23044
rect 11564 22988 15148 23044
rect 15204 22988 15214 23044
rect 16594 22988 16604 23044
rect 16660 22988 26236 23044
rect 26292 22988 26302 23044
rect 0 22932 112 22960
rect 10108 22932 10164 22988
rect 0 22876 5516 22932
rect 5572 22876 5582 22932
rect 7746 22876 7756 22932
rect 7812 22876 8092 22932
rect 8148 22876 8158 22932
rect 10108 22876 25900 22932
rect 25956 22876 25966 22932
rect 0 22848 112 22876
rect 6066 22764 6076 22820
rect 6132 22764 6412 22820
rect 6468 22764 10332 22820
rect 10388 22764 10398 22820
rect 10994 22764 11004 22820
rect 11060 22764 11340 22820
rect 11396 22764 11406 22820
rect 13346 22764 13356 22820
rect 13412 22764 20692 22820
rect 4454 22708 4464 22764
rect 4520 22708 4568 22764
rect 4624 22708 4672 22764
rect 4728 22708 4738 22764
rect 10994 22652 11004 22708
rect 11060 22652 11116 22708
rect 11172 22652 11182 22708
rect 20636 22596 20692 22764
rect 24454 22708 24464 22764
rect 24520 22708 24568 22764
rect 24624 22708 24672 22764
rect 24728 22708 24738 22764
rect 28448 22708 28560 22736
rect 27234 22652 27244 22708
rect 27300 22652 28560 22708
rect 28448 22624 28560 22652
rect 5618 22540 5628 22596
rect 5684 22540 10444 22596
rect 10500 22540 11788 22596
rect 11844 22540 11854 22596
rect 13346 22540 13356 22596
rect 13412 22540 18172 22596
rect 18228 22540 18238 22596
rect 20636 22540 26236 22596
rect 26292 22540 26302 22596
rect 11442 22428 11452 22484
rect 11508 22428 14812 22484
rect 14868 22428 14878 22484
rect 18050 22428 18060 22484
rect 18116 22428 21868 22484
rect 21924 22428 22876 22484
rect 22932 22428 22942 22484
rect 2594 22316 2604 22372
rect 2660 22316 5628 22372
rect 5684 22316 5694 22372
rect 10882 22316 10892 22372
rect 10948 22316 11676 22372
rect 11732 22316 12236 22372
rect 12292 22316 12302 22372
rect 15362 22316 15372 22372
rect 15428 22316 20076 22372
rect 20132 22316 21420 22372
rect 21476 22316 21486 22372
rect 28448 22260 28560 22288
rect 2818 22204 2828 22260
rect 2884 22204 3164 22260
rect 3220 22204 3230 22260
rect 19282 22204 19292 22260
rect 19348 22204 20636 22260
rect 20692 22204 20702 22260
rect 27122 22204 27132 22260
rect 27188 22204 28560 22260
rect 28448 22176 28560 22204
rect 5170 22092 5180 22148
rect 5236 22092 5628 22148
rect 5684 22092 6076 22148
rect 6132 22092 6142 22148
rect 11890 22092 11900 22148
rect 11956 22092 14140 22148
rect 14196 22092 14206 22148
rect 16034 22092 16044 22148
rect 16100 22092 19068 22148
rect 19124 22092 19628 22148
rect 19684 22092 19694 22148
rect 0 22036 112 22064
rect 0 21980 1484 22036
rect 1540 21980 1550 22036
rect 5730 21980 5740 22036
rect 5796 21980 7532 22036
rect 7588 21980 7598 22036
rect 11218 21980 11228 22036
rect 11284 21980 14700 22036
rect 14756 21980 14766 22036
rect 19730 21980 19740 22036
rect 19796 21980 19806 22036
rect 23426 21980 23436 22036
rect 23492 21980 23660 22036
rect 23716 21980 23726 22036
rect 0 21952 112 21980
rect 3794 21924 3804 21980
rect 3860 21924 3908 21980
rect 3964 21924 4012 21980
rect 4068 21924 4078 21980
rect 9538 21868 9548 21924
rect 9604 21868 10892 21924
rect 10948 21868 10958 21924
rect 13346 21868 13356 21924
rect 13412 21868 15372 21924
rect 15428 21868 15438 21924
rect 19740 21812 19796 21980
rect 23794 21924 23804 21980
rect 23860 21924 23908 21980
rect 23964 21924 24012 21980
rect 24068 21924 24078 21980
rect 28448 21812 28560 21840
rect 578 21756 588 21812
rect 644 21756 1596 21812
rect 1652 21756 3164 21812
rect 3220 21756 4172 21812
rect 4228 21756 4238 21812
rect 11106 21756 11116 21812
rect 11172 21756 12348 21812
rect 12404 21756 12414 21812
rect 15138 21756 15148 21812
rect 15204 21756 16156 21812
rect 16212 21756 16222 21812
rect 19740 21756 21980 21812
rect 22036 21756 22046 21812
rect 25666 21756 25676 21812
rect 25732 21756 28560 21812
rect 28448 21728 28560 21756
rect 2930 21644 2940 21700
rect 2996 21644 4956 21700
rect 5012 21644 6972 21700
rect 7028 21644 7038 21700
rect 13990 21644 14028 21700
rect 14084 21644 14094 21700
rect 17266 21644 17276 21700
rect 17332 21644 18508 21700
rect 18564 21644 18956 21700
rect 19012 21644 20748 21700
rect 20804 21644 20814 21700
rect 21186 21644 21196 21700
rect 21252 21644 25788 21700
rect 25844 21644 25854 21700
rect 5394 21532 5404 21588
rect 5460 21532 6748 21588
rect 6804 21532 6814 21588
rect 10546 21532 10556 21588
rect 10612 21532 11228 21588
rect 11284 21532 11294 21588
rect 12114 21532 12124 21588
rect 12180 21532 14812 21588
rect 14868 21532 14878 21588
rect 16146 21532 16156 21588
rect 16212 21532 16828 21588
rect 16884 21532 16894 21588
rect 17378 21532 17388 21588
rect 17444 21532 19292 21588
rect 19348 21532 19358 21588
rect 19506 21532 19516 21588
rect 19572 21532 21084 21588
rect 21140 21532 21150 21588
rect 5170 21420 5180 21476
rect 5236 21420 8540 21476
rect 8596 21420 9212 21476
rect 9268 21420 9278 21476
rect 14018 21420 14028 21476
rect 14084 21420 15148 21476
rect 15204 21420 15214 21476
rect 15362 21420 15372 21476
rect 15428 21420 16492 21476
rect 16548 21420 16558 21476
rect 19842 21420 19852 21476
rect 19908 21420 26236 21476
rect 26292 21420 26302 21476
rect 28448 21364 28560 21392
rect 4274 21308 4284 21364
rect 4340 21308 7308 21364
rect 7364 21308 7374 21364
rect 10994 21308 11004 21364
rect 11060 21308 16828 21364
rect 16884 21308 16894 21364
rect 17602 21308 17612 21364
rect 17668 21308 18284 21364
rect 18340 21308 18350 21364
rect 19618 21308 19628 21364
rect 19684 21308 20636 21364
rect 20692 21308 20702 21364
rect 20962 21308 20972 21364
rect 21028 21308 28560 21364
rect 28448 21280 28560 21308
rect 6738 21196 6748 21252
rect 6804 21196 7084 21252
rect 7140 21196 7150 21252
rect 15138 21196 15148 21252
rect 15204 21196 23548 21252
rect 0 21140 112 21168
rect 4454 21140 4464 21196
rect 4520 21140 4568 21196
rect 4624 21140 4672 21196
rect 4728 21140 4738 21196
rect 0 21084 3108 21140
rect 3602 21084 3612 21140
rect 3668 21084 4172 21140
rect 4228 21084 4238 21140
rect 8306 21084 8316 21140
rect 8372 21084 19796 21140
rect 19954 21084 19964 21140
rect 20020 21084 20188 21140
rect 20244 21084 20254 21140
rect 0 21056 112 21084
rect 3052 21028 3108 21084
rect 3052 20972 5292 21028
rect 5348 20972 5358 21028
rect 10210 20972 10220 21028
rect 10276 20972 15148 21028
rect 17938 20972 17948 21028
rect 18004 20972 18844 21028
rect 18900 20972 18910 21028
rect 19058 20972 19068 21028
rect 19124 20972 19292 21028
rect 19348 20972 19358 21028
rect 15092 20916 15148 20972
rect 19740 20916 19796 21084
rect 23492 21028 23548 21196
rect 24454 21140 24464 21196
rect 24520 21140 24568 21196
rect 24624 21140 24672 21196
rect 24728 21140 24738 21196
rect 23492 20972 25228 21028
rect 25284 20972 25294 21028
rect 28448 20916 28560 20944
rect 1810 20860 1820 20916
rect 1876 20860 3164 20916
rect 3220 20860 3230 20916
rect 13570 20860 13580 20916
rect 13636 20860 14812 20916
rect 14868 20860 14878 20916
rect 15092 20860 19516 20916
rect 19572 20860 19582 20916
rect 19740 20860 25564 20916
rect 25620 20860 25630 20916
rect 27318 20860 27356 20916
rect 27412 20860 27422 20916
rect 28130 20860 28140 20916
rect 28196 20860 28560 20916
rect 28448 20832 28560 20860
rect 4386 20748 4396 20804
rect 4452 20748 6524 20804
rect 6580 20748 6590 20804
rect 6738 20748 6748 20804
rect 6804 20748 12348 20804
rect 12404 20748 15148 20804
rect 16034 20748 16044 20804
rect 16100 20748 16828 20804
rect 16884 20748 16894 20804
rect 19282 20748 19292 20804
rect 19348 20748 20188 20804
rect 20244 20748 20254 20804
rect 21746 20748 21756 20804
rect 21812 20748 21980 20804
rect 22036 20748 22046 20804
rect 7186 20636 7196 20692
rect 7252 20636 8428 20692
rect 8484 20636 8494 20692
rect 15092 20580 15148 20748
rect 15250 20636 15260 20692
rect 15316 20636 19068 20692
rect 19124 20636 19134 20692
rect 5842 20524 5852 20580
rect 5908 20524 6524 20580
rect 6580 20524 6590 20580
rect 12562 20524 12572 20580
rect 12628 20524 13356 20580
rect 13412 20524 13422 20580
rect 15092 20524 20748 20580
rect 20804 20524 21196 20580
rect 21252 20524 21262 20580
rect 23202 20524 23212 20580
rect 23268 20524 24388 20580
rect 25778 20524 25788 20580
rect 25844 20524 26348 20580
rect 26404 20524 26414 20580
rect 24332 20468 24388 20524
rect 28448 20468 28560 20496
rect 1922 20412 1932 20468
rect 1988 20412 2828 20468
rect 2884 20412 2894 20468
rect 24332 20412 28560 20468
rect 3794 20356 3804 20412
rect 3860 20356 3908 20412
rect 3964 20356 4012 20412
rect 4068 20356 4078 20412
rect 23794 20356 23804 20412
rect 23860 20356 23908 20412
rect 23964 20356 24012 20412
rect 24068 20356 24078 20412
rect 28448 20384 28560 20412
rect 19506 20300 19516 20356
rect 19572 20300 19628 20356
rect 19684 20300 19694 20356
rect 20290 20300 20300 20356
rect 20356 20300 20524 20356
rect 20580 20300 20590 20356
rect 0 20244 112 20272
rect 0 20188 2716 20244
rect 2772 20188 2782 20244
rect 2930 20188 2940 20244
rect 2996 20188 9100 20244
rect 9156 20188 9772 20244
rect 9828 20188 11116 20244
rect 11172 20188 11182 20244
rect 14578 20188 14588 20244
rect 14644 20188 14924 20244
rect 14980 20188 14990 20244
rect 18050 20188 18060 20244
rect 18116 20188 18620 20244
rect 18676 20188 18686 20244
rect 0 20160 112 20188
rect 6178 20076 6188 20132
rect 6244 20076 7980 20132
rect 8036 20076 8046 20132
rect 8754 20076 8764 20132
rect 8820 20076 11340 20132
rect 11396 20076 11406 20132
rect 13020 20076 20748 20132
rect 20804 20076 20814 20132
rect 20962 20076 20972 20132
rect 21028 20076 22204 20132
rect 22260 20076 22270 20132
rect 7858 19964 7868 20020
rect 7924 19964 9604 20020
rect 9986 19964 9996 20020
rect 10052 19964 12796 20020
rect 12852 19964 12862 20020
rect 9548 19908 9604 19964
rect 13020 19908 13076 20076
rect 28448 20020 28560 20048
rect 13570 19964 13580 20020
rect 13636 19964 14700 20020
rect 14756 19964 14766 20020
rect 14914 19964 14924 20020
rect 14980 19964 16492 20020
rect 16548 19964 16558 20020
rect 19954 19964 19964 20020
rect 20020 19964 20860 20020
rect 20916 19964 20926 20020
rect 28354 19964 28364 20020
rect 28420 19964 28560 20020
rect 28448 19936 28560 19964
rect 7970 19852 7980 19908
rect 8036 19852 8876 19908
rect 8932 19852 8942 19908
rect 9548 19852 13076 19908
rect 14802 19852 14812 19908
rect 14868 19852 17612 19908
rect 17668 19852 17678 19908
rect 17826 19852 17836 19908
rect 17892 19852 18620 19908
rect 18676 19852 18686 19908
rect 17612 19796 17668 19852
rect 2118 19740 2156 19796
rect 2212 19740 2492 19796
rect 2548 19740 2558 19796
rect 10882 19740 10892 19796
rect 10948 19740 13468 19796
rect 13524 19740 13916 19796
rect 13972 19740 13982 19796
rect 17612 19740 17948 19796
rect 18004 19740 18014 19796
rect 19730 19740 19740 19796
rect 19796 19740 20860 19796
rect 20916 19740 20926 19796
rect 6738 19628 6748 19684
rect 6804 19628 6972 19684
rect 7028 19628 15148 19684
rect 4454 19572 4464 19628
rect 4520 19572 4568 19628
rect 4624 19572 4672 19628
rect 4728 19572 4738 19628
rect 15092 19572 15148 19628
rect 24454 19572 24464 19628
rect 24520 19572 24568 19628
rect 24624 19572 24672 19628
rect 24728 19572 24738 19628
rect 28448 19572 28560 19600
rect 8194 19516 8204 19572
rect 8260 19516 14476 19572
rect 14532 19516 14812 19572
rect 14868 19516 14878 19572
rect 15092 19516 24220 19572
rect 24276 19516 24286 19572
rect 25106 19516 25116 19572
rect 25172 19516 28560 19572
rect 28448 19488 28560 19516
rect 12786 19404 12796 19460
rect 12852 19404 12862 19460
rect 16258 19404 16268 19460
rect 16324 19404 25900 19460
rect 25956 19404 25966 19460
rect 0 19348 112 19376
rect 0 19292 1148 19348
rect 1204 19292 1214 19348
rect 2230 19292 2268 19348
rect 2324 19292 2334 19348
rect 9846 19292 9884 19348
rect 9940 19292 9950 19348
rect 12002 19292 12012 19348
rect 12068 19292 12572 19348
rect 12628 19292 12638 19348
rect 0 19264 112 19292
rect 4610 19180 4620 19236
rect 4676 19180 5404 19236
rect 5460 19180 5470 19236
rect 7298 19180 7308 19236
rect 7364 19180 7868 19236
rect 7924 19180 7934 19236
rect 12796 19124 12852 19404
rect 15474 19292 15484 19348
rect 15540 19292 15932 19348
rect 15988 19292 16716 19348
rect 16772 19292 16782 19348
rect 26450 19292 26460 19348
rect 26516 19292 27244 19348
rect 27300 19292 27310 19348
rect 13234 19180 13244 19236
rect 13300 19180 13580 19236
rect 13636 19180 13646 19236
rect 17378 19180 17388 19236
rect 17444 19180 19628 19236
rect 19684 19180 19694 19236
rect 28448 19124 28560 19152
rect 3042 19068 3052 19124
rect 3108 19068 3612 19124
rect 3668 19068 7420 19124
rect 7476 19068 11116 19124
rect 11172 19068 11182 19124
rect 12450 19068 12460 19124
rect 12516 19068 15932 19124
rect 15988 19068 15998 19124
rect 16146 19068 16156 19124
rect 16212 19068 17276 19124
rect 17332 19068 17342 19124
rect 26852 19068 28560 19124
rect 26852 19012 26908 19068
rect 28448 19040 28560 19068
rect 5730 18956 5740 19012
rect 5796 18956 5964 19012
rect 6020 18956 26908 19012
rect 12114 18844 12124 18900
rect 12180 18844 13020 18900
rect 13076 18844 13086 18900
rect 16034 18844 16044 18900
rect 16100 18844 18620 18900
rect 18676 18844 18686 18900
rect 3794 18788 3804 18844
rect 3860 18788 3908 18844
rect 3964 18788 4012 18844
rect 4068 18788 4078 18844
rect 23794 18788 23804 18844
rect 23860 18788 23908 18844
rect 23964 18788 24012 18844
rect 24068 18788 24078 18844
rect 5030 18732 5068 18788
rect 5124 18732 5134 18788
rect 5506 18732 5516 18788
rect 5572 18732 5964 18788
rect 6020 18732 6030 18788
rect 14018 18732 14028 18788
rect 14084 18732 23324 18788
rect 23380 18732 23390 18788
rect 28448 18676 28560 18704
rect 1362 18620 1372 18676
rect 1428 18620 6076 18676
rect 6132 18620 6142 18676
rect 10546 18620 10556 18676
rect 10612 18620 10780 18676
rect 10836 18620 13020 18676
rect 13076 18620 13086 18676
rect 16706 18620 16716 18676
rect 16772 18620 20412 18676
rect 20468 18620 20478 18676
rect 20738 18620 20748 18676
rect 20804 18620 28560 18676
rect 5058 18508 5068 18564
rect 5124 18508 16604 18564
rect 16660 18508 16670 18564
rect 0 18452 112 18480
rect 0 18396 700 18452
rect 756 18396 766 18452
rect 2146 18396 2156 18452
rect 2212 18396 2380 18452
rect 2436 18396 2446 18452
rect 3938 18396 3948 18452
rect 4004 18396 4844 18452
rect 4900 18396 4910 18452
rect 5394 18396 5404 18452
rect 5460 18396 6188 18452
rect 6244 18396 6254 18452
rect 14690 18396 14700 18452
rect 14756 18396 16716 18452
rect 16772 18396 16782 18452
rect 17602 18396 17612 18452
rect 17668 18396 17948 18452
rect 18004 18396 18014 18452
rect 0 18368 112 18396
rect 4834 18284 4844 18340
rect 4900 18284 6524 18340
rect 6580 18284 6590 18340
rect 7970 18284 7980 18340
rect 8036 18284 8764 18340
rect 8820 18284 9324 18340
rect 9380 18284 9390 18340
rect 10994 18284 11004 18340
rect 11060 18284 11452 18340
rect 11508 18284 14028 18340
rect 14084 18284 14094 18340
rect 17378 18284 17388 18340
rect 17444 18284 18172 18340
rect 18228 18284 18238 18340
rect 1698 18172 1708 18228
rect 1764 18172 3500 18228
rect 3556 18172 13580 18228
rect 13636 18172 13646 18228
rect 18396 18116 18452 18620
rect 28448 18592 28560 18620
rect 18834 18508 18844 18564
rect 18900 18508 18910 18564
rect 22082 18508 22092 18564
rect 22148 18508 23436 18564
rect 23492 18508 23502 18564
rect 18582 18284 18620 18340
rect 18676 18284 18686 18340
rect 18844 18116 18900 18508
rect 21522 18396 21532 18452
rect 21588 18396 21756 18452
rect 21812 18396 22148 18452
rect 22306 18396 22316 18452
rect 22372 18396 23660 18452
rect 23716 18396 23726 18452
rect 22092 18340 22148 18396
rect 20290 18284 20300 18340
rect 20356 18284 21420 18340
rect 21476 18284 21486 18340
rect 22092 18284 22652 18340
rect 22708 18284 22718 18340
rect 28448 18228 28560 18256
rect 19058 18172 19068 18228
rect 19124 18172 28560 18228
rect 28448 18144 28560 18172
rect 5926 18060 5964 18116
rect 6020 18060 6030 18116
rect 10994 18060 11004 18116
rect 11060 18060 11564 18116
rect 11620 18060 11630 18116
rect 17826 18060 17836 18116
rect 17892 18060 18060 18116
rect 18116 18060 18126 18116
rect 18396 18060 18620 18116
rect 18676 18060 18686 18116
rect 18844 18060 19516 18116
rect 19572 18060 19582 18116
rect 20598 18060 20636 18116
rect 20692 18060 20702 18116
rect 4454 18004 4464 18060
rect 4520 18004 4568 18060
rect 4624 18004 4672 18060
rect 4728 18004 4738 18060
rect 24454 18004 24464 18060
rect 24520 18004 24568 18060
rect 24624 18004 24672 18060
rect 24728 18004 24738 18060
rect 7298 17948 7308 18004
rect 7364 17948 21812 18004
rect 3378 17836 3388 17892
rect 3444 17836 3724 17892
rect 3780 17836 3790 17892
rect 4274 17836 4284 17892
rect 4340 17836 6524 17892
rect 6580 17836 6590 17892
rect 12674 17836 12684 17892
rect 12740 17836 13356 17892
rect 13412 17836 13422 17892
rect 16818 17836 16828 17892
rect 16884 17836 19516 17892
rect 19572 17836 19582 17892
rect 3826 17724 3836 17780
rect 3892 17724 5852 17780
rect 5908 17724 5918 17780
rect 6066 17724 6076 17780
rect 6132 17724 8876 17780
rect 8932 17724 8942 17780
rect 9874 17724 9884 17780
rect 9940 17724 16716 17780
rect 16772 17724 16782 17780
rect 17490 17724 17500 17780
rect 17556 17724 18844 17780
rect 18900 17724 18910 17780
rect 19058 17724 19068 17780
rect 19124 17724 19162 17780
rect 21756 17668 21812 17948
rect 22978 17836 22988 17892
rect 23044 17836 26908 17892
rect 26852 17780 26908 17836
rect 28448 17780 28560 17808
rect 22754 17724 22764 17780
rect 22820 17724 24556 17780
rect 24612 17724 24622 17780
rect 26852 17724 28560 17780
rect 28448 17696 28560 17724
rect 2930 17612 2940 17668
rect 2996 17612 4284 17668
rect 4340 17612 4350 17668
rect 4722 17612 4732 17668
rect 4788 17612 7308 17668
rect 7364 17612 7374 17668
rect 8194 17612 8204 17668
rect 8260 17612 9100 17668
rect 9156 17612 9166 17668
rect 18498 17612 18508 17668
rect 18564 17612 19292 17668
rect 19348 17612 20412 17668
rect 20468 17612 20860 17668
rect 20916 17612 21532 17668
rect 21588 17612 21598 17668
rect 21756 17612 25116 17668
rect 25172 17612 25182 17668
rect 0 17556 112 17584
rect 0 17500 1036 17556
rect 1092 17500 1102 17556
rect 2706 17500 2716 17556
rect 2772 17500 5068 17556
rect 5124 17500 5852 17556
rect 5908 17500 5918 17556
rect 10098 17500 10108 17556
rect 10164 17500 14924 17556
rect 14980 17500 14990 17556
rect 17378 17500 17388 17556
rect 17444 17500 17948 17556
rect 18004 17500 18014 17556
rect 18162 17500 18172 17556
rect 18228 17500 19404 17556
rect 19460 17500 22092 17556
rect 22148 17500 22158 17556
rect 0 17472 112 17500
rect 1250 17388 1260 17444
rect 1316 17388 1708 17444
rect 1764 17388 5236 17444
rect 5394 17388 5404 17444
rect 5460 17388 6412 17444
rect 6468 17388 6478 17444
rect 7522 17388 7532 17444
rect 7588 17388 11004 17444
rect 11060 17388 11070 17444
rect 11554 17388 11564 17444
rect 11620 17388 16156 17444
rect 16212 17388 16222 17444
rect 18050 17388 18060 17444
rect 18116 17388 18126 17444
rect 20178 17388 20188 17444
rect 20244 17388 26908 17444
rect 5180 17332 5236 17388
rect 18060 17332 18116 17388
rect 26852 17332 26908 17388
rect 28448 17332 28560 17360
rect 5180 17276 9996 17332
rect 10052 17276 10332 17332
rect 10388 17276 11116 17332
rect 11172 17276 12124 17332
rect 12180 17276 12190 17332
rect 15586 17276 15596 17332
rect 15652 17276 16940 17332
rect 16996 17276 20972 17332
rect 21028 17276 21038 17332
rect 26852 17276 28560 17332
rect 3794 17220 3804 17276
rect 3860 17220 3908 17276
rect 3964 17220 4012 17276
rect 4068 17220 4078 17276
rect 23794 17220 23804 17276
rect 23860 17220 23908 17276
rect 23964 17220 24012 17276
rect 24068 17220 24078 17276
rect 28448 17248 28560 17276
rect 5842 17164 5852 17220
rect 5908 17164 16940 17220
rect 16996 17164 17006 17220
rect 17154 17164 17164 17220
rect 17220 17164 19740 17220
rect 19796 17164 19806 17220
rect 1810 17052 1820 17108
rect 1876 17052 7812 17108
rect 9090 17052 9100 17108
rect 9156 17052 14700 17108
rect 14756 17052 14766 17108
rect 14914 17052 14924 17108
rect 14980 17052 19796 17108
rect 19954 17052 19964 17108
rect 20020 17052 21644 17108
rect 21700 17052 21710 17108
rect 7756 16996 7812 17052
rect 19740 16996 19796 17052
rect 2146 16940 2156 16996
rect 2212 16940 7532 16996
rect 7588 16940 7598 16996
rect 7746 16940 7756 16996
rect 7812 16940 8988 16996
rect 9044 16940 9054 16996
rect 9650 16940 9660 16996
rect 9716 16940 10108 16996
rect 10164 16940 10174 16996
rect 14354 16940 14364 16996
rect 14420 16940 19068 16996
rect 19124 16940 19134 16996
rect 19740 16940 26908 16996
rect 26852 16884 26908 16940
rect 28448 16884 28560 16912
rect 3350 16828 3388 16884
rect 3444 16828 3454 16884
rect 3826 16828 3836 16884
rect 3892 16828 4956 16884
rect 5012 16828 5022 16884
rect 8194 16828 8204 16884
rect 8260 16828 9324 16884
rect 9380 16828 9390 16884
rect 9874 16828 9884 16884
rect 9940 16828 10444 16884
rect 10500 16828 10510 16884
rect 12786 16828 12796 16884
rect 12852 16828 15036 16884
rect 15092 16828 15102 16884
rect 16930 16828 16940 16884
rect 16996 16828 22540 16884
rect 22596 16828 22988 16884
rect 23044 16828 23054 16884
rect 26852 16828 28560 16884
rect 28448 16800 28560 16828
rect 1586 16716 1596 16772
rect 1652 16716 2044 16772
rect 2100 16716 2268 16772
rect 2324 16716 2334 16772
rect 5058 16716 5068 16772
rect 5124 16716 6412 16772
rect 6468 16716 6478 16772
rect 6626 16716 6636 16772
rect 6692 16716 10108 16772
rect 10164 16716 10174 16772
rect 11218 16716 11228 16772
rect 11284 16716 13020 16772
rect 13076 16716 13468 16772
rect 13524 16716 13534 16772
rect 17266 16716 17276 16772
rect 17332 16716 18060 16772
rect 18116 16716 18126 16772
rect 18284 16716 19964 16772
rect 20020 16716 20030 16772
rect 20514 16716 20524 16772
rect 20580 16716 24892 16772
rect 24948 16716 24958 16772
rect 0 16660 112 16688
rect 18284 16660 18340 16716
rect 0 16604 5292 16660
rect 5348 16604 5358 16660
rect 15922 16604 15932 16660
rect 15988 16604 18340 16660
rect 18610 16604 18620 16660
rect 18676 16604 20860 16660
rect 20916 16604 20926 16660
rect 0 16576 112 16604
rect 6178 16492 6188 16548
rect 6244 16492 6636 16548
rect 6692 16492 6702 16548
rect 12114 16492 12124 16548
rect 12180 16492 18732 16548
rect 18788 16492 19068 16548
rect 19124 16492 19134 16548
rect 19366 16492 19404 16548
rect 19460 16492 19470 16548
rect 19702 16492 19740 16548
rect 19796 16492 19806 16548
rect 19954 16492 19964 16548
rect 20020 16492 24332 16548
rect 24388 16492 24398 16548
rect 4454 16436 4464 16492
rect 4520 16436 4568 16492
rect 4624 16436 4672 16492
rect 4728 16436 4738 16492
rect 24454 16436 24464 16492
rect 24520 16436 24568 16492
rect 24624 16436 24672 16492
rect 24728 16436 24738 16492
rect 28448 16436 28560 16464
rect 10098 16380 10108 16436
rect 10164 16380 11676 16436
rect 11732 16380 11742 16436
rect 17602 16380 17612 16436
rect 17668 16380 18060 16436
rect 18116 16380 20636 16436
rect 20692 16380 21308 16436
rect 21364 16380 21374 16436
rect 26852 16380 28560 16436
rect 26852 16324 26908 16380
rect 28448 16352 28560 16380
rect 1782 16268 1820 16324
rect 1876 16268 1886 16324
rect 2706 16268 2716 16324
rect 2772 16268 5516 16324
rect 5572 16268 5582 16324
rect 7074 16268 7084 16324
rect 7140 16268 9660 16324
rect 9716 16268 9726 16324
rect 10322 16268 10332 16324
rect 10388 16268 15932 16324
rect 15988 16268 15998 16324
rect 16146 16268 16156 16324
rect 16212 16268 26908 16324
rect 1820 16212 1876 16268
rect 1820 16156 2716 16212
rect 2772 16156 2782 16212
rect 3574 16156 3612 16212
rect 3668 16156 3678 16212
rect 4050 16156 4060 16212
rect 4116 16156 4172 16212
rect 4228 16156 4238 16212
rect 8950 16156 8988 16212
rect 9044 16156 9054 16212
rect 10406 16156 10444 16212
rect 10500 16156 10510 16212
rect 16034 16156 16044 16212
rect 16100 16156 19404 16212
rect 19460 16156 19470 16212
rect 19618 16156 19628 16212
rect 19684 16156 19740 16212
rect 19796 16156 19806 16212
rect 15922 16044 15932 16100
rect 15988 16044 16380 16100
rect 16436 16044 16446 16100
rect 16930 16044 16940 16100
rect 16996 16044 18284 16100
rect 18340 16044 18350 16100
rect 21942 16044 21980 16100
rect 22036 16044 22046 16100
rect 28448 15988 28560 16016
rect 6626 15932 6636 15988
rect 6692 15932 8204 15988
rect 8260 15932 8270 15988
rect 8530 15932 8540 15988
rect 8596 15932 9100 15988
rect 9156 15932 9166 15988
rect 16380 15932 28560 15988
rect 3378 15820 3388 15876
rect 3444 15820 5852 15876
rect 5908 15820 7532 15876
rect 7588 15820 8876 15876
rect 8932 15820 8942 15876
rect 10098 15820 10108 15876
rect 10164 15820 14364 15876
rect 14420 15820 14532 15876
rect 15026 15820 15036 15876
rect 15092 15820 16156 15876
rect 16212 15820 16222 15876
rect 0 15764 112 15792
rect 14476 15764 14532 15820
rect 0 15708 2828 15764
rect 2884 15708 2894 15764
rect 14476 15708 16156 15764
rect 16212 15708 16222 15764
rect 0 15680 112 15708
rect 3794 15652 3804 15708
rect 3860 15652 3908 15708
rect 3964 15652 4012 15708
rect 4068 15652 4078 15708
rect 6402 15596 6412 15652
rect 6468 15596 15148 15652
rect 15092 15540 15148 15596
rect 16380 15540 16436 15932
rect 28448 15904 28560 15932
rect 18050 15820 18060 15876
rect 18116 15820 18844 15876
rect 18900 15820 18910 15876
rect 19394 15820 19404 15876
rect 19460 15820 25452 15876
rect 25508 15820 25518 15876
rect 17490 15708 17500 15764
rect 17556 15708 21532 15764
rect 21588 15708 21598 15764
rect 23794 15652 23804 15708
rect 23860 15652 23908 15708
rect 23964 15652 24012 15708
rect 24068 15652 24078 15708
rect 17266 15596 17276 15652
rect 17332 15596 18396 15652
rect 18452 15596 18462 15652
rect 18610 15596 18620 15652
rect 18676 15596 18956 15652
rect 19012 15596 19022 15652
rect 19730 15596 19740 15652
rect 19796 15596 20188 15652
rect 20244 15596 20254 15652
rect 2146 15484 2156 15540
rect 2212 15484 8092 15540
rect 8148 15484 8158 15540
rect 8306 15484 8316 15540
rect 8372 15484 9996 15540
rect 10052 15484 10556 15540
rect 10612 15484 13244 15540
rect 13300 15484 14924 15540
rect 14980 15484 14990 15540
rect 15092 15484 16436 15540
rect 18956 15540 19012 15596
rect 28448 15540 28560 15568
rect 18956 15484 21420 15540
rect 21476 15484 21486 15540
rect 22530 15484 22540 15540
rect 22596 15484 28560 15540
rect 8316 15428 8372 15484
rect 28448 15456 28560 15484
rect 4274 15372 4284 15428
rect 4340 15372 5180 15428
rect 5236 15372 8372 15428
rect 19842 15372 19852 15428
rect 19908 15372 20076 15428
rect 20132 15372 20142 15428
rect 1698 15260 1708 15316
rect 1764 15260 3164 15316
rect 3220 15260 5740 15316
rect 5796 15260 5806 15316
rect 6738 15260 6748 15316
rect 6804 15260 7084 15316
rect 7140 15260 7868 15316
rect 7924 15260 7934 15316
rect 10966 15260 11004 15316
rect 11060 15260 11070 15316
rect 12450 15260 12460 15316
rect 12516 15260 15148 15316
rect 15204 15260 15214 15316
rect 17938 15260 17948 15316
rect 18004 15260 19180 15316
rect 19236 15260 19246 15316
rect 2594 15148 2604 15204
rect 2660 15148 3388 15204
rect 3444 15148 3454 15204
rect 6748 15092 6804 15260
rect 7718 15148 7756 15204
rect 7812 15148 7822 15204
rect 9650 15148 9660 15204
rect 9716 15148 13804 15204
rect 13860 15148 13870 15204
rect 17490 15148 17500 15204
rect 17556 15148 18396 15204
rect 18452 15148 18462 15204
rect 20066 15148 20076 15204
rect 20132 15148 21644 15204
rect 21700 15148 21710 15204
rect 28448 15092 28560 15120
rect 4274 15036 4284 15092
rect 4340 15036 6804 15092
rect 12786 15036 12796 15092
rect 12852 15036 15148 15092
rect 17042 15036 17052 15092
rect 17108 15036 21308 15092
rect 21364 15036 22092 15092
rect 22148 15036 22158 15092
rect 22642 15036 22652 15092
rect 22708 15036 23324 15092
rect 23380 15036 23390 15092
rect 24210 15036 24220 15092
rect 24276 15036 28560 15092
rect 15092 14980 15148 15036
rect 28448 15008 28560 15036
rect 7074 14924 7084 14980
rect 7140 14924 7756 14980
rect 7812 14924 7822 14980
rect 14326 14924 14364 14980
rect 14420 14924 14430 14980
rect 15092 14924 24220 14980
rect 24276 14924 24286 14980
rect 0 14868 112 14896
rect 4454 14868 4464 14924
rect 4520 14868 4568 14924
rect 4624 14868 4672 14924
rect 4728 14868 4738 14924
rect 24454 14868 24464 14924
rect 24520 14868 24568 14924
rect 24624 14868 24672 14924
rect 24728 14868 24738 14924
rect 0 14812 2436 14868
rect 6178 14812 6188 14868
rect 6244 14812 9324 14868
rect 9380 14812 9390 14868
rect 13794 14812 13804 14868
rect 13860 14812 22540 14868
rect 22596 14812 23324 14868
rect 23380 14812 23390 14868
rect 0 14784 112 14812
rect 2380 14756 2436 14812
rect 2380 14700 6412 14756
rect 6468 14700 6478 14756
rect 7634 14700 7644 14756
rect 7700 14700 9100 14756
rect 9156 14700 9166 14756
rect 9986 14700 9996 14756
rect 10052 14700 10062 14756
rect 16818 14700 16828 14756
rect 16884 14700 18508 14756
rect 18564 14700 18574 14756
rect 19954 14700 19964 14756
rect 20020 14700 20860 14756
rect 20916 14700 20926 14756
rect 6850 14588 6860 14644
rect 6916 14588 7868 14644
rect 7924 14588 8876 14644
rect 8932 14588 8942 14644
rect 1362 14476 1372 14532
rect 1428 14476 1596 14532
rect 1652 14476 1662 14532
rect 4162 14476 4172 14532
rect 4228 14476 6748 14532
rect 6804 14476 6814 14532
rect 8194 14476 8204 14532
rect 8260 14476 8764 14532
rect 8820 14476 8830 14532
rect 8390 14364 8428 14420
rect 8484 14364 8494 14420
rect 9996 14308 10052 14700
rect 28448 14644 28560 14672
rect 14690 14588 14700 14644
rect 14756 14588 17276 14644
rect 17332 14588 18620 14644
rect 18676 14588 19180 14644
rect 19236 14588 19246 14644
rect 23762 14588 23772 14644
rect 23828 14588 24780 14644
rect 24836 14588 25004 14644
rect 25060 14588 25070 14644
rect 26852 14588 28560 14644
rect 16706 14476 16716 14532
rect 16772 14476 17948 14532
rect 18004 14476 18014 14532
rect 18498 14476 18508 14532
rect 18564 14476 18844 14532
rect 18900 14476 18910 14532
rect 19842 14476 19852 14532
rect 19908 14476 19964 14532
rect 20020 14476 22876 14532
rect 22932 14476 22942 14532
rect 23538 14476 23548 14532
rect 23604 14476 24668 14532
rect 24724 14476 24734 14532
rect 14690 14364 14700 14420
rect 14756 14364 15036 14420
rect 15092 14364 15102 14420
rect 16818 14364 16828 14420
rect 16884 14364 18284 14420
rect 18340 14364 20748 14420
rect 20804 14364 21084 14420
rect 21140 14364 23660 14420
rect 23716 14364 24332 14420
rect 24388 14364 24398 14420
rect 26852 14308 26908 14588
rect 28448 14560 28560 14588
rect 3490 14252 3500 14308
rect 3556 14252 3668 14308
rect 4722 14252 4732 14308
rect 4788 14252 7308 14308
rect 7364 14252 7374 14308
rect 8194 14252 8204 14308
rect 8260 14252 8652 14308
rect 8708 14252 8718 14308
rect 9874 14252 9884 14308
rect 9940 14252 10052 14308
rect 12114 14252 12124 14308
rect 12180 14252 19964 14308
rect 20020 14252 20030 14308
rect 23492 14252 26908 14308
rect 0 13972 112 14000
rect 3612 13972 3668 14252
rect 23492 14196 23548 14252
rect 28448 14196 28560 14224
rect 7298 14140 7308 14196
rect 7364 14140 12572 14196
rect 12628 14140 12638 14196
rect 13122 14140 13132 14196
rect 13188 14140 13468 14196
rect 13524 14140 13534 14196
rect 14466 14140 14476 14196
rect 14532 14140 23548 14196
rect 24210 14140 24220 14196
rect 24276 14140 28560 14196
rect 3794 14084 3804 14140
rect 3860 14084 3908 14140
rect 3964 14084 4012 14140
rect 4068 14084 4078 14140
rect 23794 14084 23804 14140
rect 23860 14084 23908 14140
rect 23964 14084 24012 14140
rect 24068 14084 24078 14140
rect 28448 14112 28560 14140
rect 4162 14028 4172 14084
rect 4228 14028 15260 14084
rect 15316 14028 15326 14084
rect 17154 14028 17164 14084
rect 17220 14028 19068 14084
rect 19124 14028 19134 14084
rect 19506 14028 19516 14084
rect 19572 14028 20972 14084
rect 21028 14028 21420 14084
rect 21476 14028 21486 14084
rect 4172 13972 4228 14028
rect 0 13916 1372 13972
rect 1428 13916 1438 13972
rect 3612 13916 3724 13972
rect 3780 13916 3790 13972
rect 3938 13916 3948 13972
rect 4004 13916 4228 13972
rect 4386 13916 4396 13972
rect 4452 13916 14252 13972
rect 14308 13916 14318 13972
rect 16594 13916 16604 13972
rect 16660 13916 17388 13972
rect 17444 13916 17454 13972
rect 17602 13916 17612 13972
rect 17668 13916 17724 13972
rect 17780 13916 17790 13972
rect 23650 13916 23660 13972
rect 23716 13916 23726 13972
rect 0 13888 112 13916
rect 23660 13860 23716 13916
rect 7298 13804 7308 13860
rect 7364 13804 14924 13860
rect 14980 13804 14990 13860
rect 15250 13804 15260 13860
rect 15316 13804 23716 13860
rect 24770 13804 24780 13860
rect 24836 13804 24846 13860
rect 24780 13748 24836 13804
rect 28448 13748 28560 13776
rect 3602 13692 3612 13748
rect 3668 13692 6972 13748
rect 7028 13692 7038 13748
rect 8530 13692 8540 13748
rect 8596 13692 9324 13748
rect 9380 13692 9390 13748
rect 10070 13692 10108 13748
rect 10164 13692 10174 13748
rect 14802 13692 14812 13748
rect 14868 13692 15428 13748
rect 18386 13692 18396 13748
rect 18452 13692 19516 13748
rect 19572 13692 19582 13748
rect 20850 13692 20860 13748
rect 20916 13692 21420 13748
rect 21476 13692 21644 13748
rect 21700 13692 21710 13748
rect 24210 13692 24220 13748
rect 24276 13692 25340 13748
rect 25396 13692 25406 13748
rect 26002 13692 26012 13748
rect 26068 13692 28560 13748
rect 15372 13636 15428 13692
rect 28448 13664 28560 13692
rect 3378 13580 3388 13636
rect 3444 13580 4956 13636
rect 5012 13580 5022 13636
rect 6738 13580 6748 13636
rect 6804 13580 8764 13636
rect 8820 13580 8830 13636
rect 8978 13580 8988 13636
rect 9044 13580 9082 13636
rect 13794 13580 13804 13636
rect 13860 13580 15148 13636
rect 15204 13580 15214 13636
rect 15372 13580 17836 13636
rect 17892 13580 18284 13636
rect 18340 13580 18350 13636
rect 19954 13580 19964 13636
rect 20020 13580 20972 13636
rect 21028 13580 21038 13636
rect 5842 13468 5852 13524
rect 5908 13468 6636 13524
rect 6692 13468 6702 13524
rect 7410 13468 7420 13524
rect 7476 13468 8204 13524
rect 8260 13468 10108 13524
rect 10164 13468 11340 13524
rect 11396 13468 11406 13524
rect 13458 13468 13468 13524
rect 13524 13468 15036 13524
rect 15092 13468 15102 13524
rect 19730 13468 19740 13524
rect 19796 13468 20748 13524
rect 20804 13468 20814 13524
rect 20972 13468 21308 13524
rect 21364 13468 21374 13524
rect 20972 13412 21028 13468
rect 9090 13356 9100 13412
rect 9156 13356 13580 13412
rect 13636 13356 13646 13412
rect 20850 13356 20860 13412
rect 20916 13356 21028 13412
rect 4454 13300 4464 13356
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4728 13300 4738 13356
rect 24454 13300 24464 13356
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24728 13300 24738 13356
rect 28448 13300 28560 13328
rect 10658 13244 10668 13300
rect 10724 13244 11004 13300
rect 11060 13244 11070 13300
rect 12898 13244 12908 13300
rect 12964 13244 17164 13300
rect 17220 13244 17612 13300
rect 17668 13244 17678 13300
rect 26852 13244 28560 13300
rect 26852 13188 26908 13244
rect 28448 13216 28560 13244
rect 2258 13132 2268 13188
rect 2324 13132 4620 13188
rect 4676 13132 4686 13188
rect 4946 13132 4956 13188
rect 5012 13132 14924 13188
rect 14980 13132 14990 13188
rect 20962 13132 20972 13188
rect 21028 13132 26908 13188
rect 0 13076 112 13104
rect 0 13020 2940 13076
rect 2996 13020 3006 13076
rect 3126 13020 3164 13076
rect 3220 13020 3230 13076
rect 11442 13020 11452 13076
rect 11508 13020 12572 13076
rect 12628 13020 12638 13076
rect 20178 13020 20188 13076
rect 20244 13020 20636 13076
rect 20692 13020 20702 13076
rect 0 12992 112 13020
rect 7186 12908 7196 12964
rect 7252 12908 7756 12964
rect 7812 12908 7822 12964
rect 10546 12908 10556 12964
rect 10612 12908 11564 12964
rect 11620 12908 11630 12964
rect 13458 12908 13468 12964
rect 13524 12908 14028 12964
rect 14084 12908 14364 12964
rect 14420 12908 14430 12964
rect 16034 12908 16044 12964
rect 16100 12908 17388 12964
rect 17444 12908 18396 12964
rect 18452 12908 18462 12964
rect 28448 12852 28560 12880
rect 5730 12796 5740 12852
rect 5796 12796 19628 12852
rect 19684 12796 19694 12852
rect 26852 12796 28560 12852
rect 26852 12740 26908 12796
rect 28448 12768 28560 12796
rect 7410 12684 7420 12740
rect 7476 12684 7868 12740
rect 7924 12684 7934 12740
rect 8194 12684 8204 12740
rect 8260 12684 9324 12740
rect 9380 12684 9390 12740
rect 13682 12684 13692 12740
rect 13748 12684 26908 12740
rect 8306 12572 8316 12628
rect 8372 12572 13412 12628
rect 18946 12572 18956 12628
rect 19012 12572 19292 12628
rect 19348 12572 19358 12628
rect 19506 12572 19516 12628
rect 19572 12572 20188 12628
rect 20244 12572 20254 12628
rect 3794 12516 3804 12572
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 4068 12516 4078 12572
rect 10070 12460 10108 12516
rect 10164 12460 10174 12516
rect 11890 12460 11900 12516
rect 11956 12460 12572 12516
rect 12628 12460 12638 12516
rect 13356 12404 13412 12572
rect 23794 12516 23804 12572
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 24068 12516 24078 12572
rect 13570 12460 13580 12516
rect 13636 12460 20972 12516
rect 21028 12460 21038 12516
rect 28448 12404 28560 12432
rect 6962 12348 6972 12404
rect 7028 12348 9436 12404
rect 9492 12348 12236 12404
rect 12292 12348 12302 12404
rect 13356 12348 28560 12404
rect 28448 12320 28560 12348
rect 3714 12236 3724 12292
rect 3780 12236 4956 12292
rect 5012 12236 5022 12292
rect 11862 12236 11900 12292
rect 11956 12236 11966 12292
rect 16146 12236 16156 12292
rect 16212 12236 17612 12292
rect 17668 12236 19628 12292
rect 19684 12236 19694 12292
rect 23090 12236 23100 12292
rect 23156 12236 23436 12292
rect 23492 12236 23502 12292
rect 0 12180 112 12208
rect 0 12124 812 12180
rect 868 12124 878 12180
rect 2146 12124 2156 12180
rect 2212 12124 2604 12180
rect 2660 12124 5516 12180
rect 5572 12124 5582 12180
rect 14018 12124 14028 12180
rect 14084 12124 14812 12180
rect 14868 12124 14878 12180
rect 16482 12124 16492 12180
rect 16548 12124 18508 12180
rect 18564 12124 19964 12180
rect 20020 12124 20030 12180
rect 20850 12124 20860 12180
rect 20916 12124 21532 12180
rect 21588 12124 21598 12180
rect 0 12096 112 12124
rect 2482 12012 2492 12068
rect 2548 12012 5628 12068
rect 5684 12012 5694 12068
rect 8530 12012 8540 12068
rect 8596 12012 8988 12068
rect 9044 12012 9054 12068
rect 17714 12012 17724 12068
rect 17780 12012 18060 12068
rect 18116 12012 18126 12068
rect 18508 12012 24108 12068
rect 24164 12012 24174 12068
rect 18508 11956 18564 12012
rect 28448 11956 28560 11984
rect 2492 11900 2716 11956
rect 2772 11900 2782 11956
rect 4162 11900 4172 11956
rect 4228 11900 6748 11956
rect 6804 11900 6814 11956
rect 9314 11900 9324 11956
rect 9380 11900 9884 11956
rect 9940 11900 9950 11956
rect 11078 11900 11116 11956
rect 11172 11900 11182 11956
rect 15092 11900 18508 11956
rect 18564 11900 18574 11956
rect 18722 11900 18732 11956
rect 18788 11900 18798 11956
rect 19730 11900 19740 11956
rect 19796 11900 21084 11956
rect 21140 11900 21150 11956
rect 24994 11900 25004 11956
rect 25060 11900 28560 11956
rect 2492 11844 2548 11900
rect 15092 11844 15148 11900
rect 2482 11788 2492 11844
rect 2548 11788 2558 11844
rect 5506 11788 5516 11844
rect 5572 11788 5964 11844
rect 6020 11788 6300 11844
rect 6356 11788 6366 11844
rect 7298 11788 7308 11844
rect 7364 11788 8428 11844
rect 8484 11788 8764 11844
rect 8820 11788 15148 11844
rect 4454 11732 4464 11788
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4728 11732 4738 11788
rect 7308 11732 7364 11788
rect 18732 11732 18788 11900
rect 28448 11872 28560 11900
rect 19506 11788 19516 11844
rect 19572 11788 20636 11844
rect 20692 11788 20702 11844
rect 24454 11732 24464 11788
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24728 11732 24738 11788
rect 1810 11676 1820 11732
rect 1876 11676 2044 11732
rect 2100 11676 3276 11732
rect 3332 11676 3342 11732
rect 6514 11676 6524 11732
rect 6580 11676 7364 11732
rect 11106 11676 11116 11732
rect 11172 11676 13020 11732
rect 13076 11676 13086 11732
rect 15586 11676 15596 11732
rect 15652 11676 16940 11732
rect 16996 11676 17006 11732
rect 17602 11676 17612 11732
rect 17668 11676 18788 11732
rect 1586 11564 1596 11620
rect 1652 11564 2268 11620
rect 2324 11564 2334 11620
rect 3332 11564 20804 11620
rect 23202 11564 23212 11620
rect 23268 11564 23772 11620
rect 23828 11564 23838 11620
rect 3332 11396 3388 11564
rect 20748 11508 20804 11564
rect 28448 11508 28560 11536
rect 3602 11452 3612 11508
rect 3668 11452 5068 11508
rect 5124 11452 5134 11508
rect 8194 11452 8204 11508
rect 8260 11452 9212 11508
rect 9268 11452 9278 11508
rect 9874 11452 9884 11508
rect 9940 11452 12908 11508
rect 12964 11452 12974 11508
rect 18246 11452 18284 11508
rect 18340 11452 18350 11508
rect 18834 11452 18844 11508
rect 18900 11452 19404 11508
rect 19460 11452 19470 11508
rect 20748 11452 26348 11508
rect 26404 11452 26414 11508
rect 26852 11452 28560 11508
rect 8204 11396 8260 11452
rect 2258 11340 2268 11396
rect 2324 11340 3388 11396
rect 4274 11340 4284 11396
rect 4340 11340 6188 11396
rect 6244 11340 6254 11396
rect 6626 11340 6636 11396
rect 6692 11340 8260 11396
rect 11106 11340 11116 11396
rect 11172 11340 11452 11396
rect 11508 11340 11518 11396
rect 12674 11340 12684 11396
rect 12740 11340 13020 11396
rect 13076 11340 13086 11396
rect 17266 11340 17276 11396
rect 17332 11340 18396 11396
rect 18452 11340 19180 11396
rect 19236 11340 19246 11396
rect 19954 11340 19964 11396
rect 20020 11340 21196 11396
rect 21252 11340 21262 11396
rect 0 11284 112 11312
rect 7084 11284 7140 11340
rect 26852 11284 26908 11452
rect 28448 11424 28560 11452
rect 0 11228 3052 11284
rect 3108 11228 3118 11284
rect 3266 11228 3276 11284
rect 3332 11228 6748 11284
rect 6804 11228 6814 11284
rect 7074 11228 7084 11284
rect 7140 11228 7150 11284
rect 9538 11228 9548 11284
rect 9604 11228 26908 11284
rect 0 11200 112 11228
rect 3276 11116 7644 11172
rect 7700 11116 7710 11172
rect 8642 11116 8652 11172
rect 8708 11116 16268 11172
rect 16324 11116 16334 11172
rect 16716 11116 26908 11172
rect 3276 11060 3332 11116
rect 16716 11060 16772 11116
rect 26852 11060 26908 11116
rect 28448 11060 28560 11088
rect 3266 11004 3276 11060
rect 3332 11004 3342 11060
rect 9062 11004 9100 11060
rect 9156 11004 9166 11060
rect 12002 11004 12012 11060
rect 12068 11004 12796 11060
rect 12852 11004 12862 11060
rect 13010 11004 13020 11060
rect 13076 11004 13748 11060
rect 15474 11004 15484 11060
rect 15540 11004 16772 11060
rect 17042 11004 17052 11060
rect 17108 11004 18956 11060
rect 19012 11004 19022 11060
rect 26852 11004 28560 11060
rect 3794 10948 3804 11004
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 4068 10948 4078 11004
rect 7186 10892 7196 10948
rect 7252 10892 7756 10948
rect 7812 10892 7822 10948
rect 8754 10892 8764 10948
rect 8820 10892 9212 10948
rect 9268 10892 9278 10948
rect 10882 10892 10892 10948
rect 10948 10892 11564 10948
rect 11620 10892 11630 10948
rect 5170 10780 5180 10836
rect 5236 10780 8260 10836
rect 11106 10780 11116 10836
rect 11172 10780 11340 10836
rect 11396 10780 13244 10836
rect 13300 10780 13310 10836
rect 8204 10724 8260 10780
rect 2594 10668 2604 10724
rect 2660 10668 7980 10724
rect 8036 10668 8046 10724
rect 8194 10668 8204 10724
rect 8260 10668 8764 10724
rect 8820 10668 8830 10724
rect 10098 10668 10108 10724
rect 10164 10668 10668 10724
rect 10724 10668 10734 10724
rect 13692 10612 13748 11004
rect 23794 10948 23804 11004
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 24068 10948 24078 11004
rect 28448 10976 28560 11004
rect 18722 10892 18732 10948
rect 18788 10892 20076 10948
rect 20132 10892 20142 10948
rect 18274 10780 18284 10836
rect 18340 10780 19628 10836
rect 19684 10780 21308 10836
rect 21364 10780 21374 10836
rect 14802 10668 14812 10724
rect 14868 10668 19964 10724
rect 20020 10668 22988 10724
rect 23044 10668 23054 10724
rect 28448 10612 28560 10640
rect 2034 10556 2044 10612
rect 2100 10556 6524 10612
rect 6580 10556 6590 10612
rect 7858 10556 7868 10612
rect 7924 10556 9436 10612
rect 9492 10556 9502 10612
rect 11442 10556 11452 10612
rect 11508 10556 12348 10612
rect 12404 10556 12414 10612
rect 13692 10556 15148 10612
rect 18274 10556 18284 10612
rect 18340 10556 18620 10612
rect 18676 10556 18686 10612
rect 22642 10556 22652 10612
rect 22708 10556 28560 10612
rect 15092 10500 15148 10556
rect 28448 10528 28560 10556
rect 6738 10444 6748 10500
rect 6804 10444 7756 10500
rect 7812 10444 9660 10500
rect 9716 10444 9726 10500
rect 11004 10444 11564 10500
rect 11620 10444 11630 10500
rect 12226 10444 12236 10500
rect 12292 10444 13020 10500
rect 13076 10444 13086 10500
rect 15092 10444 19404 10500
rect 19460 10444 25116 10500
rect 25172 10444 25182 10500
rect 0 10388 112 10416
rect 0 10332 3164 10388
rect 3220 10332 3230 10388
rect 7074 10332 7084 10388
rect 7140 10332 7644 10388
rect 7700 10332 7710 10388
rect 8082 10332 8092 10388
rect 8148 10332 9548 10388
rect 9604 10332 9614 10388
rect 0 10304 112 10332
rect 11004 10276 11060 10444
rect 11218 10332 11228 10388
rect 11284 10332 13692 10388
rect 13748 10332 13758 10388
rect 15586 10332 15596 10388
rect 15652 10332 17612 10388
rect 17668 10332 17678 10388
rect 6178 10220 6188 10276
rect 6244 10220 8204 10276
rect 8260 10220 11060 10276
rect 4454 10164 4464 10220
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4728 10164 4738 10220
rect 24454 10164 24464 10220
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24728 10164 24738 10220
rect 28448 10164 28560 10192
rect 6962 10108 6972 10164
rect 7028 10108 7038 10164
rect 10098 10108 10108 10164
rect 10164 10108 10174 10164
rect 11666 10108 11676 10164
rect 11732 10108 15148 10164
rect 15204 10108 16044 10164
rect 16100 10108 16110 10164
rect 16258 10108 16268 10164
rect 16324 10108 18172 10164
rect 18228 10108 19404 10164
rect 19460 10108 19470 10164
rect 19618 10108 19628 10164
rect 19684 10108 19852 10164
rect 19908 10108 19918 10164
rect 24882 10108 24892 10164
rect 24948 10108 28560 10164
rect 6972 10052 7028 10108
rect 10108 10052 10164 10108
rect 28448 10080 28560 10108
rect 2482 9996 2492 10052
rect 2548 9996 5404 10052
rect 5460 9996 5470 10052
rect 6738 9996 6748 10052
rect 6804 9996 7028 10052
rect 9762 9996 9772 10052
rect 9828 9996 10164 10052
rect 11106 9996 11116 10052
rect 11172 9996 11452 10052
rect 11508 9996 11518 10052
rect 11890 9996 11900 10052
rect 11956 9996 12124 10052
rect 12180 9996 13132 10052
rect 13188 9996 13198 10052
rect 13682 9996 13692 10052
rect 13748 9996 15036 10052
rect 15092 9996 15102 10052
rect 16482 9996 16492 10052
rect 16548 9996 17276 10052
rect 17332 9996 17342 10052
rect 17826 9996 17836 10052
rect 17892 9996 18956 10052
rect 19012 9996 19022 10052
rect 20850 9996 20860 10052
rect 20916 9996 22092 10052
rect 22148 9996 22158 10052
rect 6514 9884 6524 9940
rect 6580 9884 6972 9940
rect 7028 9884 7532 9940
rect 7588 9884 8988 9940
rect 9044 9884 9054 9940
rect 12226 9884 12236 9940
rect 12292 9884 16156 9940
rect 16212 9884 17948 9940
rect 18004 9884 18014 9940
rect 20860 9828 20916 9996
rect 7858 9772 7868 9828
rect 7924 9772 8876 9828
rect 8932 9772 8942 9828
rect 13122 9772 13132 9828
rect 13188 9772 13804 9828
rect 13860 9772 13870 9828
rect 15250 9772 15260 9828
rect 15316 9772 17052 9828
rect 17108 9772 17118 9828
rect 17266 9772 17276 9828
rect 17332 9772 20916 9828
rect 28448 9716 28560 9744
rect 3826 9660 3836 9716
rect 3892 9660 16940 9716
rect 16996 9660 17006 9716
rect 17938 9660 17948 9716
rect 18004 9660 19516 9716
rect 19572 9660 19582 9716
rect 26852 9660 28560 9716
rect 26852 9604 26908 9660
rect 28448 9632 28560 9660
rect 11330 9548 11340 9604
rect 11396 9548 26908 9604
rect 0 9492 112 9520
rect 0 9436 2716 9492
rect 2772 9436 2782 9492
rect 10546 9436 10556 9492
rect 10612 9436 10892 9492
rect 10948 9436 15148 9492
rect 15362 9436 15372 9492
rect 15428 9436 15708 9492
rect 15764 9436 16604 9492
rect 16660 9436 16670 9492
rect 0 9408 112 9436
rect 3794 9380 3804 9436
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 4068 9380 4078 9436
rect 15092 9380 15148 9436
rect 23794 9380 23804 9436
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 24068 9380 24078 9436
rect 12114 9324 12124 9380
rect 12180 9324 12348 9380
rect 12404 9324 14028 9380
rect 14084 9324 14094 9380
rect 15092 9324 18172 9380
rect 18228 9324 18238 9380
rect 28448 9268 28560 9296
rect 690 9212 700 9268
rect 756 9212 1260 9268
rect 1316 9212 1326 9268
rect 9314 9212 9324 9268
rect 9380 9212 10556 9268
rect 10612 9212 12460 9268
rect 12516 9212 12796 9268
rect 12852 9212 12862 9268
rect 13794 9212 13804 9268
rect 13860 9212 14812 9268
rect 14868 9212 14878 9268
rect 15092 9212 17164 9268
rect 17220 9212 17230 9268
rect 21970 9212 21980 9268
rect 22036 9212 25564 9268
rect 25620 9212 25630 9268
rect 26852 9212 28560 9268
rect 15092 9156 15148 9212
rect 26852 9156 26908 9212
rect 28448 9184 28560 9212
rect 6374 9100 6412 9156
rect 6468 9100 6478 9156
rect 7410 9100 7420 9156
rect 7476 9100 9884 9156
rect 9940 9100 9950 9156
rect 11554 9100 11564 9156
rect 11620 9100 15148 9156
rect 15810 9100 15820 9156
rect 15876 9100 16044 9156
rect 16100 9100 26908 9156
rect 2034 8988 2044 9044
rect 2100 8988 21868 9044
rect 21924 8988 21934 9044
rect 6738 8876 6748 8932
rect 6804 8876 7308 8932
rect 7364 8876 17724 8932
rect 17780 8876 19292 8932
rect 19348 8876 19628 8932
rect 19684 8876 19694 8932
rect 28448 8820 28560 8848
rect 1820 8764 2380 8820
rect 2436 8764 2446 8820
rect 13244 8764 15372 8820
rect 15428 8764 15438 8820
rect 20066 8764 20076 8820
rect 20132 8764 28560 8820
rect 0 8596 112 8624
rect 0 8540 1596 8596
rect 1652 8540 1662 8596
rect 0 8512 112 8540
rect 1820 8428 1876 8764
rect 13244 8708 13300 8764
rect 28448 8736 28560 8764
rect 2156 8652 2604 8708
rect 2660 8652 2670 8708
rect 7186 8652 7196 8708
rect 7252 8652 8540 8708
rect 8596 8652 9772 8708
rect 9828 8652 13300 8708
rect 2156 8428 2212 8652
rect 4454 8596 4464 8652
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4728 8596 4738 8652
rect 24454 8596 24464 8652
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24728 8596 24738 8652
rect 8082 8540 8092 8596
rect 8148 8540 9324 8596
rect 9380 8540 11452 8596
rect 11508 8540 12852 8596
rect 12796 8484 12852 8540
rect 8418 8428 8428 8484
rect 8484 8428 10220 8484
rect 10276 8428 10286 8484
rect 12786 8428 12796 8484
rect 12852 8428 13132 8484
rect 13188 8428 13198 8484
rect 13906 8428 13916 8484
rect 13972 8428 14924 8484
rect 14980 8428 14990 8484
rect 21074 8428 21084 8484
rect 21140 8428 21252 8484
rect 1810 8372 1820 8428
rect 1876 8372 1886 8428
rect 2146 8372 2156 8428
rect 2212 8372 2222 8428
rect 21196 8372 21252 8428
rect 28448 8372 28560 8400
rect 6290 8316 6300 8372
rect 6356 8316 6748 8372
rect 6804 8316 10108 8372
rect 10164 8316 10174 8372
rect 10322 8316 10332 8372
rect 10388 8316 11116 8372
rect 11172 8316 11182 8372
rect 15092 8316 16716 8372
rect 16772 8316 16782 8372
rect 17826 8316 17836 8372
rect 17892 8316 18508 8372
rect 18564 8316 18574 8372
rect 20178 8316 20188 8372
rect 20244 8316 20972 8372
rect 21028 8316 21038 8372
rect 21196 8316 21308 8372
rect 21364 8316 22316 8372
rect 22372 8316 22540 8372
rect 22596 8316 22606 8372
rect 26852 8316 28560 8372
rect 15092 8260 15148 8316
rect 26852 8260 26908 8316
rect 28448 8288 28560 8316
rect 3602 8204 3612 8260
rect 3668 8204 15148 8260
rect 15474 8204 15484 8260
rect 15540 8204 16940 8260
rect 16996 8204 17006 8260
rect 17164 8204 18844 8260
rect 18900 8204 18910 8260
rect 19618 8204 19628 8260
rect 19684 8204 26908 8260
rect 17164 8148 17220 8204
rect 3826 8092 3836 8148
rect 3892 8092 7588 8148
rect 7746 8092 7756 8148
rect 7812 8092 15932 8148
rect 15988 8092 15998 8148
rect 16156 8092 17220 8148
rect 2258 7980 2268 8036
rect 2324 7980 5068 8036
rect 5124 7980 5134 8036
rect 7532 7924 7588 8092
rect 16156 8036 16212 8092
rect 13458 7980 13468 8036
rect 13524 7980 15596 8036
rect 15652 7980 16212 8036
rect 18834 7980 18844 8036
rect 18900 7980 20300 8036
rect 20356 7980 20366 8036
rect 21186 7980 21196 8036
rect 21252 7980 26908 8036
rect 26852 7924 26908 7980
rect 28448 7924 28560 7952
rect 7532 7868 19740 7924
rect 19796 7868 19806 7924
rect 19954 7868 19964 7924
rect 20020 7868 21756 7924
rect 21812 7868 21822 7924
rect 26852 7868 28560 7924
rect 3794 7812 3804 7868
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 4068 7812 4078 7868
rect 23794 7812 23804 7868
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 24068 7812 24078 7868
rect 28448 7840 28560 7868
rect 7074 7756 7084 7812
rect 7140 7756 14252 7812
rect 14308 7756 16604 7812
rect 16660 7756 17052 7812
rect 17108 7756 17118 7812
rect 0 7700 112 7728
rect 0 7644 1708 7700
rect 1764 7644 1774 7700
rect 12226 7644 12236 7700
rect 12292 7644 13244 7700
rect 13300 7644 13310 7700
rect 16706 7644 16716 7700
rect 16772 7644 17388 7700
rect 17444 7644 17454 7700
rect 21858 7644 21868 7700
rect 21924 7644 26124 7700
rect 26180 7644 26190 7700
rect 0 7616 112 7644
rect 7270 7532 7308 7588
rect 7364 7532 7374 7588
rect 15586 7532 15596 7588
rect 15652 7532 16380 7588
rect 16436 7532 16446 7588
rect 28448 7476 28560 7504
rect 3826 7420 3836 7476
rect 3892 7420 13580 7476
rect 13636 7420 13646 7476
rect 14578 7420 14588 7476
rect 14644 7420 15484 7476
rect 15540 7420 16156 7476
rect 16212 7420 16222 7476
rect 16930 7420 16940 7476
rect 16996 7420 17388 7476
rect 17444 7420 21308 7476
rect 21364 7420 21374 7476
rect 22082 7420 22092 7476
rect 22148 7420 28560 7476
rect 28448 7392 28560 7420
rect 9762 7308 9772 7364
rect 9828 7308 10444 7364
rect 10500 7308 11004 7364
rect 11060 7308 11070 7364
rect 12226 7308 12236 7364
rect 12292 7308 13356 7364
rect 13412 7308 13422 7364
rect 14914 7308 14924 7364
rect 14980 7308 15596 7364
rect 15652 7308 15662 7364
rect 16258 7308 16268 7364
rect 16324 7308 22764 7364
rect 22820 7308 22830 7364
rect 11218 7196 11228 7252
rect 11284 7196 15708 7252
rect 15764 7196 19964 7252
rect 20020 7196 20030 7252
rect 20290 7196 20300 7252
rect 20356 7196 26908 7252
rect 4454 7028 4464 7084
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4728 7028 4738 7084
rect 24454 7028 24464 7084
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 24728 7028 24738 7084
rect 26852 7028 26908 7196
rect 28448 7028 28560 7056
rect 26852 6972 28560 7028
rect 28448 6944 28560 6972
rect 914 6860 924 6916
rect 980 6860 2044 6916
rect 2100 6860 2110 6916
rect 2370 6860 2380 6916
rect 2436 6860 22652 6916
rect 22708 6860 22718 6916
rect 0 6804 112 6832
rect 0 6748 1484 6804
rect 1540 6748 1550 6804
rect 6066 6748 6076 6804
rect 6132 6748 7756 6804
rect 7812 6748 7822 6804
rect 10994 6748 11004 6804
rect 11060 6748 12684 6804
rect 12740 6748 12750 6804
rect 20850 6748 20860 6804
rect 20916 6748 27132 6804
rect 27188 6748 27198 6804
rect 0 6720 112 6748
rect 19506 6636 19516 6692
rect 19572 6636 26572 6692
rect 26628 6636 26638 6692
rect 28448 6580 28560 6608
rect 20962 6524 20972 6580
rect 21028 6524 22428 6580
rect 22484 6524 22494 6580
rect 26852 6524 28560 6580
rect 3042 6412 3052 6468
rect 3108 6412 15764 6468
rect 15922 6412 15932 6468
rect 15988 6412 25788 6468
rect 25844 6412 25854 6468
rect 15708 6356 15764 6412
rect 26852 6356 26908 6524
rect 28448 6496 28560 6524
rect 15708 6300 20860 6356
rect 20916 6300 20926 6356
rect 24220 6300 26908 6356
rect 3794 6244 3804 6300
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 4068 6244 4078 6300
rect 23794 6244 23804 6300
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 24068 6244 24078 6300
rect 9762 6188 9772 6244
rect 9828 6188 21868 6244
rect 21924 6188 21934 6244
rect 24220 6132 24276 6300
rect 28448 6132 28560 6160
rect 2258 6076 2268 6132
rect 2324 6076 14140 6132
rect 14196 6076 14206 6132
rect 21746 6076 21756 6132
rect 21812 6076 24276 6132
rect 24332 6076 28560 6132
rect 24332 6020 24388 6076
rect 28448 6048 28560 6076
rect 3154 5964 3164 6020
rect 3220 5964 16268 6020
rect 16324 5964 16334 6020
rect 19506 5964 19516 6020
rect 19572 5964 24388 6020
rect 0 5908 112 5936
rect 0 5852 2828 5908
rect 2884 5852 2894 5908
rect 11666 5852 11676 5908
rect 11732 5852 13692 5908
rect 13748 5852 13758 5908
rect 15138 5852 15148 5908
rect 15204 5852 26012 5908
rect 26068 5852 26078 5908
rect 0 5824 112 5852
rect 12114 5740 12124 5796
rect 12180 5740 26684 5796
rect 26740 5740 26750 5796
rect 26852 5684 26964 6020
rect 28448 5684 28560 5712
rect 7746 5628 7756 5684
rect 7812 5628 8876 5684
rect 8932 5628 11116 5684
rect 11172 5628 11182 5684
rect 14802 5628 14812 5684
rect 14868 5628 15372 5684
rect 15428 5628 15438 5684
rect 22530 5628 22540 5684
rect 22596 5628 28560 5684
rect 28448 5600 28560 5628
rect 4454 5460 4464 5516
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4728 5460 4738 5516
rect 24454 5460 24464 5516
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24728 5460 24738 5516
rect 9324 5404 17556 5460
rect 9324 5348 9380 5404
rect 3602 5292 3612 5348
rect 3668 5292 9380 5348
rect 12786 5292 12796 5348
rect 12852 5292 15148 5348
rect 15204 5292 15214 5348
rect 8306 5180 8316 5236
rect 8372 5180 9212 5236
rect 9268 5180 9278 5236
rect 17500 5124 17556 5404
rect 28448 5236 28560 5264
rect 17714 5180 17724 5236
rect 17780 5180 28560 5236
rect 28448 5152 28560 5180
rect 17500 5068 27580 5124
rect 27636 5068 27646 5124
rect 0 5012 112 5040
rect 0 4956 1932 5012
rect 1988 4956 1998 5012
rect 0 4928 112 4956
rect 18050 4844 18060 4900
rect 18116 4844 26908 4900
rect 26852 4788 26908 4844
rect 28448 4788 28560 4816
rect 26852 4732 28560 4788
rect 3794 4676 3804 4732
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 4068 4676 4078 4732
rect 23794 4676 23804 4732
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 24068 4676 24078 4732
rect 28448 4704 28560 4732
rect 16818 4508 16828 4564
rect 16884 4508 27020 4564
rect 27076 4508 27086 4564
rect 15474 4396 15484 4452
rect 15540 4396 27020 4452
rect 27076 4396 27086 4452
rect 28448 4340 28560 4368
rect 18834 4284 18844 4340
rect 18900 4284 28560 4340
rect 28448 4256 28560 4284
rect 2258 4172 2268 4228
rect 2324 4172 17500 4228
rect 17556 4172 17566 4228
rect 0 4116 112 4144
rect 0 4060 1484 4116
rect 1540 4060 1550 4116
rect 16930 4060 16940 4116
rect 16996 4060 26908 4116
rect 0 4032 112 4060
rect 4454 3892 4464 3948
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4728 3892 4738 3948
rect 24454 3892 24464 3948
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24728 3892 24738 3948
rect 26852 3892 26908 4060
rect 28448 3892 28560 3920
rect 10098 3836 10108 3892
rect 10164 3836 17948 3892
rect 18004 3836 18014 3892
rect 26852 3836 28560 3892
rect 28448 3808 28560 3836
rect 2258 3500 2268 3556
rect 2324 3500 23100 3556
rect 23156 3500 23166 3556
rect 28448 3444 28560 3472
rect 19058 3388 19068 3444
rect 19124 3388 28560 3444
rect 28448 3360 28560 3388
rect 0 3220 112 3248
rect 0 3164 1260 3220
rect 1316 3164 1326 3220
rect 0 3136 112 3164
rect 3794 3108 3804 3164
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 4068 3108 4078 3164
rect 23794 3108 23804 3164
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 24068 3108 24078 3164
rect 28448 2996 28560 3024
rect 21074 2940 21084 2996
rect 21140 2940 28560 2996
rect 28448 2912 28560 2940
rect 28448 2548 28560 2576
rect 22642 2492 22652 2548
rect 22708 2492 28560 2548
rect 28448 2464 28560 2492
rect 0 2324 112 2352
rect 4454 2324 4464 2380
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4728 2324 4738 2380
rect 24454 2324 24464 2380
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24728 2324 24738 2380
rect 0 2268 1820 2324
rect 1876 2268 1886 2324
rect 0 2240 112 2268
rect 11442 2156 11452 2212
rect 11508 2156 17724 2212
rect 17780 2156 17790 2212
rect 21298 2156 21308 2212
rect 21364 2156 27468 2212
rect 27524 2156 27534 2212
rect 28448 2100 28560 2128
rect 13234 2044 13244 2100
rect 13300 2044 20972 2100
rect 21028 2044 21038 2100
rect 24322 2044 24332 2100
rect 24388 2044 28560 2100
rect 28448 2016 28560 2044
rect 13794 1932 13804 1988
rect 13860 1932 22204 1988
rect 22260 1932 22270 1988
rect 12002 1708 12012 1764
rect 12068 1708 26236 1764
rect 26292 1708 26302 1764
rect 28448 1652 28560 1680
rect 466 1596 476 1652
rect 532 1596 3388 1652
rect 3444 1596 3454 1652
rect 24882 1596 24892 1652
rect 24948 1596 26908 1652
rect 26964 1596 26974 1652
rect 27132 1596 28560 1652
rect 3794 1540 3804 1596
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 4068 1540 4078 1596
rect 23794 1540 23804 1596
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 24068 1540 24078 1596
rect 27132 1428 27188 1596
rect 28448 1568 28560 1596
rect 22530 1372 22540 1428
rect 22596 1372 27188 1428
rect 28448 1204 28560 1232
rect 28354 1148 28364 1204
rect 28420 1148 28560 1204
rect 28448 1120 28560 1148
rect 12114 1036 12124 1092
rect 12180 1036 25956 1092
rect 14130 924 14140 980
rect 14196 924 25676 980
rect 25732 924 25742 980
rect 4454 756 4464 812
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4728 756 4738 812
rect 24454 756 24464 812
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24728 756 24738 812
rect 25900 756 25956 1036
rect 28448 756 28560 784
rect 25900 700 28560 756
rect 28448 672 28560 700
rect 690 588 700 644
rect 756 588 10892 644
rect 10948 588 10958 644
rect 18162 588 18172 644
rect 18228 588 26012 644
rect 26068 588 26078 644
rect 242 476 252 532
rect 308 476 4732 532
rect 4788 476 4798 532
rect 16706 476 16716 532
rect 16772 476 23548 532
rect 23604 476 23614 532
rect 19506 364 19516 420
rect 19572 364 26908 420
rect 26964 364 26974 420
rect 28448 308 28560 336
rect 18498 252 18508 308
rect 18564 252 28560 308
rect 28448 224 28560 252
rect 6850 140 6860 196
rect 6916 140 7420 196
rect 7476 140 7486 196
rect 11442 140 11452 196
rect 11508 140 21980 196
rect 22036 140 22046 196
<< via3 >>
rect 3804 56420 3860 56476
rect 3908 56420 3964 56476
rect 4012 56420 4068 56476
rect 23804 56420 23860 56476
rect 23908 56420 23964 56476
rect 24012 56420 24068 56476
rect 19516 55916 19572 55972
rect 21308 55916 21364 55972
rect 4464 55636 4520 55692
rect 4568 55636 4624 55692
rect 4672 55636 4728 55692
rect 24464 55636 24520 55692
rect 24568 55636 24624 55692
rect 24672 55636 24728 55692
rect 20860 55244 20916 55300
rect 22428 55244 22484 55300
rect 3164 55132 3220 55188
rect 27020 55132 27076 55188
rect 3804 54852 3860 54908
rect 3908 54852 3964 54908
rect 4012 54852 4068 54908
rect 23804 54852 23860 54908
rect 23908 54852 23964 54908
rect 24012 54852 24068 54908
rect 19068 54236 19124 54292
rect 17724 54124 17780 54180
rect 4464 54068 4520 54124
rect 4568 54068 4624 54124
rect 4672 54068 4728 54124
rect 24464 54068 24520 54124
rect 24568 54068 24624 54124
rect 24672 54068 24728 54124
rect 20076 53900 20132 53956
rect 17948 53788 18004 53844
rect 16716 53676 16772 53732
rect 3804 53284 3860 53340
rect 3908 53284 3964 53340
rect 4012 53284 4068 53340
rect 23804 53284 23860 53340
rect 23908 53284 23964 53340
rect 24012 53284 24068 53340
rect 12572 52668 12628 52724
rect 4464 52500 4520 52556
rect 4568 52500 4624 52556
rect 4672 52500 4728 52556
rect 24464 52500 24520 52556
rect 24568 52500 24624 52556
rect 24672 52500 24728 52556
rect 27132 52332 27188 52388
rect 22764 52108 22820 52164
rect 3804 51716 3860 51772
rect 3908 51716 3964 51772
rect 4012 51716 4068 51772
rect 23804 51716 23860 51772
rect 23908 51716 23964 51772
rect 24012 51716 24068 51772
rect 9212 51436 9268 51492
rect 11340 51212 11396 51268
rect 4464 50932 4520 50988
rect 4568 50932 4624 50988
rect 4672 50932 4728 50988
rect 24464 50932 24520 50988
rect 24568 50932 24624 50988
rect 24672 50932 24728 50988
rect 26908 50540 26964 50596
rect 3804 50148 3860 50204
rect 3908 50148 3964 50204
rect 4012 50148 4068 50204
rect 23804 50148 23860 50204
rect 23908 50148 23964 50204
rect 24012 50148 24068 50204
rect 6188 49868 6244 49924
rect 14252 49644 14308 49700
rect 4464 49364 4520 49420
rect 4568 49364 4624 49420
rect 4672 49364 4728 49420
rect 24464 49364 24520 49420
rect 24568 49364 24624 49420
rect 24672 49364 24728 49420
rect 2380 48972 2436 49028
rect 3804 48580 3860 48636
rect 3908 48580 3964 48636
rect 4012 48580 4068 48636
rect 23804 48580 23860 48636
rect 23908 48580 23964 48636
rect 24012 48580 24068 48636
rect 15932 48076 15988 48132
rect 4464 47796 4520 47852
rect 4568 47796 4624 47852
rect 4672 47796 4728 47852
rect 24464 47796 24520 47852
rect 24568 47796 24624 47852
rect 24672 47796 24728 47852
rect 3804 47012 3860 47068
rect 3908 47012 3964 47068
rect 4012 47012 4068 47068
rect 23804 47012 23860 47068
rect 23908 47012 23964 47068
rect 24012 47012 24068 47068
rect 4464 46228 4520 46284
rect 4568 46228 4624 46284
rect 4672 46228 4728 46284
rect 24464 46228 24520 46284
rect 24568 46228 24624 46284
rect 24672 46228 24728 46284
rect 3804 45444 3860 45500
rect 3908 45444 3964 45500
rect 4012 45444 4068 45500
rect 23804 45444 23860 45500
rect 23908 45444 23964 45500
rect 24012 45444 24068 45500
rect 4464 44660 4520 44716
rect 4568 44660 4624 44716
rect 4672 44660 4728 44716
rect 24464 44660 24520 44716
rect 24568 44660 24624 44716
rect 24672 44660 24728 44716
rect 3804 43876 3860 43932
rect 3908 43876 3964 43932
rect 4012 43876 4068 43932
rect 23804 43876 23860 43932
rect 23908 43876 23964 43932
rect 24012 43876 24068 43932
rect 4464 43092 4520 43148
rect 4568 43092 4624 43148
rect 4672 43092 4728 43148
rect 24464 43092 24520 43148
rect 24568 43092 24624 43148
rect 24672 43092 24728 43148
rect 3804 42308 3860 42364
rect 3908 42308 3964 42364
rect 4012 42308 4068 42364
rect 23804 42308 23860 42364
rect 23908 42308 23964 42364
rect 24012 42308 24068 42364
rect 6412 41580 6468 41636
rect 4464 41524 4520 41580
rect 4568 41524 4624 41580
rect 4672 41524 4728 41580
rect 24464 41524 24520 41580
rect 24568 41524 24624 41580
rect 24672 41524 24728 41580
rect 27244 41244 27300 41300
rect 3804 40740 3860 40796
rect 3908 40740 3964 40796
rect 4012 40740 4068 40796
rect 23804 40740 23860 40796
rect 23908 40740 23964 40796
rect 24012 40740 24068 40796
rect 4464 39956 4520 40012
rect 4568 39956 4624 40012
rect 4672 39956 4728 40012
rect 24464 39956 24520 40012
rect 24568 39956 24624 40012
rect 24672 39956 24728 40012
rect 10444 39228 10500 39284
rect 3804 39172 3860 39228
rect 3908 39172 3964 39228
rect 4012 39172 4068 39228
rect 23804 39172 23860 39228
rect 23908 39172 23964 39228
rect 24012 39172 24068 39228
rect 4464 38388 4520 38444
rect 4568 38388 4624 38444
rect 4672 38388 4728 38444
rect 24464 38388 24520 38444
rect 24568 38388 24624 38444
rect 24672 38388 24728 38444
rect 27356 37772 27412 37828
rect 1820 37660 1876 37716
rect 3804 37604 3860 37660
rect 3908 37604 3964 37660
rect 4012 37604 4068 37660
rect 23804 37604 23860 37660
rect 23908 37604 23964 37660
rect 24012 37604 24068 37660
rect 8092 37100 8148 37156
rect 8540 37100 8596 37156
rect 4464 36820 4520 36876
rect 4568 36820 4624 36876
rect 4672 36820 4728 36876
rect 24464 36820 24520 36876
rect 24568 36820 24624 36876
rect 24672 36820 24728 36876
rect 1820 36204 1876 36260
rect 3804 36036 3860 36092
rect 3908 36036 3964 36092
rect 4012 36036 4068 36092
rect 23804 36036 23860 36092
rect 23908 36036 23964 36092
rect 24012 36036 24068 36092
rect 4464 35252 4520 35308
rect 4568 35252 4624 35308
rect 4672 35252 4728 35308
rect 24464 35252 24520 35308
rect 24568 35252 24624 35308
rect 24672 35252 24728 35308
rect 10892 34860 10948 34916
rect 4844 34636 4900 34692
rect 18396 34636 18452 34692
rect 3804 34468 3860 34524
rect 3908 34468 3964 34524
rect 4012 34468 4068 34524
rect 23804 34468 23860 34524
rect 23908 34468 23964 34524
rect 24012 34468 24068 34524
rect 9100 34412 9156 34468
rect 4284 34188 4340 34244
rect 13580 34076 13636 34132
rect 8204 33964 8260 34020
rect 8988 33740 9044 33796
rect 4464 33684 4520 33740
rect 4568 33684 4624 33740
rect 4672 33684 4728 33740
rect 24464 33684 24520 33740
rect 24568 33684 24624 33740
rect 24672 33684 24728 33740
rect 4284 33628 4340 33684
rect 8204 33180 8260 33236
rect 3804 32900 3860 32956
rect 3908 32900 3964 32956
rect 4012 32900 4068 32956
rect 23804 32900 23860 32956
rect 23908 32900 23964 32956
rect 24012 32900 24068 32956
rect 12348 32844 12404 32900
rect 11676 32172 11732 32228
rect 4464 32116 4520 32172
rect 4568 32116 4624 32172
rect 4672 32116 4728 32172
rect 24464 32116 24520 32172
rect 24568 32116 24624 32172
rect 24672 32116 24728 32172
rect 9100 31724 9156 31780
rect 10220 31612 10276 31668
rect 2268 31500 2324 31556
rect 3804 31332 3860 31388
rect 3908 31332 3964 31388
rect 4012 31332 4068 31388
rect 23804 31332 23860 31388
rect 23908 31332 23964 31388
rect 24012 31332 24068 31388
rect 10220 31052 10276 31108
rect 1820 30716 1876 30772
rect 3164 30716 3220 30772
rect 13244 30716 13300 30772
rect 13468 30716 13524 30772
rect 4464 30548 4520 30604
rect 4568 30548 4624 30604
rect 4672 30548 4728 30604
rect 24464 30548 24520 30604
rect 24568 30548 24624 30604
rect 24672 30548 24728 30604
rect 22652 30492 22708 30548
rect 15260 30044 15316 30100
rect 13468 29820 13524 29876
rect 3804 29764 3860 29820
rect 3908 29764 3964 29820
rect 4012 29764 4068 29820
rect 23804 29764 23860 29820
rect 23908 29764 23964 29820
rect 24012 29764 24068 29820
rect 8316 29708 8372 29764
rect 18396 29708 18452 29764
rect 12348 29484 12404 29540
rect 15260 29372 15316 29428
rect 8316 29260 8372 29316
rect 4464 28980 4520 29036
rect 4568 28980 4624 29036
rect 4672 28980 4728 29036
rect 24464 28980 24520 29036
rect 24568 28980 24624 29036
rect 24672 28980 24728 29036
rect 8988 28924 9044 28980
rect 20076 28364 20132 28420
rect 22988 28252 23044 28308
rect 3804 28196 3860 28252
rect 3908 28196 3964 28252
rect 4012 28196 4068 28252
rect 23804 28196 23860 28252
rect 23908 28196 23964 28252
rect 24012 28196 24068 28252
rect 13244 27804 13300 27860
rect 15372 27804 15428 27860
rect 28364 27804 28420 27860
rect 4464 27412 4520 27468
rect 4568 27412 4624 27468
rect 4672 27412 4728 27468
rect 24464 27412 24520 27468
rect 24568 27412 24624 27468
rect 24672 27412 24728 27468
rect 7868 27132 7924 27188
rect 5292 27020 5348 27076
rect 9436 26908 9492 26964
rect 19068 26908 19124 26964
rect 12348 26684 12404 26740
rect 3804 26628 3860 26684
rect 3908 26628 3964 26684
rect 4012 26628 4068 26684
rect 23804 26628 23860 26684
rect 23908 26628 23964 26684
rect 24012 26628 24068 26684
rect 2156 26124 2212 26180
rect 9436 26012 9492 26068
rect 4464 25844 4520 25900
rect 4568 25844 4624 25900
rect 4672 25844 4728 25900
rect 24464 25844 24520 25900
rect 24568 25844 24624 25900
rect 24672 25844 24728 25900
rect 7196 25676 7252 25732
rect 11676 25564 11732 25620
rect 3804 25060 3860 25116
rect 3908 25060 3964 25116
rect 4012 25060 4068 25116
rect 23804 25060 23860 25116
rect 23908 25060 23964 25116
rect 24012 25060 24068 25116
rect 3500 24668 3556 24724
rect 7868 24556 7924 24612
rect 15372 24556 15428 24612
rect 3164 24444 3220 24500
rect 11340 24444 11396 24500
rect 17836 24444 17892 24500
rect 3500 24332 3556 24388
rect 9884 24332 9940 24388
rect 4464 24276 4520 24332
rect 4568 24276 4624 24332
rect 4672 24276 4728 24332
rect 24464 24276 24520 24332
rect 24568 24276 24624 24332
rect 24672 24276 24728 24332
rect 7196 24108 7252 24164
rect 26012 24108 26068 24164
rect 8988 23996 9044 24052
rect 5292 23884 5348 23940
rect 13580 23884 13636 23940
rect 17836 23884 17892 23940
rect 8988 23772 9044 23828
rect 24892 23772 24948 23828
rect 9100 23660 9156 23716
rect 20188 23548 20244 23604
rect 3804 23492 3860 23548
rect 3908 23492 3964 23548
rect 4012 23492 4068 23548
rect 23804 23492 23860 23548
rect 23908 23492 23964 23548
rect 24012 23492 24068 23548
rect 10108 23324 10164 23380
rect 19852 23324 19908 23380
rect 4464 22708 4520 22764
rect 4568 22708 4624 22764
rect 4672 22708 4728 22764
rect 11004 22652 11060 22708
rect 24464 22708 24520 22764
rect 24568 22708 24624 22764
rect 24672 22708 24728 22764
rect 20636 22204 20692 22260
rect 11900 22092 11956 22148
rect 3804 21924 3860 21980
rect 3908 21924 3964 21980
rect 4012 21924 4068 21980
rect 23804 21924 23860 21980
rect 23908 21924 23964 21980
rect 24012 21924 24068 21980
rect 14028 21644 14084 21700
rect 6748 21532 6804 21588
rect 15148 21420 15204 21476
rect 19852 21420 19908 21476
rect 15148 21196 15204 21252
rect 4464 21140 4520 21196
rect 4568 21140 4624 21196
rect 4672 21140 4728 21196
rect 4172 21084 4228 21140
rect 24464 21140 24520 21196
rect 24568 21140 24624 21196
rect 24672 21140 24728 21196
rect 27356 20860 27412 20916
rect 6748 20748 6804 20804
rect 21980 20748 22036 20804
rect 19068 20636 19124 20692
rect 3804 20356 3860 20412
rect 3908 20356 3964 20412
rect 4012 20356 4068 20412
rect 23804 20356 23860 20412
rect 23908 20356 23964 20412
rect 24012 20356 24068 20412
rect 19628 20300 19684 20356
rect 2716 20188 2772 20244
rect 14924 20188 14980 20244
rect 18060 20188 18116 20244
rect 20748 20076 20804 20132
rect 14924 19964 14980 20020
rect 2156 19740 2212 19796
rect 13468 19740 13524 19796
rect 4464 19572 4520 19628
rect 4568 19572 4624 19628
rect 4672 19572 4728 19628
rect 24464 19572 24520 19628
rect 24568 19572 24624 19628
rect 24672 19572 24728 19628
rect 2268 19292 2324 19348
rect 9884 19292 9940 19348
rect 27244 19292 27300 19348
rect 3612 19068 3668 19124
rect 5964 18956 6020 19012
rect 18620 18844 18676 18900
rect 3804 18788 3860 18844
rect 3908 18788 3964 18844
rect 4012 18788 4068 18844
rect 23804 18788 23860 18844
rect 23908 18788 23964 18844
rect 24012 18788 24068 18844
rect 5068 18732 5124 18788
rect 14028 18732 14084 18788
rect 20748 18620 20804 18676
rect 2380 18396 2436 18452
rect 17612 18396 17668 18452
rect 4844 18284 4900 18340
rect 14028 18284 14084 18340
rect 18620 18284 18676 18340
rect 19068 18172 19124 18228
rect 5964 18060 6020 18116
rect 18060 18060 18116 18116
rect 18620 18060 18676 18116
rect 20636 18060 20692 18116
rect 4464 18004 4520 18060
rect 4568 18004 4624 18060
rect 4672 18004 4728 18060
rect 24464 18004 24520 18060
rect 24568 18004 24624 18060
rect 24672 18004 24728 18060
rect 3388 17836 3444 17892
rect 19068 17724 19124 17780
rect 22988 17836 23044 17892
rect 14924 17500 14980 17556
rect 19404 17500 19460 17556
rect 20188 17388 20244 17444
rect 3804 17220 3860 17276
rect 3908 17220 3964 17276
rect 4012 17220 4068 17276
rect 23804 17220 23860 17276
rect 23908 17220 23964 17276
rect 24012 17220 24068 17276
rect 16940 17164 16996 17220
rect 19740 17164 19796 17220
rect 14924 17052 14980 17108
rect 3388 16828 3444 16884
rect 16940 16828 16996 16884
rect 5068 16716 5124 16772
rect 19964 16716 20020 16772
rect 19068 16492 19124 16548
rect 19404 16492 19460 16548
rect 19740 16492 19796 16548
rect 19964 16492 20020 16548
rect 4464 16436 4520 16492
rect 4568 16436 4624 16492
rect 4672 16436 4728 16492
rect 24464 16436 24520 16492
rect 24568 16436 24624 16492
rect 24672 16436 24728 16492
rect 18060 16380 18116 16436
rect 1820 16268 1876 16324
rect 2716 16268 2772 16324
rect 16156 16268 16212 16324
rect 3612 16156 3668 16212
rect 4172 16156 4228 16212
rect 8988 16156 9044 16212
rect 10444 16156 10500 16212
rect 19404 16156 19460 16212
rect 19628 16156 19684 16212
rect 21980 16044 22036 16100
rect 10108 15820 10164 15876
rect 14364 15820 14420 15876
rect 16156 15708 16212 15764
rect 3804 15652 3860 15708
rect 3908 15652 3964 15708
rect 4012 15652 4068 15708
rect 19404 15820 19460 15876
rect 23804 15652 23860 15708
rect 23908 15652 23964 15708
rect 24012 15652 24068 15708
rect 18620 15596 18676 15652
rect 19852 15372 19908 15428
rect 7868 15260 7924 15316
rect 11004 15260 11060 15316
rect 7756 15148 7812 15204
rect 7756 14924 7812 14980
rect 14364 14924 14420 14980
rect 24220 14924 24276 14980
rect 4464 14868 4520 14924
rect 4568 14868 4624 14924
rect 4672 14868 4728 14924
rect 24464 14868 24520 14924
rect 24568 14868 24624 14924
rect 24672 14868 24728 14924
rect 6748 14476 6804 14532
rect 8428 14364 8484 14420
rect 19852 14476 19908 14532
rect 7308 14140 7364 14196
rect 12572 14140 12628 14196
rect 24220 14140 24276 14196
rect 3804 14084 3860 14140
rect 3908 14084 3964 14140
rect 4012 14084 4068 14140
rect 23804 14084 23860 14140
rect 23908 14084 23964 14140
rect 24012 14084 24068 14140
rect 4172 14028 4228 14084
rect 14252 13916 14308 13972
rect 17612 13916 17668 13972
rect 14924 13804 14980 13860
rect 15260 13804 15316 13860
rect 3612 13692 3668 13748
rect 10108 13692 10164 13748
rect 26012 13692 26068 13748
rect 6748 13580 6804 13636
rect 8988 13580 9044 13636
rect 13468 13468 13524 13524
rect 9100 13356 9156 13412
rect 13580 13356 13636 13412
rect 4464 13300 4520 13356
rect 4568 13300 4624 13356
rect 4672 13300 4728 13356
rect 24464 13300 24520 13356
rect 24568 13300 24624 13356
rect 24672 13300 24728 13356
rect 11004 13244 11060 13300
rect 17612 13244 17668 13300
rect 20972 13132 21028 13188
rect 3164 13020 3220 13076
rect 7868 12684 7924 12740
rect 3804 12516 3860 12572
rect 3908 12516 3964 12572
rect 4012 12516 4068 12572
rect 10108 12460 10164 12516
rect 23804 12516 23860 12572
rect 23908 12516 23964 12572
rect 24012 12516 24068 12572
rect 13580 12460 13636 12516
rect 20972 12460 21028 12516
rect 11900 12236 11956 12292
rect 11116 11900 11172 11956
rect 8428 11788 8484 11844
rect 4464 11732 4520 11788
rect 4568 11732 4624 11788
rect 4672 11732 4728 11788
rect 20636 11788 20692 11844
rect 24464 11732 24520 11788
rect 24568 11732 24624 11788
rect 24672 11732 24728 11788
rect 18284 11452 18340 11508
rect 6188 11340 6244 11396
rect 9100 11004 9156 11060
rect 3804 10948 3860 11004
rect 3908 10948 3964 11004
rect 4012 10948 4068 11004
rect 8204 10668 8260 10724
rect 10108 10668 10164 10724
rect 23804 10948 23860 11004
rect 23908 10948 23964 11004
rect 24012 10948 24068 11004
rect 18284 10556 18340 10612
rect 22652 10556 22708 10612
rect 4464 10164 4520 10220
rect 4568 10164 4624 10220
rect 4672 10164 4728 10220
rect 24464 10164 24520 10220
rect 24568 10164 24624 10220
rect 24672 10164 24728 10220
rect 24892 10108 24948 10164
rect 11116 9996 11172 10052
rect 3804 9380 3860 9436
rect 3908 9380 3964 9436
rect 4012 9380 4068 9436
rect 23804 9380 23860 9436
rect 23908 9380 23964 9436
rect 24012 9380 24068 9436
rect 6412 9100 6468 9156
rect 4464 8596 4520 8652
rect 4568 8596 4624 8652
rect 4672 8596 4728 8652
rect 24464 8596 24520 8652
rect 24568 8596 24624 8652
rect 24672 8596 24728 8652
rect 10108 8316 10164 8372
rect 17836 8316 17892 8372
rect 15932 8092 15988 8148
rect 3804 7812 3860 7868
rect 3908 7812 3964 7868
rect 4012 7812 4068 7868
rect 23804 7812 23860 7868
rect 23908 7812 23964 7868
rect 24012 7812 24068 7868
rect 7308 7532 7364 7588
rect 22764 7308 22820 7364
rect 4464 7028 4520 7084
rect 4568 7028 4624 7084
rect 4672 7028 4728 7084
rect 24464 7028 24520 7084
rect 24568 7028 24624 7084
rect 24672 7028 24728 7084
rect 27132 6748 27188 6804
rect 19516 6636 19572 6692
rect 22428 6524 22484 6580
rect 20860 6300 20916 6356
rect 3804 6244 3860 6300
rect 3908 6244 3964 6300
rect 4012 6244 4068 6300
rect 23804 6244 23860 6300
rect 23908 6244 23964 6300
rect 24012 6244 24068 6300
rect 15148 5852 15204 5908
rect 4464 5460 4520 5516
rect 4568 5460 4624 5516
rect 4672 5460 4728 5516
rect 24464 5460 24520 5516
rect 24568 5460 24624 5516
rect 24672 5460 24728 5516
rect 15148 5292 15204 5348
rect 9212 5180 9268 5236
rect 3804 4676 3860 4732
rect 3908 4676 3964 4732
rect 4012 4676 4068 4732
rect 23804 4676 23860 4732
rect 23908 4676 23964 4732
rect 24012 4676 24068 4732
rect 27020 4508 27076 4564
rect 18844 4284 18900 4340
rect 4464 3892 4520 3948
rect 4568 3892 4624 3948
rect 4672 3892 4728 3948
rect 24464 3892 24520 3948
rect 24568 3892 24624 3948
rect 24672 3892 24728 3948
rect 17948 3836 18004 3892
rect 3804 3108 3860 3164
rect 3908 3108 3964 3164
rect 4012 3108 4068 3164
rect 23804 3108 23860 3164
rect 23908 3108 23964 3164
rect 24012 3108 24068 3164
rect 4464 2324 4520 2380
rect 4568 2324 4624 2380
rect 4672 2324 4728 2380
rect 24464 2324 24520 2380
rect 24568 2324 24624 2380
rect 24672 2324 24728 2380
rect 17724 2156 17780 2212
rect 21308 2156 21364 2212
rect 26908 1596 26964 1652
rect 3804 1540 3860 1596
rect 3908 1540 3964 1596
rect 4012 1540 4068 1596
rect 23804 1540 23860 1596
rect 23908 1540 23964 1596
rect 24012 1540 24068 1596
rect 28364 1148 28420 1204
rect 4464 756 4520 812
rect 4568 756 4624 812
rect 4672 756 4728 812
rect 24464 756 24520 812
rect 24568 756 24624 812
rect 24672 756 24728 812
rect 10892 588 10948 644
rect 16716 476 16772 532
<< metal4 >>
rect 3776 56476 4096 57456
rect 3776 56420 3804 56476
rect 3860 56420 3908 56476
rect 3964 56420 4012 56476
rect 4068 56420 4096 56476
rect 3164 55188 3220 55198
rect 2380 49028 2436 49038
rect 1820 37716 1876 37726
rect 1820 36260 1876 37660
rect 1820 36194 1876 36204
rect 2268 31556 2324 31566
rect 1820 30772 1876 30782
rect 1820 16324 1876 30716
rect 2156 26180 2212 26190
rect 2156 19796 2212 26124
rect 2156 19730 2212 19740
rect 2268 19348 2324 31500
rect 2268 19282 2324 19292
rect 2380 18452 2436 48972
rect 3164 30772 3220 55132
rect 3164 30706 3220 30716
rect 3776 54908 4096 56420
rect 3776 54852 3804 54908
rect 3860 54852 3908 54908
rect 3964 54852 4012 54908
rect 4068 54852 4096 54908
rect 3776 53340 4096 54852
rect 3776 53284 3804 53340
rect 3860 53284 3908 53340
rect 3964 53284 4012 53340
rect 4068 53284 4096 53340
rect 3776 51772 4096 53284
rect 3776 51716 3804 51772
rect 3860 51716 3908 51772
rect 3964 51716 4012 51772
rect 4068 51716 4096 51772
rect 3776 50204 4096 51716
rect 3776 50148 3804 50204
rect 3860 50148 3908 50204
rect 3964 50148 4012 50204
rect 4068 50148 4096 50204
rect 3776 48636 4096 50148
rect 3776 48580 3804 48636
rect 3860 48580 3908 48636
rect 3964 48580 4012 48636
rect 4068 48580 4096 48636
rect 3776 47068 4096 48580
rect 3776 47012 3804 47068
rect 3860 47012 3908 47068
rect 3964 47012 4012 47068
rect 4068 47012 4096 47068
rect 3776 45500 4096 47012
rect 3776 45444 3804 45500
rect 3860 45444 3908 45500
rect 3964 45444 4012 45500
rect 4068 45444 4096 45500
rect 3776 43932 4096 45444
rect 3776 43876 3804 43932
rect 3860 43876 3908 43932
rect 3964 43876 4012 43932
rect 4068 43876 4096 43932
rect 3776 42364 4096 43876
rect 3776 42308 3804 42364
rect 3860 42308 3908 42364
rect 3964 42308 4012 42364
rect 4068 42308 4096 42364
rect 3776 40796 4096 42308
rect 3776 40740 3804 40796
rect 3860 40740 3908 40796
rect 3964 40740 4012 40796
rect 4068 40740 4096 40796
rect 3776 39228 4096 40740
rect 3776 39172 3804 39228
rect 3860 39172 3908 39228
rect 3964 39172 4012 39228
rect 4068 39172 4096 39228
rect 3776 37660 4096 39172
rect 3776 37604 3804 37660
rect 3860 37604 3908 37660
rect 3964 37604 4012 37660
rect 4068 37604 4096 37660
rect 3776 36092 4096 37604
rect 3776 36036 3804 36092
rect 3860 36036 3908 36092
rect 3964 36036 4012 36092
rect 4068 36036 4096 36092
rect 3776 34524 4096 36036
rect 3776 34468 3804 34524
rect 3860 34468 3908 34524
rect 3964 34468 4012 34524
rect 4068 34468 4096 34524
rect 3776 32956 4096 34468
rect 4436 55692 4756 57456
rect 23776 56476 24096 57456
rect 23776 56420 23804 56476
rect 23860 56420 23908 56476
rect 23964 56420 24012 56476
rect 24068 56420 24096 56476
rect 4436 55636 4464 55692
rect 4520 55636 4568 55692
rect 4624 55636 4672 55692
rect 4728 55636 4756 55692
rect 4436 54124 4756 55636
rect 19516 55972 19572 55982
rect 19068 54292 19124 54302
rect 4436 54068 4464 54124
rect 4520 54068 4568 54124
rect 4624 54068 4672 54124
rect 4728 54068 4756 54124
rect 4436 52556 4756 54068
rect 17724 54180 17780 54190
rect 16716 53732 16772 53742
rect 4436 52500 4464 52556
rect 4520 52500 4568 52556
rect 4624 52500 4672 52556
rect 4728 52500 4756 52556
rect 4436 50988 4756 52500
rect 12572 52724 12628 52734
rect 4436 50932 4464 50988
rect 4520 50932 4568 50988
rect 4624 50932 4672 50988
rect 4728 50932 4756 50988
rect 4436 49420 4756 50932
rect 9212 51492 9268 51502
rect 4436 49364 4464 49420
rect 4520 49364 4568 49420
rect 4624 49364 4672 49420
rect 4728 49364 4756 49420
rect 4436 47852 4756 49364
rect 4436 47796 4464 47852
rect 4520 47796 4568 47852
rect 4624 47796 4672 47852
rect 4728 47796 4756 47852
rect 4436 46284 4756 47796
rect 4436 46228 4464 46284
rect 4520 46228 4568 46284
rect 4624 46228 4672 46284
rect 4728 46228 4756 46284
rect 4436 44716 4756 46228
rect 4436 44660 4464 44716
rect 4520 44660 4568 44716
rect 4624 44660 4672 44716
rect 4728 44660 4756 44716
rect 4436 43148 4756 44660
rect 4436 43092 4464 43148
rect 4520 43092 4568 43148
rect 4624 43092 4672 43148
rect 4728 43092 4756 43148
rect 4436 41580 4756 43092
rect 4436 41524 4464 41580
rect 4520 41524 4568 41580
rect 4624 41524 4672 41580
rect 4728 41524 4756 41580
rect 4436 40012 4756 41524
rect 4436 39956 4464 40012
rect 4520 39956 4568 40012
rect 4624 39956 4672 40012
rect 4728 39956 4756 40012
rect 4436 38444 4756 39956
rect 4436 38388 4464 38444
rect 4520 38388 4568 38444
rect 4624 38388 4672 38444
rect 4728 38388 4756 38444
rect 4436 36876 4756 38388
rect 4436 36820 4464 36876
rect 4520 36820 4568 36876
rect 4624 36820 4672 36876
rect 4728 36820 4756 36876
rect 4436 35308 4756 36820
rect 4436 35252 4464 35308
rect 4520 35252 4568 35308
rect 4624 35252 4672 35308
rect 4728 35252 4756 35308
rect 4284 34244 4340 34254
rect 4284 33684 4340 34188
rect 4284 33618 4340 33628
rect 4436 33740 4756 35252
rect 6188 49924 6244 49934
rect 4436 33684 4464 33740
rect 4520 33684 4568 33740
rect 4624 33684 4672 33740
rect 4728 33684 4756 33740
rect 3776 32900 3804 32956
rect 3860 32900 3908 32956
rect 3964 32900 4012 32956
rect 4068 32900 4096 32956
rect 3776 31388 4096 32900
rect 3776 31332 3804 31388
rect 3860 31332 3908 31388
rect 3964 31332 4012 31388
rect 4068 31332 4096 31388
rect 3776 29820 4096 31332
rect 3776 29764 3804 29820
rect 3860 29764 3908 29820
rect 3964 29764 4012 29820
rect 4068 29764 4096 29820
rect 3776 28252 4096 29764
rect 3776 28196 3804 28252
rect 3860 28196 3908 28252
rect 3964 28196 4012 28252
rect 4068 28196 4096 28252
rect 3776 26684 4096 28196
rect 3776 26628 3804 26684
rect 3860 26628 3908 26684
rect 3964 26628 4012 26684
rect 4068 26628 4096 26684
rect 3776 25116 4096 26628
rect 3776 25060 3804 25116
rect 3860 25060 3908 25116
rect 3964 25060 4012 25116
rect 4068 25060 4096 25116
rect 3500 24724 3556 24734
rect 3164 24500 3220 24510
rect 2380 18386 2436 18396
rect 2716 20244 2772 20254
rect 1820 16258 1876 16268
rect 2716 16324 2772 20188
rect 2716 16258 2772 16268
rect 3164 13076 3220 24444
rect 3500 24388 3556 24668
rect 3500 24322 3556 24332
rect 3776 23548 4096 25060
rect 3776 23492 3804 23548
rect 3860 23492 3908 23548
rect 3964 23492 4012 23548
rect 4068 23492 4096 23548
rect 3776 21980 4096 23492
rect 3776 21924 3804 21980
rect 3860 21924 3908 21980
rect 3964 21924 4012 21980
rect 4068 21924 4096 21980
rect 3776 20412 4096 21924
rect 4436 32172 4756 33684
rect 4436 32116 4464 32172
rect 4520 32116 4568 32172
rect 4624 32116 4672 32172
rect 4728 32116 4756 32172
rect 4436 30604 4756 32116
rect 4436 30548 4464 30604
rect 4520 30548 4568 30604
rect 4624 30548 4672 30604
rect 4728 30548 4756 30604
rect 4436 29036 4756 30548
rect 4436 28980 4464 29036
rect 4520 28980 4568 29036
rect 4624 28980 4672 29036
rect 4728 28980 4756 29036
rect 4436 27468 4756 28980
rect 4436 27412 4464 27468
rect 4520 27412 4568 27468
rect 4624 27412 4672 27468
rect 4728 27412 4756 27468
rect 4436 25900 4756 27412
rect 4436 25844 4464 25900
rect 4520 25844 4568 25900
rect 4624 25844 4672 25900
rect 4728 25844 4756 25900
rect 4436 24332 4756 25844
rect 4436 24276 4464 24332
rect 4520 24276 4568 24332
rect 4624 24276 4672 24332
rect 4728 24276 4756 24332
rect 4436 22764 4756 24276
rect 4436 22708 4464 22764
rect 4520 22708 4568 22764
rect 4624 22708 4672 22764
rect 4728 22708 4756 22764
rect 4436 21196 4756 22708
rect 3776 20356 3804 20412
rect 3860 20356 3908 20412
rect 3964 20356 4012 20412
rect 4068 20356 4096 20412
rect 3612 19124 3668 19134
rect 3388 17892 3444 17902
rect 3388 16884 3444 17836
rect 3388 16818 3444 16828
rect 3612 16212 3668 19068
rect 3612 13748 3668 16156
rect 3612 13682 3668 13692
rect 3776 18844 4096 20356
rect 3776 18788 3804 18844
rect 3860 18788 3908 18844
rect 3964 18788 4012 18844
rect 4068 18788 4096 18844
rect 3776 17276 4096 18788
rect 3776 17220 3804 17276
rect 3860 17220 3908 17276
rect 3964 17220 4012 17276
rect 4068 17220 4096 17276
rect 3776 15708 4096 17220
rect 3776 15652 3804 15708
rect 3860 15652 3908 15708
rect 3964 15652 4012 15708
rect 4068 15652 4096 15708
rect 3776 14140 4096 15652
rect 3776 14084 3804 14140
rect 3860 14084 3908 14140
rect 3964 14084 4012 14140
rect 4068 14084 4096 14140
rect 3164 13010 3220 13020
rect 3776 12572 4096 14084
rect 4172 21140 4228 21150
rect 4172 16212 4228 21084
rect 4172 14084 4228 16156
rect 4172 14018 4228 14028
rect 4436 21140 4464 21196
rect 4520 21140 4568 21196
rect 4624 21140 4672 21196
rect 4728 21140 4756 21196
rect 4436 19628 4756 21140
rect 4436 19572 4464 19628
rect 4520 19572 4568 19628
rect 4624 19572 4672 19628
rect 4728 19572 4756 19628
rect 4436 18060 4756 19572
rect 4844 34692 4900 34702
rect 4844 18340 4900 34636
rect 5292 27076 5348 27086
rect 5292 23940 5348 27020
rect 5292 23874 5348 23884
rect 5964 19012 6020 19022
rect 4844 18274 4900 18284
rect 5068 18788 5124 18798
rect 4436 18004 4464 18060
rect 4520 18004 4568 18060
rect 4624 18004 4672 18060
rect 4728 18004 4756 18060
rect 4436 16492 4756 18004
rect 5068 16772 5124 18732
rect 5964 18116 6020 18956
rect 5964 18050 6020 18060
rect 5068 16706 5124 16716
rect 4436 16436 4464 16492
rect 4520 16436 4568 16492
rect 4624 16436 4672 16492
rect 4728 16436 4756 16492
rect 4436 14924 4756 16436
rect 4436 14868 4464 14924
rect 4520 14868 4568 14924
rect 4624 14868 4672 14924
rect 4728 14868 4756 14924
rect 3776 12516 3804 12572
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 4068 12516 4096 12572
rect 3776 11004 4096 12516
rect 3776 10948 3804 11004
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 4068 10948 4096 11004
rect 3776 9436 4096 10948
rect 3776 9380 3804 9436
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 4068 9380 4096 9436
rect 3776 7868 4096 9380
rect 3776 7812 3804 7868
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 4068 7812 4096 7868
rect 3776 6300 4096 7812
rect 3776 6244 3804 6300
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 4068 6244 4096 6300
rect 3776 4732 4096 6244
rect 3776 4676 3804 4732
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 4068 4676 4096 4732
rect 3776 3164 4096 4676
rect 3776 3108 3804 3164
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 4068 3108 4096 3164
rect 3776 1596 4096 3108
rect 3776 1540 3804 1596
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 4068 1540 4096 1596
rect 3776 0 4096 1540
rect 4436 13356 4756 14868
rect 4436 13300 4464 13356
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4728 13300 4756 13356
rect 4436 11788 4756 13300
rect 4436 11732 4464 11788
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4728 11732 4756 11788
rect 4436 10220 4756 11732
rect 6188 11396 6244 49868
rect 6188 11330 6244 11340
rect 6412 41636 6468 41646
rect 4436 10164 4464 10220
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4728 10164 4756 10220
rect 4436 8652 4756 10164
rect 6412 9156 6468 41580
rect 8092 37156 8596 37198
rect 8148 37142 8540 37156
rect 8092 37090 8148 37100
rect 8540 37090 8596 37100
rect 9100 34468 9156 34478
rect 8204 34020 8260 34030
rect 8204 33236 8260 33964
rect 8204 33170 8260 33180
rect 8988 33796 9044 33806
rect 8316 29764 8372 29774
rect 8316 29316 8372 29708
rect 7868 27188 7924 27198
rect 7196 25732 7252 25742
rect 7196 24164 7252 25676
rect 7868 24612 7924 27132
rect 7868 24546 7924 24556
rect 7196 24098 7252 24108
rect 6748 21588 6804 21598
rect 6748 20804 6804 21532
rect 8316 20998 8372 29260
rect 8988 28980 9044 33740
rect 8988 28914 9044 28924
rect 9100 31780 9156 34412
rect 8988 24052 9044 24062
rect 8988 23828 9044 23996
rect 8988 23762 9044 23772
rect 9100 23716 9156 31724
rect 9100 23650 9156 23660
rect 6748 14532 6804 20748
rect 8204 20942 8372 20998
rect 7868 15316 7924 15326
rect 7756 15204 7812 15214
rect 7756 14980 7812 15148
rect 7756 14914 7812 14924
rect 6748 13636 6804 14476
rect 6748 13570 6804 13580
rect 7308 14196 7364 14206
rect 6412 9090 6468 9100
rect 4436 8596 4464 8652
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4728 8596 4756 8652
rect 4436 7084 4756 8596
rect 7308 7588 7364 14140
rect 7868 12740 7924 15260
rect 7868 12674 7924 12684
rect 8204 10724 8260 20942
rect 8988 16212 9044 16222
rect 8428 14420 8484 14430
rect 8428 11844 8484 14364
rect 8988 13636 9044 16156
rect 9044 13580 9156 13618
rect 8988 13562 9156 13580
rect 8428 11778 8484 11788
rect 9100 13412 9156 13562
rect 9100 11060 9156 13356
rect 9100 10994 9156 11004
rect 8204 10658 8260 10668
rect 7308 7522 7364 7532
rect 4436 7028 4464 7084
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4728 7028 4756 7084
rect 4436 5516 4756 7028
rect 4436 5460 4464 5516
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4728 5460 4756 5516
rect 4436 3948 4756 5460
rect 9212 5236 9268 51436
rect 11340 51268 11396 51278
rect 10444 39284 10500 39294
rect 10220 31668 10276 31678
rect 10220 31108 10276 31612
rect 10220 31042 10276 31052
rect 9436 26964 9492 26974
rect 9436 26068 9492 26908
rect 9436 26002 9492 26012
rect 9884 24388 9940 24398
rect 9884 19348 9940 24332
rect 9884 19282 9940 19292
rect 10108 23380 10164 23390
rect 10108 15876 10164 23324
rect 10444 16212 10500 39228
rect 10444 16146 10500 16156
rect 10892 34916 10948 34926
rect 10108 15810 10164 15820
rect 10108 13748 10164 13758
rect 10108 12516 10164 13692
rect 10108 12450 10164 12460
rect 10108 10724 10164 10734
rect 10108 8372 10164 10668
rect 10108 8306 10164 8316
rect 9212 5170 9268 5180
rect 4436 3892 4464 3948
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4728 3892 4756 3948
rect 4436 2380 4756 3892
rect 4436 2324 4464 2380
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4728 2324 4756 2380
rect 4436 812 4756 2324
rect 4436 756 4464 812
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4728 756 4756 812
rect 4436 0 4756 756
rect 10892 644 10948 34860
rect 11340 24500 11396 51212
rect 12348 32900 12404 32910
rect 11676 32228 11732 32238
rect 11676 25620 11732 32172
rect 12348 29540 12404 32844
rect 12348 26740 12404 29484
rect 12348 26674 12404 26684
rect 11676 25554 11732 25564
rect 11340 24434 11396 24444
rect 11004 22708 11060 22718
rect 11004 15316 11060 22652
rect 11004 13300 11060 15260
rect 11004 13234 11060 13244
rect 11900 22148 11956 22158
rect 11900 12292 11956 22092
rect 12572 14196 12628 52668
rect 14252 49700 14308 49710
rect 13580 34132 13636 34142
rect 13244 30772 13300 30782
rect 13244 27860 13300 30716
rect 13468 30772 13524 30782
rect 13468 29876 13524 30716
rect 13468 29810 13524 29820
rect 13244 27794 13300 27804
rect 13580 23940 13636 34076
rect 13580 23874 13636 23884
rect 14028 21700 14084 21710
rect 12572 14130 12628 14140
rect 13468 19796 13524 19806
rect 13468 13524 13524 19740
rect 14028 18788 14084 21644
rect 14028 18340 14084 18732
rect 14028 18274 14084 18284
rect 14252 13972 14308 49644
rect 15932 48132 15988 48142
rect 15260 30100 15316 30110
rect 15260 29428 15316 30044
rect 15260 29362 15316 29372
rect 15372 27860 15428 27870
rect 15372 24612 15428 27804
rect 15372 24546 15428 24556
rect 15148 21476 15204 21486
rect 15148 21252 15204 21420
rect 15148 21186 15204 21196
rect 14924 20244 14980 20254
rect 14924 20020 14980 20188
rect 14924 19954 14980 19964
rect 14924 17556 14980 17566
rect 14924 17108 14980 17500
rect 14924 17042 14980 17052
rect 14364 15876 14420 15886
rect 14364 14980 14420 15820
rect 14364 14914 14420 14924
rect 14252 13906 14308 13916
rect 14924 13860 14980 13870
rect 14924 13798 14980 13804
rect 15260 13860 15316 13870
rect 15260 13798 15316 13804
rect 14924 13742 15316 13798
rect 13468 13458 13524 13468
rect 13580 13412 13636 13422
rect 13580 12516 13636 13356
rect 13580 12450 13636 12460
rect 11900 12226 11956 12236
rect 11116 11956 11172 11966
rect 11116 10052 11172 11900
rect 11116 9986 11172 9996
rect 15932 8148 15988 48076
rect 16156 16324 16212 16334
rect 16156 15764 16212 16268
rect 16156 15698 16212 15708
rect 15932 8082 15988 8092
rect 15148 5908 15204 5918
rect 15148 5348 15204 5852
rect 15148 5282 15204 5292
rect 10892 578 10948 588
rect 16716 532 16772 53676
rect 17612 18452 17668 18462
rect 16940 17220 16996 17230
rect 16940 16884 16996 17164
rect 16940 16818 16996 16828
rect 17612 13972 17668 18396
rect 17612 13300 17668 13916
rect 17612 13234 17668 13244
rect 17724 2212 17780 54124
rect 17948 53844 18004 53854
rect 17836 24500 17892 24510
rect 17836 23940 17892 24444
rect 17836 8372 17892 23884
rect 17836 8306 17892 8316
rect 17948 3892 18004 53788
rect 18396 34692 18452 34702
rect 18396 29764 18452 34636
rect 18396 29698 18452 29708
rect 19068 26964 19124 54236
rect 19068 26898 19124 26908
rect 19068 20692 19124 20702
rect 18060 20244 18116 20254
rect 18060 18116 18116 20188
rect 18620 18900 18676 18910
rect 18620 18340 18676 18844
rect 18676 18284 18900 18298
rect 18620 18242 18900 18284
rect 18060 16436 18116 18060
rect 18060 16370 18116 16380
rect 18620 18116 18676 18126
rect 18620 15652 18676 18060
rect 18620 15586 18676 15596
rect 18284 11508 18340 11518
rect 18284 10612 18340 11452
rect 18284 10546 18340 10556
rect 18844 4340 18900 18242
rect 19068 18228 19124 20636
rect 19068 18162 19124 18172
rect 19068 17780 19124 17790
rect 19068 16548 19124 17724
rect 19068 16482 19124 16492
rect 19404 17556 19460 17566
rect 19404 16548 19460 17500
rect 19404 16482 19460 16492
rect 19404 16212 19460 16222
rect 19404 15876 19460 16156
rect 19404 15810 19460 15820
rect 19516 6692 19572 55916
rect 21308 55972 21364 55982
rect 20860 55300 20916 55310
rect 20076 53956 20132 53966
rect 20076 28420 20132 53900
rect 20076 28354 20132 28364
rect 20188 23604 20244 23614
rect 19852 23380 19908 23390
rect 19852 21476 19908 23324
rect 19852 21410 19908 21420
rect 19628 20356 19684 20366
rect 19628 16212 19684 20300
rect 20188 17444 20244 23548
rect 20188 17378 20244 17388
rect 20636 22260 20692 22270
rect 20636 18116 20692 22204
rect 20748 20132 20804 20142
rect 20748 18676 20804 20076
rect 20748 18610 20804 18620
rect 19740 17220 19796 17230
rect 19740 16548 19796 17164
rect 19740 16482 19796 16492
rect 19964 16772 20020 16782
rect 19964 16548 20020 16716
rect 19964 16482 20020 16492
rect 19628 16146 19684 16156
rect 19852 15428 19908 15438
rect 19852 14532 19908 15372
rect 19852 14466 19908 14476
rect 20636 11844 20692 18060
rect 20636 11778 20692 11788
rect 19516 6626 19572 6636
rect 20860 6356 20916 55244
rect 20972 13188 21028 13198
rect 20972 12516 21028 13132
rect 20972 12450 21028 12460
rect 20860 6290 20916 6300
rect 18844 4274 18900 4284
rect 17948 3826 18004 3836
rect 17724 2146 17780 2156
rect 21308 2212 21364 55916
rect 22428 55300 22484 55310
rect 21980 20804 22036 20814
rect 21980 16100 22036 20748
rect 21980 16034 22036 16044
rect 22428 6580 22484 55244
rect 23776 54908 24096 56420
rect 23776 54852 23804 54908
rect 23860 54852 23908 54908
rect 23964 54852 24012 54908
rect 24068 54852 24096 54908
rect 23776 53340 24096 54852
rect 23776 53284 23804 53340
rect 23860 53284 23908 53340
rect 23964 53284 24012 53340
rect 24068 53284 24096 53340
rect 22764 52164 22820 52174
rect 22652 30548 22708 30558
rect 22652 10612 22708 30492
rect 22652 10546 22708 10556
rect 22764 7364 22820 52108
rect 23776 51772 24096 53284
rect 23776 51716 23804 51772
rect 23860 51716 23908 51772
rect 23964 51716 24012 51772
rect 24068 51716 24096 51772
rect 23776 50204 24096 51716
rect 23776 50148 23804 50204
rect 23860 50148 23908 50204
rect 23964 50148 24012 50204
rect 24068 50148 24096 50204
rect 23776 48636 24096 50148
rect 23776 48580 23804 48636
rect 23860 48580 23908 48636
rect 23964 48580 24012 48636
rect 24068 48580 24096 48636
rect 23776 47068 24096 48580
rect 23776 47012 23804 47068
rect 23860 47012 23908 47068
rect 23964 47012 24012 47068
rect 24068 47012 24096 47068
rect 23776 45500 24096 47012
rect 23776 45444 23804 45500
rect 23860 45444 23908 45500
rect 23964 45444 24012 45500
rect 24068 45444 24096 45500
rect 23776 43932 24096 45444
rect 23776 43876 23804 43932
rect 23860 43876 23908 43932
rect 23964 43876 24012 43932
rect 24068 43876 24096 43932
rect 23776 42364 24096 43876
rect 23776 42308 23804 42364
rect 23860 42308 23908 42364
rect 23964 42308 24012 42364
rect 24068 42308 24096 42364
rect 23776 40796 24096 42308
rect 23776 40740 23804 40796
rect 23860 40740 23908 40796
rect 23964 40740 24012 40796
rect 24068 40740 24096 40796
rect 23776 39228 24096 40740
rect 23776 39172 23804 39228
rect 23860 39172 23908 39228
rect 23964 39172 24012 39228
rect 24068 39172 24096 39228
rect 23776 37660 24096 39172
rect 23776 37604 23804 37660
rect 23860 37604 23908 37660
rect 23964 37604 24012 37660
rect 24068 37604 24096 37660
rect 23776 36092 24096 37604
rect 23776 36036 23804 36092
rect 23860 36036 23908 36092
rect 23964 36036 24012 36092
rect 24068 36036 24096 36092
rect 23776 34524 24096 36036
rect 23776 34468 23804 34524
rect 23860 34468 23908 34524
rect 23964 34468 24012 34524
rect 24068 34468 24096 34524
rect 23776 32956 24096 34468
rect 23776 32900 23804 32956
rect 23860 32900 23908 32956
rect 23964 32900 24012 32956
rect 24068 32900 24096 32956
rect 23776 31388 24096 32900
rect 23776 31332 23804 31388
rect 23860 31332 23908 31388
rect 23964 31332 24012 31388
rect 24068 31332 24096 31388
rect 23776 29820 24096 31332
rect 23776 29764 23804 29820
rect 23860 29764 23908 29820
rect 23964 29764 24012 29820
rect 24068 29764 24096 29820
rect 22988 28308 23044 28318
rect 22988 17892 23044 28252
rect 22988 17826 23044 17836
rect 23776 28252 24096 29764
rect 23776 28196 23804 28252
rect 23860 28196 23908 28252
rect 23964 28196 24012 28252
rect 24068 28196 24096 28252
rect 23776 26684 24096 28196
rect 23776 26628 23804 26684
rect 23860 26628 23908 26684
rect 23964 26628 24012 26684
rect 24068 26628 24096 26684
rect 23776 25116 24096 26628
rect 23776 25060 23804 25116
rect 23860 25060 23908 25116
rect 23964 25060 24012 25116
rect 24068 25060 24096 25116
rect 23776 23548 24096 25060
rect 23776 23492 23804 23548
rect 23860 23492 23908 23548
rect 23964 23492 24012 23548
rect 24068 23492 24096 23548
rect 23776 21980 24096 23492
rect 23776 21924 23804 21980
rect 23860 21924 23908 21980
rect 23964 21924 24012 21980
rect 24068 21924 24096 21980
rect 23776 20412 24096 21924
rect 23776 20356 23804 20412
rect 23860 20356 23908 20412
rect 23964 20356 24012 20412
rect 24068 20356 24096 20412
rect 23776 18844 24096 20356
rect 23776 18788 23804 18844
rect 23860 18788 23908 18844
rect 23964 18788 24012 18844
rect 24068 18788 24096 18844
rect 22764 7298 22820 7308
rect 23776 17276 24096 18788
rect 23776 17220 23804 17276
rect 23860 17220 23908 17276
rect 23964 17220 24012 17276
rect 24068 17220 24096 17276
rect 23776 15708 24096 17220
rect 23776 15652 23804 15708
rect 23860 15652 23908 15708
rect 23964 15652 24012 15708
rect 24068 15652 24096 15708
rect 23776 14140 24096 15652
rect 24436 55692 24756 57456
rect 24436 55636 24464 55692
rect 24520 55636 24568 55692
rect 24624 55636 24672 55692
rect 24728 55636 24756 55692
rect 24436 54124 24756 55636
rect 24436 54068 24464 54124
rect 24520 54068 24568 54124
rect 24624 54068 24672 54124
rect 24728 54068 24756 54124
rect 24436 52556 24756 54068
rect 24436 52500 24464 52556
rect 24520 52500 24568 52556
rect 24624 52500 24672 52556
rect 24728 52500 24756 52556
rect 24436 50988 24756 52500
rect 24436 50932 24464 50988
rect 24520 50932 24568 50988
rect 24624 50932 24672 50988
rect 24728 50932 24756 50988
rect 24436 49420 24756 50932
rect 27020 55188 27076 55198
rect 24436 49364 24464 49420
rect 24520 49364 24568 49420
rect 24624 49364 24672 49420
rect 24728 49364 24756 49420
rect 24436 47852 24756 49364
rect 24436 47796 24464 47852
rect 24520 47796 24568 47852
rect 24624 47796 24672 47852
rect 24728 47796 24756 47852
rect 24436 46284 24756 47796
rect 24436 46228 24464 46284
rect 24520 46228 24568 46284
rect 24624 46228 24672 46284
rect 24728 46228 24756 46284
rect 24436 44716 24756 46228
rect 24436 44660 24464 44716
rect 24520 44660 24568 44716
rect 24624 44660 24672 44716
rect 24728 44660 24756 44716
rect 24436 43148 24756 44660
rect 24436 43092 24464 43148
rect 24520 43092 24568 43148
rect 24624 43092 24672 43148
rect 24728 43092 24756 43148
rect 24436 41580 24756 43092
rect 24436 41524 24464 41580
rect 24520 41524 24568 41580
rect 24624 41524 24672 41580
rect 24728 41524 24756 41580
rect 24436 40012 24756 41524
rect 24436 39956 24464 40012
rect 24520 39956 24568 40012
rect 24624 39956 24672 40012
rect 24728 39956 24756 40012
rect 24436 38444 24756 39956
rect 24436 38388 24464 38444
rect 24520 38388 24568 38444
rect 24624 38388 24672 38444
rect 24728 38388 24756 38444
rect 24436 36876 24756 38388
rect 24436 36820 24464 36876
rect 24520 36820 24568 36876
rect 24624 36820 24672 36876
rect 24728 36820 24756 36876
rect 24436 35308 24756 36820
rect 24436 35252 24464 35308
rect 24520 35252 24568 35308
rect 24624 35252 24672 35308
rect 24728 35252 24756 35308
rect 24436 33740 24756 35252
rect 24436 33684 24464 33740
rect 24520 33684 24568 33740
rect 24624 33684 24672 33740
rect 24728 33684 24756 33740
rect 24436 32172 24756 33684
rect 24436 32116 24464 32172
rect 24520 32116 24568 32172
rect 24624 32116 24672 32172
rect 24728 32116 24756 32172
rect 24436 30604 24756 32116
rect 24436 30548 24464 30604
rect 24520 30548 24568 30604
rect 24624 30548 24672 30604
rect 24728 30548 24756 30604
rect 24436 29036 24756 30548
rect 24436 28980 24464 29036
rect 24520 28980 24568 29036
rect 24624 28980 24672 29036
rect 24728 28980 24756 29036
rect 24436 27468 24756 28980
rect 24436 27412 24464 27468
rect 24520 27412 24568 27468
rect 24624 27412 24672 27468
rect 24728 27412 24756 27468
rect 24436 25900 24756 27412
rect 24436 25844 24464 25900
rect 24520 25844 24568 25900
rect 24624 25844 24672 25900
rect 24728 25844 24756 25900
rect 24436 24332 24756 25844
rect 24436 24276 24464 24332
rect 24520 24276 24568 24332
rect 24624 24276 24672 24332
rect 24728 24276 24756 24332
rect 24436 22764 24756 24276
rect 26908 50596 26964 50606
rect 26012 24164 26068 24174
rect 24436 22708 24464 22764
rect 24520 22708 24568 22764
rect 24624 22708 24672 22764
rect 24728 22708 24756 22764
rect 24436 21196 24756 22708
rect 24436 21140 24464 21196
rect 24520 21140 24568 21196
rect 24624 21140 24672 21196
rect 24728 21140 24756 21196
rect 24436 19628 24756 21140
rect 24436 19572 24464 19628
rect 24520 19572 24568 19628
rect 24624 19572 24672 19628
rect 24728 19572 24756 19628
rect 24436 18060 24756 19572
rect 24436 18004 24464 18060
rect 24520 18004 24568 18060
rect 24624 18004 24672 18060
rect 24728 18004 24756 18060
rect 24436 16492 24756 18004
rect 24436 16436 24464 16492
rect 24520 16436 24568 16492
rect 24624 16436 24672 16492
rect 24728 16436 24756 16492
rect 23776 14084 23804 14140
rect 23860 14084 23908 14140
rect 23964 14084 24012 14140
rect 24068 14084 24096 14140
rect 24220 14980 24276 14990
rect 24220 14196 24276 14924
rect 24220 14130 24276 14140
rect 24436 14924 24756 16436
rect 24436 14868 24464 14924
rect 24520 14868 24568 14924
rect 24624 14868 24672 14924
rect 24728 14868 24756 14924
rect 23776 12572 24096 14084
rect 23776 12516 23804 12572
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 24068 12516 24096 12572
rect 23776 11004 24096 12516
rect 23776 10948 23804 11004
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 24068 10948 24096 11004
rect 23776 9436 24096 10948
rect 23776 9380 23804 9436
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 24068 9380 24096 9436
rect 23776 7868 24096 9380
rect 23776 7812 23804 7868
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 24068 7812 24096 7868
rect 22428 6514 22484 6524
rect 21308 2146 21364 2156
rect 23776 6300 24096 7812
rect 23776 6244 23804 6300
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 24068 6244 24096 6300
rect 23776 4732 24096 6244
rect 23776 4676 23804 4732
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 24068 4676 24096 4732
rect 23776 3164 24096 4676
rect 23776 3108 23804 3164
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 24068 3108 24096 3164
rect 16716 466 16772 476
rect 23776 1596 24096 3108
rect 23776 1540 23804 1596
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 24068 1540 24096 1596
rect 23776 0 24096 1540
rect 24436 13356 24756 14868
rect 24436 13300 24464 13356
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24728 13300 24756 13356
rect 24436 11788 24756 13300
rect 24436 11732 24464 11788
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24728 11732 24756 11788
rect 24436 10220 24756 11732
rect 24436 10164 24464 10220
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24728 10164 24756 10220
rect 24436 8652 24756 10164
rect 24892 23828 24948 23838
rect 24892 10164 24948 23772
rect 26012 13748 26068 24108
rect 26012 13682 26068 13692
rect 24892 10098 24948 10108
rect 24436 8596 24464 8652
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24728 8596 24756 8652
rect 24436 7084 24756 8596
rect 24436 7028 24464 7084
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 24728 7028 24756 7084
rect 24436 5516 24756 7028
rect 24436 5460 24464 5516
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24728 5460 24756 5516
rect 24436 3948 24756 5460
rect 24436 3892 24464 3948
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24728 3892 24756 3948
rect 24436 2380 24756 3892
rect 24436 2324 24464 2380
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24728 2324 24756 2380
rect 24436 812 24756 2324
rect 26908 1652 26964 50540
rect 27020 4564 27076 55132
rect 27132 52388 27188 52398
rect 27132 6804 27188 52332
rect 27244 41300 27300 41310
rect 27244 19348 27300 41244
rect 27356 37828 27412 37838
rect 27356 20916 27412 37772
rect 27356 20850 27412 20860
rect 28364 27860 28420 27870
rect 27244 19282 27300 19292
rect 27132 6738 27188 6748
rect 27020 4498 27076 4508
rect 26908 1586 26964 1596
rect 28364 1204 28420 27804
rect 28364 1138 28420 1148
rect 24436 756 24464 812
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24728 756 24756 812
rect 24436 0 24756 756
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _078_
timestamp 1486834041
transform 1 0 15904 0 -1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _079_
timestamp 1486834041
transform -1 0 10080 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _080_
timestamp 1486834041
transform -1 0 17584 0 1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _081_
timestamp 1486834041
transform -1 0 16352 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _082_
timestamp 1486834041
transform 1 0 14784 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _083_
timestamp 1486834041
transform 1 0 3360 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _084_
timestamp 1486834041
transform 1 0 11984 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _085_
timestamp 1486834041
transform 1 0 8064 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _086_
timestamp 1486834041
transform -1 0 21840 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _087_
timestamp 1486834041
transform 1 0 16576 0 -1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _088_
timestamp 1486834041
transform 1 0 15904 0 -1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _089_
timestamp 1486834041
transform -1 0 20272 0 1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _090_
timestamp 1486834041
transform 1 0 6832 0 1 19600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _091_
timestamp 1486834041
transform 1 0 4928 0 -1 18032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _092_
timestamp 1486834041
transform 1 0 4928 0 -1 19600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _093_
timestamp 1486834041
transform 1 0 13440 0 1 27440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _094_
timestamp 1486834041
transform 1 0 11088 0 -1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _095_
timestamp 1486834041
transform 1 0 18144 0 -1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _096_
timestamp 1486834041
transform 1 0 11312 0 -1 32144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _097_
timestamp 1486834041
transform 1 0 15232 0 -1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _098_
timestamp 1486834041
transform 1 0 14784 0 -1 10192
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _099_
timestamp 1486834041
transform 1 0 15232 0 -1 8624
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _100_
timestamp 1486834041
transform 1 0 16016 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _101_
timestamp 1486834041
transform -1 0 17472 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _102_
timestamp 1486834041
transform 1 0 15456 0 1 7056
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _103_
timestamp 1486834041
transform 1 0 16576 0 1 10192
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _104_
timestamp 1486834041
transform 1 0 16576 0 -1 8624
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _105_
timestamp 1486834041
transform 1 0 8736 0 -1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _106_
timestamp 1486834041
transform 1 0 6944 0 -1 11760
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _107_
timestamp 1486834041
transform 1 0 3808 0 -1 14896
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _108_
timestamp 1486834041
transform 1 0 7616 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _109_
timestamp 1486834041
transform -1 0 7952 0 1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _110_
timestamp 1486834041
transform 1 0 5712 0 -1 16464
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _111_
timestamp 1486834041
transform -1 0 9520 0 -1 14896
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _112_
timestamp 1486834041
transform 1 0 7168 0 -1 14896
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _113_
timestamp 1486834041
transform -1 0 13328 0 1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _114_
timestamp 1486834041
transform 1 0 11312 0 1 10192
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _115_
timestamp 1486834041
transform -1 0 13664 0 -1 10192
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _116_
timestamp 1486834041
transform 1 0 13664 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _117_
timestamp 1486834041
transform 1 0 11312 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _118_
timestamp 1486834041
transform -1 0 11312 0 -1 11760
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _119_
timestamp 1486834041
transform 1 0 10528 0 1 10192
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _120_
timestamp 1486834041
transform 1 0 12656 0 1 10192
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _121_
timestamp 1486834041
transform -1 0 9408 0 -1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _122_
timestamp 1486834041
transform 1 0 6944 0 -1 10192
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _123_
timestamp 1486834041
transform -1 0 9072 0 1 11760
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _124_
timestamp 1486834041
transform 1 0 8736 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _125_
timestamp 1486834041
transform -1 0 7728 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _126_
timestamp 1486834041
transform 1 0 7952 0 -1 8624
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _127_
timestamp 1486834041
transform -1 0 10304 0 1 10192
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _128_
timestamp 1486834041
transform 1 0 7056 0 1 10192
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _129_
timestamp 1486834041
transform 1 0 19376 0 -1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _130_
timestamp 1486834041
transform 1 0 20496 0 1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _131_
timestamp 1486834041
transform 1 0 19040 0 -1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _132_
timestamp 1486834041
transform 1 0 20496 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _133_
timestamp 1486834041
transform 1 0 20496 0 1 14896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _134_
timestamp 1486834041
transform -1 0 20272 0 1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _135_
timestamp 1486834041
transform 1 0 17136 0 1 13328
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _136_
timestamp 1486834041
transform -1 0 21168 0 1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _137_
timestamp 1486834041
transform 1 0 17696 0 -1 16464
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _138_
timestamp 1486834041
transform 1 0 16576 0 -1 16464
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _139_
timestamp 1486834041
transform 1 0 18928 0 1 13328
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _140_
timestamp 1486834041
transform 1 0 20496 0 1 18032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _141_
timestamp 1486834041
transform -1 0 20160 0 1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _142_
timestamp 1486834041
transform 1 0 18816 0 -1 16464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _143_
timestamp 1486834041
transform -1 0 19936 0 1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _144_
timestamp 1486834041
transform -1 0 19040 0 1 18032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _145_
timestamp 1486834041
transform 1 0 18480 0 1 19600
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _146_
timestamp 1486834041
transform 1 0 17696 0 -1 18032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _147_
timestamp 1486834041
transform -1 0 17696 0 -1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _148_
timestamp 1486834041
transform 1 0 18144 0 1 16464
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _149_
timestamp 1486834041
transform 1 0 17808 0 -1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _150_
timestamp 1486834041
transform -1 0 18032 0 1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _151_
timestamp 1486834041
transform 1 0 17584 0 -1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _152_
timestamp 1486834041
transform 1 0 19264 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _153_
timestamp 1486834041
transform 1 0 17584 0 -1 14896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _154_
timestamp 1486834041
transform -1 0 18928 0 -1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _155_
timestamp 1486834041
transform 1 0 16576 0 -1 13328
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _156_
timestamp 1486834041
transform 1 0 16576 0 -1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _157_
timestamp 1486834041
transform -1 0 19376 0 1 14896
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _158_
timestamp 1486834041
transform 1 0 16800 0 1 11760
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _159_
timestamp 1486834041
transform 1 0 17920 0 1 11760
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _160_
timestamp 1486834041
transform 1 0 19152 0 -1 22736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _161_
timestamp 1486834041
transform 1 0 20496 0 1 19600
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _162_
timestamp 1486834041
transform 1 0 18592 0 -1 21168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _163_
timestamp 1486834041
transform -1 0 20272 0 1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _164_
timestamp 1486834041
transform -1 0 21504 0 -1 19600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _165_
timestamp 1486834041
transform -1 0 20272 0 1 19600
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _166_
timestamp 1486834041
transform -1 0 18256 0 -1 21168
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _167_
timestamp 1486834041
transform -1 0 18704 0 1 21168
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _168_
timestamp 1486834041
transform 1 0 16800 0 -1 19600
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _169_
timestamp 1486834041
transform 1 0 18704 0 1 21168
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _170_
timestamp 1486834041
transform 1 0 20496 0 1 21168
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _171_
timestamp 1486834041
transform 1 0 15008 0 1 36848
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _172_
timestamp 1486834041
transform 1 0 8624 0 1 33712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _173_
timestamp 1486834041
transform 1 0 12432 0 -1 30576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _174_
timestamp 1486834041
transform 1 0 2016 0 -1 21168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _175_
timestamp 1486834041
transform 1 0 14448 0 1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _176_
timestamp 1486834041
transform 1 0 8848 0 1 16464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _177_
timestamp 1486834041
transform 1 0 19264 0 -1 29008
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _178_
timestamp 1486834041
transform -1 0 12432 0 1 30576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _179_
timestamp 1486834041
transform 1 0 20496 0 1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _180_
timestamp 1486834041
transform 1 0 2240 0 -1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _181_
timestamp 1486834041
transform 1 0 15344 0 1 30576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _182_
timestamp 1486834041
transform 1 0 3360 0 -1 30576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _183_
timestamp 1486834041
transform 1 0 12320 0 -1 19600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _184_
timestamp 1486834041
transform 1 0 14560 0 1 16464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _185_
timestamp 1486834041
transform 1 0 20496 0 1 30576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _186_
timestamp 1486834041
transform 1 0 7840 0 1 38416
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _187_
timestamp 1486834041
transform 1 0 2688 0 -1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _188_
timestamp 1486834041
transform 1 0 6832 0 1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _189_
timestamp 1486834041
transform 1 0 4928 0 -1 32144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _190_
timestamp 1486834041
transform 1 0 2128 0 -1 33712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _191_
timestamp 1486834041
transform 1 0 12656 0 1 19600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _192_
timestamp 1486834041
transform 1 0 14560 0 1 14896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _193_
timestamp 1486834041
transform 1 0 10192 0 -1 21168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _194_
timestamp 1486834041
transform 1 0 8848 0 1 25872
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _195_
timestamp 1486834041
transform 1 0 20048 0 -1 32144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _196_
timestamp 1486834041
transform 1 0 5936 0 1 39984
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _197_
timestamp 1486834041
transform 1 0 1008 0 1 33712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _198_
timestamp 1486834041
transform 1 0 2464 0 -1 25872
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _199_
timestamp 1486834041
transform 1 0 13664 0 1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _200_
timestamp 1486834041
transform 1 0 8960 0 -1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _201_
timestamp 1486834041
transform 1 0 17248 0 -1 27440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _202_
timestamp 1486834041
transform 1 0 12656 0 1 38416
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _203_
timestamp 1486834041
transform 1 0 14224 0 1 29008
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _204_
timestamp 1486834041
transform -1 0 8736 0 1 21168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _205_
timestamp 1486834041
transform -1 0 4928 0 -1 18032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _206_
timestamp 1486834041
transform 1 0 3136 0 -1 27440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _207_
timestamp 1486834041
transform 1 0 13552 0 1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _208_
timestamp 1486834041
transform 1 0 8848 0 1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _209_
timestamp 1486834041
transform 1 0 16576 0 -1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _210_
timestamp 1486834041
transform 1 0 11424 0 -1 29008
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _211_
timestamp 1486834041
transform 1 0 14336 0 1 21168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _212_
timestamp 1486834041
transform -1 0 8848 0 1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _213_
timestamp 1486834041
transform -1 0 7056 0 -1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _214_
timestamp 1486834041
transform -1 0 25648 0 1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _215_
timestamp 1486834041
transform -1 0 19040 0 1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _216_
timestamp 1486834041
transform -1 0 9744 0 1 5488
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _217_
timestamp 1486834041
transform -1 0 24528 0 1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _218_
timestamp 1486834041
transform 1 0 24416 0 -1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _219_
timestamp 1486834041
transform -1 0 24192 0 1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _220_
timestamp 1486834041
transform 1 0 1456 0 1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _221_
timestamp 1486834041
transform 1 0 1680 0 1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _222_
timestamp 1486834041
transform -1 0 3584 0 -1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _223_
timestamp 1486834041
transform 1 0 1680 0 1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _224_
timestamp 1486834041
transform -1 0 8512 0 -1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _225_
timestamp 1486834041
transform -1 0 8624 0 1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _226_
timestamp 1486834041
transform 1 0 1904 0 1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _227_
timestamp 1486834041
transform -1 0 7280 0 -1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _228_
timestamp 1486834041
transform 1 0 10080 0 -1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _229_
timestamp 1486834041
transform 1 0 9520 0 1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _230_
timestamp 1486834041
transform 1 0 17024 0 1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _231_
timestamp 1486834041
transform 1 0 17472 0 -1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _232_
timestamp 1486834041
transform 1 0 5712 0 1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _233_
timestamp 1486834041
transform 1 0 10976 0 -1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _234_
timestamp 1486834041
transform 1 0 11200 0 -1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _235_
timestamp 1486834041
transform 1 0 13440 0 -1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _236_
timestamp 1486834041
transform 1 0 2688 0 -1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _237_
timestamp 1486834041
transform -1 0 7840 0 -1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _238_
timestamp 1486834041
transform 1 0 3248 0 -1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _239_
timestamp 1486834041
transform 1 0 2352 0 1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _240_
timestamp 1486834041
transform 1 0 2352 0 1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _241_
timestamp 1486834041
transform 1 0 5264 0 -1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _242_
timestamp 1486834041
transform 1 0 10192 0 1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _243_
timestamp 1486834041
transform -1 0 18816 0 -1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _244_
timestamp 1486834041
transform 1 0 9184 0 -1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _245_
timestamp 1486834041
transform 1 0 10192 0 1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _246_
timestamp 1486834041
transform 1 0 14336 0 1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _247_
timestamp 1486834041
transform 1 0 11424 0 -1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _248_
timestamp 1486834041
transform 1 0 6608 0 1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _249_
timestamp 1486834041
transform 1 0 9072 0 1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _250_
timestamp 1486834041
transform 1 0 12208 0 -1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _251_
timestamp 1486834041
transform 1 0 11872 0 -1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _252_
timestamp 1486834041
transform 1 0 2016 0 1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _253_
timestamp 1486834041
transform 1 0 1680 0 1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _254_
timestamp 1486834041
transform 1 0 1344 0 -1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _255_
timestamp 1486834041
transform 1 0 1008 0 -1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _256_
timestamp 1486834041
transform 1 0 5824 0 -1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _257_
timestamp 1486834041
transform -1 0 9744 0 1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _258_
timestamp 1486834041
transform 1 0 12768 0 1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _259_
timestamp 1486834041
transform 1 0 13888 0 1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _260_
timestamp 1486834041
transform 1 0 6272 0 -1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _261_
timestamp 1486834041
transform 1 0 10192 0 1 39984
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _262_
timestamp 1486834041
transform 1 0 16688 0 -1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _263_
timestamp 1486834041
transform 1 0 17024 0 -1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _264_
timestamp 1486834041
transform 1 0 7728 0 1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _265_
timestamp 1486834041
transform 1 0 8960 0 1 7056
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _266_
timestamp 1486834041
transform 1 0 12544 0 -1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _267_
timestamp 1486834041
transform 1 0 12992 0 -1 5488
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _268_
timestamp 1486834041
transform 1 0 896 0 -1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _269_
timestamp 1486834041
transform 1 0 1568 0 1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _270_
timestamp 1486834041
transform -1 0 3136 0 1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _271_
timestamp 1486834041
transform 1 0 1008 0 -1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _272_
timestamp 1486834041
transform 1 0 4032 0 -1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _273_
timestamp 1486834041
transform 1 0 5040 0 1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _274_
timestamp 1486834041
transform 1 0 18928 0 -1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _275_
timestamp 1486834041
transform 1 0 21168 0 -1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _276_
timestamp 1486834041
transform -1 0 10976 0 -1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _277_
timestamp 1486834041
transform 1 0 8736 0 -1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _278_
timestamp 1486834041
transform 1 0 9184 0 -1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _279_
timestamp 1486834041
transform 1 0 10080 0 1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _280_
timestamp 1486834041
transform 1 0 10528 0 -1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _281_
timestamp 1486834041
transform 1 0 13104 0 -1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _282_
timestamp 1486834041
transform 1 0 12656 0 1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _283_
timestamp 1486834041
transform 1 0 10192 0 1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _284_
timestamp 1486834041
transform 1 0 896 0 1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _285_
timestamp 1486834041
transform 1 0 1344 0 -1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _286_
timestamp 1486834041
transform 1 0 5264 0 1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _287_
timestamp 1486834041
transform 1 0 2352 0 1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _288_
timestamp 1486834041
transform 1 0 6048 0 1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _289_
timestamp 1486834041
transform 1 0 6272 0 -1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _290_
timestamp 1486834041
transform -1 0 5040 0 -1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _291_
timestamp 1486834041
transform 1 0 2352 0 1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _292_
timestamp 1486834041
transform 1 0 6160 0 1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _293_
timestamp 1486834041
transform -1 0 10976 0 -1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _294_
timestamp 1486834041
transform 1 0 18032 0 -1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _295_
timestamp 1486834041
transform 1 0 17808 0 -1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _296_
timestamp 1486834041
transform 1 0 10864 0 -1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _297_
timestamp 1486834041
transform 1 0 9632 0 -1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _298_
timestamp 1486834041
transform 1 0 11872 0 -1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _299_
timestamp 1486834041
transform 1 0 10080 0 -1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _300_
timestamp 1486834041
transform 1 0 2352 0 1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _301_
timestamp 1486834041
transform 1 0 1680 0 -1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _302_
timestamp 1486834041
transform 1 0 13104 0 1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _303_
timestamp 1486834041
transform 1 0 6944 0 1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _304_
timestamp 1486834041
transform 1 0 896 0 -1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _305_
timestamp 1486834041
transform 1 0 1904 0 1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _306_
timestamp 1486834041
transform 1 0 20160 0 -1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _307_
timestamp 1486834041
transform 1 0 20496 0 1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _308_
timestamp 1486834041
transform 1 0 8176 0 1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _309_
timestamp 1486834041
transform 1 0 7840 0 1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _310_
timestamp 1486834041
transform 1 0 19376 0 -1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _311_
timestamp 1486834041
transform 1 0 18032 0 1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _312_
timestamp 1486834041
transform 1 0 7952 0 1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _313_
timestamp 1486834041
transform 1 0 6272 0 -1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _314_
timestamp 1486834041
transform 1 0 14112 0 -1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _315_
timestamp 1486834041
transform 1 0 12880 0 1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _316_
timestamp 1486834041
transform 1 0 896 0 1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _317_
timestamp 1486834041
transform 1 0 1344 0 1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _318_
timestamp 1486834041
transform 1 0 6608 0 1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _319_
timestamp 1486834041
transform 1 0 10192 0 -1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _320_
timestamp 1486834041
transform 1 0 6160 0 1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _321_
timestamp 1486834041
transform 1 0 6272 0 -1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _322_
timestamp 1486834041
transform 1 0 14112 0 1 39984
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _323_
timestamp 1486834041
transform 1 0 13552 0 -1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _324_
timestamp 1486834041
transform 1 0 14112 0 -1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _325_
timestamp 1486834041
transform 1 0 14112 0 -1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _326_
timestamp 1486834041
transform 1 0 17808 0 1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _327_
timestamp 1486834041
transform 1 0 17808 0 1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _328_
timestamp 1486834041
transform 1 0 14560 0 1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _329_
timestamp 1486834041
transform 1 0 11984 0 -1 7056
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _330_
timestamp 1486834041
transform 1 0 12656 0 1 7056
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _331_
timestamp 1486834041
transform 1 0 14336 0 1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _332_
timestamp 1486834041
transform 1 0 12768 0 -1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _333_
timestamp 1486834041
transform 1 0 14112 0 -1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _334_
timestamp 1486834041
transform 1 0 14560 0 1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _335_
timestamp 1486834041
transform 1 0 4928 0 -1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _336_
timestamp 1486834041
transform -1 0 4592 0 1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _337_
timestamp 1486834041
transform 1 0 4816 0 1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _338_
timestamp 1486834041
transform 1 0 16240 0 1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _339_
timestamp 1486834041
transform -1 0 23520 0 -1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _340_
timestamp 1486834041
transform 1 0 7952 0 1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _341_
timestamp 1486834041
transform 1 0 10192 0 1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _342_
timestamp 1486834041
transform 1 0 9632 0 -1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _343_
timestamp 1486834041
transform 1 0 10192 0 1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _344_
timestamp 1486834041
transform 1 0 10304 0 -1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _345_
timestamp 1486834041
transform -1 0 23408 0 -1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _346_
timestamp 1486834041
transform -1 0 20272 0 1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _347_
timestamp 1486834041
transform -1 0 23408 0 1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _348_
timestamp 1486834041
transform 1 0 3808 0 -1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _349_
timestamp 1486834041
transform 1 0 4816 0 1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _350_
timestamp 1486834041
transform 1 0 4704 0 -1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _351_
timestamp 1486834041
transform 1 0 4592 0 -1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_4  _352_
timestamp 1486834041
transform 1 0 12320 0 -1 33712
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_4  _353_
timestamp 1486834041
transform 1 0 8400 0 1 36848
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_4  _354_
timestamp 1486834041
transform 1 0 12656 0 1 33712
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_4  _355_
timestamp 1486834041
transform 1 0 8400 0 1 35280
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _356_
timestamp 1486834041
transform -1 0 11312 0 -1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _357_
timestamp 1486834041
transform 1 0 19376 0 1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _358_
timestamp 1486834041
transform 1 0 12656 0 1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _359_
timestamp 1486834041
transform 1 0 15120 0 1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _360_
timestamp 1486834041
transform -1 0 5712 0 1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _361_
timestamp 1486834041
transform 1 0 8736 0 -1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _362_
timestamp 1486834041
transform 1 0 8736 0 -1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _363_
timestamp 1486834041
transform 1 0 15344 0 -1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _364_
timestamp 1486834041
transform -1 0 12432 0 1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _365_
timestamp 1486834041
transform 1 0 18032 0 1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _366_
timestamp 1486834041
transform 1 0 9632 0 -1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _367_
timestamp 1486834041
transform 1 0 15008 0 -1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _368_
timestamp 1486834041
transform 1 0 4816 0 1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _369_
timestamp 1486834041
transform 1 0 3136 0 1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _370_
timestamp 1486834041
transform -1 0 5936 0 1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _371_
timestamp 1486834041
transform 1 0 15344 0 -1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _372_
timestamp 1486834041
transform -1 0 13552 0 1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _373_
timestamp 1486834041
transform 1 0 18480 0 -1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _374_
timestamp 1486834041
transform -1 0 10416 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _375_
timestamp 1486834041
transform 1 0 15232 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _376_
timestamp 1486834041
transform 1 0 4816 0 1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _377_
timestamp 1486834041
transform 1 0 16576 0 -1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _378_
timestamp 1486834041
transform -1 0 1904 0 1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _379_
timestamp 1486834041
transform 1 0 21616 0 -1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _380_
timestamp 1486834041
transform -1 0 10416 0 -1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _381_
timestamp 1486834041
transform 1 0 20496 0 1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _382_
timestamp 1486834041
transform 1 0 9744 0 -1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _383_
timestamp 1486834041
transform 1 0 16576 0 -1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _384_
timestamp 1486834041
transform -1 0 2016 0 -1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _385_
timestamp 1486834041
transform 1 0 13328 0 1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _386_
timestamp 1486834041
transform 1 0 9408 0 -1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _387_
timestamp 1486834041
transform 1 0 16576 0 -1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _388_
timestamp 1486834041
transform 1 0 4816 0 1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _389_
timestamp 1486834041
transform 1 0 1792 0 -1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _390_
timestamp 1486834041
transform -1 0 7168 0 -1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _391_
timestamp 1486834041
transform 1 0 21392 0 1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _392_
timestamp 1486834041
transform 1 0 10416 0 1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _393_
timestamp 1486834041
transform -1 0 11088 0 -1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _394_
timestamp 1486834041
transform 1 0 15344 0 -1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _395_
timestamp 1486834041
transform -1 0 14000 0 1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _396_
timestamp 1486834041
transform 1 0 3136 0 1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _397_
timestamp 1486834041
transform 1 0 5712 0 1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _398_
timestamp 1486834041
transform 1 0 7616 0 -1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _399_
timestamp 1486834041
transform -1 0 2800 0 -1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _400_
timestamp 1486834041
transform 1 0 8848 0 -1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _401_
timestamp 1486834041
transform -1 0 21392 0 1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _402_
timestamp 1486834041
transform -1 0 15904 0 -1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _403_
timestamp 1486834041
transform 1 0 13328 0 1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _404_
timestamp 1486834041
transform 1 0 8736 0 -1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _405_
timestamp 1486834041
transform 1 0 5264 0 1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _406_
timestamp 1486834041
transform 1 0 3696 0 1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _407_
timestamp 1486834041
transform 1 0 11536 0 1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _408_
timestamp 1486834041
transform 1 0 16240 0 1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _409_
timestamp 1486834041
transform 1 0 15008 0 -1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _410_
timestamp 1486834041
transform 1 0 19040 0 1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _411_
timestamp 1486834041
transform 1 0 17248 0 -1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _412_
timestamp 1486834041
transform 1 0 7056 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _413_
timestamp 1486834041
transform 1 0 10864 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _414_
timestamp 1486834041
transform 1 0 12096 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _415_
timestamp 1486834041
transform 1 0 11424 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _416_
timestamp 1486834041
transform 1 0 1456 0 1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _417_
timestamp 1486834041
transform 1 0 3584 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _418_
timestamp 1486834041
transform 1 0 3696 0 1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _419_
timestamp 1486834041
transform 1 0 1456 0 1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _420_
timestamp 1486834041
transform 1 0 1008 0 1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _421_
timestamp 1486834041
transform 1 0 2352 0 -1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _422_
timestamp 1486834041
transform 1 0 22400 0 -1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _423_
timestamp 1486834041
transform 1 0 22736 0 -1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _424_
timestamp 1486834041
transform 1 0 9184 0 -1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _425_
timestamp 1486834041
transform 1 0 6608 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _426_
timestamp 1486834041
transform 1 0 23296 0 1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _427_
timestamp 1486834041
transform 1 0 17136 0 1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _428_
timestamp 1486834041
transform 1 0 7616 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _429_
timestamp 1486834041
transform 1 0 23072 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _430_
timestamp 1486834041
transform -1 0 25312 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _431_
timestamp 1486834041
transform 1 0 11312 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _432_
timestamp 1486834041
transform 1 0 4816 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _433_
timestamp 1486834041
transform 1 0 2464 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _434_
timestamp 1486834041
transform 1 0 5712 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _435_
timestamp 1486834041
transform 1 0 2464 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _436_
timestamp 1486834041
transform -1 0 8064 0 -1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _437_
timestamp 1486834041
transform 1 0 2464 0 -1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _438_
timestamp 1486834041
transform -1 0 20608 0 -1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _439_
timestamp 1486834041
transform 1 0 1456 0 1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _440_
timestamp 1486834041
transform -1 0 25312 0 -1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _441_
timestamp 1486834041
transform 1 0 25760 0 -1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _442_
timestamp 1486834041
transform 1 0 20496 0 1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _443_
timestamp 1486834041
transform 1 0 25200 0 1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _444_
timestamp 1486834041
transform 1 0 18928 0 1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _445_
timestamp 1486834041
transform 1 0 25760 0 -1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _446_
timestamp 1486834041
transform 1 0 26656 0 -1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _447_
timestamp 1486834041
transform 1 0 19824 0 -1 55664
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _448_
timestamp 1486834041
transform 1 0 25872 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _449_
timestamp 1486834041
transform 1 0 26768 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _450_
timestamp 1486834041
transform 1 0 21280 0 -1 52528
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _451_
timestamp 1486834041
transform -1 0 14000 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _452_
timestamp 1486834041
transform -1 0 22624 0 -1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _453_
timestamp 1486834041
transform -1 0 24192 0 -1 50960
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _454_
timestamp 1486834041
transform -1 0 12208 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _455_
timestamp 1486834041
transform -1 0 3808 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _456_
timestamp 1486834041
transform -1 0 10752 0 -1 36848
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_UserCLK_regs
timestamp 1486834041
transform 1 0 12656 0 1 35280
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_UserCLK
timestamp 1486834041
transform 1 0 10752 0 -1 35280
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_UserCLK
timestamp 1486834041
transform -1 0 15344 0 -1 39984
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_UserCLK_regs
timestamp 1486834041
transform 1 0 13440 0 1 32144
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_UserCLK_regs
timestamp 1486834041
transform -1 0 14896 0 -1 38416
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_regs_0_UserCLK
timestamp 1486834041
transform 1 0 10752 0 -1 36848
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout38
timestamp 1486834041
transform 1 0 6384 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout39
timestamp 1486834041
transform 1 0 10416 0 1 19600
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout40
timestamp 1486834041
transform 1 0 6272 0 1 27440
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout41
timestamp 1486834041
transform 1 0 6944 0 -1 29008
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout42
timestamp 1486834041
transform 1 0 8736 0 -1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout43
timestamp 1486834041
transform 1 0 5936 0 1 22736
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout44
timestamp 1486834041
transform 1 0 4816 0 1 32144
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout45
timestamp 1486834041
transform 1 0 4816 0 1 33712
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout46
timestamp 1486834041
transform -1 0 4144 0 -1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout47
timestamp 1486834041
transform -1 0 2464 0 -1 30576
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout48
timestamp 1486834041
transform 1 0 6944 0 -1 30576
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout49
timestamp 1486834041
transform -1 0 5488 0 -1 29008
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout50
timestamp 1486834041
transform -1 0 1792 0 1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout51
timestamp 1486834041
transform -1 0 14224 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout52
timestamp 1486834041
transform 1 0 12656 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout53
timestamp 1486834041
transform 1 0 8624 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout54
timestamp 1486834041
transform -1 0 8176 0 -1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout55
timestamp 1486834041
transform 1 0 11536 0 -1 41552
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2
timestamp 1486834041
transform 1 0 896 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36
timestamp 1486834041
transform 1 0 4704 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_70
timestamp 1486834041
transform 1 0 8512 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_104
timestamp 1486834041
transform 1 0 12320 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_138
timestamp 1486834041
transform 1 0 16128 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_172
timestamp 1486834041
transform 1 0 19936 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_206
timestamp 1486834041
transform 1 0 23744 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_240
timestamp 1486834041
transform 1 0 27552 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_2
timestamp 1486834041
transform 1 0 896 0 -1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_66
timestamp 1486834041
transform 1 0 8064 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_72
timestamp 1486834041
transform 1 0 8736 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_88
timestamp 1486834041
transform 1 0 10528 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_92
timestamp 1486834041
transform 1 0 10976 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_94
timestamp 1486834041
transform 1 0 11200 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_103
timestamp 1486834041
transform 1 0 12208 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_119
timestamp 1486834041
transform 1 0 14000 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_135
timestamp 1486834041
transform 1 0 15792 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_139
timestamp 1486834041
transform 1 0 16240 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_142
timestamp 1486834041
transform 1 0 16576 0 -1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_206
timestamp 1486834041
transform 1 0 23744 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_212
timestamp 1486834041
transform 1 0 24416 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_220
timestamp 1486834041
transform 1 0 25312 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_224
timestamp 1486834041
transform 1 0 25760 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_2
timestamp 1486834041
transform 1 0 896 0 1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1486834041
transform 1 0 4480 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_37
timestamp 1486834041
transform 1 0 4816 0 1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_101
timestamp 1486834041
transform 1 0 11984 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_107
timestamp 1486834041
transform 1 0 12656 0 1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_171
timestamp 1486834041
transform 1 0 19824 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_177
timestamp 1486834041
transform 1 0 20496 0 1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_16
timestamp 1486834041
transform 1 0 2464 0 -1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_48
timestamp 1486834041
transform 1 0 6048 0 -1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_64
timestamp 1486834041
transform 1 0 7840 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_68
timestamp 1486834041
transform 1 0 8288 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_72
timestamp 1486834041
transform 1 0 8736 0 -1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_136
timestamp 1486834041
transform 1 0 15904 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_142
timestamp 1486834041
transform 1 0 16576 0 -1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_206
timestamp 1486834041
transform 1 0 23744 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_212
timestamp 1486834041
transform 1 0 24416 0 -1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_228
timestamp 1486834041
transform 1 0 26208 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_236
timestamp 1486834041
transform 1 0 27104 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_240
timestamp 1486834041
transform 1 0 27552 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_16
timestamp 1486834041
transform 1 0 2464 0 1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_32
timestamp 1486834041
transform 1 0 4256 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1486834041
transform 1 0 4480 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_37
timestamp 1486834041
transform 1 0 4816 0 1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_101
timestamp 1486834041
transform 1 0 11984 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_107
timestamp 1486834041
transform 1 0 12656 0 1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_171
timestamp 1486834041
transform 1 0 19824 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_177
timestamp 1486834041
transform 1 0 20496 0 1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_16
timestamp 1486834041
transform 1 0 2464 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_28
timestamp 1486834041
transform 1 0 3808 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_60
timestamp 1486834041
transform 1 0 7392 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_72
timestamp 1486834041
transform 1 0 8736 0 -1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_88
timestamp 1486834041
transform 1 0 10528 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_96
timestamp 1486834041
transform 1 0 11424 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_100
timestamp 1486834041
transform 1 0 11872 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_138
timestamp 1486834041
transform 1 0 16128 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_142
timestamp 1486834041
transform 1 0 16576 0 -1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_206
timestamp 1486834041
transform 1 0 23744 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_212
timestamp 1486834041
transform 1 0 24416 0 -1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_228
timestamp 1486834041
transform 1 0 26208 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_236
timestamp 1486834041
transform 1 0 27104 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_240
timestamp 1486834041
transform 1 0 27552 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_24
timestamp 1486834041
transform 1 0 3360 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_32
timestamp 1486834041
transform 1 0 4256 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1486834041
transform 1 0 4480 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_37
timestamp 1486834041
transform 1 0 4816 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_53
timestamp 1486834041
transform 1 0 6608 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_81
timestamp 1486834041
transform 1 0 9744 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_89
timestamp 1486834041
transform 1 0 10640 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_93
timestamp 1486834041
transform 1 0 11088 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_95
timestamp 1486834041
transform 1 0 11312 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_104
timestamp 1486834041
transform 1 0 12320 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_107
timestamp 1486834041
transform 1 0 12656 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_115
timestamp 1486834041
transform 1 0 13552 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_148
timestamp 1486834041
transform 1 0 17248 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_164
timestamp 1486834041
transform 1 0 19040 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_172
timestamp 1486834041
transform 1 0 19936 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_174
timestamp 1486834041
transform 1 0 20160 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_177
timestamp 1486834041
transform 1 0 20496 0 1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_30
timestamp 1486834041
transform 1 0 4032 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_62
timestamp 1486834041
transform 1 0 7616 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_72
timestamp 1486834041
transform 1 0 8736 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_76
timestamp 1486834041
transform 1 0 9184 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_78
timestamp 1486834041
transform 1 0 9408 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_87
timestamp 1486834041
transform 1 0 10416 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_99
timestamp 1486834041
transform 1 0 11760 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_121
timestamp 1486834041
transform 1 0 14224 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_137
timestamp 1486834041
transform 1 0 16016 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_139
timestamp 1486834041
transform 1 0 16240 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_142
timestamp 1486834041
transform 1 0 16576 0 -1 7056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_206
timestamp 1486834041
transform 1 0 23744 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_212
timestamp 1486834041
transform 1 0 24416 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_228
timestamp 1486834041
transform 1 0 26208 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_236
timestamp 1486834041
transform 1 0 27104 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_240
timestamp 1486834041
transform 1 0 27552 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_30
timestamp 1486834041
transform 1 0 4032 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1486834041
transform 1 0 4480 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_37
timestamp 1486834041
transform 1 0 4816 0 1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_61
timestamp 1486834041
transform 1 0 7504 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_69
timestamp 1486834041
transform 1 0 8400 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_73
timestamp 1486834041
transform 1 0 8848 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_94
timestamp 1486834041
transform 1 0 11200 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_98
timestamp 1486834041
transform 1 0 11648 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_100
timestamp 1486834041
transform 1 0 11872 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_127
timestamp 1486834041
transform 1 0 14896 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_131
timestamp 1486834041
transform 1 0 15344 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_151
timestamp 1486834041
transform 1 0 17584 0 1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_167
timestamp 1486834041
transform 1 0 19376 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_177
timestamp 1486834041
transform 1 0 20496 0 1 7056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_30
timestamp 1486834041
transform 1 0 4032 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_34
timestamp 1486834041
transform 1 0 4480 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_36
timestamp 1486834041
transform 1 0 4704 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_72
timestamp 1486834041
transform 1 0 8736 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_80
timestamp 1486834041
transform 1 0 9632 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_84
timestamp 1486834041
transform 1 0 10080 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_154
timestamp 1486834041
transform 1 0 17920 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_162
timestamp 1486834041
transform 1 0 18816 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_166
timestamp 1486834041
transform 1 0 19264 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_199
timestamp 1486834041
transform 1 0 22960 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_207
timestamp 1486834041
transform 1 0 23856 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_209
timestamp 1486834041
transform 1 0 24080 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_212
timestamp 1486834041
transform 1 0 24416 0 -1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_228
timestamp 1486834041
transform 1 0 26208 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_236
timestamp 1486834041
transform 1 0 27104 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_240
timestamp 1486834041
transform 1 0 27552 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_30
timestamp 1486834041
transform 1 0 4032 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1486834041
transform 1 0 4480 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_53
timestamp 1486834041
transform 1 0 6608 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_83
timestamp 1486834041
transform 1 0 9968 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_121
timestamp 1486834041
transform 1 0 14224 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_123
timestamp 1486834041
transform 1 0 14448 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_164
timestamp 1486834041
transform 1 0 19040 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_172
timestamp 1486834041
transform 1 0 19936 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_174
timestamp 1486834041
transform 1 0 20160 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_177
timestamp 1486834041
transform 1 0 20496 0 1 8624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_30
timestamp 1486834041
transform 1 0 4032 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_34
timestamp 1486834041
transform 1 0 4480 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_55
timestamp 1486834041
transform 1 0 6832 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_66
timestamp 1486834041
transform 1 0 8064 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_72
timestamp 1486834041
transform 1 0 8736 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_124
timestamp 1486834041
transform 1 0 14560 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_150
timestamp 1486834041
transform 1 0 17472 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_152
timestamp 1486834041
transform 1 0 17696 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_185
timestamp 1486834041
transform 1 0 21392 0 -1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_201
timestamp 1486834041
transform 1 0 23184 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_209
timestamp 1486834041
transform 1 0 24080 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_212
timestamp 1486834041
transform 1 0 24416 0 -1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_228
timestamp 1486834041
transform 1 0 26208 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_236
timestamp 1486834041
transform 1 0 27104 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_240
timestamp 1486834041
transform 1 0 27552 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_2
timestamp 1486834041
transform 1 0 896 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_6
timestamp 1486834041
transform 1 0 1344 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_8
timestamp 1486834041
transform 1 0 1568 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_29
timestamp 1486834041
transform 1 0 3920 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_33
timestamp 1486834041
transform 1 0 4368 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_69
timestamp 1486834041
transform 1 0 8400 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_86
timestamp 1486834041
transform 1 0 10304 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_119
timestamp 1486834041
transform 1 0 14000 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_121
timestamp 1486834041
transform 1 0 14224 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_177
timestamp 1486834041
transform 1 0 20496 0 1 10192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_2
timestamp 1486834041
transform 1 0 896 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_34
timestamp 1486834041
transform 1 0 4480 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_84
timestamp 1486834041
transform 1 0 10080 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_88
timestamp 1486834041
transform 1 0 10528 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_123
timestamp 1486834041
transform 1 0 14448 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_127
timestamp 1486834041
transform 1 0 14896 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_129
timestamp 1486834041
transform 1 0 15120 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_136
timestamp 1486834041
transform 1 0 15904 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_148
timestamp 1486834041
transform 1 0 17248 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_150
timestamp 1486834041
transform 1 0 17472 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_183
timestamp 1486834041
transform 1 0 21168 0 -1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_199
timestamp 1486834041
transform 1 0 22960 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_208
timestamp 1486834041
transform 1 0 23968 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_212
timestamp 1486834041
transform 1 0 24416 0 -1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_228
timestamp 1486834041
transform 1 0 26208 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_236
timestamp 1486834041
transform 1 0 27104 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_240
timestamp 1486834041
transform 1 0 27552 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_2
timestamp 1486834041
transform 1 0 896 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_6
timestamp 1486834041
transform 1 0 1344 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_8
timestamp 1486834041
transform 1 0 1568 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_29
timestamp 1486834041
transform 1 0 3920 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_33
timestamp 1486834041
transform 1 0 4368 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_103
timestamp 1486834041
transform 1 0 12208 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_121
timestamp 1486834041
transform 1 0 14224 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_123
timestamp 1486834041
transform 1 0 14448 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_174
timestamp 1486834041
transform 1 0 20160 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_189
timestamp 1486834041
transform 1 0 21840 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_213
timestamp 1486834041
transform 1 0 24528 0 1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_229
timestamp 1486834041
transform 1 0 26320 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_237
timestamp 1486834041
transform 1 0 27216 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_78
timestamp 1486834041
transform 1 0 9408 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_163
timestamp 1486834041
transform 1 0 18928 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_196
timestamp 1486834041
transform 1 0 22624 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_204
timestamp 1486834041
transform 1 0 23520 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_208
timestamp 1486834041
transform 1 0 23968 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_220
timestamp 1486834041
transform 1 0 25312 0 -1 13328
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_236
timestamp 1486834041
transform 1 0 27104 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_240
timestamp 1486834041
transform 1 0 27552 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_2
timestamp 1486834041
transform 1 0 896 0 1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_6
timestamp 1486834041
transform 1 0 1344 0 1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_51
timestamp 1486834041
transform 1 0 6384 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_113
timestamp 1486834041
transform 1 0 13328 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_162
timestamp 1486834041
transform 1 0 18816 0 1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_223
timestamp 1486834041
transform 1 0 25648 0 1 13328
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_239
timestamp 1486834041
transform 1 0 27440 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_2
timestamp 1486834041
transform 1 0 896 0 -1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_26
timestamp 1486834041
transform 1 0 3584 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_79
timestamp 1486834041
transform 1 0 9520 0 -1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_148
timestamp 1486834041
transform 1 0 17248 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_150
timestamp 1486834041
transform 1 0 17472 0 -1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_203
timestamp 1486834041
transform 1 0 23408 0 -1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_207
timestamp 1486834041
transform 1 0 23856 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_209
timestamp 1486834041
transform 1 0 24080 0 -1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_232
timestamp 1486834041
transform 1 0 26656 0 -1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_240
timestamp 1486834041
transform 1 0 27552 0 -1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_2
timestamp 1486834041
transform 1 0 896 0 1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_6
timestamp 1486834041
transform 1 0 1344 0 1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_107
timestamp 1486834041
transform 1 0 12656 0 1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_115
timestamp 1486834041
transform 1 0 13552 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_117
timestamp 1486834041
transform 1 0 13776 0 1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_156
timestamp 1486834041
transform 1 0 18144 0 1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_167
timestamp 1486834041
transform 1 0 19376 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_209
timestamp 1486834041
transform 1 0 24080 0 1 14896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_2
timestamp 1486834041
transform 1 0 896 0 -1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_43
timestamp 1486834041
transform 1 0 5488 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_78
timestamp 1486834041
transform 1 0 9408 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_80
timestamp 1486834041
transform 1 0 9632 0 -1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_89
timestamp 1486834041
transform 1 0 10640 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_139
timestamp 1486834041
transform 1 0 16240 0 -1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_194
timestamp 1486834041
transform 1 0 22400 0 -1 16464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_212
timestamp 1486834041
transform 1 0 24416 0 -1 16464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_228
timestamp 1486834041
transform 1 0 26208 0 -1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_236
timestamp 1486834041
transform 1 0 27104 0 -1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_240
timestamp 1486834041
transform 1 0 27552 0 -1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_30
timestamp 1486834041
transform 1 0 4032 0 1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_34
timestamp 1486834041
transform 1 0 4480 0 1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_51
timestamp 1486834041
transform 1 0 6384 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_107
timestamp 1486834041
transform 1 0 12656 0 1 16464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_123
timestamp 1486834041
transform 1 0 14448 0 1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_174
timestamp 1486834041
transform 1 0 20160 0 1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_183
timestamp 1486834041
transform 1 0 21168 0 1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_187
timestamp 1486834041
transform 1 0 21616 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_189
timestamp 1486834041
transform 1 0 21840 0 1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_210
timestamp 1486834041
transform 1 0 24192 0 1 16464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_226
timestamp 1486834041
transform 1 0 25984 0 1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_234
timestamp 1486834041
transform 1 0 26880 0 1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_238
timestamp 1486834041
transform 1 0 27328 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_240
timestamp 1486834041
transform 1 0 27552 0 1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_2
timestamp 1486834041
transform 1 0 896 0 -1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_120
timestamp 1486834041
transform 1 0 14112 0 -1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_136
timestamp 1486834041
transform 1 0 15904 0 -1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_204
timestamp 1486834041
transform 1 0 23520 0 -1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_208
timestamp 1486834041
transform 1 0 23968 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_220
timestamp 1486834041
transform 1 0 25312 0 -1 18032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_236
timestamp 1486834041
transform 1 0 27104 0 -1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_240
timestamp 1486834041
transform 1 0 27552 0 -1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_2
timestamp 1486834041
transform 1 0 896 0 1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_6
timestamp 1486834041
transform 1 0 1344 0 1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_127
timestamp 1486834041
transform 1 0 14896 0 1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_131
timestamp 1486834041
transform 1 0 15344 0 1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_172
timestamp 1486834041
transform 1 0 19936 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_174
timestamp 1486834041
transform 1 0 20160 0 1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_209
timestamp 1486834041
transform 1 0 24080 0 1 18032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_16
timestamp 1486834041
transform 1 0 2464 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_72
timestamp 1486834041
transform 1 0 8736 0 -1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_142
timestamp 1486834041
transform 1 0 16576 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_186
timestamp 1486834041
transform 1 0 21504 0 -1 19600
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_202
timestamp 1486834041
transform 1 0 23296 0 -1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_212
timestamp 1486834041
transform 1 0 24416 0 -1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_220
timestamp 1486834041
transform 1 0 25312 0 -1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_232
timestamp 1486834041
transform 1 0 26656 0 -1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_240
timestamp 1486834041
transform 1 0 27552 0 -1 19600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_2
timestamp 1486834041
transform 1 0 896 0 1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_26
timestamp 1486834041
transform 1 0 3584 0 1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_34
timestamp 1486834041
transform 1 0 4480 0 1 19600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_51
timestamp 1486834041
transform 1 0 6384 0 1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_101
timestamp 1486834041
transform 1 0 11984 0 1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_165
timestamp 1486834041
transform 1 0 19152 0 1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_183
timestamp 1486834041
transform 1 0 21168 0 1 19600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_215
timestamp 1486834041
transform 1 0 24752 0 1 19600
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_231
timestamp 1486834041
transform 1 0 26544 0 1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_239
timestamp 1486834041
transform 1 0 27440 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_2
timestamp 1486834041
transform 1 0 896 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_64
timestamp 1486834041
transform 1 0 7840 0 -1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_68
timestamp 1486834041
transform 1 0 8288 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_80
timestamp 1486834041
transform 1 0 9632 0 -1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_84
timestamp 1486834041
transform 1 0 10080 0 -1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_117
timestamp 1486834041
transform 1 0 13776 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_119
timestamp 1486834041
transform 1 0 14000 0 -1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_157
timestamp 1486834041
transform 1 0 18256 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_159
timestamp 1486834041
transform 1 0 18480 0 -1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_192
timestamp 1486834041
transform 1 0 22176 0 -1 21168
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_208
timestamp 1486834041
transform 1 0 23968 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_212
timestamp 1486834041
transform 1 0 24416 0 -1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_220
timestamp 1486834041
transform 1 0 25312 0 -1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_240
timestamp 1486834041
transform 1 0 27552 0 -1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_2
timestamp 1486834041
transform 1 0 896 0 1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_10
timestamp 1486834041
transform 1 0 1792 0 1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_14
timestamp 1486834041
transform 1 0 2240 0 1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_37
timestamp 1486834041
transform 1 0 4816 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_39
timestamp 1486834041
transform 1 0 5040 0 1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_72
timestamp 1486834041
transform 1 0 8736 0 1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_80
timestamp 1486834041
transform 1 0 9632 0 1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_84
timestamp 1486834041
transform 1 0 10080 0 1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_107
timestamp 1486834041
transform 1 0 12656 0 1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_111
timestamp 1486834041
transform 1 0 13104 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_121
timestamp 1486834041
transform 1 0 14224 0 1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_154
timestamp 1486834041
transform 1 0 17920 0 1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_200
timestamp 1486834041
transform 1 0 23072 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_210
timestamp 1486834041
transform 1 0 24192 0 1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_218
timestamp 1486834041
transform 1 0 25088 0 1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_36
timestamp 1486834041
transform 1 0 4704 0 -1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_40
timestamp 1486834041
transform 1 0 5152 0 -1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_61
timestamp 1486834041
transform 1 0 7504 0 -1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_69
timestamp 1486834041
transform 1 0 8400 0 -1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_72
timestamp 1486834041
transform 1 0 8736 0 -1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_116
timestamp 1486834041
transform 1 0 13664 0 -1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_162
timestamp 1486834041
transform 1 0 18816 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_164
timestamp 1486834041
transform 1 0 19040 0 -1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_205
timestamp 1486834041
transform 1 0 23632 0 -1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_209
timestamp 1486834041
transform 1 0 24080 0 -1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_212
timestamp 1486834041
transform 1 0 24416 0 -1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_2
timestamp 1486834041
transform 1 0 896 0 1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_31
timestamp 1486834041
transform 1 0 4144 0 1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_37
timestamp 1486834041
transform 1 0 4816 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_81
timestamp 1486834041
transform 1 0 9744 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_83
timestamp 1486834041
transform 1 0 9968 0 1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_104
timestamp 1486834041
transform 1 0 12320 0 1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_107
timestamp 1486834041
transform 1 0 12656 0 1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_119
timestamp 1486834041
transform 1 0 14000 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_121
timestamp 1486834041
transform 1 0 14224 0 1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_142
timestamp 1486834041
transform 1 0 16576 0 1 22736
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_158
timestamp 1486834041
transform 1 0 18368 0 1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_166
timestamp 1486834041
transform 1 0 19264 0 1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_177
timestamp 1486834041
transform 1 0 20496 0 1 22736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_209
timestamp 1486834041
transform 1 0 24080 0 1 22736
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_225
timestamp 1486834041
transform 1 0 25872 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_2
timestamp 1486834041
transform 1 0 896 0 -1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_10
timestamp 1486834041
transform 1 0 1792 0 -1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_66
timestamp 1486834041
transform 1 0 8064 0 -1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_72
timestamp 1486834041
transform 1 0 8736 0 -1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_80
timestamp 1486834041
transform 1 0 9632 0 -1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_84
timestamp 1486834041
transform 1 0 10080 0 -1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_125
timestamp 1486834041
transform 1 0 14672 0 -1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_129
timestamp 1486834041
transform 1 0 15120 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_139
timestamp 1486834041
transform 1 0 16240 0 -1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_202
timestamp 1486834041
transform 1 0 23296 0 -1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_212
timestamp 1486834041
transform 1 0 24416 0 -1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_2
timestamp 1486834041
transform 1 0 896 0 1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_6
timestamp 1486834041
transform 1 0 1344 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_28
timestamp 1486834041
transform 1 0 3808 0 1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_32
timestamp 1486834041
transform 1 0 4256 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_34
timestamp 1486834041
transform 1 0 4480 0 1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_51
timestamp 1486834041
transform 1 0 6384 0 1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_95
timestamp 1486834041
transform 1 0 11312 0 1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_103
timestamp 1486834041
transform 1 0 12208 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_115
timestamp 1486834041
transform 1 0 13552 0 1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_163
timestamp 1486834041
transform 1 0 18928 0 1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_171
timestamp 1486834041
transform 1 0 19824 0 1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_209
timestamp 1486834041
transform 1 0 24080 0 1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_48
timestamp 1486834041
transform 1 0 6048 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_112
timestamp 1486834041
transform 1 0 13216 0 -1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_150
timestamp 1486834041
transform 1 0 17472 0 -1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_158
timestamp 1486834041
transform 1 0 18368 0 -1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_195
timestamp 1486834041
transform 1 0 22512 0 -1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_203
timestamp 1486834041
transform 1 0 23408 0 -1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_207
timestamp 1486834041
transform 1 0 23856 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_209
timestamp 1486834041
transform 1 0 24080 0 -1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_212
timestamp 1486834041
transform 1 0 24416 0 -1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_2
timestamp 1486834041
transform 1 0 896 0 1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_6
timestamp 1486834041
transform 1 0 1344 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_8
timestamp 1486834041
transform 1 0 1568 0 1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_29
timestamp 1486834041
transform 1 0 3920 0 1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_33
timestamp 1486834041
transform 1 0 4368 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_45
timestamp 1486834041
transform 1 0 5712 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_47
timestamp 1486834041
transform 1 0 5936 0 1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_68
timestamp 1486834041
transform 1 0 8288 0 1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_72
timestamp 1486834041
transform 1 0 8736 0 1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_107
timestamp 1486834041
transform 1 0 12656 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_137
timestamp 1486834041
transform 1 0 16016 0 1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_145
timestamp 1486834041
transform 1 0 16912 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_197
timestamp 1486834041
transform 1 0 22736 0 1 25872
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_213
timestamp 1486834041
transform 1 0 24528 0 1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_221
timestamp 1486834041
transform 1 0 25424 0 1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_225
timestamp 1486834041
transform 1 0 25872 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_54
timestamp 1486834041
transform 1 0 6720 0 -1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_92
timestamp 1486834041
transform 1 0 10976 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_134
timestamp 1486834041
transform 1 0 15680 0 -1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_138
timestamp 1486834041
transform 1 0 16128 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_142
timestamp 1486834041
transform 1 0 16576 0 -1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_146
timestamp 1486834041
transform 1 0 17024 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_180
timestamp 1486834041
transform 1 0 20832 0 -1 27440
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_196
timestamp 1486834041
transform 1 0 22624 0 -1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_204
timestamp 1486834041
transform 1 0 23520 0 -1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_208
timestamp 1486834041
transform 1 0 23968 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_212
timestamp 1486834041
transform 1 0 24416 0 -1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_2
timestamp 1486834041
transform 1 0 896 0 1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_10
timestamp 1486834041
transform 1 0 1792 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_32
timestamp 1486834041
transform 1 0 4256 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_34
timestamp 1486834041
transform 1 0 4480 0 1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_45
timestamp 1486834041
transform 1 0 5712 0 1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_49
timestamp 1486834041
transform 1 0 6160 0 1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_84
timestamp 1486834041
transform 1 0 10080 0 1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_107
timestamp 1486834041
transform 1 0 12656 0 1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_111
timestamp 1486834041
transform 1 0 13104 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_113
timestamp 1486834041
transform 1 0 13328 0 1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_146
timestamp 1486834041
transform 1 0 17024 0 1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_150
timestamp 1486834041
transform 1 0 17472 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_152
timestamp 1486834041
transform 1 0 17696 0 1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_173
timestamp 1486834041
transform 1 0 20048 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_185
timestamp 1486834041
transform 1 0 21392 0 1 27440
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_201
timestamp 1486834041
transform 1 0 23184 0 1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_209
timestamp 1486834041
transform 1 0 24080 0 1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_2
timestamp 1486834041
transform 1 0 896 0 -1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_6
timestamp 1486834041
transform 1 0 1344 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_8
timestamp 1486834041
transform 1 0 1568 0 -1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_43
timestamp 1486834041
transform 1 0 5488 0 -1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_51
timestamp 1486834041
transform 1 0 6384 0 -1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_55
timestamp 1486834041
transform 1 0 6832 0 -1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_72
timestamp 1486834041
transform 1 0 8736 0 -1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_128
timestamp 1486834041
transform 1 0 15008 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_130
timestamp 1486834041
transform 1 0 15232 0 -1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_139
timestamp 1486834041
transform 1 0 16240 0 -1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_142
timestamp 1486834041
transform 1 0 16576 0 -1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_198
timestamp 1486834041
transform 1 0 22848 0 -1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_206
timestamp 1486834041
transform 1 0 23744 0 -1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_212
timestamp 1486834041
transform 1 0 24416 0 -1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_220
timestamp 1486834041
transform 1 0 25312 0 -1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_224
timestamp 1486834041
transform 1 0 25760 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_226
timestamp 1486834041
transform 1 0 25984 0 -1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_10
timestamp 1486834041
transform 1 0 1792 0 1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_14
timestamp 1486834041
transform 1 0 2240 0 1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_37
timestamp 1486834041
transform 1 0 4816 0 1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_61
timestamp 1486834041
transform 1 0 7504 0 1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_65
timestamp 1486834041
transform 1 0 7952 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_87
timestamp 1486834041
transform 1 0 10416 0 1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_95
timestamp 1486834041
transform 1 0 11312 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_107
timestamp 1486834041
transform 1 0 12656 0 1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_111
timestamp 1486834041
transform 1 0 13104 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_173
timestamp 1486834041
transform 1 0 20048 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_177
timestamp 1486834041
transform 1 0 20496 0 1 29008
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_209
timestamp 1486834041
transform 1 0 24080 0 1 29008
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_225
timestamp 1486834041
transform 1 0 25872 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_80
timestamp 1486834041
transform 1 0 9632 0 -1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_84
timestamp 1486834041
transform 1 0 10080 0 -1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_137
timestamp 1486834041
transform 1 0 16016 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_139
timestamp 1486834041
transform 1 0 16240 0 -1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_142
timestamp 1486834041
transform 1 0 16576 0 -1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_203
timestamp 1486834041
transform 1 0 23408 0 -1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_207
timestamp 1486834041
transform 1 0 23856 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_209
timestamp 1486834041
transform 1 0 24080 0 -1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_212
timestamp 1486834041
transform 1 0 24416 0 -1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_220
timestamp 1486834041
transform 1 0 25312 0 -1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_224
timestamp 1486834041
transform 1 0 25760 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_226
timestamp 1486834041
transform 1 0 25984 0 -1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_2
timestamp 1486834041
transform 1 0 896 0 1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_10
timestamp 1486834041
transform 1 0 1792 0 1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_14
timestamp 1486834041
transform 1 0 2240 0 1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_107
timestamp 1486834041
transform 1 0 12656 0 1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_163
timestamp 1486834041
transform 1 0 18928 0 1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_171
timestamp 1486834041
transform 1 0 19824 0 1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_209
timestamp 1486834041
transform 1 0 24080 0 1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_2
timestamp 1486834041
transform 1 0 896 0 -1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_26
timestamp 1486834041
transform 1 0 3584 0 -1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_34
timestamp 1486834041
transform 1 0 4480 0 -1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_72
timestamp 1486834041
transform 1 0 8736 0 -1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_76
timestamp 1486834041
transform 1 0 9184 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_78
timestamp 1486834041
transform 1 0 9408 0 -1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_127
timestamp 1486834041
transform 1 0 14896 0 -1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_135
timestamp 1486834041
transform 1 0 15792 0 -1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_139
timestamp 1486834041
transform 1 0 16240 0 -1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_150
timestamp 1486834041
transform 1 0 17472 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_152
timestamp 1486834041
transform 1 0 17696 0 -1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_205
timestamp 1486834041
transform 1 0 23632 0 -1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_209
timestamp 1486834041
transform 1 0 24080 0 -1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_212
timestamp 1486834041
transform 1 0 24416 0 -1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_30
timestamp 1486834041
transform 1 0 4032 0 1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_34
timestamp 1486834041
transform 1 0 4480 0 1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_51
timestamp 1486834041
transform 1 0 6384 0 1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_55
timestamp 1486834041
transform 1 0 6832 0 1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_76
timestamp 1486834041
transform 1 0 9184 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_78
timestamp 1486834041
transform 1 0 9408 0 1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_99
timestamp 1486834041
transform 1 0 11760 0 1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_103
timestamp 1486834041
transform 1 0 12208 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_107
timestamp 1486834041
transform 1 0 12656 0 1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_111
timestamp 1486834041
transform 1 0 13104 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_113
timestamp 1486834041
transform 1 0 13328 0 1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_172
timestamp 1486834041
transform 1 0 19936 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_174
timestamp 1486834041
transform 1 0 20160 0 1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_193
timestamp 1486834041
transform 1 0 22288 0 1 32144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_225
timestamp 1486834041
transform 1 0 25872 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_2
timestamp 1486834041
transform 1 0 896 0 -1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_10
timestamp 1486834041
transform 1 0 1792 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_12
timestamp 1486834041
transform 1 0 2016 0 -1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_45
timestamp 1486834041
transform 1 0 5712 0 -1 33712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_49
timestamp 1486834041
transform 1 0 6160 0 -1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_80
timestamp 1486834041
transform 1 0 9632 0 -1 33712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_142
timestamp 1486834041
transform 1 0 16576 0 -1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_150
timestamp 1486834041
transform 1 0 17472 0 -1 33712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_154
timestamp 1486834041
transform 1 0 17920 0 -1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_41_175
timestamp 1486834041
transform 1 0 20272 0 -1 33712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_207
timestamp 1486834041
transform 1 0 23856 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_209
timestamp 1486834041
transform 1 0 24080 0 -1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_212
timestamp 1486834041
transform 1 0 24416 0 -1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_2
timestamp 1486834041
transform 1 0 896 0 1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_103
timestamp 1486834041
transform 1 0 12208 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_143
timestamp 1486834041
transform 1 0 16688 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_145
timestamp 1486834041
transform 1 0 16912 0 1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_166
timestamp 1486834041
transform 1 0 19264 0 1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_177
timestamp 1486834041
transform 1 0 20496 0 1 33712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_209
timestamp 1486834041
transform 1 0 24080 0 1 33712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_2
timestamp 1486834041
transform 1 0 896 0 -1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_72
timestamp 1486834041
transform 1 0 8736 0 -1 35280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_76
timestamp 1486834041
transform 1 0 9184 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_86
timestamp 1486834041
transform 1 0 10304 0 -1 35280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_142
timestamp 1486834041
transform 1 0 16576 0 -1 35280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_146
timestamp 1486834041
transform 1 0 17024 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_188
timestamp 1486834041
transform 1 0 21728 0 -1 35280
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_204
timestamp 1486834041
transform 1 0 23520 0 -1 35280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_208
timestamp 1486834041
transform 1 0 23968 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_212
timestamp 1486834041
transform 1 0 24416 0 -1 35280
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_22
timestamp 1486834041
transform 1 0 3136 0 1 35280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_26
timestamp 1486834041
transform 1 0 3584 0 1 35280
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_37
timestamp 1486834041
transform 1 0 4816 0 1 35280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_157
timestamp 1486834041
transform 1 0 18256 0 1 35280
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_173
timestamp 1486834041
transform 1 0 20048 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_177
timestamp 1486834041
transform 1 0 20496 0 1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_209
timestamp 1486834041
transform 1 0 24080 0 1 35280
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_225
timestamp 1486834041
transform 1 0 25872 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_2
timestamp 1486834041
transform 1 0 896 0 -1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_10
timestamp 1486834041
transform 1 0 1792 0 -1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_67
timestamp 1486834041
transform 1 0 8176 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_69
timestamp 1486834041
transform 1 0 8400 0 -1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_72
timestamp 1486834041
transform 1 0 8736 0 -1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_80
timestamp 1486834041
transform 1 0 9632 0 -1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_45_178
timestamp 1486834041
transform 1 0 20608 0 -1 36848
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_212
timestamp 1486834041
transform 1 0 24416 0 -1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_2
timestamp 1486834041
transform 1 0 896 0 1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_6
timestamp 1486834041
transform 1 0 1344 0 1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_37
timestamp 1486834041
transform 1 0 4816 0 1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_45
timestamp 1486834041
transform 1 0 5712 0 1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_107
timestamp 1486834041
transform 1 0 12656 0 1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_160
timestamp 1486834041
transform 1 0 18592 0 1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_168
timestamp 1486834041
transform 1 0 19488 0 1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_172
timestamp 1486834041
transform 1 0 19936 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_174
timestamp 1486834041
transform 1 0 20160 0 1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_46_177
timestamp 1486834041
transform 1 0 20496 0 1 36848
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_209
timestamp 1486834041
transform 1 0 24080 0 1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_2
timestamp 1486834041
transform 1 0 896 0 -1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_23
timestamp 1486834041
transform 1 0 3248 0 -1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_27
timestamp 1486834041
transform 1 0 3696 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_29
timestamp 1486834041
transform 1 0 3920 0 -1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_72
timestamp 1486834041
transform 1 0 8736 0 -1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_76
timestamp 1486834041
transform 1 0 9184 0 -1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_127
timestamp 1486834041
transform 1 0 14896 0 -1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_136
timestamp 1486834041
transform 1 0 15904 0 -1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_142
timestamp 1486834041
transform 1 0 16576 0 -1 38416
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_206
timestamp 1486834041
transform 1 0 23744 0 -1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_212
timestamp 1486834041
transform 1 0 24416 0 -1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_2
timestamp 1486834041
transform 1 0 896 0 1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_31
timestamp 1486834041
transform 1 0 4144 0 1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_37
timestamp 1486834041
transform 1 0 4816 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_59
timestamp 1486834041
transform 1 0 7280 0 1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_63
timestamp 1486834041
transform 1 0 7728 0 1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_96
timestamp 1486834041
transform 1 0 11424 0 1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_147
timestamp 1486834041
transform 1 0 17136 0 1 38416
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_163
timestamp 1486834041
transform 1 0 18928 0 1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_171
timestamp 1486834041
transform 1 0 19824 0 1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_48_177
timestamp 1486834041
transform 1 0 20496 0 1 38416
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_209
timestamp 1486834041
transform 1 0 24080 0 1 38416
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_225
timestamp 1486834041
transform 1 0 25872 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_2
timestamp 1486834041
transform 1 0 896 0 -1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_10
timestamp 1486834041
transform 1 0 1792 0 -1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_14
timestamp 1486834041
transform 1 0 2240 0 -1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_31
timestamp 1486834041
transform 1 0 4144 0 -1 39984
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_47
timestamp 1486834041
transform 1 0 5936 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_49
timestamp 1486834041
transform 1 0 6160 0 -1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_66
timestamp 1486834041
transform 1 0 8064 0 -1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_72
timestamp 1486834041
transform 1 0 8736 0 -1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_131
timestamp 1486834041
transform 1 0 15344 0 -1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_139
timestamp 1486834041
transform 1 0 16240 0 -1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_142
timestamp 1486834041
transform 1 0 16576 0 -1 39984
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_206
timestamp 1486834041
transform 1 0 23744 0 -1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_212
timestamp 1486834041
transform 1 0 24416 0 -1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_2
timestamp 1486834041
transform 1 0 896 0 1 39984
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_34
timestamp 1486834041
transform 1 0 4480 0 1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_37
timestamp 1486834041
transform 1 0 4816 0 1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_45
timestamp 1486834041
transform 1 0 5712 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_79
timestamp 1486834041
transform 1 0 9520 0 1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_83
timestamp 1486834041
transform 1 0 9968 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_115
timestamp 1486834041
transform 1 0 13552 0 1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_119
timestamp 1486834041
transform 1 0 14000 0 1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_140
timestamp 1486834041
transform 1 0 16352 0 1 39984
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_172
timestamp 1486834041
transform 1 0 19936 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_174
timestamp 1486834041
transform 1 0 20160 0 1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_177
timestamp 1486834041
transform 1 0 20496 0 1 39984
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_209
timestamp 1486834041
transform 1 0 24080 0 1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_2
timestamp 1486834041
transform 1 0 896 0 -1 41552
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_66
timestamp 1486834041
transform 1 0 8064 0 -1 41552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_92
timestamp 1486834041
transform 1 0 10976 0 -1 41552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_96
timestamp 1486834041
transform 1 0 11424 0 -1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_105
timestamp 1486834041
transform 1 0 12432 0 -1 41552
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_113
timestamp 1486834041
transform 1 0 13328 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_135
timestamp 1486834041
transform 1 0 15792 0 -1 41552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_139
timestamp 1486834041
transform 1 0 16240 0 -1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_142
timestamp 1486834041
transform 1 0 16576 0 -1 41552
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_206
timestamp 1486834041
transform 1 0 23744 0 -1 41552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_212
timestamp 1486834041
transform 1 0 24416 0 -1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_52_2
timestamp 1486834041
transform 1 0 896 0 1 41552
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_34
timestamp 1486834041
transform 1 0 4480 0 1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_37
timestamp 1486834041
transform 1 0 4816 0 1 41552
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_101
timestamp 1486834041
transform 1 0 11984 0 1 41552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_107
timestamp 1486834041
transform 1 0 12656 0 1 41552
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_115
timestamp 1486834041
transform 1 0 13552 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_117
timestamp 1486834041
transform 1 0 13776 0 1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_52_138
timestamp 1486834041
transform 1 0 16128 0 1 41552
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_170
timestamp 1486834041
transform 1 0 19712 0 1 41552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_174
timestamp 1486834041
transform 1 0 20160 0 1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_52_177
timestamp 1486834041
transform 1 0 20496 0 1 41552
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_209
timestamp 1486834041
transform 1 0 24080 0 1 41552
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_225
timestamp 1486834041
transform 1 0 25872 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_2
timestamp 1486834041
transform 1 0 896 0 -1 43120
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_66
timestamp 1486834041
transform 1 0 8064 0 -1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_72
timestamp 1486834041
transform 1 0 8736 0 -1 43120
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_136
timestamp 1486834041
transform 1 0 15904 0 -1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_142
timestamp 1486834041
transform 1 0 16576 0 -1 43120
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_206
timestamp 1486834041
transform 1 0 23744 0 -1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_212
timestamp 1486834041
transform 1 0 24416 0 -1 43120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_2
timestamp 1486834041
transform 1 0 896 0 1 43120
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_34
timestamp 1486834041
transform 1 0 4480 0 1 43120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_37
timestamp 1486834041
transform 1 0 4816 0 1 43120
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_101
timestamp 1486834041
transform 1 0 11984 0 1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_107
timestamp 1486834041
transform 1 0 12656 0 1 43120
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_171
timestamp 1486834041
transform 1 0 19824 0 1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_177
timestamp 1486834041
transform 1 0 20496 0 1 43120
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_209
timestamp 1486834041
transform 1 0 24080 0 1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_2
timestamp 1486834041
transform 1 0 896 0 -1 44688
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_66
timestamp 1486834041
transform 1 0 8064 0 -1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_72
timestamp 1486834041
transform 1 0 8736 0 -1 44688
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_136
timestamp 1486834041
transform 1 0 15904 0 -1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_142
timestamp 1486834041
transform 1 0 16576 0 -1 44688
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_206
timestamp 1486834041
transform 1 0 23744 0 -1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_212
timestamp 1486834041
transform 1 0 24416 0 -1 44688
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_56_2
timestamp 1486834041
transform 1 0 896 0 1 44688
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_34
timestamp 1486834041
transform 1 0 4480 0 1 44688
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_37
timestamp 1486834041
transform 1 0 4816 0 1 44688
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_101
timestamp 1486834041
transform 1 0 11984 0 1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_107
timestamp 1486834041
transform 1 0 12656 0 1 44688
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_171
timestamp 1486834041
transform 1 0 19824 0 1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_56_177
timestamp 1486834041
transform 1 0 20496 0 1 44688
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_56_209
timestamp 1486834041
transform 1 0 24080 0 1 44688
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_225
timestamp 1486834041
transform 1 0 25872 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_2
timestamp 1486834041
transform 1 0 896 0 -1 46256
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_66
timestamp 1486834041
transform 1 0 8064 0 -1 46256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_72
timestamp 1486834041
transform 1 0 8736 0 -1 46256
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_136
timestamp 1486834041
transform 1 0 15904 0 -1 46256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_142
timestamp 1486834041
transform 1 0 16576 0 -1 46256
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_206
timestamp 1486834041
transform 1 0 23744 0 -1 46256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_212
timestamp 1486834041
transform 1 0 24416 0 -1 46256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_58_2
timestamp 1486834041
transform 1 0 896 0 1 46256
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_34
timestamp 1486834041
transform 1 0 4480 0 1 46256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_37
timestamp 1486834041
transform 1 0 4816 0 1 46256
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_101
timestamp 1486834041
transform 1 0 11984 0 1 46256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_107
timestamp 1486834041
transform 1 0 12656 0 1 46256
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_171
timestamp 1486834041
transform 1 0 19824 0 1 46256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_58_177
timestamp 1486834041
transform 1 0 20496 0 1 46256
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_209
timestamp 1486834041
transform 1 0 24080 0 1 46256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_2
timestamp 1486834041
transform 1 0 896 0 -1 47824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_66
timestamp 1486834041
transform 1 0 8064 0 -1 47824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_72
timestamp 1486834041
transform 1 0 8736 0 -1 47824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_136
timestamp 1486834041
transform 1 0 15904 0 -1 47824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_142
timestamp 1486834041
transform 1 0 16576 0 -1 47824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_206
timestamp 1486834041
transform 1 0 23744 0 -1 47824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_212
timestamp 1486834041
transform 1 0 24416 0 -1 47824
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_2
timestamp 1486834041
transform 1 0 896 0 1 47824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_34
timestamp 1486834041
transform 1 0 4480 0 1 47824
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_37
timestamp 1486834041
transform 1 0 4816 0 1 47824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_101
timestamp 1486834041
transform 1 0 11984 0 1 47824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_107
timestamp 1486834041
transform 1 0 12656 0 1 47824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_171
timestamp 1486834041
transform 1 0 19824 0 1 47824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_177
timestamp 1486834041
transform 1 0 20496 0 1 47824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_60_209
timestamp 1486834041
transform 1 0 24080 0 1 47824
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_225
timestamp 1486834041
transform 1 0 25872 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_2
timestamp 1486834041
transform 1 0 896 0 -1 49392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_66
timestamp 1486834041
transform 1 0 8064 0 -1 49392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_72
timestamp 1486834041
transform 1 0 8736 0 -1 49392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_136
timestamp 1486834041
transform 1 0 15904 0 -1 49392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_142
timestamp 1486834041
transform 1 0 16576 0 -1 49392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_206
timestamp 1486834041
transform 1 0 23744 0 -1 49392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_212
timestamp 1486834041
transform 1 0 24416 0 -1 49392
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_62_2
timestamp 1486834041
transform 1 0 896 0 1 49392
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_34
timestamp 1486834041
transform 1 0 4480 0 1 49392
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_37
timestamp 1486834041
transform 1 0 4816 0 1 49392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_101
timestamp 1486834041
transform 1 0 11984 0 1 49392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_107
timestamp 1486834041
transform 1 0 12656 0 1 49392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_171
timestamp 1486834041
transform 1 0 19824 0 1 49392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_62_177
timestamp 1486834041
transform 1 0 20496 0 1 49392
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_209
timestamp 1486834041
transform 1 0 24080 0 1 49392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_2
timestamp 1486834041
transform 1 0 896 0 -1 50960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_66
timestamp 1486834041
transform 1 0 8064 0 -1 50960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_72
timestamp 1486834041
transform 1 0 8736 0 -1 50960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_136
timestamp 1486834041
transform 1 0 15904 0 -1 50960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_63_142
timestamp 1486834041
transform 1 0 16576 0 -1 50960
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_63_174
timestamp 1486834041
transform 1 0 20160 0 -1 50960
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_190
timestamp 1486834041
transform 1 0 21952 0 -1 50960
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_198
timestamp 1486834041
transform 1 0 22848 0 -1 50960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_212
timestamp 1486834041
transform 1 0 24416 0 -1 50960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_64_2
timestamp 1486834041
transform 1 0 896 0 1 50960
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_34
timestamp 1486834041
transform 1 0 4480 0 1 50960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_37
timestamp 1486834041
transform 1 0 4816 0 1 50960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_101
timestamp 1486834041
transform 1 0 11984 0 1 50960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_107
timestamp 1486834041
transform 1 0 12656 0 1 50960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_171
timestamp 1486834041
transform 1 0 19824 0 1 50960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_64_177
timestamp 1486834041
transform 1 0 20496 0 1 50960
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_209
timestamp 1486834041
transform 1 0 24080 0 1 50960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_2
timestamp 1486834041
transform 1 0 896 0 -1 52528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_66
timestamp 1486834041
transform 1 0 8064 0 -1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_72
timestamp 1486834041
transform 1 0 8736 0 -1 52528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_136
timestamp 1486834041
transform 1 0 15904 0 -1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_65_142
timestamp 1486834041
transform 1 0 16576 0 -1 52528
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_174
timestamp 1486834041
transform 1 0 20160 0 -1 52528
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_182
timestamp 1486834041
transform 1 0 21056 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_192
timestamp 1486834041
transform 1 0 22176 0 -1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_212
timestamp 1486834041
transform 1 0 24416 0 -1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_66_2
timestamp 1486834041
transform 1 0 896 0 1 52528
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_34
timestamp 1486834041
transform 1 0 4480 0 1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_37
timestamp 1486834041
transform 1 0 4816 0 1 52528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_101
timestamp 1486834041
transform 1 0 11984 0 1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_107
timestamp 1486834041
transform 1 0 12656 0 1 52528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_171
timestamp 1486834041
transform 1 0 19824 0 1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_177
timestamp 1486834041
transform 1 0 20496 0 1 52528
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_193
timestamp 1486834041
transform 1 0 22288 0 1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_197
timestamp 1486834041
transform 1 0 22736 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_2
timestamp 1486834041
transform 1 0 896 0 -1 54096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_66
timestamp 1486834041
transform 1 0 8064 0 -1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_72
timestamp 1486834041
transform 1 0 8736 0 -1 54096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_136
timestamp 1486834041
transform 1 0 15904 0 -1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_142
timestamp 1486834041
transform 1 0 16576 0 -1 54096
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_174
timestamp 1486834041
transform 1 0 20160 0 -1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_182
timestamp 1486834041
transform 1 0 21056 0 -1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_186
timestamp 1486834041
transform 1 0 21504 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_212
timestamp 1486834041
transform 1 0 24416 0 -1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_68_2
timestamp 1486834041
transform 1 0 896 0 1 54096
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_34
timestamp 1486834041
transform 1 0 4480 0 1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_37
timestamp 1486834041
transform 1 0 4816 0 1 54096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_101
timestamp 1486834041
transform 1 0 11984 0 1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_68_107
timestamp 1486834041
transform 1 0 12656 0 1 54096
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_68_139
timestamp 1486834041
transform 1 0 16240 0 1 54096
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_68_155
timestamp 1486834041
transform 1 0 18032 0 1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_171
timestamp 1486834041
transform 1 0 19824 0 1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_69_2
timestamp 1486834041
transform 1 0 896 0 -1 55664
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_10
timestamp 1486834041
transform 1 0 1792 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_12
timestamp 1486834041
transform 1 0 2016 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_69_27
timestamp 1486834041
transform 1 0 3696 0 -1 55664
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_43
timestamp 1486834041
transform 1 0 5488 0 -1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_47
timestamp 1486834041
transform 1 0 5936 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_63
timestamp 1486834041
transform 1 0 7728 0 -1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_67
timestamp 1486834041
transform 1 0 8176 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_69
timestamp 1486834041
transform 1 0 8400 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_69_72
timestamp 1486834041
transform 1 0 8736 0 -1 55664
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_69_88
timestamp 1486834041
transform 1 0 10528 0 -1 55664
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_96
timestamp 1486834041
transform 1 0 11424 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_69_111
timestamp 1486834041
transform 1 0 13104 0 -1 55664
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_69_127
timestamp 1486834041
transform 1 0 14896 0 -1 55664
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_135
timestamp 1486834041
transform 1 0 15792 0 -1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_139
timestamp 1486834041
transform 1 0 16240 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_142
timestamp 1486834041
transform 1 0 16576 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_144
timestamp 1486834041
transform 1 0 16800 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_69_159
timestamp 1486834041
transform 1 0 18480 0 -1 55664
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_167
timestamp 1486834041
transform 1 0 19376 0 -1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_207
timestamp 1486834041
transform 1 0 23856 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_209
timestamp 1486834041
transform 1 0 24080 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_212
timestamp 1486834041
transform 1 0 24416 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_70_8
timestamp 1486834041
transform 1 0 1568 0 1 55664
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_16
timestamp 1486834041
transform 1 0 2464 0 1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_36
timestamp 1486834041
transform 1 0 4704 0 1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_51
timestamp 1486834041
transform 1 0 6384 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_53
timestamp 1486834041
transform 1 0 6608 0 1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_70
timestamp 1486834041
transform 1 0 8512 0 1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_99
timestamp 1486834041
transform 1 0 11760 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_101
timestamp 1486834041
transform 1 0 11984 0 1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_104
timestamp 1486834041
transform 1 0 12320 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_106
timestamp 1486834041
transform 1 0 12544 0 1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_135
timestamp 1486834041
transform 1 0 15792 0 1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_152
timestamp 1486834041
transform 1 0 17696 0 1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_200
timestamp 1486834041
transform 1 0 23072 0 1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_234
timestamp 1486834041
transform 1 0 26880 0 1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_240
timestamp 1486834041
transform 1 0 27552 0 1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output1
timestamp 1486834041
transform -1 0 2464 0 -1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output2
timestamp 1486834041
transform -1 0 2464 0 1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output3
timestamp 1486834041
transform -1 0 4032 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output4
timestamp 1486834041
transform -1 0 2464 0 1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output5
timestamp 1486834041
transform -1 0 7616 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output6
timestamp 1486834041
transform -1 0 4032 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output7
timestamp 1486834041
transform -1 0 4032 0 -1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output8
timestamp 1486834041
transform -1 0 2464 0 -1 5488
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output9
timestamp 1486834041
transform -1 0 6384 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output10
timestamp 1486834041
transform -1 0 2464 0 -1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output11
timestamp 1486834041
transform -1 0 2464 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output12
timestamp 1486834041
transform -1 0 2464 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output13
timestamp 1486834041
transform -1 0 2464 0 1 5488
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output14
timestamp 1486834041
transform -1 0 4032 0 1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output15
timestamp 1486834041
transform 1 0 4816 0 1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output16
timestamp 1486834041
transform 1 0 4816 0 1 16464
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output17
timestamp 1486834041
transform -1 0 2464 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output18
timestamp 1486834041
transform 1 0 4816 0 1 19600
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output19
timestamp 1486834041
transform -1 0 4032 0 -1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output20
timestamp 1486834041
transform -1 0 2464 0 -1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output21
timestamp 1486834041
transform -1 0 2464 0 -1 19600
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output22
timestamp 1486834041
transform -1 0 4704 0 -1 22736
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output23
timestamp 1486834041
transform 1 0 4816 0 1 24304
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output24
timestamp 1486834041
transform -1 0 2464 0 -1 25872
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output25
timestamp 1486834041
transform 1 0 24528 0 -1 22736
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output26
timestamp 1486834041
transform 1 0 26096 0 1 21168
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output27
timestamp 1486834041
transform 1 0 26096 0 -1 22736
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output28
timestamp 1486834041
transform 1 0 24528 0 -1 24304
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output29
timestamp 1486834041
transform 1 0 26096 0 1 22736
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output30
timestamp 1486834041
transform 1 0 24528 0 1 24304
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output31
timestamp 1486834041
transform 1 0 26096 0 -1 24304
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output32
timestamp 1486834041
transform 1 0 24528 0 -1 25872
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output33
timestamp 1486834041
transform 1 0 26096 0 1 24304
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output34
timestamp 1486834041
transform 1 0 26096 0 -1 25872
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output35
timestamp 1486834041
transform 1 0 24528 0 -1 27440
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output36
timestamp 1486834041
transform 1 0 26096 0 1 25872
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output37
timestamp 1486834041
transform 1 0 24528 0 1 27440
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output38
timestamp 1486834041
transform 1 0 26096 0 -1 27440
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output39
timestamp 1486834041
transform 1 0 26096 0 1 27440
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output40
timestamp 1486834041
transform 1 0 26096 0 -1 29008
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output41
timestamp 1486834041
transform 1 0 26096 0 1 29008
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output42
timestamp 1486834041
transform 1 0 26096 0 -1 30576
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output43
timestamp 1486834041
transform 1 0 26096 0 1 30576
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output44
timestamp 1486834041
transform 1 0 26096 0 -1 32144
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output45
timestamp 1486834041
transform 1 0 24528 0 -1 38416
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output46
timestamp 1486834041
transform 1 0 24528 0 -1 43120
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output47
timestamp 1486834041
transform 1 0 26096 0 -1 44688
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output48
timestamp 1486834041
transform 1 0 26096 0 -1 39984
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output49
timestamp 1486834041
transform 1 0 26096 0 1 39984
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output50
timestamp 1486834041
transform 1 0 24528 0 -1 39984
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output51
timestamp 1486834041
transform 1 0 26096 0 -1 41552
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output52
timestamp 1486834041
transform 1 0 24528 0 1 39984
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output53
timestamp 1486834041
transform 1 0 26096 0 1 41552
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output54
timestamp 1486834041
transform 1 0 24528 0 -1 41552
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output55
timestamp 1486834041
transform 1 0 26096 0 -1 43120
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output56
timestamp 1486834041
transform 1 0 26096 0 1 43120
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output57
timestamp 1486834041
transform 1 0 24528 0 1 30576
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output58
timestamp 1486834041
transform 1 0 26096 0 -1 36848
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output59
timestamp 1486834041
transform 1 0 26096 0 1 36848
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output60
timestamp 1486834041
transform 1 0 24528 0 -1 36848
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output61
timestamp 1486834041
transform 1 0 26096 0 -1 38416
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output62
timestamp 1486834041
transform 1 0 24528 0 1 36848
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output63
timestamp 1486834041
transform 1 0 26096 0 1 38416
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output64
timestamp 1486834041
transform 1 0 26096 0 1 32144
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output65
timestamp 1486834041
transform 1 0 24528 0 -1 32144
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output66
timestamp 1486834041
transform 1 0 26096 0 -1 33712
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output67
timestamp 1486834041
transform 1 0 26096 0 1 33712
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output68
timestamp 1486834041
transform 1 0 24528 0 -1 33712
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output69
timestamp 1486834041
transform 1 0 26096 0 -1 35280
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output70
timestamp 1486834041
transform 1 0 24528 0 1 33712
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output71
timestamp 1486834041
transform 1 0 26096 0 1 35280
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output72
timestamp 1486834041
transform 1 0 24528 0 -1 35280
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output73
timestamp 1486834041
transform 1 0 24528 0 1 43120
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output74
timestamp 1486834041
transform 1 0 26096 0 -1 49392
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output75
timestamp 1486834041
transform 1 0 26096 0 1 49392
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output76
timestamp 1486834041
transform 1 0 24528 0 -1 49392
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output77
timestamp 1486834041
transform 1 0 26096 0 -1 50960
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output78
timestamp 1486834041
transform 1 0 24528 0 1 49392
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output79
timestamp 1486834041
transform 1 0 26096 0 1 50960
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output80
timestamp 1486834041
transform 1 0 24528 0 -1 50960
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output81
timestamp 1486834041
transform 1 0 26096 0 -1 52528
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output82
timestamp 1486834041
transform 1 0 26096 0 1 52528
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output83
timestamp 1486834041
transform 1 0 24528 0 -1 52528
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output84
timestamp 1486834041
transform 1 0 26096 0 1 44688
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output85
timestamp 1486834041
transform 1 0 26096 0 -1 54096
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output86
timestamp 1486834041
transform 1 0 24528 0 1 52528
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output87
timestamp 1486834041
transform 1 0 26096 0 1 54096
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output88
timestamp 1486834041
transform 1 0 24528 0 -1 54096
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output89
timestamp 1486834041
transform 1 0 26096 0 -1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output90
timestamp 1486834041
transform 1 0 24528 0 -1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output91
timestamp 1486834041
transform -1 0 24528 0 1 54096
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output92
timestamp 1486834041
transform 1 0 22624 0 -1 54096
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output93
timestamp 1486834041
transform 1 0 21392 0 1 54096
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output94
timestamp 1486834041
transform 1 0 24528 0 1 50960
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output95
timestamp 1486834041
transform 1 0 24528 0 -1 44688
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output96
timestamp 1486834041
transform 1 0 22960 0 1 52528
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output97
timestamp 1486834041
transform 1 0 22624 0 -1 52528
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output98
timestamp 1486834041
transform 1 0 26096 0 -1 46256
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output99
timestamp 1486834041
transform 1 0 26096 0 1 46256
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output100
timestamp 1486834041
transform 1 0 24528 0 -1 46256
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output101
timestamp 1486834041
transform 1 0 26096 0 -1 47824
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output102
timestamp 1486834041
transform 1 0 24528 0 1 46256
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output103
timestamp 1486834041
transform 1 0 26096 0 1 47824
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output104
timestamp 1486834041
transform 1 0 24528 0 -1 47824
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output105
timestamp 1486834041
transform -1 0 3696 0 -1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output106
timestamp 1486834041
transform -1 0 17696 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output107
timestamp 1486834041
transform -1 0 18480 0 -1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output108
timestamp 1486834041
transform -1 0 19712 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output109
timestamp 1486834041
transform -1 0 21504 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output110
timestamp 1486834041
transform 1 0 21504 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output111
timestamp 1486834041
transform 1 0 22288 0 -1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output112
timestamp 1486834041
transform 1 0 23744 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output113
timestamp 1486834041
transform 1 0 25312 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output114
timestamp 1486834041
transform 1 0 24528 0 1 54096
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output115
timestamp 1486834041
transform 1 0 20720 0 -1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output116
timestamp 1486834041
transform 1 0 2912 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output117
timestamp 1486834041
transform -1 0 6384 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output118
timestamp 1486834041
transform 1 0 6160 0 -1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output119
timestamp 1486834041
transform -1 0 8288 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output120
timestamp 1486834041
transform -1 0 10192 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output121
timestamp 1486834041
transform -1 0 11760 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output122
timestamp 1486834041
transform -1 0 13104 0 -1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output123
timestamp 1486834041
transform -1 0 14224 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output124
timestamp 1486834041
transform -1 0 15792 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output125
timestamp 1486834041
transform -1 0 1568 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_71
timestamp 1486834041
transform 1 0 672 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1486834041
transform -1 0 27888 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_72
timestamp 1486834041
transform 1 0 672 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1486834041
transform -1 0 27888 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_73
timestamp 1486834041
transform 1 0 672 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1486834041
transform -1 0 27888 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_74
timestamp 1486834041
transform 1 0 672 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1486834041
transform -1 0 27888 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_75
timestamp 1486834041
transform 1 0 672 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1486834041
transform -1 0 27888 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_76
timestamp 1486834041
transform 1 0 672 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1486834041
transform -1 0 27888 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_77
timestamp 1486834041
transform 1 0 672 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1486834041
transform -1 0 27888 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_78
timestamp 1486834041
transform 1 0 672 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1486834041
transform -1 0 27888 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_79
timestamp 1486834041
transform 1 0 672 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1486834041
transform -1 0 27888 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_80
timestamp 1486834041
transform 1 0 672 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1486834041
transform -1 0 27888 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_81
timestamp 1486834041
transform 1 0 672 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1486834041
transform -1 0 27888 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_82
timestamp 1486834041
transform 1 0 672 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1486834041
transform -1 0 27888 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_83
timestamp 1486834041
transform 1 0 672 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1486834041
transform -1 0 27888 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_84
timestamp 1486834041
transform 1 0 672 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1486834041
transform -1 0 27888 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_85
timestamp 1486834041
transform 1 0 672 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1486834041
transform -1 0 27888 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_86
timestamp 1486834041
transform 1 0 672 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1486834041
transform -1 0 27888 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_87
timestamp 1486834041
transform 1 0 672 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1486834041
transform -1 0 27888 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_88
timestamp 1486834041
transform 1 0 672 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1486834041
transform -1 0 27888 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_89
timestamp 1486834041
transform 1 0 672 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1486834041
transform -1 0 27888 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_90
timestamp 1486834041
transform 1 0 672 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1486834041
transform -1 0 27888 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_91
timestamp 1486834041
transform 1 0 672 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1486834041
transform -1 0 27888 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_92
timestamp 1486834041
transform 1 0 672 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1486834041
transform -1 0 27888 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_93
timestamp 1486834041
transform 1 0 672 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1486834041
transform -1 0 27888 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_94
timestamp 1486834041
transform 1 0 672 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1486834041
transform -1 0 27888 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_95
timestamp 1486834041
transform 1 0 672 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1486834041
transform -1 0 27888 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_96
timestamp 1486834041
transform 1 0 672 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1486834041
transform -1 0 27888 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_97
timestamp 1486834041
transform 1 0 672 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1486834041
transform -1 0 27888 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_98
timestamp 1486834041
transform 1 0 672 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1486834041
transform -1 0 27888 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_99
timestamp 1486834041
transform 1 0 672 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1486834041
transform -1 0 27888 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_100
timestamp 1486834041
transform 1 0 672 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1486834041
transform -1 0 27888 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_101
timestamp 1486834041
transform 1 0 672 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1486834041
transform -1 0 27888 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_102
timestamp 1486834041
transform 1 0 672 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1486834041
transform -1 0 27888 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_103
timestamp 1486834041
transform 1 0 672 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1486834041
transform -1 0 27888 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_104
timestamp 1486834041
transform 1 0 672 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1486834041
transform -1 0 27888 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_105
timestamp 1486834041
transform 1 0 672 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1486834041
transform -1 0 27888 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_106
timestamp 1486834041
transform 1 0 672 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1486834041
transform -1 0 27888 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_107
timestamp 1486834041
transform 1 0 672 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1486834041
transform -1 0 27888 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_108
timestamp 1486834041
transform 1 0 672 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1486834041
transform -1 0 27888 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_109
timestamp 1486834041
transform 1 0 672 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1486834041
transform -1 0 27888 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_110
timestamp 1486834041
transform 1 0 672 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1486834041
transform -1 0 27888 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_111
timestamp 1486834041
transform 1 0 672 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1486834041
transform -1 0 27888 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_112
timestamp 1486834041
transform 1 0 672 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1486834041
transform -1 0 27888 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_113
timestamp 1486834041
transform 1 0 672 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1486834041
transform -1 0 27888 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_114
timestamp 1486834041
transform 1 0 672 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1486834041
transform -1 0 27888 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_115
timestamp 1486834041
transform 1 0 672 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1486834041
transform -1 0 27888 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_116
timestamp 1486834041
transform 1 0 672 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1486834041
transform -1 0 27888 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_117
timestamp 1486834041
transform 1 0 672 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1486834041
transform -1 0 27888 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_118
timestamp 1486834041
transform 1 0 672 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1486834041
transform -1 0 27888 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_119
timestamp 1486834041
transform 1 0 672 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1486834041
transform -1 0 27888 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_120
timestamp 1486834041
transform 1 0 672 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1486834041
transform -1 0 27888 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_121
timestamp 1486834041
transform 1 0 672 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1486834041
transform -1 0 27888 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_122
timestamp 1486834041
transform 1 0 672 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1486834041
transform -1 0 27888 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_123
timestamp 1486834041
transform 1 0 672 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1486834041
transform -1 0 27888 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_124
timestamp 1486834041
transform 1 0 672 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1486834041
transform -1 0 27888 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_125
timestamp 1486834041
transform 1 0 672 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1486834041
transform -1 0 27888 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_126
timestamp 1486834041
transform 1 0 672 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1486834041
transform -1 0 27888 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_127
timestamp 1486834041
transform 1 0 672 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1486834041
transform -1 0 27888 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_128
timestamp 1486834041
transform 1 0 672 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1486834041
transform -1 0 27888 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_129
timestamp 1486834041
transform 1 0 672 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1486834041
transform -1 0 27888 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_130
timestamp 1486834041
transform 1 0 672 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1486834041
transform -1 0 27888 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_131
timestamp 1486834041
transform 1 0 672 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1486834041
transform -1 0 27888 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_132
timestamp 1486834041
transform 1 0 672 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1486834041
transform -1 0 27888 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Left_133
timestamp 1486834041
transform 1 0 672 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Right_62
timestamp 1486834041
transform -1 0 27888 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Left_134
timestamp 1486834041
transform 1 0 672 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Right_63
timestamp 1486834041
transform -1 0 27888 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Left_135
timestamp 1486834041
transform 1 0 672 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Right_64
timestamp 1486834041
transform -1 0 27888 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Left_136
timestamp 1486834041
transform 1 0 672 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Right_65
timestamp 1486834041
transform -1 0 27888 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Left_137
timestamp 1486834041
transform 1 0 672 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Right_66
timestamp 1486834041
transform -1 0 27888 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Left_138
timestamp 1486834041
transform 1 0 672 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Right_67
timestamp 1486834041
transform -1 0 27888 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Left_139
timestamp 1486834041
transform 1 0 672 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Right_68
timestamp 1486834041
transform -1 0 27888 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Left_140
timestamp 1486834041
transform 1 0 672 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Right_69
timestamp 1486834041
transform -1 0 27888 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Left_141
timestamp 1486834041
transform 1 0 672 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Right_70
timestamp 1486834041
transform -1 0 27888 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_142
timestamp 1486834041
transform 1 0 4480 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_143
timestamp 1486834041
transform 1 0 8288 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_144
timestamp 1486834041
transform 1 0 12096 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_145
timestamp 1486834041
transform 1 0 15904 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_146
timestamp 1486834041
transform 1 0 19712 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_147
timestamp 1486834041
transform 1 0 23520 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_148
timestamp 1486834041
transform 1 0 27328 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_149
timestamp 1486834041
transform 1 0 8512 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_150
timestamp 1486834041
transform 1 0 16352 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_151
timestamp 1486834041
transform 1 0 24192 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_152
timestamp 1486834041
transform 1 0 4592 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_153
timestamp 1486834041
transform 1 0 12432 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_154
timestamp 1486834041
transform 1 0 20272 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_155
timestamp 1486834041
transform 1 0 8512 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_156
timestamp 1486834041
transform 1 0 16352 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_157
timestamp 1486834041
transform 1 0 24192 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_158
timestamp 1486834041
transform 1 0 4592 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_159
timestamp 1486834041
transform 1 0 12432 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_160
timestamp 1486834041
transform 1 0 20272 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_161
timestamp 1486834041
transform 1 0 8512 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_162
timestamp 1486834041
transform 1 0 16352 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_163
timestamp 1486834041
transform 1 0 24192 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_164
timestamp 1486834041
transform 1 0 4592 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_165
timestamp 1486834041
transform 1 0 12432 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_166
timestamp 1486834041
transform 1 0 20272 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_167
timestamp 1486834041
transform 1 0 8512 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_168
timestamp 1486834041
transform 1 0 16352 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_169
timestamp 1486834041
transform 1 0 24192 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_170
timestamp 1486834041
transform 1 0 4592 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_171
timestamp 1486834041
transform 1 0 12432 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_172
timestamp 1486834041
transform 1 0 20272 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_173
timestamp 1486834041
transform 1 0 8512 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_174
timestamp 1486834041
transform 1 0 16352 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_175
timestamp 1486834041
transform 1 0 24192 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_176
timestamp 1486834041
transform 1 0 4592 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_177
timestamp 1486834041
transform 1 0 12432 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_178
timestamp 1486834041
transform 1 0 20272 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_179
timestamp 1486834041
transform 1 0 8512 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_180
timestamp 1486834041
transform 1 0 16352 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_181
timestamp 1486834041
transform 1 0 24192 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_182
timestamp 1486834041
transform 1 0 4592 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_183
timestamp 1486834041
transform 1 0 12432 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_184
timestamp 1486834041
transform 1 0 20272 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_185
timestamp 1486834041
transform 1 0 8512 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_186
timestamp 1486834041
transform 1 0 16352 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_187
timestamp 1486834041
transform 1 0 24192 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_188
timestamp 1486834041
transform 1 0 4592 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_189
timestamp 1486834041
transform 1 0 12432 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_190
timestamp 1486834041
transform 1 0 20272 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_191
timestamp 1486834041
transform 1 0 8512 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_192
timestamp 1486834041
transform 1 0 16352 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_193
timestamp 1486834041
transform 1 0 24192 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_194
timestamp 1486834041
transform 1 0 4592 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_195
timestamp 1486834041
transform 1 0 12432 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_196
timestamp 1486834041
transform 1 0 20272 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_197
timestamp 1486834041
transform 1 0 8512 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_198
timestamp 1486834041
transform 1 0 16352 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_199
timestamp 1486834041
transform 1 0 24192 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_200
timestamp 1486834041
transform 1 0 4592 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_201
timestamp 1486834041
transform 1 0 12432 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_202
timestamp 1486834041
transform 1 0 20272 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_203
timestamp 1486834041
transform 1 0 8512 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_204
timestamp 1486834041
transform 1 0 16352 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_205
timestamp 1486834041
transform 1 0 24192 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_206
timestamp 1486834041
transform 1 0 4592 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_207
timestamp 1486834041
transform 1 0 12432 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_208
timestamp 1486834041
transform 1 0 20272 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_209
timestamp 1486834041
transform 1 0 8512 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_210
timestamp 1486834041
transform 1 0 16352 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_211
timestamp 1486834041
transform 1 0 24192 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_212
timestamp 1486834041
transform 1 0 4592 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_213
timestamp 1486834041
transform 1 0 12432 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_214
timestamp 1486834041
transform 1 0 20272 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_215
timestamp 1486834041
transform 1 0 8512 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_216
timestamp 1486834041
transform 1 0 16352 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_217
timestamp 1486834041
transform 1 0 24192 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_218
timestamp 1486834041
transform 1 0 4592 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_219
timestamp 1486834041
transform 1 0 12432 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_220
timestamp 1486834041
transform 1 0 20272 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_221
timestamp 1486834041
transform 1 0 8512 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_222
timestamp 1486834041
transform 1 0 16352 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_223
timestamp 1486834041
transform 1 0 24192 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_224
timestamp 1486834041
transform 1 0 4592 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_225
timestamp 1486834041
transform 1 0 12432 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_226
timestamp 1486834041
transform 1 0 20272 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_227
timestamp 1486834041
transform 1 0 8512 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_228
timestamp 1486834041
transform 1 0 16352 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_229
timestamp 1486834041
transform 1 0 24192 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_230
timestamp 1486834041
transform 1 0 4592 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_231
timestamp 1486834041
transform 1 0 12432 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_232
timestamp 1486834041
transform 1 0 20272 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_233
timestamp 1486834041
transform 1 0 8512 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_234
timestamp 1486834041
transform 1 0 16352 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_235
timestamp 1486834041
transform 1 0 24192 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_236
timestamp 1486834041
transform 1 0 4592 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_237
timestamp 1486834041
transform 1 0 12432 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_238
timestamp 1486834041
transform 1 0 20272 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_239
timestamp 1486834041
transform 1 0 8512 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_240
timestamp 1486834041
transform 1 0 16352 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_241
timestamp 1486834041
transform 1 0 24192 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1486834041
transform 1 0 4592 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1486834041
transform 1 0 12432 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_244
timestamp 1486834041
transform 1 0 20272 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1486834041
transform 1 0 8512 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1486834041
transform 1 0 16352 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1486834041
transform 1 0 24192 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1486834041
transform 1 0 4592 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1486834041
transform 1 0 12432 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1486834041
transform 1 0 20272 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_251
timestamp 1486834041
transform 1 0 8512 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_252
timestamp 1486834041
transform 1 0 16352 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1486834041
transform 1 0 24192 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_254
timestamp 1486834041
transform 1 0 4592 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_255
timestamp 1486834041
transform 1 0 12432 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_256
timestamp 1486834041
transform 1 0 20272 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_257
timestamp 1486834041
transform 1 0 8512 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_258
timestamp 1486834041
transform 1 0 16352 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_259
timestamp 1486834041
transform 1 0 24192 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_260
timestamp 1486834041
transform 1 0 4592 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_261
timestamp 1486834041
transform 1 0 12432 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_262
timestamp 1486834041
transform 1 0 20272 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_263
timestamp 1486834041
transform 1 0 8512 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_264
timestamp 1486834041
transform 1 0 16352 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_265
timestamp 1486834041
transform 1 0 24192 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_266
timestamp 1486834041
transform 1 0 4592 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_267
timestamp 1486834041
transform 1 0 12432 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_268
timestamp 1486834041
transform 1 0 20272 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_269
timestamp 1486834041
transform 1 0 8512 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_270
timestamp 1486834041
transform 1 0 16352 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_271
timestamp 1486834041
transform 1 0 24192 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_272
timestamp 1486834041
transform 1 0 4592 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_273
timestamp 1486834041
transform 1 0 12432 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_274
timestamp 1486834041
transform 1 0 20272 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_275
timestamp 1486834041
transform 1 0 8512 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_276
timestamp 1486834041
transform 1 0 16352 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_277
timestamp 1486834041
transform 1 0 24192 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_278
timestamp 1486834041
transform 1 0 4592 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_279
timestamp 1486834041
transform 1 0 12432 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_280
timestamp 1486834041
transform 1 0 20272 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_281
timestamp 1486834041
transform 1 0 8512 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_282
timestamp 1486834041
transform 1 0 16352 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_283
timestamp 1486834041
transform 1 0 24192 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_284
timestamp 1486834041
transform 1 0 4592 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_285
timestamp 1486834041
transform 1 0 12432 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_286
timestamp 1486834041
transform 1 0 20272 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_287
timestamp 1486834041
transform 1 0 8512 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_288
timestamp 1486834041
transform 1 0 16352 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_289
timestamp 1486834041
transform 1 0 24192 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_290
timestamp 1486834041
transform 1 0 4592 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_291
timestamp 1486834041
transform 1 0 12432 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_292
timestamp 1486834041
transform 1 0 20272 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_293
timestamp 1486834041
transform 1 0 8512 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_294
timestamp 1486834041
transform 1 0 16352 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_295
timestamp 1486834041
transform 1 0 24192 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_296
timestamp 1486834041
transform 1 0 4592 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_297
timestamp 1486834041
transform 1 0 12432 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_298
timestamp 1486834041
transform 1 0 20272 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_299
timestamp 1486834041
transform 1 0 8512 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_300
timestamp 1486834041
transform 1 0 16352 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_301
timestamp 1486834041
transform 1 0 24192 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_302
timestamp 1486834041
transform 1 0 4592 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_303
timestamp 1486834041
transform 1 0 12432 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_304
timestamp 1486834041
transform 1 0 20272 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_305
timestamp 1486834041
transform 1 0 8512 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_306
timestamp 1486834041
transform 1 0 16352 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_307
timestamp 1486834041
transform 1 0 24192 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_308
timestamp 1486834041
transform 1 0 4592 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_309
timestamp 1486834041
transform 1 0 12432 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_310
timestamp 1486834041
transform 1 0 20272 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_311
timestamp 1486834041
transform 1 0 8512 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_312
timestamp 1486834041
transform 1 0 16352 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_313
timestamp 1486834041
transform 1 0 24192 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_314
timestamp 1486834041
transform 1 0 4592 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_315
timestamp 1486834041
transform 1 0 12432 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_316
timestamp 1486834041
transform 1 0 20272 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_317
timestamp 1486834041
transform 1 0 8512 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_318
timestamp 1486834041
transform 1 0 16352 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_319
timestamp 1486834041
transform 1 0 24192 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_320
timestamp 1486834041
transform 1 0 4592 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_321
timestamp 1486834041
transform 1 0 12432 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_322
timestamp 1486834041
transform 1 0 20272 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_323
timestamp 1486834041
transform 1 0 8512 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_324
timestamp 1486834041
transform 1 0 16352 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_325
timestamp 1486834041
transform 1 0 24192 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_326
timestamp 1486834041
transform 1 0 4592 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_327
timestamp 1486834041
transform 1 0 12432 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_328
timestamp 1486834041
transform 1 0 20272 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_329
timestamp 1486834041
transform 1 0 8512 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_330
timestamp 1486834041
transform 1 0 16352 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_331
timestamp 1486834041
transform 1 0 24192 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_332
timestamp 1486834041
transform 1 0 4592 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_333
timestamp 1486834041
transform 1 0 12432 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_334
timestamp 1486834041
transform 1 0 20272 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_335
timestamp 1486834041
transform 1 0 8512 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_336
timestamp 1486834041
transform 1 0 16352 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_337
timestamp 1486834041
transform 1 0 24192 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_338
timestamp 1486834041
transform 1 0 4592 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_339
timestamp 1486834041
transform 1 0 12432 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_340
timestamp 1486834041
transform 1 0 20272 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_341
timestamp 1486834041
transform 1 0 8512 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_342
timestamp 1486834041
transform 1 0 16352 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_343
timestamp 1486834041
transform 1 0 24192 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_344
timestamp 1486834041
transform 1 0 4592 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_345
timestamp 1486834041
transform 1 0 12432 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_346
timestamp 1486834041
transform 1 0 20272 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_347
timestamp 1486834041
transform 1 0 8512 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_348
timestamp 1486834041
transform 1 0 16352 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_349
timestamp 1486834041
transform 1 0 24192 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_350
timestamp 1486834041
transform 1 0 4592 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_351
timestamp 1486834041
transform 1 0 12432 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_352
timestamp 1486834041
transform 1 0 20272 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_353
timestamp 1486834041
transform 1 0 8512 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_354
timestamp 1486834041
transform 1 0 16352 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_355
timestamp 1486834041
transform 1 0 24192 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_356
timestamp 1486834041
transform 1 0 4480 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_357
timestamp 1486834041
transform 1 0 8288 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_358
timestamp 1486834041
transform 1 0 12096 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_359
timestamp 1486834041
transform 1 0 15904 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_360
timestamp 1486834041
transform 1 0 19712 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_361
timestamp 1486834041
transform 1 0 23520 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_362
timestamp 1486834041
transform 1 0 27328 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  wire126
timestamp 1486834041
transform -1 0 17248 0 -1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  wire127
timestamp 1486834041
transform -1 0 14560 0 1 14896
box -86 -86 758 870
<< labels >>
flabel metal3 s 0 3136 112 3248 0 FreeSans 448 0 0 0 A_I_top
port 0 nsew signal output
flabel metal3 s 0 2240 112 2352 0 FreeSans 448 0 0 0 A_O_top
port 1 nsew signal input
flabel metal3 s 0 4032 112 4144 0 FreeSans 448 0 0 0 A_T_top
port 2 nsew signal output
flabel metal3 s 0 12992 112 13104 0 FreeSans 448 0 0 0 A_config_C_bit0
port 3 nsew signal output
flabel metal3 s 0 13888 112 14000 0 FreeSans 448 0 0 0 A_config_C_bit1
port 4 nsew signal output
flabel metal3 s 0 14784 112 14896 0 FreeSans 448 0 0 0 A_config_C_bit2
port 5 nsew signal output
flabel metal3 s 0 15680 112 15792 0 FreeSans 448 0 0 0 A_config_C_bit3
port 6 nsew signal output
flabel metal3 s 0 5824 112 5936 0 FreeSans 448 0 0 0 B_I_top
port 7 nsew signal output
flabel metal3 s 0 4928 112 5040 0 FreeSans 448 0 0 0 B_O_top
port 8 nsew signal input
flabel metal3 s 0 6720 112 6832 0 FreeSans 448 0 0 0 B_T_top
port 9 nsew signal output
flabel metal3 s 0 16576 112 16688 0 FreeSans 448 0 0 0 B_config_C_bit0
port 10 nsew signal output
flabel metal3 s 0 17472 112 17584 0 FreeSans 448 0 0 0 B_config_C_bit1
port 11 nsew signal output
flabel metal3 s 0 18368 112 18480 0 FreeSans 448 0 0 0 B_config_C_bit2
port 12 nsew signal output
flabel metal3 s 0 19264 112 19376 0 FreeSans 448 0 0 0 B_config_C_bit3
port 13 nsew signal output
flabel metal3 s 0 8512 112 8624 0 FreeSans 448 0 0 0 C_I_top
port 14 nsew signal output
flabel metal3 s 0 7616 112 7728 0 FreeSans 448 0 0 0 C_O_top
port 15 nsew signal input
flabel metal3 s 0 9408 112 9520 0 FreeSans 448 0 0 0 C_T_top
port 16 nsew signal output
flabel metal3 s 0 20160 112 20272 0 FreeSans 448 0 0 0 C_config_C_bit0
port 17 nsew signal output
flabel metal3 s 0 21056 112 21168 0 FreeSans 448 0 0 0 C_config_C_bit1
port 18 nsew signal output
flabel metal3 s 0 21952 112 22064 0 FreeSans 448 0 0 0 C_config_C_bit2
port 19 nsew signal output
flabel metal3 s 0 22848 112 22960 0 FreeSans 448 0 0 0 C_config_C_bit3
port 20 nsew signal output
flabel metal3 s 0 11200 112 11312 0 FreeSans 448 0 0 0 D_I_top
port 21 nsew signal output
flabel metal3 s 0 10304 112 10416 0 FreeSans 448 0 0 0 D_O_top
port 22 nsew signal input
flabel metal3 s 0 12096 112 12208 0 FreeSans 448 0 0 0 D_T_top
port 23 nsew signal output
flabel metal3 s 0 23744 112 23856 0 FreeSans 448 0 0 0 D_config_C_bit0
port 24 nsew signal output
flabel metal3 s 0 24640 112 24752 0 FreeSans 448 0 0 0 D_config_C_bit1
port 25 nsew signal output
flabel metal3 s 0 25536 112 25648 0 FreeSans 448 0 0 0 D_config_C_bit2
port 26 nsew signal output
flabel metal3 s 0 26432 112 26544 0 FreeSans 448 0 0 0 D_config_C_bit3
port 27 nsew signal output
flabel metal3 s 28448 21728 28560 21840 0 FreeSans 448 0 0 0 E1BEG[0]
port 28 nsew signal output
flabel metal3 s 28448 22176 28560 22288 0 FreeSans 448 0 0 0 E1BEG[1]
port 29 nsew signal output
flabel metal3 s 28448 22624 28560 22736 0 FreeSans 448 0 0 0 E1BEG[2]
port 30 nsew signal output
flabel metal3 s 28448 23072 28560 23184 0 FreeSans 448 0 0 0 E1BEG[3]
port 31 nsew signal output
flabel metal3 s 28448 23520 28560 23632 0 FreeSans 448 0 0 0 E2BEG[0]
port 32 nsew signal output
flabel metal3 s 28448 23968 28560 24080 0 FreeSans 448 0 0 0 E2BEG[1]
port 33 nsew signal output
flabel metal3 s 28448 24416 28560 24528 0 FreeSans 448 0 0 0 E2BEG[2]
port 34 nsew signal output
flabel metal3 s 28448 24864 28560 24976 0 FreeSans 448 0 0 0 E2BEG[3]
port 35 nsew signal output
flabel metal3 s 28448 25312 28560 25424 0 FreeSans 448 0 0 0 E2BEG[4]
port 36 nsew signal output
flabel metal3 s 28448 25760 28560 25872 0 FreeSans 448 0 0 0 E2BEG[5]
port 37 nsew signal output
flabel metal3 s 28448 26208 28560 26320 0 FreeSans 448 0 0 0 E2BEG[6]
port 38 nsew signal output
flabel metal3 s 28448 26656 28560 26768 0 FreeSans 448 0 0 0 E2BEG[7]
port 39 nsew signal output
flabel metal3 s 28448 27104 28560 27216 0 FreeSans 448 0 0 0 E2BEGb[0]
port 40 nsew signal output
flabel metal3 s 28448 27552 28560 27664 0 FreeSans 448 0 0 0 E2BEGb[1]
port 41 nsew signal output
flabel metal3 s 28448 28000 28560 28112 0 FreeSans 448 0 0 0 E2BEGb[2]
port 42 nsew signal output
flabel metal3 s 28448 28448 28560 28560 0 FreeSans 448 0 0 0 E2BEGb[3]
port 43 nsew signal output
flabel metal3 s 28448 28896 28560 29008 0 FreeSans 448 0 0 0 E2BEGb[4]
port 44 nsew signal output
flabel metal3 s 28448 29344 28560 29456 0 FreeSans 448 0 0 0 E2BEGb[5]
port 45 nsew signal output
flabel metal3 s 28448 29792 28560 29904 0 FreeSans 448 0 0 0 E2BEGb[6]
port 46 nsew signal output
flabel metal3 s 28448 30240 28560 30352 0 FreeSans 448 0 0 0 E2BEGb[7]
port 47 nsew signal output
flabel metal3 s 28448 37856 28560 37968 0 FreeSans 448 0 0 0 E6BEG[0]
port 48 nsew signal output
flabel metal3 s 28448 42336 28560 42448 0 FreeSans 448 0 0 0 E6BEG[10]
port 49 nsew signal output
flabel metal3 s 28448 42784 28560 42896 0 FreeSans 448 0 0 0 E6BEG[11]
port 50 nsew signal output
flabel metal3 s 28448 38304 28560 38416 0 FreeSans 448 0 0 0 E6BEG[1]
port 51 nsew signal output
flabel metal3 s 28448 38752 28560 38864 0 FreeSans 448 0 0 0 E6BEG[2]
port 52 nsew signal output
flabel metal3 s 28448 39200 28560 39312 0 FreeSans 448 0 0 0 E6BEG[3]
port 53 nsew signal output
flabel metal3 s 28448 39648 28560 39760 0 FreeSans 448 0 0 0 E6BEG[4]
port 54 nsew signal output
flabel metal3 s 28448 40096 28560 40208 0 FreeSans 448 0 0 0 E6BEG[5]
port 55 nsew signal output
flabel metal3 s 28448 40544 28560 40656 0 FreeSans 448 0 0 0 E6BEG[6]
port 56 nsew signal output
flabel metal3 s 28448 40992 28560 41104 0 FreeSans 448 0 0 0 E6BEG[7]
port 57 nsew signal output
flabel metal3 s 28448 41440 28560 41552 0 FreeSans 448 0 0 0 E6BEG[8]
port 58 nsew signal output
flabel metal3 s 28448 41888 28560 42000 0 FreeSans 448 0 0 0 E6BEG[9]
port 59 nsew signal output
flabel metal3 s 28448 30688 28560 30800 0 FreeSans 448 0 0 0 EE4BEG[0]
port 60 nsew signal output
flabel metal3 s 28448 35168 28560 35280 0 FreeSans 448 0 0 0 EE4BEG[10]
port 61 nsew signal output
flabel metal3 s 28448 35616 28560 35728 0 FreeSans 448 0 0 0 EE4BEG[11]
port 62 nsew signal output
flabel metal3 s 28448 36064 28560 36176 0 FreeSans 448 0 0 0 EE4BEG[12]
port 63 nsew signal output
flabel metal3 s 28448 36512 28560 36624 0 FreeSans 448 0 0 0 EE4BEG[13]
port 64 nsew signal output
flabel metal3 s 28448 36960 28560 37072 0 FreeSans 448 0 0 0 EE4BEG[14]
port 65 nsew signal output
flabel metal3 s 28448 37408 28560 37520 0 FreeSans 448 0 0 0 EE4BEG[15]
port 66 nsew signal output
flabel metal3 s 28448 31136 28560 31248 0 FreeSans 448 0 0 0 EE4BEG[1]
port 67 nsew signal output
flabel metal3 s 28448 31584 28560 31696 0 FreeSans 448 0 0 0 EE4BEG[2]
port 68 nsew signal output
flabel metal3 s 28448 32032 28560 32144 0 FreeSans 448 0 0 0 EE4BEG[3]
port 69 nsew signal output
flabel metal3 s 28448 32480 28560 32592 0 FreeSans 448 0 0 0 EE4BEG[4]
port 70 nsew signal output
flabel metal3 s 28448 32928 28560 33040 0 FreeSans 448 0 0 0 EE4BEG[5]
port 71 nsew signal output
flabel metal3 s 28448 33376 28560 33488 0 FreeSans 448 0 0 0 EE4BEG[6]
port 72 nsew signal output
flabel metal3 s 28448 33824 28560 33936 0 FreeSans 448 0 0 0 EE4BEG[7]
port 73 nsew signal output
flabel metal3 s 28448 34272 28560 34384 0 FreeSans 448 0 0 0 EE4BEG[8]
port 74 nsew signal output
flabel metal3 s 28448 34720 28560 34832 0 FreeSans 448 0 0 0 EE4BEG[9]
port 75 nsew signal output
flabel metal3 s 0 27328 112 27440 0 FreeSans 448 0 0 0 FrameData[0]
port 76 nsew signal input
flabel metal3 s 0 36288 112 36400 0 FreeSans 448 0 0 0 FrameData[10]
port 77 nsew signal input
flabel metal3 s 0 37184 112 37296 0 FreeSans 448 0 0 0 FrameData[11]
port 78 nsew signal input
flabel metal3 s 0 38080 112 38192 0 FreeSans 448 0 0 0 FrameData[12]
port 79 nsew signal input
flabel metal3 s 0 38976 112 39088 0 FreeSans 448 0 0 0 FrameData[13]
port 80 nsew signal input
flabel metal3 s 0 39872 112 39984 0 FreeSans 448 0 0 0 FrameData[14]
port 81 nsew signal input
flabel metal3 s 0 40768 112 40880 0 FreeSans 448 0 0 0 FrameData[15]
port 82 nsew signal input
flabel metal3 s 0 41664 112 41776 0 FreeSans 448 0 0 0 FrameData[16]
port 83 nsew signal input
flabel metal3 s 0 42560 112 42672 0 FreeSans 448 0 0 0 FrameData[17]
port 84 nsew signal input
flabel metal3 s 0 43456 112 43568 0 FreeSans 448 0 0 0 FrameData[18]
port 85 nsew signal input
flabel metal3 s 0 44352 112 44464 0 FreeSans 448 0 0 0 FrameData[19]
port 86 nsew signal input
flabel metal3 s 0 28224 112 28336 0 FreeSans 448 0 0 0 FrameData[1]
port 87 nsew signal input
flabel metal3 s 0 45248 112 45360 0 FreeSans 448 0 0 0 FrameData[20]
port 88 nsew signal input
flabel metal3 s 0 46144 112 46256 0 FreeSans 448 0 0 0 FrameData[21]
port 89 nsew signal input
flabel metal3 s 0 47040 112 47152 0 FreeSans 448 0 0 0 FrameData[22]
port 90 nsew signal input
flabel metal3 s 0 47936 112 48048 0 FreeSans 448 0 0 0 FrameData[23]
port 91 nsew signal input
flabel metal3 s 0 48832 112 48944 0 FreeSans 448 0 0 0 FrameData[24]
port 92 nsew signal input
flabel metal3 s 0 49728 112 49840 0 FreeSans 448 0 0 0 FrameData[25]
port 93 nsew signal input
flabel metal3 s 0 50624 112 50736 0 FreeSans 448 0 0 0 FrameData[26]
port 94 nsew signal input
flabel metal3 s 0 51520 112 51632 0 FreeSans 448 0 0 0 FrameData[27]
port 95 nsew signal input
flabel metal3 s 0 52416 112 52528 0 FreeSans 448 0 0 0 FrameData[28]
port 96 nsew signal input
flabel metal3 s 0 53312 112 53424 0 FreeSans 448 0 0 0 FrameData[29]
port 97 nsew signal input
flabel metal3 s 0 29120 112 29232 0 FreeSans 448 0 0 0 FrameData[2]
port 98 nsew signal input
flabel metal3 s 0 54208 112 54320 0 FreeSans 448 0 0 0 FrameData[30]
port 99 nsew signal input
flabel metal3 s 0 55104 112 55216 0 FreeSans 448 0 0 0 FrameData[31]
port 100 nsew signal input
flabel metal3 s 0 30016 112 30128 0 FreeSans 448 0 0 0 FrameData[3]
port 101 nsew signal input
flabel metal3 s 0 30912 112 31024 0 FreeSans 448 0 0 0 FrameData[4]
port 102 nsew signal input
flabel metal3 s 0 31808 112 31920 0 FreeSans 448 0 0 0 FrameData[5]
port 103 nsew signal input
flabel metal3 s 0 32704 112 32816 0 FreeSans 448 0 0 0 FrameData[6]
port 104 nsew signal input
flabel metal3 s 0 33600 112 33712 0 FreeSans 448 0 0 0 FrameData[7]
port 105 nsew signal input
flabel metal3 s 0 34496 112 34608 0 FreeSans 448 0 0 0 FrameData[8]
port 106 nsew signal input
flabel metal3 s 0 35392 112 35504 0 FreeSans 448 0 0 0 FrameData[9]
port 107 nsew signal input
flabel metal3 s 28448 43232 28560 43344 0 FreeSans 448 0 0 0 FrameData_O[0]
port 108 nsew signal output
flabel metal3 s 28448 47712 28560 47824 0 FreeSans 448 0 0 0 FrameData_O[10]
port 109 nsew signal output
flabel metal3 s 28448 48160 28560 48272 0 FreeSans 448 0 0 0 FrameData_O[11]
port 110 nsew signal output
flabel metal3 s 28448 48608 28560 48720 0 FreeSans 448 0 0 0 FrameData_O[12]
port 111 nsew signal output
flabel metal3 s 28448 49056 28560 49168 0 FreeSans 448 0 0 0 FrameData_O[13]
port 112 nsew signal output
flabel metal3 s 28448 49504 28560 49616 0 FreeSans 448 0 0 0 FrameData_O[14]
port 113 nsew signal output
flabel metal3 s 28448 49952 28560 50064 0 FreeSans 448 0 0 0 FrameData_O[15]
port 114 nsew signal output
flabel metal3 s 28448 50400 28560 50512 0 FreeSans 448 0 0 0 FrameData_O[16]
port 115 nsew signal output
flabel metal3 s 28448 50848 28560 50960 0 FreeSans 448 0 0 0 FrameData_O[17]
port 116 nsew signal output
flabel metal3 s 28448 51296 28560 51408 0 FreeSans 448 0 0 0 FrameData_O[18]
port 117 nsew signal output
flabel metal3 s 28448 51744 28560 51856 0 FreeSans 448 0 0 0 FrameData_O[19]
port 118 nsew signal output
flabel metal3 s 28448 43680 28560 43792 0 FreeSans 448 0 0 0 FrameData_O[1]
port 119 nsew signal output
flabel metal3 s 28448 52192 28560 52304 0 FreeSans 448 0 0 0 FrameData_O[20]
port 120 nsew signal output
flabel metal3 s 28448 52640 28560 52752 0 FreeSans 448 0 0 0 FrameData_O[21]
port 121 nsew signal output
flabel metal3 s 28448 53088 28560 53200 0 FreeSans 448 0 0 0 FrameData_O[22]
port 122 nsew signal output
flabel metal3 s 28448 53536 28560 53648 0 FreeSans 448 0 0 0 FrameData_O[23]
port 123 nsew signal output
flabel metal3 s 28448 53984 28560 54096 0 FreeSans 448 0 0 0 FrameData_O[24]
port 124 nsew signal output
flabel metal3 s 28448 54432 28560 54544 0 FreeSans 448 0 0 0 FrameData_O[25]
port 125 nsew signal output
flabel metal3 s 28448 54880 28560 54992 0 FreeSans 448 0 0 0 FrameData_O[26]
port 126 nsew signal output
flabel metal3 s 28448 55328 28560 55440 0 FreeSans 448 0 0 0 FrameData_O[27]
port 127 nsew signal output
flabel metal3 s 28448 55776 28560 55888 0 FreeSans 448 0 0 0 FrameData_O[28]
port 128 nsew signal output
flabel metal3 s 28448 56224 28560 56336 0 FreeSans 448 0 0 0 FrameData_O[29]
port 129 nsew signal output
flabel metal3 s 28448 44128 28560 44240 0 FreeSans 448 0 0 0 FrameData_O[2]
port 130 nsew signal output
flabel metal3 s 28448 56672 28560 56784 0 FreeSans 448 0 0 0 FrameData_O[30]
port 131 nsew signal output
flabel metal3 s 28448 57120 28560 57232 0 FreeSans 448 0 0 0 FrameData_O[31]
port 132 nsew signal output
flabel metal3 s 28448 44576 28560 44688 0 FreeSans 448 0 0 0 FrameData_O[3]
port 133 nsew signal output
flabel metal3 s 28448 45024 28560 45136 0 FreeSans 448 0 0 0 FrameData_O[4]
port 134 nsew signal output
flabel metal3 s 28448 45472 28560 45584 0 FreeSans 448 0 0 0 FrameData_O[5]
port 135 nsew signal output
flabel metal3 s 28448 45920 28560 46032 0 FreeSans 448 0 0 0 FrameData_O[6]
port 136 nsew signal output
flabel metal3 s 28448 46368 28560 46480 0 FreeSans 448 0 0 0 FrameData_O[7]
port 137 nsew signal output
flabel metal3 s 28448 46816 28560 46928 0 FreeSans 448 0 0 0 FrameData_O[8]
port 138 nsew signal output
flabel metal3 s 28448 47264 28560 47376 0 FreeSans 448 0 0 0 FrameData_O[9]
port 139 nsew signal output
flabel metal2 s 2016 0 2128 112 0 FreeSans 448 0 0 0 FrameStrobe[0]
port 140 nsew signal input
flabel metal2 s 15456 0 15568 112 0 FreeSans 448 0 0 0 FrameStrobe[10]
port 141 nsew signal input
flabel metal2 s 16800 0 16912 112 0 FreeSans 448 0 0 0 FrameStrobe[11]
port 142 nsew signal input
flabel metal2 s 18144 0 18256 112 0 FreeSans 448 0 0 0 FrameStrobe[12]
port 143 nsew signal input
flabel metal2 s 19488 0 19600 112 0 FreeSans 448 0 0 0 FrameStrobe[13]
port 144 nsew signal input
flabel metal2 s 20832 0 20944 112 0 FreeSans 448 0 0 0 FrameStrobe[14]
port 145 nsew signal input
flabel metal2 s 22176 0 22288 112 0 FreeSans 448 0 0 0 FrameStrobe[15]
port 146 nsew signal input
flabel metal2 s 23520 0 23632 112 0 FreeSans 448 0 0 0 FrameStrobe[16]
port 147 nsew signal input
flabel metal2 s 24864 0 24976 112 0 FreeSans 448 0 0 0 FrameStrobe[17]
port 148 nsew signal input
flabel metal2 s 26208 0 26320 112 0 FreeSans 448 0 0 0 FrameStrobe[18]
port 149 nsew signal input
flabel metal2 s 27552 0 27664 112 0 FreeSans 448 0 0 0 FrameStrobe[19]
port 150 nsew signal input
flabel metal2 s 3360 0 3472 112 0 FreeSans 448 0 0 0 FrameStrobe[1]
port 151 nsew signal input
flabel metal2 s 4704 0 4816 112 0 FreeSans 448 0 0 0 FrameStrobe[2]
port 152 nsew signal input
flabel metal2 s 6048 0 6160 112 0 FreeSans 448 0 0 0 FrameStrobe[3]
port 153 nsew signal input
flabel metal2 s 7392 0 7504 112 0 FreeSans 448 0 0 0 FrameStrobe[4]
port 154 nsew signal input
flabel metal2 s 8736 0 8848 112 0 FreeSans 448 0 0 0 FrameStrobe[5]
port 155 nsew signal input
flabel metal2 s 10080 0 10192 112 0 FreeSans 448 0 0 0 FrameStrobe[6]
port 156 nsew signal input
flabel metal2 s 11424 0 11536 112 0 FreeSans 448 0 0 0 FrameStrobe[7]
port 157 nsew signal input
flabel metal2 s 12768 0 12880 112 0 FreeSans 448 0 0 0 FrameStrobe[8]
port 158 nsew signal input
flabel metal2 s 14112 0 14224 112 0 FreeSans 448 0 0 0 FrameStrobe[9]
port 159 nsew signal input
flabel metal2 s 2016 57344 2128 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[0]
port 160 nsew signal output
flabel metal2 s 15456 57344 15568 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[10]
port 161 nsew signal output
flabel metal2 s 16800 57344 16912 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[11]
port 162 nsew signal output
flabel metal2 s 18144 57344 18256 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[12]
port 163 nsew signal output
flabel metal2 s 19488 57344 19600 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[13]
port 164 nsew signal output
flabel metal2 s 20832 57344 20944 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[14]
port 165 nsew signal output
flabel metal2 s 22176 57344 22288 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[15]
port 166 nsew signal output
flabel metal2 s 23520 57344 23632 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[16]
port 167 nsew signal output
flabel metal2 s 24864 57344 24976 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[17]
port 168 nsew signal output
flabel metal2 s 26208 57344 26320 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[18]
port 169 nsew signal output
flabel metal2 s 27552 57344 27664 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[19]
port 170 nsew signal output
flabel metal2 s 3360 57344 3472 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[1]
port 171 nsew signal output
flabel metal2 s 4704 57344 4816 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[2]
port 172 nsew signal output
flabel metal2 s 6048 57344 6160 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[3]
port 173 nsew signal output
flabel metal2 s 7392 57344 7504 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[4]
port 174 nsew signal output
flabel metal2 s 8736 57344 8848 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[5]
port 175 nsew signal output
flabel metal2 s 10080 57344 10192 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[6]
port 176 nsew signal output
flabel metal2 s 11424 57344 11536 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[7]
port 177 nsew signal output
flabel metal2 s 12768 57344 12880 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[8]
port 178 nsew signal output
flabel metal2 s 14112 57344 14224 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[9]
port 179 nsew signal output
flabel metal2 s 672 0 784 112 0 FreeSans 448 0 0 0 UserCLK
port 180 nsew signal input
flabel metal2 s 672 57344 784 57456 0 FreeSans 448 0 0 0 UserCLKo
port 181 nsew signal output
flabel metal4 s 3776 0 4096 57456 0 FreeSans 1472 90 0 0 VDD
port 182 nsew power bidirectional
flabel metal4 s 3776 0 4096 56 0 FreeSans 368 0 0 0 VDD
port 182 nsew power bidirectional
flabel metal4 s 3776 57400 4096 57456 0 FreeSans 368 0 0 0 VDD
port 182 nsew power bidirectional
flabel metal4 s 23776 0 24096 57456 0 FreeSans 1472 90 0 0 VDD
port 182 nsew power bidirectional
flabel metal4 s 23776 0 24096 56 0 FreeSans 368 0 0 0 VDD
port 182 nsew power bidirectional
flabel metal4 s 23776 57400 24096 57456 0 FreeSans 368 0 0 0 VDD
port 182 nsew power bidirectional
flabel metal4 s 4436 0 4756 57456 0 FreeSans 1472 90 0 0 VSS
port 183 nsew ground bidirectional
flabel metal4 s 4436 0 4756 56 0 FreeSans 368 0 0 0 VSS
port 183 nsew ground bidirectional
flabel metal4 s 4436 57400 4756 57456 0 FreeSans 368 0 0 0 VSS
port 183 nsew ground bidirectional
flabel metal4 s 24436 0 24756 57456 0 FreeSans 1472 90 0 0 VSS
port 183 nsew ground bidirectional
flabel metal4 s 24436 0 24756 56 0 FreeSans 368 0 0 0 VSS
port 183 nsew ground bidirectional
flabel metal4 s 24436 57400 24756 57456 0 FreeSans 368 0 0 0 VSS
port 183 nsew ground bidirectional
flabel metal3 s 28448 224 28560 336 0 FreeSans 448 0 0 0 W1END[0]
port 184 nsew signal input
flabel metal3 s 28448 672 28560 784 0 FreeSans 448 0 0 0 W1END[1]
port 185 nsew signal input
flabel metal3 s 28448 1120 28560 1232 0 FreeSans 448 0 0 0 W1END[2]
port 186 nsew signal input
flabel metal3 s 28448 1568 28560 1680 0 FreeSans 448 0 0 0 W1END[3]
port 187 nsew signal input
flabel metal3 s 28448 5600 28560 5712 0 FreeSans 448 0 0 0 W2END[0]
port 188 nsew signal input
flabel metal3 s 28448 6048 28560 6160 0 FreeSans 448 0 0 0 W2END[1]
port 189 nsew signal input
flabel metal3 s 28448 6496 28560 6608 0 FreeSans 448 0 0 0 W2END[2]
port 190 nsew signal input
flabel metal3 s 28448 6944 28560 7056 0 FreeSans 448 0 0 0 W2END[3]
port 191 nsew signal input
flabel metal3 s 28448 7392 28560 7504 0 FreeSans 448 0 0 0 W2END[4]
port 192 nsew signal input
flabel metal3 s 28448 7840 28560 7952 0 FreeSans 448 0 0 0 W2END[5]
port 193 nsew signal input
flabel metal3 s 28448 8288 28560 8400 0 FreeSans 448 0 0 0 W2END[6]
port 194 nsew signal input
flabel metal3 s 28448 8736 28560 8848 0 FreeSans 448 0 0 0 W2END[7]
port 195 nsew signal input
flabel metal3 s 28448 2016 28560 2128 0 FreeSans 448 0 0 0 W2MID[0]
port 196 nsew signal input
flabel metal3 s 28448 2464 28560 2576 0 FreeSans 448 0 0 0 W2MID[1]
port 197 nsew signal input
flabel metal3 s 28448 2912 28560 3024 0 FreeSans 448 0 0 0 W2MID[2]
port 198 nsew signal input
flabel metal3 s 28448 3360 28560 3472 0 FreeSans 448 0 0 0 W2MID[3]
port 199 nsew signal input
flabel metal3 s 28448 3808 28560 3920 0 FreeSans 448 0 0 0 W2MID[4]
port 200 nsew signal input
flabel metal3 s 28448 4256 28560 4368 0 FreeSans 448 0 0 0 W2MID[5]
port 201 nsew signal input
flabel metal3 s 28448 4704 28560 4816 0 FreeSans 448 0 0 0 W2MID[6]
port 202 nsew signal input
flabel metal3 s 28448 5152 28560 5264 0 FreeSans 448 0 0 0 W2MID[7]
port 203 nsew signal input
flabel metal3 s 28448 16352 28560 16464 0 FreeSans 448 0 0 0 W6END[0]
port 204 nsew signal input
flabel metal3 s 28448 20832 28560 20944 0 FreeSans 448 0 0 0 W6END[10]
port 205 nsew signal input
flabel metal3 s 28448 21280 28560 21392 0 FreeSans 448 0 0 0 W6END[11]
port 206 nsew signal input
flabel metal3 s 28448 16800 28560 16912 0 FreeSans 448 0 0 0 W6END[1]
port 207 nsew signal input
flabel metal3 s 28448 17248 28560 17360 0 FreeSans 448 0 0 0 W6END[2]
port 208 nsew signal input
flabel metal3 s 28448 17696 28560 17808 0 FreeSans 448 0 0 0 W6END[3]
port 209 nsew signal input
flabel metal3 s 28448 18144 28560 18256 0 FreeSans 448 0 0 0 W6END[4]
port 210 nsew signal input
flabel metal3 s 28448 18592 28560 18704 0 FreeSans 448 0 0 0 W6END[5]
port 211 nsew signal input
flabel metal3 s 28448 19040 28560 19152 0 FreeSans 448 0 0 0 W6END[6]
port 212 nsew signal input
flabel metal3 s 28448 19488 28560 19600 0 FreeSans 448 0 0 0 W6END[7]
port 213 nsew signal input
flabel metal3 s 28448 19936 28560 20048 0 FreeSans 448 0 0 0 W6END[8]
port 214 nsew signal input
flabel metal3 s 28448 20384 28560 20496 0 FreeSans 448 0 0 0 W6END[9]
port 215 nsew signal input
flabel metal3 s 28448 9184 28560 9296 0 FreeSans 448 0 0 0 WW4END[0]
port 216 nsew signal input
flabel metal3 s 28448 13664 28560 13776 0 FreeSans 448 0 0 0 WW4END[10]
port 217 nsew signal input
flabel metal3 s 28448 14112 28560 14224 0 FreeSans 448 0 0 0 WW4END[11]
port 218 nsew signal input
flabel metal3 s 28448 14560 28560 14672 0 FreeSans 448 0 0 0 WW4END[12]
port 219 nsew signal input
flabel metal3 s 28448 15008 28560 15120 0 FreeSans 448 0 0 0 WW4END[13]
port 220 nsew signal input
flabel metal3 s 28448 15456 28560 15568 0 FreeSans 448 0 0 0 WW4END[14]
port 221 nsew signal input
flabel metal3 s 28448 15904 28560 16016 0 FreeSans 448 0 0 0 WW4END[15]
port 222 nsew signal input
flabel metal3 s 28448 9632 28560 9744 0 FreeSans 448 0 0 0 WW4END[1]
port 223 nsew signal input
flabel metal3 s 28448 10080 28560 10192 0 FreeSans 448 0 0 0 WW4END[2]
port 224 nsew signal input
flabel metal3 s 28448 10528 28560 10640 0 FreeSans 448 0 0 0 WW4END[3]
port 225 nsew signal input
flabel metal3 s 28448 10976 28560 11088 0 FreeSans 448 0 0 0 WW4END[4]
port 226 nsew signal input
flabel metal3 s 28448 11424 28560 11536 0 FreeSans 448 0 0 0 WW4END[5]
port 227 nsew signal input
flabel metal3 s 28448 11872 28560 11984 0 FreeSans 448 0 0 0 WW4END[6]
port 228 nsew signal input
flabel metal3 s 28448 12320 28560 12432 0 FreeSans 448 0 0 0 WW4END[7]
port 229 nsew signal input
flabel metal3 s 28448 12768 28560 12880 0 FreeSans 448 0 0 0 WW4END[8]
port 230 nsew signal input
flabel metal3 s 28448 13216 28560 13328 0 FreeSans 448 0 0 0 WW4END[9]
port 231 nsew signal input
rlabel metal1 14280 56448 14280 56448 0 VDD
rlabel metal1 14280 55664 14280 55664 0 VSS
rlabel metal3 686 3192 686 3192 0 A_I_top
rlabel metal3 966 2296 966 2296 0 A_O_top
rlabel metal3 798 4088 798 4088 0 A_T_top
rlabel metal2 2968 11088 2968 11088 0 A_config_C_bit0
rlabel metal3 742 13944 742 13944 0 A_config_C_bit1
rlabel metal3 1246 14840 1246 14840 0 A_config_C_bit2
rlabel metal3 1470 15736 1470 15736 0 A_config_C_bit3
rlabel metal3 1470 5880 1470 5880 0 B_I_top
rlabel metal3 1022 4984 1022 4984 0 B_O_top
rlabel metal3 798 6776 798 6776 0 B_T_top
rlabel metal3 2702 16632 2702 16632 0 B_config_C_bit0
rlabel metal2 1288 8260 1288 8260 0 B_config_C_bit1
rlabel metal3 1008 9240 1008 9240 0 B_config_C_bit2
rlabel metal3 630 19320 630 19320 0 B_config_C_bit3
rlabel metal3 854 8568 854 8568 0 C_I_top
rlabel metal3 910 7672 910 7672 0 C_O_top
rlabel metal2 2800 7672 2800 7672 0 C_T_top
rlabel metal3 1414 20216 1414 20216 0 C_config_C_bit0
rlabel metal3 1582 21112 1582 21112 0 C_config_C_bit1
rlabel metal3 798 22008 798 22008 0 C_config_C_bit2
rlabel metal2 5544 21560 5544 21560 0 C_config_C_bit3
rlabel metal3 1582 11256 1582 11256 0 D_I_top
rlabel metal2 2968 20496 2968 20496 0 D_O_top
rlabel metal2 1064 6552 1064 6552 0 D_T_top
rlabel metal3 742 23800 742 23800 0 D_config_C_bit0
rlabel metal4 3528 24528 3528 24528 0 D_config_C_bit1
rlabel metal2 5544 25256 5544 25256 0 D_config_C_bit2
rlabel metal3 686 26488 686 26488 0 D_config_C_bit3
rlabel metal2 25704 21952 25704 21952 0 E1BEG[0]
rlabel metal2 27160 21952 27160 21952 0 E1BEG[1]
rlabel metal2 27272 22456 27272 22456 0 E1BEG[2]
rlabel metal2 25704 23408 25704 23408 0 E1BEG[3]
rlabel metal2 27272 23464 27272 23464 0 E2BEG[0]
rlabel metal2 25704 24416 25704 24416 0 E2BEG[1]
rlabel metal2 27272 24136 27272 24136 0 E2BEG[2]
rlabel metal3 27706 24920 27706 24920 0 E2BEG[3]
rlabel metal2 27160 25088 27160 25088 0 E2BEG[4]
rlabel metal2 27272 25592 27272 25592 0 E2BEG[5]
rlabel metal3 27090 26264 27090 26264 0 E2BEG[6]
rlabel metal2 27272 26600 27272 26600 0 E2BEG[7]
rlabel metal2 25704 27552 25704 27552 0 E2BEGb[0]
rlabel metal2 27048 27384 27048 27384 0 E2BEGb[1]
rlabel metal3 27874 28056 27874 28056 0 E2BEGb[2]
rlabel metal3 27874 28504 27874 28504 0 E2BEGb[3]
rlabel metal3 27874 28952 27874 28952 0 E2BEGb[4]
rlabel metal3 27818 29400 27818 29400 0 E2BEGb[5]
rlabel metal3 27762 29848 27762 29848 0 E2BEGb[6]
rlabel metal3 27874 30296 27874 30296 0 E2BEGb[7]
rlabel metal3 27090 37912 27090 37912 0 E6BEG[0]
rlabel metal3 27090 42392 27090 42392 0 E6BEG[10]
rlabel metal3 27874 42840 27874 42840 0 E6BEG[11]
rlabel metal3 27874 38360 27874 38360 0 E6BEG[1]
rlabel metal3 27818 38808 27818 38808 0 E6BEG[2]
rlabel metal3 27090 39256 27090 39256 0 E6BEG[3]
rlabel metal3 27874 39704 27874 39704 0 E6BEG[4]
rlabel metal3 27090 40152 27090 40152 0 E6BEG[5]
rlabel metal3 27762 40600 27762 40600 0 E6BEG[6]
rlabel metal3 27090 41048 27090 41048 0 E6BEG[7]
rlabel metal3 27874 41496 27874 41496 0 E6BEG[8]
rlabel metal3 27818 41944 27818 41944 0 E6BEG[9]
rlabel metal2 25480 30800 25480 30800 0 EE4BEG[0]
rlabel metal3 27874 35224 27874 35224 0 EE4BEG[10]
rlabel metal3 27818 35672 27818 35672 0 EE4BEG[11]
rlabel metal2 25704 36176 25704 36176 0 EE4BEG[12]
rlabel metal3 27874 36568 27874 36568 0 EE4BEG[13]
rlabel metal2 25480 37072 25480 37072 0 EE4BEG[14]
rlabel metal3 27762 37464 27762 37464 0 EE4BEG[15]
rlabel metal3 27762 31192 27762 31192 0 EE4BEG[1]
rlabel metal3 27090 31640 27090 31640 0 EE4BEG[2]
rlabel metal3 27874 32088 27874 32088 0 EE4BEG[3]
rlabel metal3 27818 32536 27818 32536 0 EE4BEG[4]
rlabel metal2 25704 33040 25704 33040 0 EE4BEG[5]
rlabel metal3 27874 33432 27874 33432 0 EE4BEG[6]
rlabel metal2 25704 34048 25704 34048 0 EE4BEG[7]
rlabel metal3 27762 34328 27762 34328 0 EE4BEG[8]
rlabel metal3 27090 34776 27090 34776 0 EE4BEG[9]
rlabel metal2 6720 26152 6720 26152 0 FrameData[0]
rlabel metal2 12712 18424 12712 18424 0 FrameData[10]
rlabel metal2 10920 19600 10920 19600 0 FrameData[11]
rlabel metal2 1848 24472 1848 24472 0 FrameData[12]
rlabel metal2 2464 24584 2464 24584 0 FrameData[13]
rlabel metal3 1134 39928 1134 39928 0 FrameData[14]
rlabel metal2 3024 26040 3024 26040 0 FrameData[15]
rlabel metal2 1624 22120 1624 22120 0 FrameData[16]
rlabel metal2 2744 23072 2744 23072 0 FrameData[17]
rlabel metal2 17080 20608 17080 20608 0 FrameData[18]
rlabel metal2 17752 44044 17752 44044 0 FrameData[19]
rlabel metal3 8064 23464 8064 23464 0 FrameData[1]
rlabel metal2 9352 20160 9352 20160 0 FrameData[20]
rlabel metal2 10976 25816 10976 25816 0 FrameData[21]
rlabel metal3 574 47096 574 47096 0 FrameData[22]
rlabel metal2 17304 25928 17304 25928 0 FrameData[23]
rlabel metal3 1526 48888 1526 48888 0 FrameData[24]
rlabel metal2 22568 14784 22568 14784 0 FrameData[25]
rlabel metal3 5446 50680 5446 50680 0 FrameData[26]
rlabel metal3 6902 51576 6902 51576 0 FrameData[27]
rlabel metal3 2408 25256 2408 25256 0 FrameData[28]
rlabel metal3 2296 26152 2296 26152 0 FrameData[29]
rlabel metal2 2744 39256 2744 39256 0 FrameData[2]
rlabel metal3 3038 54264 3038 54264 0 FrameData[30]
rlabel metal3 1638 55160 1638 55160 0 FrameData[31]
rlabel metal2 2856 36008 2856 36008 0 FrameData[3]
rlabel metal2 16408 38136 16408 38136 0 FrameData[4]
rlabel metal3 13160 22456 13160 22456 0 FrameData[5]
rlabel metal2 17864 33320 17864 33320 0 FrameData[6]
rlabel metal3 18200 28728 18200 28728 0 FrameData[7]
rlabel metal3 5712 18312 5712 18312 0 FrameData[8]
rlabel metal2 10528 17752 10528 17752 0 FrameData[9]
rlabel metal3 27090 43288 27090 43288 0 FrameData_O[0]
rlabel metal3 27874 47768 27874 47768 0 FrameData_O[10]
rlabel metal3 27818 48216 27818 48216 0 FrameData_O[11]
rlabel metal3 27090 48664 27090 48664 0 FrameData_O[12]
rlabel metal3 27874 49112 27874 49112 0 FrameData_O[13]
rlabel metal3 27090 49560 27090 49560 0 FrameData_O[14]
rlabel metal3 27762 50008 27762 50008 0 FrameData_O[15]
rlabel metal3 27090 50456 27090 50456 0 FrameData_O[16]
rlabel metal3 27874 50904 27874 50904 0 FrameData_O[17]
rlabel metal3 27818 51352 27818 51352 0 FrameData_O[18]
rlabel metal3 27090 51800 27090 51800 0 FrameData_O[19]
rlabel metal3 27762 43736 27762 43736 0 FrameData_O[1]
rlabel metal3 27874 52248 27874 52248 0 FrameData_O[20]
rlabel metal3 26978 52696 26978 52696 0 FrameData_O[21]
rlabel metal3 27762 53144 27762 53144 0 FrameData_O[22]
rlabel metal3 27090 53592 27090 53592 0 FrameData_O[23]
rlabel metal3 27874 54040 27874 54040 0 FrameData_O[24]
rlabel metal3 27090 54488 27090 54488 0 FrameData_O[25]
rlabel metal3 27314 54936 27314 54936 0 FrameData_O[26]
rlabel metal2 23800 53984 23800 53984 0 FrameData_O[27]
rlabel metal3 25522 55832 25522 55832 0 FrameData_O[28]
rlabel metal2 25760 51576 25760 51576 0 FrameData_O[29]
rlabel metal3 27090 44184 27090 44184 0 FrameData_O[2]
rlabel metal2 24192 53144 24192 53144 0 FrameData_O[30]
rlabel metal2 23688 53312 23688 53312 0 FrameData_O[31]
rlabel metal3 27874 44632 27874 44632 0 FrameData_O[3]
rlabel metal3 27818 45080 27818 45080 0 FrameData_O[4]
rlabel metal3 27090 45528 27090 45528 0 FrameData_O[5]
rlabel metal3 27874 45976 27874 45976 0 FrameData_O[6]
rlabel metal3 27090 46424 27090 46424 0 FrameData_O[7]
rlabel metal3 27762 46872 27762 46872 0 FrameData_O[8]
rlabel metal3 27090 47320 27090 47320 0 FrameData_O[9]
rlabel metal2 2072 3486 2072 3486 0 FrameStrobe[0]
rlabel metal2 26936 20468 26936 20468 0 FrameStrobe[10]
rlabel metal4 27048 29848 27048 29848 0 FrameStrobe[11]
rlabel metal2 26040 1288 26040 1288 0 FrameStrobe[12]
rlabel metal2 26936 1176 26936 1176 0 FrameStrobe[13]
rlabel metal3 25760 52360 25760 52360 0 FrameStrobe[14]
rlabel metal2 22232 1022 22232 1022 0 FrameStrobe[15]
rlabel metal2 23576 294 23576 294 0 FrameStrobe[16]
rlabel metal2 24920 854 24920 854 0 FrameStrobe[17]
rlabel metal2 26264 910 26264 910 0 FrameStrobe[18]
rlabel metal2 27608 2590 27608 2590 0 FrameStrobe[19]
rlabel metal2 3416 854 3416 854 0 FrameStrobe[1]
rlabel metal2 4760 294 4760 294 0 FrameStrobe[2]
rlabel metal2 6104 182 6104 182 0 FrameStrobe[3]
rlabel metal2 7448 126 7448 126 0 FrameStrobe[4]
rlabel metal3 21112 19432 21112 19432 0 FrameStrobe[5]
rlabel metal2 20664 54040 20664 54040 0 FrameStrobe[6]
rlabel metal2 11480 126 11480 126 0 FrameStrobe[7]
rlabel metal4 19096 40600 19096 40600 0 FrameStrobe[8]
rlabel metal2 14168 518 14168 518 0 FrameStrobe[9]
rlabel metal2 2520 55300 2520 55300 0 FrameStrobe_O[0]
rlabel metal3 16016 56280 16016 56280 0 FrameStrobe_O[10]
rlabel metal2 17304 55300 17304 55300 0 FrameStrobe_O[11]
rlabel metal2 18368 56280 18368 56280 0 FrameStrobe_O[12]
rlabel metal2 20328 56840 20328 56840 0 FrameStrobe_O[13]
rlabel metal2 20888 56826 20888 56826 0 FrameStrobe_O[14]
rlabel metal2 23016 56448 23016 56448 0 FrameStrobe_O[15]
rlabel metal2 23576 56826 23576 56826 0 FrameStrobe_O[16]
rlabel metal2 24920 56826 24920 56826 0 FrameStrobe_O[17]
rlabel metal2 26264 57330 26264 57330 0 FrameStrobe_O[18]
rlabel metal2 27608 56994 27608 56994 0 FrameStrobe_O[19]
rlabel metal2 3416 56826 3416 56826 0 FrameStrobe_O[1]
rlabel metal2 5208 56448 5208 56448 0 FrameStrobe_O[2]
rlabel metal3 6496 55160 6496 55160 0 FrameStrobe_O[3]
rlabel metal2 7448 56770 7448 56770 0 FrameStrobe_O[4]
rlabel metal2 9016 56448 9016 56448 0 FrameStrobe_O[5]
rlabel metal2 10584 56504 10584 56504 0 FrameStrobe_O[6]
rlabel metal3 11704 55160 11704 55160 0 FrameStrobe_O[7]
rlabel metal2 13048 56448 13048 56448 0 FrameStrobe_O[8]
rlabel metal2 14616 56504 14616 56504 0 FrameStrobe_O[9]
rlabel metal3 21168 24808 21168 24808 0 Inst_A_IO_1_bidirectional_frame_config_pass.Q
rlabel metal2 21392 30968 21392 30968 0 Inst_B_IO_1_bidirectional_frame_config_pass.Q
rlabel metal2 15512 16072 15512 16072 0 Inst_C_IO_1_bidirectional_frame_config_pass.Q
rlabel metal3 14168 19992 14168 19992 0 Inst_D_IO_1_bidirectional_frame_config_pass.Q
rlabel metal3 9184 34104 9184 34104 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit0.Q
rlabel metal2 9128 34384 9128 34384 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit1.Q
rlabel metal2 15400 9520 15400 9520 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit10.Q
rlabel metal3 18592 15288 18592 15288 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit11.Q
rlabel metal3 18928 14616 18928 14616 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit12.Q
rlabel metal2 16072 13832 16072 13832 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit13.Q
rlabel metal3 17528 12152 17528 12152 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit14.Q
rlabel metal2 7896 14560 7896 14560 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit15.Q
rlabel metal2 7560 15568 7560 15568 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit16.Q
rlabel metal2 7504 11368 7504 11368 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit17.Q
rlabel metal2 18200 17584 18200 17584 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit18.Q
rlabel metal3 18928 17640 18928 17640 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit19.Q
rlabel metal2 16352 40152 16352 40152 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit2.Q
rlabel metal2 17192 17416 17192 17416 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit20.Q
rlabel metal2 18760 16688 18760 16688 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit21.Q
rlabel metal2 11144 10640 11144 10640 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit22.Q
rlabel metal2 11144 11592 11144 11592 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit23.Q
rlabel metal2 11928 11144 11928 11144 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit24.Q
rlabel metal2 21000 15456 21000 15456 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit25.Q
rlabel metal3 17640 16072 17640 16072 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit26.Q
rlabel metal2 20888 14168 20888 14168 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit27.Q
rlabel metal2 19656 13272 19656 13272 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit28.Q
rlabel metal2 7784 10528 7784 10528 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit29.Q
rlabel metal2 15512 39088 15512 39088 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit3.Q
rlabel metal3 8736 11480 8736 11480 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit30.Q
rlabel metal2 9016 11704 9016 11704 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit31.Q
rlabel metal3 19656 21672 19656 21672 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit4.Q
rlabel metal2 19096 21840 19096 21840 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit5.Q
rlabel metal2 19432 29176 19432 29176 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit6.Q
rlabel metal3 20328 21560 20328 21560 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit7.Q
rlabel metal2 16520 9632 16520 9632 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit8.Q
rlabel metal2 15624 7504 15624 7504 0 Inst_W_IO4_ConfigMem.Inst_frame0_bit9.Q
rlabel metal2 7448 25368 7448 25368 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit0.Q
rlabel metal2 8400 24696 8400 24696 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit1.Q
rlabel metal2 13888 19208 13888 19208 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit10.Q
rlabel metal3 12320 19320 12320 19320 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit11.Q
rlabel metal2 4984 29904 4984 29904 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit12.Q
rlabel metal2 3640 29512 3640 29512 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit13.Q
rlabel metal3 16016 30856 16016 30856 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit14.Q
rlabel metal2 8904 31640 8904 31640 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit15.Q
rlabel metal2 2856 23240 2856 23240 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit16.Q
rlabel metal2 4032 23352 4032 23352 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit17.Q
rlabel metal3 21616 24136 21616 24136 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit18.Q
rlabel metal2 22400 24696 22400 24696 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit19.Q
rlabel metal2 3136 34888 3136 34888 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit2.Q
rlabel metal2 10136 29792 10136 29792 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit20.Q
rlabel metal2 9800 28896 9800 28896 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit21.Q
rlabel metal2 21280 25704 21280 25704 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit22.Q
rlabel metal2 19936 26488 19936 26488 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit23.Q
rlabel metal2 9912 16184 9912 16184 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit24.Q
rlabel metal2 8232 16576 8232 16576 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit25.Q
rlabel metal2 16072 24976 16072 24976 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit26.Q
rlabel metal2 14896 24696 14896 24696 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit27.Q
rlabel metal2 2856 17696 2856 17696 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit28.Q
rlabel metal2 3304 20132 3304 20132 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit29.Q
rlabel metal2 4312 36008 4312 36008 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit3.Q
rlabel metal2 12936 30128 12936 30128 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit30.Q
rlabel metal3 14280 30128 14280 30128 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit31.Q
rlabel metal2 8176 38920 8176 38920 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit4.Q
rlabel metal2 9464 39872 9464 39872 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit5.Q
rlabel metal2 21000 31080 21000 31080 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit6.Q
rlabel metal3 20944 30968 20944 30968 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit7.Q
rlabel metal2 12824 16576 12824 16576 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit8.Q
rlabel metal2 16184 17136 16184 17136 0 Inst_W_IO4_ConfigMem.Inst_frame1_bit9.Q
rlabel metal2 7112 22624 7112 22624 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit0.Q
rlabel metal2 8120 22232 8120 22232 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit1.Q
rlabel metal2 14392 5880 14392 5880 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit10.Q
rlabel metal2 14952 5544 14952 5544 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit11.Q
rlabel metal2 2912 25480 2912 25480 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit12.Q
rlabel metal2 4200 25144 4200 25144 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit13.Q
rlabel metal2 1512 34776 1512 34776 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit14.Q
rlabel metal2 2912 34104 2912 34104 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit15.Q
rlabel metal3 6272 38248 6272 38248 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit16.Q
rlabel metal2 7000 39256 7000 39256 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit17.Q
rlabel metal2 20888 31080 20888 31080 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit18.Q
rlabel metal3 22456 30184 22456 30184 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit19.Q
rlabel metal2 14728 33208 14728 33208 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit2.Q
rlabel metal2 9072 26824 9072 26824 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit20.Q
rlabel metal2 10696 25984 10696 25984 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit21.Q
rlabel metal2 10808 21448 10808 21448 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit22.Q
rlabel metal2 12040 21840 12040 21840 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit23.Q
rlabel metal3 13832 15288 13832 15288 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit24.Q
rlabel metal2 16184 15568 16184 15568 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit25.Q
rlabel metal2 14616 19320 14616 19320 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit26.Q
rlabel metal2 12152 18760 12152 18760 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit27.Q
rlabel metal2 2800 32760 2800 32760 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit28.Q
rlabel metal2 3304 32536 3304 32536 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit29.Q
rlabel metal2 15904 41720 15904 41720 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit3.Q
rlabel metal3 6944 29624 6944 29624 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit30.Q
rlabel metal3 4872 31192 4872 31192 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit31.Q
rlabel metal3 10696 38696 10696 38696 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit4.Q
rlabel metal3 13216 38808 13216 38808 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit5.Q
rlabel metal2 17752 28504 17752 28504 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit6.Q
rlabel metal2 18984 27720 18984 27720 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit7.Q
rlabel metal2 9632 9240 9632 9240 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit8.Q
rlabel metal2 10864 7672 10864 7672 0 Inst_W_IO4_ConfigMem.Inst_frame2_bit9.Q
rlabel metal3 13552 27272 13552 27272 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit10.Q
rlabel metal2 15344 27272 15344 27272 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit11.Q
rlabel metal3 5040 19208 5040 19208 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit12.Q
rlabel metal2 6552 19936 6552 19936 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit13.Q
rlabel metal2 5208 16968 5208 16968 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit14.Q
rlabel metal2 6552 17808 6552 17808 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit15.Q
rlabel metal2 7336 20664 7336 20664 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit16.Q
rlabel metal2 8456 20328 8456 20328 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit17.Q
rlabel metal3 13496 21560 13496 21560 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit18.Q
rlabel metal3 16520 21560 16520 21560 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit19.Q
rlabel metal3 11536 28616 11536 28616 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit20.Q
rlabel metal2 13048 28336 13048 28336 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit21.Q
rlabel metal3 16688 23352 16688 23352 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit22.Q
rlabel metal2 18200 23240 18200 23240 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit23.Q
rlabel metal3 8960 13720 8960 13720 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit24.Q
rlabel metal2 10976 12376 10976 12376 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit25.Q
rlabel metal2 14168 12656 14168 12656 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit26.Q
rlabel metal2 13832 13384 13832 13384 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit27.Q
rlabel metal3 4368 27048 4368 27048 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit28.Q
rlabel metal2 3640 26768 3640 26768 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit29.Q
rlabel metal2 3304 16184 3304 16184 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit30.Q
rlabel metal2 2968 16968 2968 16968 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit31.Q
rlabel metal2 12936 31920 12936 31920 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit4.Q
rlabel metal2 11592 31808 11592 31808 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit5.Q
rlabel metal2 18984 34608 18984 34608 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit6.Q
rlabel metal2 19880 35560 19880 35560 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit7.Q
rlabel metal2 7672 19040 7672 19040 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit8.Q
rlabel metal2 12936 24584 12936 24584 0 Inst_W_IO4_ConfigMem.Inst_frame3_bit9.Q
rlabel metal2 12488 32032 12488 32032 0 Inst_W_IO4_switch_matrix.E1BEG0
rlabel metal2 19544 34552 19544 34552 0 Inst_W_IO4_switch_matrix.E1BEG1
rlabel metal2 12264 24304 12264 24304 0 Inst_W_IO4_switch_matrix.E1BEG2
rlabel metal3 14952 26264 14952 26264 0 Inst_W_IO4_switch_matrix.E1BEG3
rlabel metal2 5544 18592 5544 18592 0 Inst_W_IO4_switch_matrix.E2BEG0
rlabel metal3 7504 17752 7504 17752 0 Inst_W_IO4_switch_matrix.E2BEG1
rlabel metal3 8456 19880 8456 19880 0 Inst_W_IO4_switch_matrix.E2BEG2
rlabel metal2 15512 22680 15512 22680 0 Inst_W_IO4_switch_matrix.E2BEG3
rlabel metal3 12432 28840 12432 28840 0 Inst_W_IO4_switch_matrix.E2BEG4
rlabel metal2 17752 24304 17752 24304 0 Inst_W_IO4_switch_matrix.E2BEG5
rlabel metal2 10024 14056 10024 14056 0 Inst_W_IO4_switch_matrix.E2BEG6
rlabel metal2 15148 14504 15148 14504 0 Inst_W_IO4_switch_matrix.E2BEG7
rlabel metal3 4648 27272 4648 27272 0 Inst_W_IO4_switch_matrix.E2BEGb0
rlabel metal4 3416 17360 3416 17360 0 Inst_W_IO4_switch_matrix.E2BEGb1
rlabel metal2 7560 21728 7560 21728 0 Inst_W_IO4_switch_matrix.E2BEGb2
rlabel metal2 15456 29176 15456 29176 0 Inst_W_IO4_switch_matrix.E2BEGb3
rlabel metal3 13608 38696 13608 38696 0 Inst_W_IO4_switch_matrix.E2BEGb4
rlabel metal2 18536 27160 18536 27160 0 Inst_W_IO4_switch_matrix.E2BEGb5
rlabel metal2 10136 8288 10136 8288 0 Inst_W_IO4_switch_matrix.E2BEGb6
rlabel metal2 15400 5488 15400 5488 0 Inst_W_IO4_switch_matrix.E2BEGb7
rlabel metal2 4704 30408 4704 30408 0 Inst_W_IO4_switch_matrix.E6BEG0
rlabel metal2 16520 31304 16520 31304 0 Inst_W_IO4_switch_matrix.E6BEG1
rlabel metal2 9800 34440 9800 34440 0 Inst_W_IO4_switch_matrix.E6BEG10
rlabel metal2 16184 36848 16184 36848 0 Inst_W_IO4_switch_matrix.E6BEG11
rlabel metal2 1624 23576 1624 23576 0 Inst_W_IO4_switch_matrix.E6BEG2
rlabel metal2 21728 24584 21728 24584 0 Inst_W_IO4_switch_matrix.E6BEG3
rlabel metal2 11256 30968 11256 30968 0 Inst_W_IO4_switch_matrix.E6BEG4
rlabel metal2 20664 28280 20664 28280 0 Inst_W_IO4_switch_matrix.E6BEG5
rlabel metal2 10024 16352 10024 16352 0 Inst_W_IO4_switch_matrix.E6BEG6
rlabel metal3 16240 24584 16240 24584 0 Inst_W_IO4_switch_matrix.E6BEG7
rlabel metal3 2520 20888 2520 20888 0 Inst_W_IO4_switch_matrix.E6BEG8
rlabel metal2 13608 29848 13608 29848 0 Inst_W_IO4_switch_matrix.E6BEG9
rlabel metal3 4312 25704 4312 25704 0 Inst_W_IO4_switch_matrix.EE4BEG0
rlabel metal2 2128 33992 2128 33992 0 Inst_W_IO4_switch_matrix.EE4BEG1
rlabel metal3 7952 24584 7952 24584 0 Inst_W_IO4_switch_matrix.EE4BEG10
rlabel metal2 2632 35840 2632 35840 0 Inst_W_IO4_switch_matrix.EE4BEG11
rlabel metal2 9016 39144 9016 39144 0 Inst_W_IO4_switch_matrix.EE4BEG12
rlabel metal2 21672 31360 21672 31360 0 Inst_W_IO4_switch_matrix.EE4BEG13
rlabel metal2 15736 17192 15736 17192 0 Inst_W_IO4_switch_matrix.EE4BEG14
rlabel metal2 13496 20384 13496 20384 0 Inst_W_IO4_switch_matrix.EE4BEG15
rlabel metal2 7056 40152 7056 40152 0 Inst_W_IO4_switch_matrix.EE4BEG2
rlabel metal2 21280 31976 21280 31976 0 Inst_W_IO4_switch_matrix.EE4BEG3
rlabel metal2 10584 25368 10584 25368 0 Inst_W_IO4_switch_matrix.EE4BEG4
rlabel metal2 10976 23912 10976 23912 0 Inst_W_IO4_switch_matrix.EE4BEG5
rlabel metal2 15680 15176 15680 15176 0 Inst_W_IO4_switch_matrix.EE4BEG6
rlabel metal2 13832 21392 13832 21392 0 Inst_W_IO4_switch_matrix.EE4BEG7
rlabel metal2 3416 32984 3416 32984 0 Inst_W_IO4_switch_matrix.EE4BEG8
rlabel metal2 6048 30968 6048 30968 0 Inst_W_IO4_switch_matrix.EE4BEG9
rlabel metal2 728 350 728 350 0 UserCLK
rlabel metal2 13608 36008 13608 36008 0 UserCLK_regs
rlabel metal2 896 55944 896 55944 0 UserCLKo
rlabel metal3 23506 280 23506 280 0 W1END[0]
rlabel metal3 27202 728 27202 728 0 W1END[1]
rlabel metal3 28434 1176 28434 1176 0 W1END[2]
rlabel metal3 27818 1624 27818 1624 0 W1END[3]
rlabel metal3 26936 5824 26936 5824 0 W2END[0]
rlabel metal2 19544 7056 19544 7056 0 W2END[1]
rlabel metal3 18200 26600 18200 26600 0 W2END[2]
rlabel metal2 15400 23128 15400 23128 0 W2END[3]
rlabel metal3 19656 26488 19656 26488 0 W2END[4]
rlabel metal2 20776 20664 20776 20664 0 W2END[5]
rlabel metal2 1848 17362 1848 17362 0 W2END[6]
rlabel metal2 19544 20832 19544 20832 0 W2END[7]
rlabel metal3 26418 2072 26418 2072 0 W2MID[0]
rlabel metal3 25578 2520 25578 2520 0 W2MID[1]
rlabel metal3 24794 2968 24794 2968 0 W2MID[2]
rlabel metal2 15848 22176 15848 22176 0 W2MID[3]
rlabel metal2 16968 17080 16968 17080 0 W2MID[4]
rlabel metal3 23674 4312 23674 4312 0 W2MID[5]
rlabel metal3 27678 4760 27678 4760 0 W2MID[6]
rlabel metal2 15624 10976 15624 10976 0 W2MID[7]
rlabel metal3 27678 16408 27678 16408 0 W6END[0]
rlabel metal3 28322 20888 28322 20888 0 W6END[10]
rlabel metal2 20944 23800 20944 23800 0 W6END[11]
rlabel metal3 27678 16856 27678 16856 0 W6END[1]
rlabel metal3 27678 17304 27678 17304 0 W6END[2]
rlabel metal3 27678 17752 27678 17752 0 W6END[3]
rlabel metal2 2632 24976 2632 24976 0 W6END[4]
rlabel metal4 20776 19376 20776 19376 0 W6END[5]
rlabel metal3 27678 19096 27678 19096 0 W6END[6]
rlabel metal3 26810 19544 26810 19544 0 W6END[7]
rlabel metal3 28434 19992 28434 19992 0 W6END[8]
rlabel metal3 23800 20552 23800 20552 0 W6END[9]
rlabel metal2 15792 19768 15792 19768 0 WW4END[0]
rlabel metal2 16744 24136 16744 24136 0 WW4END[10]
rlabel metal4 24248 14560 24248 14560 0 WW4END[11]
rlabel metal3 27678 14616 27678 14616 0 WW4END[12]
rlabel metal2 24248 17304 24248 17304 0 WW4END[13]
rlabel metal2 2744 17584 2744 17584 0 WW4END[14]
rlabel metal3 16408 15736 16408 15736 0 WW4END[15]
rlabel metal3 27678 9688 27678 9688 0 WW4END[1]
rlabel metal2 18984 23856 18984 23856 0 WW4END[2]
rlabel metal3 25578 10584 25578 10584 0 WW4END[3]
rlabel metal2 16520 21504 16520 21504 0 WW4END[4]
rlabel metal3 27678 11480 27678 11480 0 WW4END[5]
rlabel metal2 25088 19208 25088 19208 0 WW4END[6]
rlabel metal3 7616 19208 7616 19208 0 WW4END[7]
rlabel metal3 27678 12824 27678 12824 0 WW4END[8]
rlabel metal3 27678 13272 27678 13272 0 WW4END[9]
rlabel metal2 18088 15960 18088 15960 0 _000_
rlabel metal2 9352 12040 9352 12040 0 _001_
rlabel metal2 16632 7728 16632 7728 0 _002_
rlabel metal2 15176 10024 15176 10024 0 _003_
rlabel metal2 15232 8232 15232 8232 0 _004_
rlabel metal2 3640 13832 3640 13832 0 _005_
rlabel metal3 12768 7672 12768 7672 0 _006_
rlabel metal2 8344 11648 8344 11648 0 _007_
rlabel metal2 17528 15904 17528 15904 0 _008_
rlabel metal2 19544 18032 19544 18032 0 _009_
rlabel metal2 17640 12208 17640 12208 0 _010_
rlabel metal2 19656 21672 19656 21672 0 _011_
rlabel metal2 15736 10472 15736 10472 0 _012_
rlabel metal3 16240 8232 16240 8232 0 _013_
rlabel metal2 16464 8008 16464 8008 0 _014_
rlabel metal3 17080 7672 17080 7672 0 _015_
rlabel metal2 17192 9968 17192 9968 0 _016_
rlabel metal2 15960 9016 15960 9016 0 _017_
rlabel metal2 17584 8344 17584 8344 0 _018_
rlabel metal2 7896 11536 7896 11536 0 _019_
rlabel metal2 7616 12600 7616 12600 0 _020_
rlabel metal3 6048 14280 6048 14280 0 _021_
rlabel metal2 7952 13160 7952 13160 0 _022_
rlabel metal2 7672 14896 7672 14896 0 _023_
rlabel metal3 7784 14840 7784 14840 0 _024_
rlabel metal3 8512 14504 8512 14504 0 _025_
rlabel metal2 12040 10808 12040 10808 0 _026_
rlabel metal2 12264 10416 12264 10416 0 _027_
rlabel metal2 12768 10024 12768 10024 0 _028_
rlabel metal2 13944 10304 13944 10304 0 _029_
rlabel metal2 10920 10752 10920 10752 0 _030_
rlabel metal2 10752 10472 10752 10472 0 _031_
rlabel metal3 12488 10360 12488 10360 0 _032_
rlabel metal3 8400 9800 8400 9800 0 _033_
rlabel metal2 7448 10304 7448 10304 0 _034_
rlabel metal2 7224 10864 7224 10864 0 _035_
rlabel metal3 8680 10584 8680 10584 0 _036_
rlabel metal3 8680 9128 8680 9128 0 _037_
rlabel metal3 9352 8456 9352 8456 0 _038_
rlabel metal3 8848 10360 8848 10360 0 _039_
rlabel metal2 20552 10976 20552 10976 0 _040_
rlabel metal3 20272 13496 20272 13496 0 _041_
rlabel metal2 20664 12600 20664 12600 0 _042_
rlabel metal2 20776 12488 20776 12488 0 _043_
rlabel metal3 20888 15176 20888 15176 0 _044_
rlabel metal2 19768 15260 19768 15260 0 _045_
rlabel metal2 16688 16072 16688 16072 0 _046_
rlabel metal2 18648 16352 18648 16352 0 _047_
rlabel metal2 17304 15736 17304 15736 0 _048_
rlabel metal2 17136 15624 17136 15624 0 _049_
rlabel metal3 20832 17080 20832 17080 0 _050_
rlabel metal2 18984 16576 18984 16576 0 _051_
rlabel metal2 19936 16296 19936 16296 0 _052_
rlabel metal2 19208 17136 19208 17136 0 _053_
rlabel metal2 17864 19096 17864 19096 0 _054_
rlabel metal2 18536 17248 18536 17248 0 _055_
rlabel metal3 18200 17752 18200 17752 0 _056_
rlabel metal2 18312 17136 18312 17136 0 _057_
rlabel metal3 18424 10024 18424 10024 0 _058_
rlabel metal2 17640 11200 17640 11200 0 _059_
rlabel metal2 18760 11536 18760 11536 0 _060_
rlabel metal2 18984 12376 18984 12376 0 _061_
rlabel metal2 18760 13832 18760 13832 0 _062_
rlabel metal2 18368 12376 18368 12376 0 _063_
rlabel metal2 16912 12152 16912 12152 0 _064_
rlabel metal3 17696 14728 17696 14728 0 _065_
rlabel metal3 17976 15176 17976 15176 0 _066_
rlabel metal2 17752 11984 17752 11984 0 _067_
rlabel metal2 20608 20104 20608 20104 0 _068_
rlabel metal3 21616 20104 21616 20104 0 _069_
rlabel metal2 19768 21056 19768 21056 0 _070_
rlabel metal2 19880 23128 19880 23128 0 _071_
rlabel metal2 20328 19656 20328 19656 0 _072_
rlabel metal3 20440 19992 20440 19992 0 _073_
rlabel metal3 18424 21000 18424 21000 0 _074_
rlabel metal2 17752 20440 17752 20440 0 _075_
rlabel metal3 18368 21560 18368 21560 0 _076_
rlabel metal3 20160 21336 20160 21336 0 _077_
rlabel metal2 14056 37296 14056 37296 0 clknet_0_UserCLK
rlabel metal2 14840 34048 14840 34048 0 clknet_0_UserCLK_regs
rlabel metal2 10584 38080 10584 38080 0 clknet_1_0__leaf_UserCLK
rlabel metal2 12600 32984 12600 32984 0 clknet_1_0__leaf_UserCLK_regs
rlabel metal3 9184 37240 9184 37240 0 clknet_1_1__leaf_UserCLK_regs
rlabel metal3 22792 18536 22792 18536 0 net1
rlabel metal2 2408 7560 2408 7560 0 net10
rlabel metal3 23184 52808 23184 52808 0 net100
rlabel metal3 23184 52248 23184 52248 0 net101
rlabel metal2 26488 40712 26488 40712 0 net102
rlabel metal2 26264 53592 26264 53592 0 net103
rlabel metal2 24696 52752 24696 52752 0 net104
rlabel metal2 26264 54152 26264 54152 0 net105
rlabel metal2 24696 53648 24696 53648 0 net106
rlabel metal2 26488 53368 26488 53368 0 net107
rlabel metal3 24024 55272 24024 55272 0 net108
rlabel metal3 22344 54152 22344 54152 0 net109
rlabel metal2 2296 10192 2296 10192 0 net11
rlabel metal2 22792 53032 22792 53032 0 net110
rlabel metal2 21560 54208 21560 54208 0 net111
rlabel metal4 3192 18760 3192 18760 0 net112
rlabel metal2 24920 43988 24920 43988 0 net113
rlabel metal2 23128 52696 23128 52696 0 net114
rlabel metal2 16296 6664 16296 6664 0 net115
rlabel metal2 12320 38920 12320 38920 0 net116
rlabel metal3 21616 46536 21616 46536 0 net117
rlabel metal2 24920 45192 24920 45192 0 net118
rlabel metal3 23016 47432 23016 47432 0 net119
rlabel metal2 2072 9408 2072 9408 0 net12
rlabel metal2 24528 46536 24528 46536 0 net120
rlabel metal3 21112 48104 21112 48104 0 net121
rlabel metal2 24696 47376 24696 47376 0 net122
rlabel metal3 5432 39704 5432 39704 0 net123
rlabel metal4 27384 29344 27384 29344 0 net124
rlabel metal3 19432 55272 19432 55272 0 net125
rlabel metal3 23072 6664 23072 6664 0 net126
rlabel metal2 27496 2128 27496 2128 0 net127
rlabel metal2 21896 52248 21896 52248 0 net128
rlabel metal3 17136 2072 17136 2072 0 net129
rlabel metal2 14392 16128 14392 16128 0 net13
rlabel metal3 22904 55720 22904 55720 0 net130
rlabel metal3 24528 55944 24528 55944 0 net131
rlabel metal2 24696 54320 24696 54320 0 net132
rlabel metal2 3080 5824 3080 5824 0 net133
rlabel metal2 2576 43680 2576 43680 0 net134
rlabel metal3 7728 55944 7728 55944 0 net135
rlabel metal3 4592 55272 4592 55272 0 net136
rlabel metal3 23688 17752 23688 17752 0 net137
rlabel metal4 27272 30296 27272 30296 0 net138
rlabel metal3 16408 54488 16408 54488 0 net139
rlabel metal3 8736 7448 8736 7448 0 net14
rlabel metal3 20580 40936 20580 40936 0 net140
rlabel metal3 16800 55720 16800 55720 0 net141
rlabel metal3 21112 41384 21112 41384 0 net142
rlabel metal2 1400 54824 1400 54824 0 net143
rlabel metal2 16744 9912 16744 9912 0 net144
rlabel metal2 2296 5992 2296 5992 0 net145
rlabel metal3 4200 13608 4200 13608 0 net15
rlabel metal2 3696 15848 3696 15848 0 net16
rlabel metal3 1960 11592 1960 11592 0 net17
rlabel metal2 5040 17304 5040 17304 0 net18
rlabel metal2 19768 9352 19768 9352 0 net19
rlabel metal2 17528 6160 17528 6160 0 net2
rlabel metal2 2184 7532 2184 7532 0 net20
rlabel metal4 2296 25424 2296 25424 0 net21
rlabel metal2 4312 24584 4312 24584 0 net22
rlabel metal2 4928 24696 4928 24696 0 net23
rlabel metal2 2016 25480 2016 25480 0 net24
rlabel metal2 25032 23632 25032 23632 0 net25
rlabel metal2 19992 25704 19992 25704 0 net26
rlabel metal3 20664 22680 20664 22680 0 net27
rlabel metal2 24696 24080 24696 24080 0 net28
rlabel metal2 16632 20776 16632 20776 0 net29
rlabel metal2 6888 15876 6888 15876 0 net3
rlabel metal2 24920 23968 24920 23968 0 net30
rlabel metal2 26264 23800 26264 23800 0 net31
rlabel metal2 16072 24248 16072 24248 0 net32
rlabel metal3 16520 24248 16520 24248 0 net33
rlabel metal2 18760 25144 18760 25144 0 net34
rlabel metal2 15960 16464 15960 16464 0 net35
rlabel metal3 16184 16072 16184 16072 0 net36
rlabel metal2 24360 27496 24360 27496 0 net37
rlabel metal2 23744 15512 23744 15512 0 net38
rlabel metal2 18424 22736 18424 22736 0 net39
rlabel metal2 2296 7728 2296 7728 0 net4
rlabel metal2 2072 26096 2072 26096 0 net40
rlabel metal2 1736 36848 1736 36848 0 net41
rlabel metal2 17304 32032 17304 32032 0 net42
rlabel metal3 8176 23240 8176 23240 0 net43
rlabel metal3 2072 35784 2072 35784 0 net44
rlabel metal2 2744 30912 2744 30912 0 net45
rlabel metal2 6104 22904 6104 22904 0 net46
rlabel metal3 1904 23240 1904 23240 0 net47
rlabel metal3 20104 25368 20104 25368 0 net48
rlabel metal2 2744 37128 2744 37128 0 net49
rlabel metal3 23688 13888 23688 13888 0 net5
rlabel metal3 1960 29512 1960 29512 0 net50
rlabel metal2 14560 20776 14560 20776 0 net51
rlabel metal2 23128 16324 23128 16324 0 net52
rlabel metal2 10584 9184 10584 9184 0 net53
rlabel metal2 18200 29344 18200 29344 0 net54
rlabel metal2 7784 39536 7784 39536 0 net55
rlabel metal2 3696 16968 3696 16968 0 net56
rlabel metal3 26096 27720 26096 27720 0 net57
rlabel metal3 21168 28616 21168 28616 0 net58
rlabel metal2 26264 29456 26264 29456 0 net59
rlabel metal2 17024 9240 17024 9240 0 net6
rlabel metal3 22680 28504 22680 28504 0 net60
rlabel metal2 21896 6944 21896 6944 0 net61
rlabel metal3 26096 20552 26096 20552 0 net62
rlabel metal2 24696 37744 24696 37744 0 net63
rlabel metal2 24696 42224 24696 42224 0 net64
rlabel metal2 26376 43624 26376 43624 0 net65
rlabel metal3 21952 39592 21952 39592 0 net66
rlabel metal3 784 23240 784 23240 0 net67
rlabel metal3 23632 35448 23632 35448 0 net68
rlabel metal3 23212 41160 23212 41160 0 net69
rlabel metal2 18704 12264 18704 12264 0 net7
rlabel metal3 23240 40376 23240 40376 0 net70
rlabel metal2 17080 40544 17080 40544 0 net71
rlabel metal2 24808 40656 24808 40656 0 net72
rlabel metal2 1288 21504 1288 21504 0 net73
rlabel metal2 14000 40824 14000 40824 0 net74
rlabel metal3 15624 26208 15624 26208 0 net75
rlabel metal4 18424 32200 18424 32200 0 net76
rlabel metal2 2016 36344 2016 36344 0 net77
rlabel metal3 19880 36736 19880 36736 0 net78
rlabel metal2 20776 35336 20776 35336 0 net79
rlabel metal2 3080 6776 3080 6776 0 net8
rlabel metal2 15176 19768 15176 19768 0 net80
rlabel metal3 25816 38696 25816 38696 0 net81
rlabel metal2 2520 34552 2520 34552 0 net82
rlabel metal2 24920 32648 24920 32648 0 net83
rlabel metal3 24192 32648 24192 32648 0 net84
rlabel metal3 25760 33992 25760 33992 0 net85
rlabel metal2 24696 33264 24696 33264 0 net86
rlabel metal3 22456 15848 22456 15848 0 net87
rlabel metal2 24696 33936 24696 33936 0 net88
rlabel metal2 26152 33992 26152 33992 0 net89
rlabel metal2 7784 6440 7784 6440 0 net9
rlabel metal2 24360 33208 24360 33208 0 net90
rlabel metal2 24920 41664 24920 41664 0 net91
rlabel metal2 26152 49000 26152 49000 0 net92
rlabel metal2 26600 49784 26600 49784 0 net93
rlabel metal3 2296 18424 2296 18424 0 net94
rlabel metal2 26264 50232 26264 50232 0 net95
rlabel metal3 19488 49672 19488 49672 0 net96
rlabel metal2 26264 47656 26264 47656 0 net97
rlabel metal2 24696 50512 24696 50512 0 net98
rlabel metal2 25928 49448 25928 49448 0 net99
<< properties >>
string FIXED_BBOX 0 0 28560 57456
<< end >>
