module S_WARMBOOT (BOOT_top,
    CONFIGURED_top,
    Co,
    RESET_top,
    SLOT_top0,
    SLOT_top1,
    SLOT_top2,
    SLOT_top3,
    UserCLK,
    UserCLKo,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N2BEG,
    N2BEGb,
    N4BEG,
    NN4BEG,
    S1END,
    S2END,
    S2MID,
    S4END,
    SS4END);
 output BOOT_top;
 input CONFIGURED_top;
 output Co;
 input RESET_top;
 output SLOT_top0;
 output SLOT_top1;
 output SLOT_top2;
 output SLOT_top3;
 input UserCLK;
 output UserCLKo;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 output [15:0] N4BEG;
 output [15:0] NN4BEG;
 input [3:0] S1END;
 input [7:0] S2END;
 input [7:0] S2MID;
 input [15:0] S4END;
 input [15:0] SS4END;

 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Inst_S_WARMBOOT_switch_matrix.N1BEG0 ;
 wire \Inst_S_WARMBOOT_switch_matrix.N1BEG1 ;
 wire \Inst_S_WARMBOOT_switch_matrix.N1BEG2 ;
 wire \Inst_S_WARMBOOT_switch_matrix.N1BEG3 ;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire net5;
 wire net6;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net166;

 gf180mcu_fd_sc_mcu7t5v0__inv_1 _043_ (.I(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit30.Q ),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _044_ (.I(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit31.Q ),
    .ZN(_010_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _045_ (.I(net1),
    .ZN(_011_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _046_ (.I(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit27.Q ),
    .ZN(_012_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _047_ (.I(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit28.Q ),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _048_ (.I(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit24.Q ),
    .ZN(_014_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _049_ (.I(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit25.Q ),
    .ZN(_015_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _050_ (.I(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit21.Q ),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _051_ (.I(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit22.Q ),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _052_ (.I(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit18.Q ),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _053_ (.I(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit19.Q ),
    .ZN(_019_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _054_ (.I0(net27),
    .I1(net39),
    .S(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit29.Q ),
    .Z(_020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _055_ (.A1(_009_),
    .A2(_020_),
    .ZN(_021_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _056_ (.I0(net31),
    .I1(net35),
    .S(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit29.Q ),
    .Z(_022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _057_ (.A1(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit30.Q ),
    .A2(_022_),
    .B(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit31.Q ),
    .ZN(_023_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _058_ (.I0(net43),
    .I1(net47),
    .S(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit29.Q ),
    .Z(_024_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _059_ (.I0(net51),
    .I1(net55),
    .S(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit29.Q ),
    .Z(_025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _060_ (.A1(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit30.Q ),
    .A2(_025_),
    .ZN(_026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _061_ (.A1(_009_),
    .A2(_024_),
    .B(_010_),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _062_ (.A1(_021_),
    .A2(_023_),
    .B1(_026_),
    .B2(_027_),
    .C(_011_),
    .ZN(net56));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _063_ (.I0(net43),
    .I1(net47),
    .S(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit26.Q ),
    .Z(_028_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _064_ (.I0(net51),
    .I1(net55),
    .S(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit26.Q ),
    .Z(_029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _065_ (.A1(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit27.Q ),
    .A2(_029_),
    .ZN(_030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _066_ (.A1(_012_),
    .A2(_028_),
    .B(_013_),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _067_ (.I0(net27),
    .I1(net39),
    .I2(net31),
    .I3(net35),
    .S0(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit26.Q ),
    .S1(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit27.Q ),
    .Z(_032_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _068_ (.A1(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit28.Q ),
    .A2(_032_),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _069_ (.A1(_030_),
    .A2(_031_),
    .B(_033_),
    .ZN(net164));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _070_ (.I0(net42),
    .I1(net46),
    .S(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit23.Q ),
    .Z(_034_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _071_ (.I0(net50),
    .I1(net54),
    .S(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit23.Q ),
    .Z(_035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _072_ (.A1(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit24.Q ),
    .A2(_035_),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _073_ (.A1(_014_),
    .A2(_034_),
    .B(_015_),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _074_ (.I0(net26),
    .I1(net38),
    .I2(net30),
    .I3(net34),
    .S0(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit23.Q ),
    .S1(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit24.Q ),
    .Z(_038_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _075_ (.A1(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit25.Q ),
    .A2(_038_),
    .ZN(_039_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _076_ (.A1(_036_),
    .A2(_037_),
    .B(_039_),
    .ZN(net163));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _077_ (.I0(net41),
    .I1(net45),
    .S(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit20.Q ),
    .Z(_040_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _078_ (.I0(net49),
    .I1(net53),
    .S(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit20.Q ),
    .Z(_041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _079_ (.A1(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit21.Q ),
    .A2(_041_),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _080_ (.A1(_016_),
    .A2(_040_),
    .B(_017_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _081_ (.I0(net25),
    .I1(net37),
    .I2(net29),
    .I3(net33),
    .S0(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit20.Q ),
    .S1(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit21.Q ),
    .Z(_001_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _082_ (.A1(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit22.Q ),
    .A2(_001_),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _083_ (.A1(_042_),
    .A2(_000_),
    .B(_002_),
    .ZN(net162));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _084_ (.I0(net40),
    .I1(net44),
    .S(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit17.Q ),
    .Z(_003_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _085_ (.I0(net48),
    .I1(net52),
    .S(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit17.Q ),
    .Z(_004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _086_ (.A1(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit18.Q ),
    .A2(_004_),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _087_ (.A1(_018_),
    .A2(_003_),
    .B(_019_),
    .ZN(_006_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _088_ (.I0(net24),
    .I1(net36),
    .I2(net28),
    .I3(net32),
    .S0(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit17.Q ),
    .S1(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit18.Q ),
    .Z(_007_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _089_ (.A1(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit19.Q ),
    .A2(_007_),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _090_ (.A1(_005_),
    .A2(_006_),
    .B(_008_),
    .ZN(net161));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _091_ (.I0(net24),
    .I1(net23),
    .S(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit16.Q ),
    .Z(\Inst_S_WARMBOOT_switch_matrix.N1BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _092_ (.I0(net25),
    .I1(net23),
    .S(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit15.Q ),
    .Z(\Inst_S_WARMBOOT_switch_matrix.N1BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _093_ (.I0(net26),
    .I1(net23),
    .S(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit14.Q ),
    .Z(\Inst_S_WARMBOOT_switch_matrix.N1BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _094_ (.I0(net27),
    .I1(net23),
    .S(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit13.Q ),
    .Z(\Inst_S_WARMBOOT_switch_matrix.N1BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _095_ (.D(net2),
    .E(net5),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _096_ (.D(net3),
    .E(net5),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _097_ (.D(net4),
    .E(net5),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _098_ (.D(net7),
    .E(net5),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _099_ (.D(net8),
    .E(net5),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _100_ (.D(net9),
    .E(net5),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _101_ (.D(net10),
    .E(net5),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _102_ (.D(net11),
    .E(net6),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _103_ (.D(net12),
    .E(net6),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _104_ (.D(net13),
    .E(net6),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _105_ (.D(net14),
    .E(net5),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _106_ (.D(net15),
    .E(net5),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _107_ (.D(net16),
    .E(net5),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _108_ (.D(net17),
    .E(net6),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _109_ (.D(net18),
    .E(net6),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _110_ (.D(net19),
    .E(net6),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _111_ (.D(net20),
    .E(net6),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _112_ (.D(net21),
    .E(net6),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _113_ (.D(net22),
    .E(net6),
    .Q(\Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _115_ (.I(FrameData[0]),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _116_ (.I(FrameData[1]),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _117_ (.I(FrameData[2]),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _118_ (.I(FrameData[3]),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _119_ (.I(FrameData[4]),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _120_ (.I(FrameData[5]),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _121_ (.I(FrameData[6]),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _122_ (.I(FrameData[7]),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _123_ (.I(FrameData[8]),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _124_ (.I(FrameData[9]),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _125_ (.I(FrameData[10]),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _126_ (.I(FrameData[11]),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _127_ (.I(FrameData[12]),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _128_ (.I(net2),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _129_ (.I(net3),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _130_ (.I(net4),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _131_ (.I(net7),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _132_ (.I(net8),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _133_ (.I(net9),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _134_ (.I(net10),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _135_ (.I(net11),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _136_ (.I(net12),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _137_ (.I(net13),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _138_ (.I(net14),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _139_ (.I(net15),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _140_ (.I(net16),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _141_ (.I(net17),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _142_ (.I(net18),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _143_ (.I(net19),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _144_ (.I(net20),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _145_ (.I(net21),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _146_ (.I(net22),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _147_ (.I(net6),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _148_ (.I(FrameStrobe[1]),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _149_ (.I(FrameStrobe[2]),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _150_ (.I(FrameStrobe[3]),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _151_ (.I(FrameStrobe[4]),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _152_ (.I(FrameStrobe[5]),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _153_ (.I(FrameStrobe[6]),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _154_ (.I(FrameStrobe[7]),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _155_ (.I(FrameStrobe[8]),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _156_ (.I(FrameStrobe[9]),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _157_ (.I(FrameStrobe[10]),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _158_ (.I(FrameStrobe[11]),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _159_ (.I(FrameStrobe[12]),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _160_ (.I(FrameStrobe[13]),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _161_ (.I(FrameStrobe[14]),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _162_ (.I(FrameStrobe[15]),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _163_ (.I(FrameStrobe[16]),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _164_ (.I(FrameStrobe[17]),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _165_ (.I(FrameStrobe[18]),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _166_ (.I(FrameStrobe[19]),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _167_ (.I(\Inst_S_WARMBOOT_switch_matrix.N1BEG0 ),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _168_ (.I(\Inst_S_WARMBOOT_switch_matrix.N1BEG1 ),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _169_ (.I(\Inst_S_WARMBOOT_switch_matrix.N1BEG2 ),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _170_ (.I(\Inst_S_WARMBOOT_switch_matrix.N1BEG3 ),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _171_ (.I(S2MID[7]),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _172_ (.I(S2MID[6]),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _173_ (.I(S2MID[5]),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _174_ (.I(S2MID[4]),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _175_ (.I(net39),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _176_ (.I(net38),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _177_ (.I(net37),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _178_ (.I(net36),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _179_ (.I(net35),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _180_ (.I(net34),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _181_ (.I(net33),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _182_ (.I(net32),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _183_ (.I(net31),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _184_ (.I(net30),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _185_ (.I(net29),
    .Z(net127));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _186_ (.I(net28),
    .Z(net128));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _187_ (.I(S4END[15]),
    .Z(net129));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _188_ (.I(S4END[14]),
    .Z(net136));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _189_ (.I(S4END[13]),
    .Z(net137));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _190_ (.I(S4END[12]),
    .Z(net138));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _191_ (.I(S4END[11]),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _192_ (.I(S4END[10]),
    .Z(net140));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _193_ (.I(S4END[9]),
    .Z(net141));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _194_ (.I(S4END[8]),
    .Z(net142));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _195_ (.I(net47),
    .Z(net143));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _196_ (.I(net46),
    .Z(net144));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _197_ (.I(net45),
    .Z(net130));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _198_ (.I(net44),
    .Z(net131));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _199_ (.I(net43),
    .Z(net132));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _200_ (.I(net42),
    .Z(net133));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _201_ (.I(net41),
    .Z(net134));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _202_ (.I(net40),
    .Z(net135));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _203_ (.I(SS4END[15]),
    .Z(net145));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _204_ (.I(SS4END[14]),
    .Z(net152));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _205_ (.I(SS4END[13]),
    .Z(net153));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _206_ (.I(SS4END[12]),
    .Z(net154));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _207_ (.I(SS4END[11]),
    .Z(net155));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _208_ (.I(SS4END[10]),
    .Z(net156));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _209_ (.I(SS4END[9]),
    .Z(net157));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _210_ (.I(SS4END[8]),
    .Z(net158));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _211_ (.I(net55),
    .Z(net159));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _212_ (.I(net54),
    .Z(net160));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _213_ (.I(net53),
    .Z(net146));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _214_ (.I(net52),
    .Z(net147));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _215_ (.I(net51),
    .Z(net148));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _216_ (.I(net50),
    .Z(net149));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _217_ (.I(net49),
    .Z(net150));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _218_ (.I(net48),
    .Z(net151));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _219_ (.I(UserCLK),
    .Z(net165));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_31 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_32 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_33 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_35 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_38 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_39 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_40 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_41 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_42 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_43 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_44 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_45 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_46 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_47 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_48 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_49 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_50 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_51 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_52 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_53 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_54 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_55 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_56 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_57 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_58 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_59 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_60 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_61 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_62 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_63 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_64 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_65 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_67 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_68 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_69 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_70 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_71 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_72 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_73 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_74 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_75 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_76 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_77 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_78 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_79 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_80 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_81 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_82 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_83 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_84 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_85 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_86 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_87 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_88 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_89 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_90 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_91 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_92 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_93 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_94 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_95 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_96 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_97 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_98 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_99 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_157 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout5 (.I(FrameStrobe[0]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout6 (.I(FrameStrobe[0]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input1 (.I(CONFIGURED_top),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input2 (.I(FrameData[13]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input3 (.I(FrameData[14]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input4 (.I(FrameData[15]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input5 (.I(FrameData[16]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input6 (.I(FrameData[17]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input7 (.I(FrameData[18]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input8 (.I(FrameData[19]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input9 (.I(FrameData[20]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input10 (.I(FrameData[21]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input11 (.I(FrameData[22]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input12 (.I(FrameData[23]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input13 (.I(FrameData[24]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input14 (.I(FrameData[25]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input15 (.I(FrameData[26]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input16 (.I(FrameData[27]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input17 (.I(FrameData[28]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input18 (.I(FrameData[29]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input19 (.I(FrameData[30]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input20 (.I(FrameData[31]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input21 (.I(RESET_top),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input22 (.I(S1END[0]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input23 (.I(S1END[1]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input24 (.I(S1END[2]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input25 (.I(S1END[3]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input26 (.I(S2END[0]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input27 (.I(S2END[1]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input28 (.I(S2END[2]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input29 (.I(S2END[3]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input30 (.I(S2END[4]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input31 (.I(S2END[5]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input32 (.I(S2END[6]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input33 (.I(S2END[7]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input34 (.I(S2MID[0]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input35 (.I(S2MID[1]),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input36 (.I(S2MID[2]),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input37 (.I(S2MID[3]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input38 (.I(S4END[0]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input39 (.I(S4END[1]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input40 (.I(S4END[2]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input41 (.I(S4END[3]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input42 (.I(S4END[4]),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input43 (.I(S4END[5]),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input44 (.I(S4END[6]),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input45 (.I(S4END[7]),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input46 (.I(SS4END[0]),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input47 (.I(SS4END[1]),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input48 (.I(SS4END[2]),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input49 (.I(SS4END[3]),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input50 (.I(SS4END[4]),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input51 (.I(SS4END[5]),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input52 (.I(SS4END[6]),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input53 (.I(SS4END[7]),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output54 (.I(net56),
    .Z(BOOT_top));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output55 (.I(net57),
    .Z(FrameData_O[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output56 (.I(net58),
    .Z(FrameData_O[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output57 (.I(net59),
    .Z(FrameData_O[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output58 (.I(net60),
    .Z(FrameData_O[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output59 (.I(net61),
    .Z(FrameData_O[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output60 (.I(net62),
    .Z(FrameData_O[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output61 (.I(net63),
    .Z(FrameData_O[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output62 (.I(net64),
    .Z(FrameData_O[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output63 (.I(net65),
    .Z(FrameData_O[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output64 (.I(net66),
    .Z(FrameData_O[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output65 (.I(net67),
    .Z(FrameData_O[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output66 (.I(net68),
    .Z(FrameData_O[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output67 (.I(net69),
    .Z(FrameData_O[20]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output68 (.I(net70),
    .Z(FrameData_O[21]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output69 (.I(net71),
    .Z(FrameData_O[22]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output70 (.I(net72),
    .Z(FrameData_O[23]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output71 (.I(net73),
    .Z(FrameData_O[24]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output72 (.I(net74),
    .Z(FrameData_O[25]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output73 (.I(net75),
    .Z(FrameData_O[26]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output74 (.I(net76),
    .Z(FrameData_O[27]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output75 (.I(net77),
    .Z(FrameData_O[28]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output76 (.I(net78),
    .Z(FrameData_O[29]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output77 (.I(net79),
    .Z(FrameData_O[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output78 (.I(net80),
    .Z(FrameData_O[30]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output79 (.I(net81),
    .Z(FrameData_O[31]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output80 (.I(net82),
    .Z(FrameData_O[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output81 (.I(net83),
    .Z(FrameData_O[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output82 (.I(net84),
    .Z(FrameData_O[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output83 (.I(net85),
    .Z(FrameData_O[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output84 (.I(net86),
    .Z(FrameData_O[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output85 (.I(net87),
    .Z(FrameData_O[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output86 (.I(net88),
    .Z(FrameData_O[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output87 (.I(net89),
    .Z(FrameStrobe_O[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output88 (.I(net90),
    .Z(FrameStrobe_O[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output89 (.I(net91),
    .Z(FrameStrobe_O[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output90 (.I(net92),
    .Z(FrameStrobe_O[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output91 (.I(net93),
    .Z(FrameStrobe_O[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output92 (.I(net94),
    .Z(FrameStrobe_O[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output93 (.I(net95),
    .Z(FrameStrobe_O[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output94 (.I(net96),
    .Z(FrameStrobe_O[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output95 (.I(net97),
    .Z(FrameStrobe_O[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output96 (.I(net98),
    .Z(FrameStrobe_O[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output97 (.I(net99),
    .Z(FrameStrobe_O[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output98 (.I(net100),
    .Z(FrameStrobe_O[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output99 (.I(net101),
    .Z(FrameStrobe_O[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output100 (.I(net102),
    .Z(FrameStrobe_O[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output101 (.I(net103),
    .Z(FrameStrobe_O[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output102 (.I(net104),
    .Z(FrameStrobe_O[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output103 (.I(net105),
    .Z(FrameStrobe_O[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output104 (.I(net106),
    .Z(FrameStrobe_O[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output105 (.I(net107),
    .Z(FrameStrobe_O[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output106 (.I(net108),
    .Z(FrameStrobe_O[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output107 (.I(net109),
    .Z(N1BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output108 (.I(net110),
    .Z(N1BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output109 (.I(net111),
    .Z(N1BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output110 (.I(net112),
    .Z(N1BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output111 (.I(net113),
    .Z(N2BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output112 (.I(net114),
    .Z(N2BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output113 (.I(net115),
    .Z(N2BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output114 (.I(net116),
    .Z(N2BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output115 (.I(net117),
    .Z(N2BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output116 (.I(net118),
    .Z(N2BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output117 (.I(net119),
    .Z(N2BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output118 (.I(net120),
    .Z(N2BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output119 (.I(net121),
    .Z(N2BEGb[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output120 (.I(net122),
    .Z(N2BEGb[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output121 (.I(net123),
    .Z(N2BEGb[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output122 (.I(net124),
    .Z(N2BEGb[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output123 (.I(net125),
    .Z(N2BEGb[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output124 (.I(net126),
    .Z(N2BEGb[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output125 (.I(net127),
    .Z(N2BEGb[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output126 (.I(net128),
    .Z(N2BEGb[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output127 (.I(net129),
    .Z(N4BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output128 (.I(net130),
    .Z(N4BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output129 (.I(net131),
    .Z(N4BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output130 (.I(net132),
    .Z(N4BEG[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output131 (.I(net133),
    .Z(N4BEG[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output132 (.I(net134),
    .Z(N4BEG[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output133 (.I(net135),
    .Z(N4BEG[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output134 (.I(net136),
    .Z(N4BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output135 (.I(net137),
    .Z(N4BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output136 (.I(net138),
    .Z(N4BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output137 (.I(net139),
    .Z(N4BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output138 (.I(net140),
    .Z(N4BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output139 (.I(net141),
    .Z(N4BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output140 (.I(net142),
    .Z(N4BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output141 (.I(net143),
    .Z(N4BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output142 (.I(net144),
    .Z(N4BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output143 (.I(net145),
    .Z(NN4BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output144 (.I(net146),
    .Z(NN4BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output145 (.I(net147),
    .Z(NN4BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output146 (.I(net148),
    .Z(NN4BEG[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output147 (.I(net149),
    .Z(NN4BEG[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output148 (.I(net150),
    .Z(NN4BEG[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output149 (.I(net151),
    .Z(NN4BEG[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output150 (.I(net152),
    .Z(NN4BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output151 (.I(net153),
    .Z(NN4BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output152 (.I(net154),
    .Z(NN4BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output153 (.I(net155),
    .Z(NN4BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output154 (.I(net156),
    .Z(NN4BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output155 (.I(net157),
    .Z(NN4BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output156 (.I(net158),
    .Z(NN4BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output157 (.I(net159),
    .Z(NN4BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output158 (.I(net160),
    .Z(NN4BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output159 (.I(net161),
    .Z(SLOT_top0));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output160 (.I(net162),
    .Z(SLOT_top1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output161 (.I(net163),
    .Z(SLOT_top2));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output162 (.I(net164),
    .Z(SLOT_top3));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output163 (.I(net165),
    .Z(UserCLKo));
 gf180mcu_fd_sc_mcu7t5v0__tiel S_WARMBOOT_164 (.ZN(net166));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_498 ();
 assign Co = net166;
endmodule
