magic
tech gf180mcuD
magscale 1 10
timestamp 1764324398
<< metal1 >>
rect 672 13354 56784 13388
rect 672 13302 4466 13354
rect 4518 13302 4570 13354
rect 4622 13302 4674 13354
rect 4726 13302 24466 13354
rect 24518 13302 24570 13354
rect 24622 13302 24674 13354
rect 24726 13302 44466 13354
rect 44518 13302 44570 13354
rect 44622 13302 44674 13354
rect 44726 13302 56784 13354
rect 672 13268 56784 13302
rect 2158 13186 2210 13198
rect 2158 13122 2210 13134
rect 3726 13186 3778 13198
rect 3726 13122 3778 13134
rect 5966 13186 6018 13198
rect 5966 13122 6018 13134
rect 7534 13186 7586 13198
rect 7534 13122 7586 13134
rect 9774 13186 9826 13198
rect 9774 13122 9826 13134
rect 11342 13186 11394 13198
rect 11342 13122 11394 13134
rect 17390 13186 17442 13198
rect 17390 13122 17442 13134
rect 18958 13186 19010 13198
rect 18958 13122 19010 13134
rect 22654 13186 22706 13198
rect 22654 13122 22706 13134
rect 26238 13186 26290 13198
rect 26238 13122 26290 13134
rect 27134 13186 27186 13198
rect 27134 13122 27186 13134
rect 27806 13186 27858 13198
rect 27806 13122 27858 13134
rect 28702 13186 28754 13198
rect 28702 13122 28754 13134
rect 30046 13186 30098 13198
rect 30046 13122 30098 13134
rect 31502 13186 31554 13198
rect 31502 13122 31554 13134
rect 34190 13186 34242 13198
rect 34190 13122 34242 13134
rect 35310 13186 35362 13198
rect 35310 13122 35362 13134
rect 36206 13186 36258 13198
rect 36206 13122 36258 13134
rect 37102 13186 37154 13198
rect 37102 13122 37154 13134
rect 37998 13186 38050 13198
rect 37998 13122 38050 13134
rect 40798 13186 40850 13198
rect 40798 13122 40850 13134
rect 41694 13186 41746 13198
rect 41694 13122 41746 13134
rect 42926 13186 42978 13198
rect 42926 13122 42978 13134
rect 43822 13186 43874 13198
rect 43822 13122 43874 13134
rect 48974 13186 49026 13198
rect 48974 13122 49026 13134
rect 51102 13186 51154 13198
rect 51102 13122 51154 13134
rect 54910 13186 54962 13198
rect 54910 13122 54962 13134
rect 33294 13074 33346 13086
rect 13346 13022 13358 13074
rect 13410 13022 13422 13074
rect 14914 13022 14926 13074
rect 14978 13022 14990 13074
rect 23874 13022 23886 13074
rect 23938 13022 23950 13074
rect 33294 13010 33346 13022
rect 41358 13074 41410 13086
rect 41358 13010 41410 13022
rect 43486 13074 43538 13086
rect 44930 13022 44942 13074
rect 44994 13022 45006 13074
rect 52882 13022 52894 13074
rect 52946 13022 52958 13074
rect 43486 13010 43538 13022
rect 32398 12962 32450 12974
rect 2706 12910 2718 12962
rect 2770 12910 2782 12962
rect 4274 12910 4286 12962
rect 4338 12910 4350 12962
rect 6514 12910 6526 12962
rect 6578 12910 6590 12962
rect 8082 12910 8094 12962
rect 8146 12910 8158 12962
rect 10210 12910 10222 12962
rect 10274 12910 10286 12962
rect 11890 12910 11902 12962
rect 11954 12910 11966 12962
rect 14130 12910 14142 12962
rect 14194 12910 14206 12962
rect 15698 12910 15710 12962
rect 15762 12910 15774 12962
rect 17826 12910 17838 12962
rect 17890 12910 17902 12962
rect 19282 12910 19294 12962
rect 19346 12910 19358 12962
rect 20514 12910 20526 12962
rect 20578 12910 20590 12962
rect 22082 12910 22094 12962
rect 22146 12910 22158 12962
rect 46834 12910 46846 12962
rect 46898 12910 46910 12962
rect 48402 12910 48414 12962
rect 48466 12910 48478 12962
rect 50642 12910 50654 12962
rect 50706 12910 50718 12962
rect 52322 12910 52334 12962
rect 52386 12910 52398 12962
rect 54338 12910 54350 12962
rect 54402 12910 54414 12962
rect 32398 12898 32450 12910
rect 21534 12850 21586 12862
rect 21534 12786 21586 12798
rect 24446 12850 24498 12862
rect 24446 12786 24498 12798
rect 25678 12850 25730 12862
rect 25678 12786 25730 12798
rect 26574 12850 26626 12862
rect 26574 12786 26626 12798
rect 28366 12850 28418 12862
rect 30606 12850 30658 12862
rect 32958 12850 33010 12862
rect 29138 12798 29150 12850
rect 29202 12798 29214 12850
rect 31938 12798 31950 12850
rect 32002 12798 32014 12850
rect 28366 12786 28418 12798
rect 30606 12786 30658 12798
rect 32958 12786 33010 12798
rect 33854 12850 33906 12862
rect 33854 12786 33906 12798
rect 34750 12850 34802 12862
rect 36766 12850 36818 12862
rect 35746 12798 35758 12850
rect 35810 12798 35822 12850
rect 34750 12786 34802 12798
rect 36766 12786 36818 12798
rect 37662 12850 37714 12862
rect 44382 12850 44434 12862
rect 38434 12798 38446 12850
rect 38498 12798 38510 12850
rect 42130 12798 42142 12850
rect 42194 12798 42206 12850
rect 37662 12786 37714 12798
rect 44382 12786 44434 12798
rect 45950 12850 46002 12862
rect 45950 12786 46002 12798
rect 47854 12850 47906 12862
rect 47854 12786 47906 12798
rect 672 12570 56784 12604
rect 672 12518 3806 12570
rect 3858 12518 3910 12570
rect 3962 12518 4014 12570
rect 4066 12518 23806 12570
rect 23858 12518 23910 12570
rect 23962 12518 24014 12570
rect 24066 12518 43806 12570
rect 43858 12518 43910 12570
rect 43962 12518 44014 12570
rect 44066 12518 56784 12570
rect 672 12484 56784 12518
rect 2270 12402 2322 12414
rect 2270 12338 2322 12350
rect 10110 12402 10162 12414
rect 10110 12338 10162 12350
rect 12014 12402 12066 12414
rect 12014 12338 12066 12350
rect 14814 12402 14866 12414
rect 14814 12338 14866 12350
rect 16382 12402 16434 12414
rect 16382 12338 16434 12350
rect 17950 12402 18002 12414
rect 17950 12338 18002 12350
rect 23550 12402 23602 12414
rect 23550 12338 23602 12350
rect 47966 12402 48018 12414
rect 47966 12338 48018 12350
rect 49086 12402 49138 12414
rect 49086 12338 49138 12350
rect 52558 12402 52610 12414
rect 52558 12338 52610 12350
rect 54126 12402 54178 12414
rect 54126 12338 54178 12350
rect 55694 12402 55746 12414
rect 55694 12338 55746 12350
rect 20862 12290 20914 12302
rect 27246 12290 27298 12302
rect 41358 12290 41410 12302
rect 3602 12238 3614 12290
rect 3666 12238 3678 12290
rect 5058 12238 5070 12290
rect 5122 12238 5134 12290
rect 8194 12238 8206 12290
rect 8258 12238 8270 12290
rect 19394 12238 19406 12290
rect 19458 12238 19470 12290
rect 22194 12238 22206 12290
rect 22258 12238 22270 12290
rect 31490 12238 31502 12290
rect 31554 12238 31566 12290
rect 33618 12238 33630 12290
rect 33682 12238 33694 12290
rect 34514 12238 34526 12290
rect 34578 12238 34590 12290
rect 44594 12238 44606 12290
rect 44658 12238 44670 12290
rect 20862 12226 20914 12238
rect 27246 12226 27298 12238
rect 41358 12226 41410 12238
rect 21422 12178 21474 12190
rect 30494 12178 30546 12190
rect 2818 12126 2830 12178
rect 2882 12126 2894 12178
rect 4386 12126 4398 12178
rect 4450 12126 4462 12178
rect 5394 12126 5406 12178
rect 5458 12126 5470 12178
rect 7298 12126 7310 12178
rect 7362 12126 7374 12178
rect 10434 12126 10446 12178
rect 10498 12126 10510 12178
rect 10994 12126 11006 12178
rect 11058 12126 11070 12178
rect 18386 12126 18398 12178
rect 18450 12126 18462 12178
rect 22978 12126 22990 12178
rect 23042 12126 23054 12178
rect 24546 12126 24558 12178
rect 24610 12126 24622 12178
rect 21422 12114 21474 12126
rect 30494 12114 30546 12126
rect 32286 12178 32338 12190
rect 32286 12114 32338 12126
rect 33182 12178 33234 12190
rect 33182 12114 33234 12126
rect 34078 12178 34130 12190
rect 34078 12114 34130 12126
rect 34974 12178 35026 12190
rect 34974 12114 35026 12126
rect 36878 12178 36930 12190
rect 44158 12178 44210 12190
rect 37762 12126 37774 12178
rect 37826 12126 37838 12178
rect 42690 12126 42702 12178
rect 42754 12126 42766 12178
rect 52210 12126 52222 12178
rect 52274 12126 52286 12178
rect 55234 12126 55246 12178
rect 55298 12126 55310 12178
rect 36878 12114 36930 12126
rect 44158 12114 44210 12126
rect 13806 12066 13858 12078
rect 25902 12066 25954 12078
rect 31054 12066 31106 12078
rect 9090 12014 9102 12066
rect 9154 12014 9166 12066
rect 15362 12014 15374 12066
rect 15426 12014 15438 12066
rect 16930 12014 16942 12066
rect 16994 12014 17006 12066
rect 20066 12014 20078 12066
rect 20130 12014 20142 12066
rect 26226 12014 26238 12066
rect 26290 12014 26302 12066
rect 13806 12002 13858 12014
rect 25902 12002 25954 12014
rect 31054 12002 31106 12014
rect 32846 12066 32898 12078
rect 32846 12002 32898 12014
rect 35534 12066 35586 12078
rect 35534 12002 35586 12014
rect 36318 12066 36370 12078
rect 36318 12002 36370 12014
rect 42254 12066 42306 12078
rect 42254 12002 42306 12014
rect 45614 12066 45666 12078
rect 45614 12002 45666 12014
rect 46510 12066 46562 12078
rect 50990 12066 51042 12078
rect 48514 12014 48526 12066
rect 48578 12014 48590 12066
rect 50082 12014 50094 12066
rect 50146 12014 50158 12066
rect 53554 12014 53566 12066
rect 53618 12014 53630 12066
rect 46510 12002 46562 12014
rect 50990 12002 51042 12014
rect 6974 11954 7026 11966
rect 6974 11890 7026 11902
rect 13246 11954 13298 11966
rect 13246 11890 13298 11902
rect 24894 11954 24946 11966
rect 24894 11890 24946 11902
rect 25342 11954 25394 11966
rect 25342 11890 25394 11902
rect 31950 11954 32002 11966
rect 39454 11954 39506 11966
rect 38322 11902 38334 11954
rect 38386 11902 38398 11954
rect 31950 11890 32002 11902
rect 39454 11890 39506 11902
rect 41918 11954 41970 11966
rect 41918 11890 41970 11902
rect 45054 11954 45106 11966
rect 45054 11890 45106 11902
rect 45950 11954 46002 11966
rect 45950 11890 46002 11902
rect 50430 11954 50482 11966
rect 50430 11890 50482 11902
rect 672 11786 56784 11820
rect 672 11734 4466 11786
rect 4518 11734 4570 11786
rect 4622 11734 4674 11786
rect 4726 11734 24466 11786
rect 24518 11734 24570 11786
rect 24622 11734 24674 11786
rect 24726 11734 44466 11786
rect 44518 11734 44570 11786
rect 44622 11734 44674 11786
rect 44726 11734 56784 11786
rect 672 11700 56784 11734
rect 4622 11618 4674 11630
rect 4622 11554 4674 11566
rect 6190 11618 6242 11630
rect 6190 11554 6242 11566
rect 7758 11618 7810 11630
rect 7758 11554 7810 11566
rect 10894 11618 10946 11630
rect 10894 11554 10946 11566
rect 14030 11618 14082 11630
rect 14030 11554 14082 11566
rect 17502 11618 17554 11630
rect 17502 11554 17554 11566
rect 19070 11618 19122 11630
rect 19070 11554 19122 11566
rect 25678 11618 25730 11630
rect 25678 11554 25730 11566
rect 27582 11618 27634 11630
rect 27582 11554 27634 11566
rect 32398 11618 32450 11630
rect 32398 11554 32450 11566
rect 36430 11618 36482 11630
rect 36430 11554 36482 11566
rect 37326 11618 37378 11630
rect 37326 11554 37378 11566
rect 42590 11618 42642 11630
rect 42590 11554 42642 11566
rect 43486 11618 43538 11630
rect 43486 11554 43538 11566
rect 44382 11618 44434 11630
rect 44382 11554 44434 11566
rect 46958 11618 47010 11630
rect 46958 11554 47010 11566
rect 50318 11618 50370 11630
rect 50318 11554 50370 11566
rect 53454 11618 53506 11630
rect 53454 11554 53506 11566
rect 25118 11506 25170 11518
rect 44942 11506 44994 11518
rect 55022 11506 55074 11518
rect 20402 11454 20414 11506
rect 20466 11454 20478 11506
rect 21970 11454 21982 11506
rect 22034 11454 22046 11506
rect 34738 11454 34750 11506
rect 34802 11454 34814 11506
rect 42018 11454 42030 11506
rect 42082 11454 42094 11506
rect 52098 11454 52110 11506
rect 52162 11454 52174 11506
rect 25118 11442 25170 11454
rect 44942 11442 44994 11454
rect 55022 11442 55074 11454
rect 1038 11394 1090 11406
rect 9214 11394 9266 11406
rect 31278 11394 31330 11406
rect 38446 11394 38498 11406
rect 3602 11342 3614 11394
rect 3666 11342 3678 11394
rect 5170 11342 5182 11394
rect 5234 11342 5246 11394
rect 6626 11342 6638 11394
rect 6690 11342 6702 11394
rect 8194 11342 8206 11394
rect 8258 11342 8270 11394
rect 11442 11342 11454 11394
rect 11506 11342 11518 11394
rect 13010 11342 13022 11394
rect 13074 11342 13086 11394
rect 14466 11342 14478 11394
rect 14530 11342 14542 11394
rect 16034 11342 16046 11394
rect 16098 11342 16110 11394
rect 17826 11342 17838 11394
rect 17890 11342 17902 11394
rect 19618 11342 19630 11394
rect 19682 11342 19694 11394
rect 21186 11342 21198 11394
rect 21250 11342 21262 11394
rect 22754 11342 22766 11394
rect 22818 11342 22830 11394
rect 23538 11342 23550 11394
rect 23602 11342 23614 11394
rect 26002 11342 26014 11394
rect 26066 11342 26078 11394
rect 26226 11342 26238 11394
rect 26290 11342 26302 11394
rect 34402 11342 34414 11394
rect 34466 11342 34478 11394
rect 1038 11330 1090 11342
rect 9214 11330 9266 11342
rect 31278 11330 31330 11342
rect 38446 11330 38498 11342
rect 41246 11394 41298 11406
rect 44046 11394 44098 11406
rect 41794 11342 41806 11394
rect 41858 11342 41870 11394
rect 41246 11330 41298 11342
rect 44046 11330 44098 11342
rect 46622 11394 46674 11406
rect 54462 11394 54514 11406
rect 48178 11342 48190 11394
rect 48242 11342 48254 11394
rect 49746 11342 49758 11394
rect 49810 11342 49822 11394
rect 51314 11342 51326 11394
rect 51378 11342 51390 11394
rect 52882 11342 52894 11394
rect 52946 11342 52958 11394
rect 46622 11330 46674 11342
rect 54462 11330 54514 11342
rect 1598 11282 1650 11294
rect 1598 11218 1650 11230
rect 2606 11282 2658 11294
rect 2606 11218 2658 11230
rect 9774 11282 9826 11294
rect 23998 11282 24050 11294
rect 12338 11230 12350 11282
rect 12402 11230 12414 11282
rect 15474 11230 15486 11282
rect 15538 11230 15550 11282
rect 9774 11218 9826 11230
rect 23998 11218 24050 11230
rect 28142 11282 28194 11294
rect 28142 11218 28194 11230
rect 31838 11282 31890 11294
rect 39006 11282 39058 11294
rect 46062 11282 46114 11294
rect 32834 11230 32846 11282
rect 32898 11230 32910 11282
rect 36866 11230 36878 11282
rect 36930 11230 36942 11282
rect 37762 11230 37774 11282
rect 37826 11230 37838 11282
rect 43026 11230 43038 11282
rect 43090 11230 43102 11282
rect 31838 11218 31890 11230
rect 39006 11218 39058 11230
rect 46062 11218 46114 11230
rect 47518 11282 47570 11294
rect 47518 11218 47570 11230
rect 49198 11282 49250 11294
rect 49198 11218 49250 11230
rect 26574 11170 26626 11182
rect 26574 11106 26626 11118
rect 35982 11170 36034 11182
rect 35982 11106 36034 11118
rect 40910 11170 40962 11182
rect 40910 11106 40962 11118
rect 672 11002 56784 11036
rect 672 10950 3806 11002
rect 3858 10950 3910 11002
rect 3962 10950 4014 11002
rect 4066 10950 23806 11002
rect 23858 10950 23910 11002
rect 23962 10950 24014 11002
rect 24066 10950 43806 11002
rect 43858 10950 43910 11002
rect 43962 10950 44014 11002
rect 44066 10950 56784 11002
rect 672 10916 56784 10950
rect 3390 10834 3442 10846
rect 3390 10770 3442 10782
rect 6414 10834 6466 10846
rect 6414 10770 6466 10782
rect 7982 10834 8034 10846
rect 7982 10770 8034 10782
rect 14814 10834 14866 10846
rect 14814 10770 14866 10782
rect 41582 10834 41634 10846
rect 41582 10770 41634 10782
rect 49646 10834 49698 10846
rect 49646 10770 49698 10782
rect 50878 10834 50930 10846
rect 50878 10770 50930 10782
rect 52558 10834 52610 10846
rect 52558 10770 52610 10782
rect 5518 10722 5570 10734
rect 18286 10722 18338 10734
rect 2034 10670 2046 10722
rect 2098 10670 2110 10722
rect 16482 10670 16494 10722
rect 16546 10670 16558 10722
rect 5518 10658 5570 10670
rect 18286 10658 18338 10670
rect 19518 10722 19570 10734
rect 34974 10722 35026 10734
rect 21858 10670 21870 10722
rect 21922 10670 21934 10722
rect 23762 10670 23774 10722
rect 23826 10670 23838 10722
rect 25554 10670 25566 10722
rect 25618 10670 25630 10722
rect 26226 10670 26238 10722
rect 26290 10670 26302 10722
rect 19518 10658 19570 10670
rect 34974 10658 35026 10670
rect 54574 10722 54626 10734
rect 54574 10658 54626 10670
rect 56142 10722 56194 10734
rect 56142 10658 56194 10670
rect 20078 10610 20130 10622
rect 2818 10558 2830 10610
rect 2882 10558 2894 10610
rect 4386 10558 4398 10610
rect 4450 10558 4462 10610
rect 5058 10558 5070 10610
rect 5122 10558 5134 10610
rect 7410 10558 7422 10610
rect 7474 10558 7486 10610
rect 8978 10558 8990 10610
rect 9042 10558 9054 10610
rect 9538 10558 9550 10610
rect 9602 10558 9614 10610
rect 13458 10558 13470 10610
rect 13522 10558 13534 10610
rect 24658 10558 24670 10610
rect 24722 10558 24734 10610
rect 25218 10558 25230 10610
rect 25282 10558 25294 10610
rect 29922 10558 29934 10610
rect 29986 10558 29998 10610
rect 42242 10558 42254 10610
rect 42306 10558 42318 10610
rect 47282 10558 47294 10610
rect 47346 10558 47358 10610
rect 48738 10558 48750 10610
rect 48802 10558 48814 10610
rect 52098 10558 52110 10610
rect 52162 10558 52174 10610
rect 55122 10558 55134 10610
rect 55186 10558 55198 10610
rect 20078 10546 20130 10558
rect 12126 10498 12178 10510
rect 9874 10446 9886 10498
rect 9938 10446 9950 10498
rect 12126 10434 12178 10446
rect 13918 10498 13970 10510
rect 24222 10498 24274 10510
rect 40686 10498 40738 10510
rect 14242 10446 14254 10498
rect 14306 10446 14318 10498
rect 15810 10446 15822 10498
rect 15874 10446 15886 10498
rect 17714 10446 17726 10498
rect 17778 10446 17790 10498
rect 17938 10446 17950 10498
rect 18002 10446 18014 10498
rect 21074 10446 21086 10498
rect 21138 10446 21150 10498
rect 26674 10446 26686 10498
rect 26738 10446 26750 10498
rect 30370 10446 30382 10498
rect 30434 10446 30446 10498
rect 13918 10434 13970 10446
rect 24222 10434 24274 10446
rect 40686 10434 40738 10446
rect 40798 10498 40850 10510
rect 40798 10434 40850 10446
rect 41246 10498 41298 10510
rect 46846 10498 46898 10510
rect 42130 10446 42142 10498
rect 42194 10446 42206 10498
rect 41246 10434 41298 10446
rect 46846 10434 46898 10446
rect 47742 10498 47794 10510
rect 47742 10434 47794 10446
rect 48302 10498 48354 10510
rect 51426 10446 51438 10498
rect 51490 10446 51502 10498
rect 53554 10446 53566 10498
rect 53618 10446 53630 10498
rect 48302 10434 48354 10446
rect 11118 10386 11170 10398
rect 11118 10322 11170 10334
rect 11566 10386 11618 10398
rect 11566 10322 11618 10334
rect 18622 10386 18674 10398
rect 18622 10322 18674 10334
rect 23326 10386 23378 10398
rect 23326 10322 23378 10334
rect 27806 10386 27858 10398
rect 27806 10322 27858 10334
rect 31614 10386 31666 10398
rect 31614 10322 31666 10334
rect 34414 10386 34466 10398
rect 34414 10322 34466 10334
rect 40462 10386 40514 10398
rect 40462 10322 40514 10334
rect 672 10218 56784 10252
rect 672 10166 4466 10218
rect 4518 10166 4570 10218
rect 4622 10166 4674 10218
rect 4726 10166 24466 10218
rect 24518 10166 24570 10218
rect 24622 10166 24674 10218
rect 24726 10166 44466 10218
rect 44518 10166 44570 10218
rect 44622 10166 44674 10218
rect 44726 10166 56784 10218
rect 672 10132 56784 10166
rect 17950 10050 18002 10062
rect 17950 9986 18002 9998
rect 21086 10050 21138 10062
rect 21086 9986 21138 9998
rect 23998 10050 24050 10062
rect 23998 9986 24050 9998
rect 25118 10050 25170 10062
rect 25118 9986 25170 9998
rect 30046 10050 30098 10062
rect 30046 9986 30098 9998
rect 46398 10050 46450 10062
rect 46398 9986 46450 9998
rect 17390 9938 17442 9950
rect 2258 9886 2270 9938
rect 2322 9886 2334 9938
rect 5282 9886 5294 9938
rect 5346 9886 5358 9938
rect 17390 9874 17442 9886
rect 18846 9938 18898 9950
rect 18846 9874 18898 9886
rect 21534 9938 21586 9950
rect 46958 9938 47010 9950
rect 27570 9886 27582 9938
rect 27634 9886 27646 9938
rect 21534 9874 21586 9886
rect 46958 9874 47010 9886
rect 49086 9938 49138 9950
rect 50194 9886 50206 9938
rect 50258 9886 50270 9938
rect 49086 9874 49138 9886
rect 12910 9826 12962 9838
rect 18286 9826 18338 9838
rect 42590 9826 42642 9838
rect 3042 9774 3054 9826
rect 3106 9774 3118 9826
rect 7522 9774 7534 9826
rect 7586 9774 7598 9826
rect 10434 9774 10446 9826
rect 10498 9774 10510 9826
rect 12002 9774 12014 9826
rect 12066 9774 12078 9826
rect 15138 9774 15150 9826
rect 15202 9774 15214 9826
rect 20962 9774 20974 9826
rect 21026 9774 21038 9826
rect 21970 9774 21982 9826
rect 22034 9774 22046 9826
rect 27794 9774 27806 9826
rect 27858 9774 27870 9826
rect 12910 9762 12962 9774
rect 18286 9762 18338 9774
rect 42590 9762 42642 9774
rect 48526 9826 48578 9838
rect 49410 9774 49422 9826
rect 49474 9774 49486 9826
rect 50978 9774 50990 9826
rect 51042 9774 51054 9826
rect 52546 9774 52558 9826
rect 52610 9774 52622 9826
rect 54114 9774 54126 9826
rect 54178 9774 54190 9826
rect 48526 9762 48578 9774
rect 4286 9714 4338 9726
rect 9438 9714 9490 9726
rect 6850 9662 6862 9714
rect 6914 9662 6926 9714
rect 4286 9650 4338 9662
rect 9438 9650 9490 9662
rect 11006 9714 11058 9726
rect 14142 9714 14194 9726
rect 25678 9714 25730 9726
rect 13346 9662 13358 9714
rect 13410 9662 13422 9714
rect 20626 9662 20638 9714
rect 20690 9662 20702 9714
rect 23538 9662 23550 9714
rect 23602 9662 23614 9714
rect 11006 9650 11058 9662
rect 14142 9650 14194 9662
rect 25678 9650 25730 9662
rect 30606 9714 30658 9726
rect 30606 9650 30658 9662
rect 51998 9714 52050 9726
rect 51998 9650 52050 9662
rect 53566 9714 53618 9726
rect 53566 9650 53618 9662
rect 26686 9602 26738 9614
rect 26686 9538 26738 9550
rect 27022 9602 27074 9614
rect 27022 9538 27074 9550
rect 42478 9602 42530 9614
rect 42478 9538 42530 9550
rect 55134 9602 55186 9614
rect 55134 9538 55186 9550
rect 672 9434 56784 9468
rect 672 9382 3806 9434
rect 3858 9382 3910 9434
rect 3962 9382 4014 9434
rect 4066 9382 23806 9434
rect 23858 9382 23910 9434
rect 23962 9382 24014 9434
rect 24066 9382 43806 9434
rect 43858 9382 43910 9434
rect 43962 9382 44014 9434
rect 44066 9382 56784 9434
rect 672 9348 56784 9382
rect 2046 9266 2098 9278
rect 2046 9202 2098 9214
rect 53006 9266 53058 9278
rect 53006 9202 53058 9214
rect 18062 9154 18114 9166
rect 18062 9090 18114 9102
rect 20974 9154 21026 9166
rect 20974 9090 21026 9102
rect 36318 9154 36370 9166
rect 46062 9154 46114 9166
rect 41346 9102 41358 9154
rect 41410 9102 41422 9154
rect 51090 9102 51102 9154
rect 51154 9102 51166 9154
rect 36318 9090 36370 9102
rect 46062 9090 46114 9102
rect 3838 9042 3890 9054
rect 5854 9042 5906 9054
rect 11342 9042 11394 9054
rect 18622 9042 18674 9054
rect 22654 9042 22706 9054
rect 26686 9042 26738 9054
rect 5058 8990 5070 9042
rect 5122 8990 5134 9042
rect 9986 8990 9998 9042
rect 10050 8990 10062 9042
rect 12114 8990 12126 9042
rect 12178 8990 12190 9042
rect 13346 8990 13358 9042
rect 13410 8990 13422 9042
rect 21298 8990 21310 9042
rect 21362 8990 21374 9042
rect 21858 8990 21870 9042
rect 21922 8990 21934 9042
rect 23202 8990 23214 9042
rect 23266 8990 23278 9042
rect 24098 8990 24110 9042
rect 24162 8990 24174 9042
rect 3838 8978 3890 8990
rect 5854 8978 5906 8990
rect 11342 8978 11394 8990
rect 18622 8978 18674 8990
rect 22654 8978 22706 8990
rect 26686 8978 26738 8990
rect 31726 9042 31778 9054
rect 34974 9042 35026 9054
rect 39902 9042 39954 9054
rect 33282 8990 33294 9042
rect 33346 8990 33358 9042
rect 36754 8990 36766 9042
rect 36818 8990 36830 9042
rect 38546 8990 38558 9042
rect 38610 8990 38622 9042
rect 31726 8978 31778 8990
rect 34974 8978 35026 8990
rect 39902 8978 39954 8990
rect 40014 9042 40066 9054
rect 40014 8978 40066 8990
rect 40686 9042 40738 9054
rect 48414 9042 48466 9054
rect 41794 8990 41806 9042
rect 41858 8990 41870 9042
rect 42242 8990 42254 9042
rect 42306 8990 42318 9042
rect 43138 8990 43150 9042
rect 43202 8990 43214 9042
rect 45602 8990 45614 9042
rect 45666 8990 45678 9042
rect 40686 8978 40738 8990
rect 48414 8978 48466 8990
rect 48974 9042 49026 9054
rect 48974 8978 49026 8990
rect 49310 9042 49362 9054
rect 51986 8990 51998 9042
rect 52050 8990 52062 9042
rect 49310 8978 49362 8990
rect 3502 8930 3554 8942
rect 2594 8878 2606 8930
rect 2658 8878 2670 8930
rect 3502 8866 3554 8878
rect 4398 8930 4450 8942
rect 4398 8866 4450 8878
rect 5518 8930 5570 8942
rect 5518 8866 5570 8878
rect 6414 8930 6466 8942
rect 6414 8866 6466 8878
rect 10446 8930 10498 8942
rect 12910 8930 12962 8942
rect 12002 8878 12014 8930
rect 12066 8878 12078 8930
rect 10446 8866 10498 8878
rect 12910 8866 12962 8878
rect 27246 8930 27298 8942
rect 38110 8930 38162 8942
rect 31938 8878 31950 8930
rect 32002 8878 32014 8930
rect 32498 8878 32510 8930
rect 32562 8878 32574 8930
rect 27246 8866 27298 8878
rect 38110 8866 38162 8878
rect 39566 8930 39618 8942
rect 49870 8930 49922 8942
rect 41458 8878 41470 8930
rect 41522 8878 41534 8930
rect 42466 8878 42478 8930
rect 42530 8878 42542 8930
rect 47730 8878 47742 8930
rect 47794 8878 47806 8930
rect 50194 8878 50206 8930
rect 50258 8878 50270 8930
rect 53554 8878 53566 8930
rect 53618 8878 53630 8930
rect 54338 8878 54350 8930
rect 54402 8878 54414 8930
rect 55122 8878 55134 8930
rect 55186 8878 55198 8930
rect 55906 8878 55918 8930
rect 55970 8878 55982 8930
rect 39566 8866 39618 8878
rect 49870 8866 49922 8878
rect 2942 8818 2994 8830
rect 2942 8754 2994 8766
rect 11006 8818 11058 8830
rect 31390 8818 31442 8830
rect 39790 8818 39842 8830
rect 21970 8766 21982 8818
rect 22034 8766 22046 8818
rect 33842 8766 33854 8818
rect 33906 8766 33918 8818
rect 11006 8754 11058 8766
rect 31390 8754 31442 8766
rect 39790 8754 39842 8766
rect 40798 8818 40850 8830
rect 40798 8754 40850 8766
rect 48078 8818 48130 8830
rect 48078 8754 48130 8766
rect 672 8650 56784 8684
rect 672 8598 4466 8650
rect 4518 8598 4570 8650
rect 4622 8598 4674 8650
rect 4726 8598 24466 8650
rect 24518 8598 24570 8650
rect 24622 8598 24674 8650
rect 24726 8598 44466 8650
rect 44518 8598 44570 8650
rect 44622 8598 44674 8650
rect 44726 8598 56784 8650
rect 672 8564 56784 8598
rect 4062 8370 4114 8382
rect 14926 8370 14978 8382
rect 2258 8318 2270 8370
rect 2322 8318 2334 8370
rect 13794 8318 13806 8370
rect 13858 8318 13870 8370
rect 4062 8306 4114 8318
rect 14926 8306 14978 8318
rect 18398 8370 18450 8382
rect 18398 8306 18450 8318
rect 18510 8370 18562 8382
rect 18510 8306 18562 8318
rect 28030 8370 28082 8382
rect 28030 8306 28082 8318
rect 28926 8370 28978 8382
rect 28926 8306 28978 8318
rect 31166 8370 31218 8382
rect 31166 8306 31218 8318
rect 34078 8370 34130 8382
rect 36654 8370 36706 8382
rect 39006 8370 39058 8382
rect 35746 8318 35758 8370
rect 35810 8318 35822 8370
rect 36082 8318 36094 8370
rect 36146 8318 36158 8370
rect 37986 8318 37998 8370
rect 38050 8318 38062 8370
rect 34078 8306 34130 8318
rect 36654 8306 36706 8318
rect 39006 8306 39058 8318
rect 41134 8370 41186 8382
rect 41134 8306 41186 8318
rect 41582 8370 41634 8382
rect 41582 8306 41634 8318
rect 41918 8370 41970 8382
rect 41918 8306 41970 8318
rect 42142 8370 42194 8382
rect 42142 8306 42194 8318
rect 42254 8370 42306 8382
rect 42254 8306 42306 8318
rect 50318 8370 50370 8382
rect 51762 8318 51774 8370
rect 51826 8318 51838 8370
rect 53330 8318 53342 8370
rect 53394 8318 53406 8370
rect 50318 8306 50370 8318
rect 2606 8258 2658 8270
rect 2606 8194 2658 8206
rect 3166 8258 3218 8270
rect 3166 8194 3218 8206
rect 4398 8258 4450 8270
rect 4398 8194 4450 8206
rect 7758 8258 7810 8270
rect 18734 8258 18786 8270
rect 13570 8206 13582 8258
rect 13634 8206 13646 8258
rect 14466 8206 14478 8258
rect 14530 8206 14542 8258
rect 7758 8194 7810 8206
rect 18734 8194 18786 8206
rect 19070 8258 19122 8270
rect 29486 8258 29538 8270
rect 35086 8258 35138 8270
rect 38670 8258 38722 8270
rect 28466 8206 28478 8258
rect 28530 8206 28542 8258
rect 31602 8206 31614 8258
rect 31666 8206 31678 8258
rect 33618 8206 33630 8258
rect 33682 8206 33694 8258
rect 37874 8206 37886 8258
rect 37938 8206 37950 8258
rect 19070 8194 19122 8206
rect 29486 8194 29538 8206
rect 35086 8194 35138 8206
rect 38670 8194 38722 8206
rect 40798 8258 40850 8270
rect 40798 8194 40850 8206
rect 41022 8258 41074 8270
rect 41022 8194 41074 8206
rect 41358 8258 41410 8270
rect 41358 8194 41410 8206
rect 49758 8258 49810 8270
rect 50978 8206 50990 8258
rect 51042 8206 51054 8258
rect 52546 8206 52558 8258
rect 52610 8206 52622 8258
rect 54114 8206 54126 8258
rect 54178 8206 54190 8258
rect 49758 8194 49810 8206
rect 1262 8146 1314 8158
rect 1262 8082 1314 8094
rect 3502 8146 3554 8158
rect 3502 8082 3554 8094
rect 4958 8146 5010 8158
rect 55134 8146 55186 8158
rect 8194 8094 8206 8146
rect 8258 8094 8270 8146
rect 34626 8094 34638 8146
rect 34690 8094 34702 8146
rect 4958 8082 5010 8094
rect 55134 8082 55186 8094
rect 12798 8034 12850 8046
rect 12798 7970 12850 7982
rect 13134 8034 13186 8046
rect 13134 7970 13186 7982
rect 18958 8034 19010 8046
rect 18958 7970 19010 7982
rect 36318 8034 36370 8046
rect 36318 7970 36370 7982
rect 41694 8034 41746 8046
rect 41694 7970 41746 7982
rect 672 7866 56784 7900
rect 672 7814 3806 7866
rect 3858 7814 3910 7866
rect 3962 7814 4014 7866
rect 4066 7814 23806 7866
rect 23858 7814 23910 7866
rect 23962 7814 24014 7866
rect 24066 7814 43806 7866
rect 43858 7814 43910 7866
rect 43962 7814 44014 7866
rect 44066 7814 56784 7866
rect 672 7780 56784 7814
rect 19966 7698 20018 7710
rect 19966 7634 20018 7646
rect 53006 7698 53058 7710
rect 53006 7634 53058 7646
rect 56142 7698 56194 7710
rect 56142 7634 56194 7646
rect 1598 7586 1650 7598
rect 14030 7586 14082 7598
rect 36318 7586 36370 7598
rect 3266 7534 3278 7586
rect 3330 7534 3342 7586
rect 16146 7534 16158 7586
rect 16210 7534 16222 7586
rect 19618 7534 19630 7586
rect 19682 7534 19694 7586
rect 1598 7522 1650 7534
rect 14030 7522 14082 7534
rect 36318 7522 36370 7534
rect 42590 7586 42642 7598
rect 42590 7522 42642 7534
rect 50542 7586 50594 7598
rect 50542 7522 50594 7534
rect 54574 7586 54626 7598
rect 54574 7522 54626 7534
rect 1038 7474 1090 7486
rect 1038 7410 1090 7422
rect 2830 7474 2882 7486
rect 2830 7410 2882 7422
rect 3726 7474 3778 7486
rect 12238 7474 12290 7486
rect 8306 7422 8318 7474
rect 8370 7422 8382 7474
rect 3726 7410 3778 7422
rect 12238 7410 12290 7422
rect 18622 7474 18674 7486
rect 18622 7410 18674 7422
rect 18958 7474 19010 7486
rect 18958 7410 19010 7422
rect 19294 7474 19346 7486
rect 19294 7410 19346 7422
rect 28926 7474 28978 7486
rect 37998 7474 38050 7486
rect 49982 7474 50034 7486
rect 36754 7422 36766 7474
rect 36818 7422 36830 7474
rect 37090 7422 37102 7474
rect 37154 7422 37166 7474
rect 38434 7422 38446 7474
rect 38498 7422 38510 7474
rect 39330 7422 39342 7474
rect 39394 7422 39406 7474
rect 43026 7422 43038 7474
rect 43090 7422 43102 7474
rect 28926 7410 28978 7422
rect 37998 7410 38050 7422
rect 49982 7410 50034 7422
rect 50878 7474 50930 7486
rect 52098 7422 52110 7474
rect 52162 7422 52174 7474
rect 55234 7422 55246 7474
rect 55298 7422 55310 7474
rect 50878 7410 50930 7422
rect 2494 7362 2546 7374
rect 2494 7298 2546 7310
rect 4286 7362 4338 7374
rect 17726 7362 17778 7374
rect 8642 7310 8654 7362
rect 8706 7310 8718 7362
rect 4286 7298 4338 7310
rect 17726 7298 17778 7310
rect 18286 7362 18338 7374
rect 18286 7298 18338 7310
rect 19742 7362 19794 7374
rect 51438 7362 51490 7374
rect 29138 7310 29150 7362
rect 29202 7310 29214 7362
rect 29474 7310 29486 7362
rect 29538 7310 29550 7362
rect 53554 7310 53566 7362
rect 53618 7310 53630 7362
rect 19742 7298 19794 7310
rect 51438 7298 51490 7310
rect 1934 7250 1986 7262
rect 1934 7186 1986 7198
rect 9886 7250 9938 7262
rect 9886 7186 9938 7198
rect 11902 7250 11954 7262
rect 11902 7186 11954 7198
rect 12126 7250 12178 7262
rect 12126 7186 12178 7198
rect 13470 7250 13522 7262
rect 18398 7250 18450 7262
rect 16594 7198 16606 7250
rect 16658 7198 16670 7250
rect 13470 7186 13522 7198
rect 18398 7186 18450 7198
rect 18846 7250 18898 7262
rect 18846 7186 18898 7198
rect 28590 7250 28642 7262
rect 37314 7198 37326 7250
rect 37378 7198 37390 7250
rect 28590 7186 28642 7198
rect 672 7082 56784 7116
rect 672 7030 4466 7082
rect 4518 7030 4570 7082
rect 4622 7030 4674 7082
rect 4726 7030 24466 7082
rect 24518 7030 24570 7082
rect 24622 7030 24674 7082
rect 24726 7030 44466 7082
rect 44518 7030 44570 7082
rect 44622 7030 44674 7082
rect 44726 7030 56784 7082
rect 672 6996 56784 7030
rect 1038 6914 1090 6926
rect 1038 6850 1090 6862
rect 2830 6914 2882 6926
rect 2830 6850 2882 6862
rect 18622 6914 18674 6926
rect 18622 6850 18674 6862
rect 22878 6914 22930 6926
rect 22878 6850 22930 6862
rect 45838 6914 45890 6926
rect 45838 6850 45890 6862
rect 16718 6802 16770 6814
rect 16718 6738 16770 6750
rect 17278 6802 17330 6814
rect 17278 6738 17330 6750
rect 18734 6802 18786 6814
rect 41134 6802 41186 6814
rect 21634 6750 21646 6802
rect 21698 6750 21710 6802
rect 25106 6750 25118 6802
rect 25170 6750 25182 6802
rect 42018 6750 42030 6802
rect 42082 6750 42094 6802
rect 43362 6750 43374 6802
rect 43426 6750 43438 6802
rect 43698 6750 43710 6802
rect 43762 6750 43774 6802
rect 18734 6738 18786 6750
rect 41134 6738 41186 6750
rect 1934 6690 1986 6702
rect 1934 6626 1986 6638
rect 10558 6690 10610 6702
rect 10558 6626 10610 6638
rect 11006 6690 11058 6702
rect 11006 6626 11058 6638
rect 11118 6690 11170 6702
rect 11118 6626 11170 6638
rect 11230 6690 11282 6702
rect 11230 6626 11282 6638
rect 11566 6690 11618 6702
rect 11566 6626 11618 6638
rect 11790 6690 11842 6702
rect 11790 6626 11842 6638
rect 12126 6690 12178 6702
rect 12126 6626 12178 6638
rect 12350 6690 12402 6702
rect 12350 6626 12402 6638
rect 18286 6690 18338 6702
rect 18286 6626 18338 6638
rect 18846 6690 18898 6702
rect 26350 6690 26402 6702
rect 21298 6638 21310 6690
rect 21362 6638 21374 6690
rect 24770 6638 24782 6690
rect 24834 6638 24846 6690
rect 18846 6626 18898 6638
rect 26350 6626 26402 6638
rect 31278 6690 31330 6702
rect 31278 6626 31330 6638
rect 31838 6690 31890 6702
rect 42814 6690 42866 6702
rect 42242 6638 42254 6690
rect 42306 6638 42318 6690
rect 31838 6626 31890 6638
rect 42814 6626 42866 6638
rect 50542 6690 50594 6702
rect 50542 6626 50594 6638
rect 51102 6690 51154 6702
rect 51102 6626 51154 6638
rect 51438 6690 51490 6702
rect 52546 6638 52558 6690
rect 52610 6638 52622 6690
rect 54114 6638 54126 6690
rect 54178 6638 54190 6690
rect 51438 6626 51490 6638
rect 3390 6578 3442 6590
rect 1474 6526 1486 6578
rect 1538 6526 1550 6578
rect 2370 6526 2382 6578
rect 2434 6526 2446 6578
rect 3390 6514 3442 6526
rect 12014 6578 12066 6590
rect 53566 6578 53618 6590
rect 46274 6526 46286 6578
rect 46338 6526 46350 6578
rect 51874 6526 51886 6578
rect 51938 6526 51950 6578
rect 12014 6514 12066 6526
rect 53566 6514 53618 6526
rect 10670 6466 10722 6478
rect 10670 6402 10722 6414
rect 41470 6466 41522 6478
rect 41470 6402 41522 6414
rect 43150 6466 43202 6478
rect 43150 6402 43202 6414
rect 55134 6466 55186 6478
rect 55134 6402 55186 6414
rect 672 6298 56784 6332
rect 672 6246 3806 6298
rect 3858 6246 3910 6298
rect 3962 6246 4014 6298
rect 4066 6246 23806 6298
rect 23858 6246 23910 6298
rect 23962 6246 24014 6298
rect 24066 6246 43806 6298
rect 43858 6246 43910 6298
rect 43962 6246 44014 6298
rect 44066 6246 56784 6298
rect 672 6212 56784 6246
rect 9438 6130 9490 6142
rect 9438 6066 9490 6078
rect 11566 6130 11618 6142
rect 11566 6066 11618 6078
rect 27022 6130 27074 6142
rect 27022 6066 27074 6078
rect 32622 6130 32674 6142
rect 32622 6066 32674 6078
rect 32958 6130 33010 6142
rect 32958 6066 33010 6078
rect 37326 6130 37378 6142
rect 37326 6066 37378 6078
rect 53006 6130 53058 6142
rect 53006 6066 53058 6078
rect 56142 6130 56194 6142
rect 56142 6066 56194 6078
rect 1598 6018 1650 6030
rect 1598 5954 1650 5966
rect 7310 6018 7362 6030
rect 22206 6018 22258 6030
rect 25678 6018 25730 6030
rect 7858 5966 7870 6018
rect 7922 5966 7934 6018
rect 25106 5966 25118 6018
rect 25170 5966 25182 6018
rect 7310 5954 7362 5966
rect 22206 5954 22258 5966
rect 25678 5954 25730 5966
rect 28478 6018 28530 6030
rect 37214 6018 37266 6030
rect 30482 5966 30494 6018
rect 30546 5966 30558 6018
rect 28478 5954 28530 5966
rect 37214 5954 37266 5966
rect 38558 6018 38610 6030
rect 38558 5954 38610 5966
rect 41806 6018 41858 6030
rect 54574 6018 54626 6030
rect 49410 5966 49422 6018
rect 49474 5966 49486 6018
rect 41806 5954 41858 5966
rect 54574 5954 54626 5966
rect 1038 5906 1090 5918
rect 1038 5842 1090 5854
rect 1934 5906 1986 5918
rect 1934 5842 1986 5854
rect 6750 5906 6802 5918
rect 6750 5842 6802 5854
rect 11678 5906 11730 5918
rect 11678 5842 11730 5854
rect 21646 5906 21698 5918
rect 21646 5842 21698 5854
rect 26238 5906 26290 5918
rect 29038 5906 29090 5918
rect 27682 5854 27694 5906
rect 27746 5854 27758 5906
rect 26238 5842 26290 5854
rect 29038 5842 29090 5854
rect 38446 5906 38498 5918
rect 38446 5842 38498 5854
rect 38782 5906 38834 5918
rect 38782 5842 38834 5854
rect 39566 5906 39618 5918
rect 48974 5906 49026 5918
rect 42242 5854 42254 5906
rect 42306 5854 42318 5906
rect 52098 5854 52110 5906
rect 52162 5854 52174 5906
rect 53666 5854 53678 5906
rect 53730 5854 53742 5906
rect 39566 5842 39618 5854
rect 48974 5842 49026 5854
rect 2494 5794 2546 5806
rect 32062 5794 32114 5806
rect 38110 5794 38162 5806
rect 8194 5742 8206 5794
rect 8258 5742 8270 5794
rect 27794 5742 27806 5794
rect 27858 5742 27870 5794
rect 30818 5742 30830 5794
rect 30882 5742 30894 5794
rect 33170 5742 33182 5794
rect 33234 5742 33246 5794
rect 33618 5742 33630 5794
rect 33682 5742 33694 5794
rect 55122 5742 55134 5794
rect 55186 5742 55198 5794
rect 2494 5730 2546 5742
rect 32062 5730 32114 5742
rect 38110 5730 38162 5742
rect 24670 5682 24722 5694
rect 24670 5618 24722 5630
rect 26686 5682 26738 5694
rect 26686 5618 26738 5630
rect 37102 5682 37154 5694
rect 37102 5618 37154 5630
rect 39230 5682 39282 5694
rect 39230 5618 39282 5630
rect 39454 5682 39506 5694
rect 39454 5618 39506 5630
rect 672 5514 56784 5548
rect 672 5462 4466 5514
rect 4518 5462 4570 5514
rect 4622 5462 4674 5514
rect 4726 5462 24466 5514
rect 24518 5462 24570 5514
rect 24622 5462 24674 5514
rect 24726 5462 44466 5514
rect 44518 5462 44570 5514
rect 44622 5462 44674 5514
rect 44726 5462 56784 5514
rect 672 5428 56784 5462
rect 30942 5346 30994 5358
rect 30942 5282 30994 5294
rect 39454 5346 39506 5358
rect 39454 5282 39506 5294
rect 53230 5346 53282 5358
rect 53230 5282 53282 5294
rect 11902 5234 11954 5246
rect 11902 5170 11954 5182
rect 12462 5234 12514 5246
rect 21310 5234 21362 5246
rect 31502 5234 31554 5246
rect 13458 5182 13470 5234
rect 13522 5182 13534 5234
rect 22978 5182 22990 5234
rect 23042 5182 23054 5234
rect 23202 5182 23214 5234
rect 23266 5182 23278 5234
rect 34514 5182 34526 5234
rect 34578 5182 34590 5234
rect 12462 5170 12514 5182
rect 21310 5170 21362 5182
rect 31502 5170 31554 5182
rect 1598 5122 1650 5134
rect 14142 5122 14194 5134
rect 21870 5122 21922 5134
rect 1138 5070 1150 5122
rect 1202 5070 1214 5122
rect 2034 5070 2046 5122
rect 2098 5070 2110 5122
rect 12898 5070 12910 5122
rect 12962 5070 12974 5122
rect 13346 5070 13358 5122
rect 13410 5070 13422 5122
rect 14690 5070 14702 5122
rect 14754 5070 14766 5122
rect 15586 5070 15598 5122
rect 15650 5070 15662 5122
rect 1598 5058 1650 5070
rect 14142 5058 14194 5070
rect 21870 5058 21922 5070
rect 22318 5122 22370 5134
rect 22318 5058 22370 5070
rect 38670 5122 38722 5134
rect 38670 5058 38722 5070
rect 38782 5122 38834 5134
rect 38782 5058 38834 5070
rect 39118 5122 39170 5134
rect 39118 5058 39170 5070
rect 39454 5122 39506 5134
rect 39454 5058 39506 5070
rect 39790 5122 39842 5134
rect 39790 5058 39842 5070
rect 51998 5122 52050 5134
rect 54114 5070 54126 5122
rect 54178 5070 54190 5122
rect 54898 5070 54910 5122
rect 54962 5070 54974 5122
rect 51998 5058 52050 5070
rect 2494 5010 2546 5022
rect 12126 5010 12178 5022
rect 11890 4958 11902 5010
rect 11954 4958 11966 5010
rect 2494 4946 2546 4958
rect 12126 4946 12178 4958
rect 22654 5010 22706 5022
rect 34178 4958 34190 5010
rect 34242 4958 34254 5010
rect 52434 4958 52446 5010
rect 52498 4958 52510 5010
rect 53666 4958 53678 5010
rect 53730 4958 53742 5010
rect 22654 4946 22706 4958
rect 35758 4898 35810 4910
rect 35758 4834 35810 4846
rect 672 4730 56784 4764
rect 672 4678 3806 4730
rect 3858 4678 3910 4730
rect 3962 4678 4014 4730
rect 4066 4678 23806 4730
rect 23858 4678 23910 4730
rect 23962 4678 24014 4730
rect 24066 4678 43806 4730
rect 43858 4678 43910 4730
rect 43962 4678 44014 4730
rect 44066 4678 56784 4730
rect 672 4644 56784 4678
rect 10894 4562 10946 4574
rect 10894 4498 10946 4510
rect 17950 4562 18002 4574
rect 17950 4498 18002 4510
rect 22990 4562 23042 4574
rect 22990 4498 23042 4510
rect 39454 4562 39506 4574
rect 39454 4498 39506 4510
rect 54574 4562 54626 4574
rect 54574 4498 54626 4510
rect 56142 4562 56194 4574
rect 56142 4498 56194 4510
rect 13470 4450 13522 4462
rect 9314 4398 9326 4450
rect 9378 4398 9390 4450
rect 11778 4398 11790 4450
rect 11842 4398 11854 4450
rect 13470 4386 13522 4398
rect 15150 4450 15202 4462
rect 15150 4386 15202 4398
rect 34974 4450 35026 4462
rect 53106 4398 53118 4450
rect 53170 4398 53182 4450
rect 34974 4386 35026 4398
rect 1038 4338 1090 4350
rect 1038 4274 1090 4286
rect 12238 4338 12290 4350
rect 12238 4274 12290 4286
rect 14030 4338 14082 4350
rect 14030 4274 14082 4286
rect 18286 4338 18338 4350
rect 27582 4338 27634 4350
rect 21298 4286 21310 4338
rect 21362 4286 21374 4338
rect 18286 4274 18338 4286
rect 27582 4274 27634 4286
rect 28478 4338 28530 4350
rect 39566 4338 39618 4350
rect 34514 4286 34526 4338
rect 34578 4286 34590 4338
rect 28478 4274 28530 4286
rect 39566 4274 39618 4286
rect 44494 4338 44546 4350
rect 44494 4274 44546 4286
rect 45054 4338 45106 4350
rect 45054 4274 45106 4286
rect 49870 4338 49922 4350
rect 53554 4286 53566 4338
rect 53618 4286 53630 4338
rect 49870 4274 49922 4286
rect 1598 4226 1650 4238
rect 27022 4226 27074 4238
rect 9650 4174 9662 4226
rect 9714 4174 9726 4226
rect 18498 4174 18510 4226
rect 18562 4174 18574 4226
rect 19058 4174 19070 4226
rect 19122 4174 19134 4226
rect 21746 4174 21758 4226
rect 21810 4174 21822 4226
rect 1598 4162 1650 4174
rect 27022 4162 27074 4174
rect 27246 4226 27298 4238
rect 27246 4162 27298 4174
rect 50430 4226 50482 4238
rect 50430 4162 50482 4174
rect 52670 4226 52722 4238
rect 55122 4174 55134 4226
rect 55186 4174 55198 4226
rect 52670 4162 52722 4174
rect 15710 4114 15762 4126
rect 15710 4050 15762 4062
rect 27470 4114 27522 4126
rect 27470 4050 27522 4062
rect 28590 4114 28642 4126
rect 28590 4050 28642 4062
rect 28814 4114 28866 4126
rect 28814 4050 28866 4062
rect 34414 4114 34466 4126
rect 34414 4050 34466 4062
rect 672 3946 56784 3980
rect 672 3894 4466 3946
rect 4518 3894 4570 3946
rect 4622 3894 4674 3946
rect 4726 3894 24466 3946
rect 24518 3894 24570 3946
rect 24622 3894 24674 3946
rect 24726 3894 44466 3946
rect 44518 3894 44570 3946
rect 44622 3894 44674 3946
rect 44726 3894 56784 3946
rect 672 3860 56784 3894
rect 19630 3778 19682 3790
rect 19630 3714 19682 3726
rect 26910 3778 26962 3790
rect 26910 3714 26962 3726
rect 27246 3778 27298 3790
rect 27246 3714 27298 3726
rect 29710 3778 29762 3790
rect 37326 3778 37378 3790
rect 36194 3726 36206 3778
rect 36258 3726 36270 3778
rect 29710 3714 29762 3726
rect 37326 3714 37378 3726
rect 51662 3778 51714 3790
rect 51662 3714 51714 3726
rect 17950 3666 18002 3678
rect 17950 3602 18002 3614
rect 26798 3666 26850 3678
rect 26798 3602 26850 3614
rect 27358 3666 27410 3678
rect 52546 3614 52558 3666
rect 52610 3614 52622 3666
rect 54114 3614 54126 3666
rect 54178 3614 54190 3666
rect 54898 3614 54910 3666
rect 54962 3614 54974 3666
rect 27358 3602 27410 3614
rect 28590 3554 28642 3566
rect 9426 3502 9438 3554
rect 9490 3502 9502 3554
rect 18386 3502 18398 3554
rect 18450 3502 18462 3554
rect 28590 3490 28642 3502
rect 28926 3554 28978 3566
rect 28926 3490 28978 3502
rect 29262 3554 29314 3566
rect 52222 3554 52274 3566
rect 35746 3502 35758 3554
rect 35810 3502 35822 3554
rect 29262 3490 29314 3502
rect 52222 3490 52274 3502
rect 9886 3442 9938 3454
rect 28814 3442 28866 3454
rect 53566 3442 53618 3454
rect 19170 3390 19182 3442
rect 19234 3390 19246 3442
rect 29586 3390 29598 3442
rect 29650 3390 29662 3442
rect 9886 3378 9938 3390
rect 28814 3378 28866 3390
rect 53566 3378 53618 3390
rect 29934 3330 29986 3342
rect 29934 3266 29986 3278
rect 672 3162 56784 3196
rect 672 3110 3806 3162
rect 3858 3110 3910 3162
rect 3962 3110 4014 3162
rect 4066 3110 23806 3162
rect 23858 3110 23910 3162
rect 23962 3110 24014 3162
rect 24066 3110 43806 3162
rect 43858 3110 43910 3162
rect 43962 3110 44014 3162
rect 44066 3110 56784 3162
rect 672 3076 56784 3110
rect 26910 2994 26962 3006
rect 26910 2930 26962 2942
rect 38222 2994 38274 3006
rect 38222 2930 38274 2942
rect 54574 2994 54626 3006
rect 54574 2930 54626 2942
rect 56142 2994 56194 3006
rect 56142 2930 56194 2942
rect 28926 2882 28978 2894
rect 25330 2830 25342 2882
rect 25394 2830 25406 2882
rect 28926 2818 28978 2830
rect 41582 2882 41634 2894
rect 41582 2818 41634 2830
rect 48414 2882 48466 2894
rect 48414 2818 48466 2830
rect 30382 2770 30434 2782
rect 40574 2770 40626 2782
rect 21634 2718 21646 2770
rect 21698 2718 21710 2770
rect 29250 2718 29262 2770
rect 29314 2718 29326 2770
rect 29810 2718 29822 2770
rect 29874 2718 29886 2770
rect 30930 2718 30942 2770
rect 30994 2718 31006 2770
rect 31938 2718 31950 2770
rect 32002 2718 32014 2770
rect 35298 2718 35310 2770
rect 35362 2718 35374 2770
rect 36530 2718 36542 2770
rect 36594 2718 36606 2770
rect 30382 2706 30434 2718
rect 40574 2706 40626 2718
rect 47854 2770 47906 2782
rect 47854 2706 47906 2718
rect 50878 2770 50930 2782
rect 51986 2718 51998 2770
rect 52050 2718 52062 2770
rect 53554 2718 53566 2770
rect 53618 2718 53630 2770
rect 55346 2718 55358 2770
rect 55410 2718 55422 2770
rect 50878 2706 50930 2718
rect 22094 2658 22146 2670
rect 33070 2658 33122 2670
rect 25666 2606 25678 2658
rect 25730 2606 25742 2658
rect 29922 2606 29934 2658
rect 29986 2606 29998 2658
rect 22094 2594 22146 2606
rect 33070 2594 33122 2606
rect 35758 2658 35810 2670
rect 51438 2658 51490 2670
rect 36978 2606 36990 2658
rect 37042 2606 37054 2658
rect 52770 2606 52782 2658
rect 52834 2606 52846 2658
rect 35758 2594 35810 2606
rect 51438 2594 51490 2606
rect 32510 2546 32562 2558
rect 32510 2482 32562 2494
rect 40014 2546 40066 2558
rect 40014 2482 40066 2494
rect 42142 2546 42194 2558
rect 42142 2482 42194 2494
rect 672 2378 56784 2412
rect 672 2326 4466 2378
rect 4518 2326 4570 2378
rect 4622 2326 4674 2378
rect 4726 2326 24466 2378
rect 24518 2326 24570 2378
rect 24622 2326 24674 2378
rect 24726 2326 44466 2378
rect 44518 2326 44570 2378
rect 44622 2326 44674 2378
rect 44726 2326 56784 2378
rect 672 2292 56784 2326
rect 26350 2210 26402 2222
rect 26350 2146 26402 2158
rect 28702 2210 28754 2222
rect 28702 2146 28754 2158
rect 30158 2210 30210 2222
rect 30158 2146 30210 2158
rect 36654 2210 36706 2222
rect 36654 2146 36706 2158
rect 41134 2210 41186 2222
rect 49870 2210 49922 2222
rect 49074 2158 49086 2210
rect 49138 2158 49150 2210
rect 41134 2146 41186 2158
rect 49870 2146 49922 2158
rect 50766 2210 50818 2222
rect 50766 2146 50818 2158
rect 23998 2098 24050 2110
rect 28142 2098 28194 2110
rect 12898 2046 12910 2098
rect 12962 2046 12974 2098
rect 25106 2046 25118 2098
rect 25170 2046 25182 2098
rect 23998 2034 24050 2046
rect 28142 2034 28194 2046
rect 29598 2098 29650 2110
rect 29598 2034 29650 2046
rect 37214 2098 37266 2110
rect 37214 2034 37266 2046
rect 37886 2098 37938 2110
rect 37886 2034 37938 2046
rect 41694 2098 41746 2110
rect 41694 2034 41746 2046
rect 51326 2098 51378 2110
rect 51326 2034 51378 2046
rect 51662 2098 51714 2110
rect 51662 2034 51714 2046
rect 52222 2098 52274 2110
rect 52546 2046 52558 2098
rect 52610 2046 52622 2098
rect 54898 2046 54910 2098
rect 54962 2046 54974 2098
rect 52222 2034 52274 2046
rect 38446 1986 38498 1998
rect 23538 1934 23550 1986
rect 23602 1934 23614 1986
rect 24770 1934 24782 1986
rect 24834 1934 24846 1986
rect 47058 1934 47070 1986
rect 47122 1934 47134 1986
rect 49298 1934 49310 1986
rect 49362 1934 49374 1986
rect 54114 1934 54126 1986
rect 54178 1934 54190 1986
rect 38446 1922 38498 1934
rect 53566 1874 53618 1886
rect 47394 1822 47406 1874
rect 47458 1822 47470 1874
rect 50306 1822 50318 1874
rect 50370 1822 50382 1874
rect 53566 1810 53618 1822
rect 11902 1762 11954 1774
rect 11902 1698 11954 1710
rect 672 1594 56784 1628
rect 672 1542 3806 1594
rect 3858 1542 3910 1594
rect 3962 1542 4014 1594
rect 4066 1542 23806 1594
rect 23858 1542 23910 1594
rect 23962 1542 24014 1594
rect 24066 1542 43806 1594
rect 43858 1542 43910 1594
rect 43962 1542 44014 1594
rect 44066 1542 56784 1594
rect 672 1508 56784 1542
rect 53566 1426 53618 1438
rect 53566 1362 53618 1374
rect 56142 1426 56194 1438
rect 56142 1362 56194 1374
rect 4174 1314 4226 1326
rect 4174 1250 4226 1262
rect 5518 1314 5570 1326
rect 51998 1314 52050 1326
rect 7410 1262 7422 1314
rect 7474 1262 7486 1314
rect 5518 1250 5570 1262
rect 51998 1250 52050 1262
rect 6514 1150 6526 1202
rect 6578 1150 6590 1202
rect 10882 1150 10894 1202
rect 10946 1150 10958 1202
rect 14914 1150 14926 1202
rect 14978 1150 14990 1202
rect 25666 1150 25678 1202
rect 25730 1150 25742 1202
rect 50978 1150 50990 1202
rect 51042 1150 51054 1202
rect 52546 1150 52558 1202
rect 52610 1150 52622 1202
rect 55122 1150 55134 1202
rect 55186 1150 55198 1202
rect 2158 1090 2210 1102
rect 26126 1090 26178 1102
rect 8082 1038 8094 1090
rect 8146 1038 8158 1090
rect 10098 1038 10110 1090
rect 10162 1038 10174 1090
rect 14130 1038 14142 1090
rect 14194 1038 14206 1090
rect 2158 1026 2210 1038
rect 26126 1026 26178 1038
rect 1598 978 1650 990
rect 1598 914 1650 926
rect 3614 978 3666 990
rect 3614 914 3666 926
rect 672 810 56784 844
rect 672 758 4466 810
rect 4518 758 4570 810
rect 4622 758 4674 810
rect 4726 758 24466 810
rect 24518 758 24570 810
rect 24622 758 24674 810
rect 24726 758 44466 810
rect 44518 758 44570 810
rect 44622 758 44674 810
rect 44726 758 56784 810
rect 672 724 56784 758
<< via1 >>
rect 4466 13302 4518 13354
rect 4570 13302 4622 13354
rect 4674 13302 4726 13354
rect 24466 13302 24518 13354
rect 24570 13302 24622 13354
rect 24674 13302 24726 13354
rect 44466 13302 44518 13354
rect 44570 13302 44622 13354
rect 44674 13302 44726 13354
rect 2158 13134 2210 13186
rect 3726 13134 3778 13186
rect 5966 13134 6018 13186
rect 7534 13134 7586 13186
rect 9774 13134 9826 13186
rect 11342 13134 11394 13186
rect 17390 13134 17442 13186
rect 18958 13134 19010 13186
rect 22654 13134 22706 13186
rect 26238 13134 26290 13186
rect 27134 13134 27186 13186
rect 27806 13134 27858 13186
rect 28702 13134 28754 13186
rect 30046 13134 30098 13186
rect 31502 13134 31554 13186
rect 34190 13134 34242 13186
rect 35310 13134 35362 13186
rect 36206 13134 36258 13186
rect 37102 13134 37154 13186
rect 37998 13134 38050 13186
rect 40798 13134 40850 13186
rect 41694 13134 41746 13186
rect 42926 13134 42978 13186
rect 43822 13134 43874 13186
rect 48974 13134 49026 13186
rect 51102 13134 51154 13186
rect 54910 13134 54962 13186
rect 13358 13022 13410 13074
rect 14926 13022 14978 13074
rect 23886 13022 23938 13074
rect 33294 13022 33346 13074
rect 41358 13022 41410 13074
rect 43486 13022 43538 13074
rect 44942 13022 44994 13074
rect 52894 13022 52946 13074
rect 2718 12910 2770 12962
rect 4286 12910 4338 12962
rect 6526 12910 6578 12962
rect 8094 12910 8146 12962
rect 10222 12910 10274 12962
rect 11902 12910 11954 12962
rect 14142 12910 14194 12962
rect 15710 12910 15762 12962
rect 17838 12910 17890 12962
rect 19294 12910 19346 12962
rect 20526 12910 20578 12962
rect 22094 12910 22146 12962
rect 32398 12910 32450 12962
rect 46846 12910 46898 12962
rect 48414 12910 48466 12962
rect 50654 12910 50706 12962
rect 52334 12910 52386 12962
rect 54350 12910 54402 12962
rect 21534 12798 21586 12850
rect 24446 12798 24498 12850
rect 25678 12798 25730 12850
rect 26574 12798 26626 12850
rect 28366 12798 28418 12850
rect 29150 12798 29202 12850
rect 30606 12798 30658 12850
rect 31950 12798 32002 12850
rect 32958 12798 33010 12850
rect 33854 12798 33906 12850
rect 34750 12798 34802 12850
rect 35758 12798 35810 12850
rect 36766 12798 36818 12850
rect 37662 12798 37714 12850
rect 38446 12798 38498 12850
rect 42142 12798 42194 12850
rect 44382 12798 44434 12850
rect 45950 12798 46002 12850
rect 47854 12798 47906 12850
rect 3806 12518 3858 12570
rect 3910 12518 3962 12570
rect 4014 12518 4066 12570
rect 23806 12518 23858 12570
rect 23910 12518 23962 12570
rect 24014 12518 24066 12570
rect 43806 12518 43858 12570
rect 43910 12518 43962 12570
rect 44014 12518 44066 12570
rect 2270 12350 2322 12402
rect 10110 12350 10162 12402
rect 12014 12350 12066 12402
rect 14814 12350 14866 12402
rect 16382 12350 16434 12402
rect 17950 12350 18002 12402
rect 23550 12350 23602 12402
rect 47966 12350 48018 12402
rect 49086 12350 49138 12402
rect 52558 12350 52610 12402
rect 54126 12350 54178 12402
rect 55694 12350 55746 12402
rect 3614 12238 3666 12290
rect 5070 12238 5122 12290
rect 8206 12238 8258 12290
rect 19406 12238 19458 12290
rect 20862 12238 20914 12290
rect 22206 12238 22258 12290
rect 27246 12238 27298 12290
rect 31502 12238 31554 12290
rect 33630 12238 33682 12290
rect 34526 12238 34578 12290
rect 41358 12238 41410 12290
rect 44606 12238 44658 12290
rect 2830 12126 2882 12178
rect 4398 12126 4450 12178
rect 5406 12126 5458 12178
rect 7310 12126 7362 12178
rect 10446 12126 10498 12178
rect 11006 12126 11058 12178
rect 18398 12126 18450 12178
rect 21422 12126 21474 12178
rect 22990 12126 23042 12178
rect 24558 12126 24610 12178
rect 30494 12126 30546 12178
rect 32286 12126 32338 12178
rect 33182 12126 33234 12178
rect 34078 12126 34130 12178
rect 34974 12126 35026 12178
rect 36878 12126 36930 12178
rect 37774 12126 37826 12178
rect 42702 12126 42754 12178
rect 44158 12126 44210 12178
rect 52222 12126 52274 12178
rect 55246 12126 55298 12178
rect 9102 12014 9154 12066
rect 13806 12014 13858 12066
rect 15374 12014 15426 12066
rect 16942 12014 16994 12066
rect 20078 12014 20130 12066
rect 25902 12014 25954 12066
rect 26238 12014 26290 12066
rect 31054 12014 31106 12066
rect 32846 12014 32898 12066
rect 35534 12014 35586 12066
rect 36318 12014 36370 12066
rect 42254 12014 42306 12066
rect 45614 12014 45666 12066
rect 46510 12014 46562 12066
rect 48526 12014 48578 12066
rect 50094 12014 50146 12066
rect 50990 12014 51042 12066
rect 53566 12014 53618 12066
rect 6974 11902 7026 11954
rect 13246 11902 13298 11954
rect 24894 11902 24946 11954
rect 25342 11902 25394 11954
rect 31950 11902 32002 11954
rect 38334 11902 38386 11954
rect 39454 11902 39506 11954
rect 41918 11902 41970 11954
rect 45054 11902 45106 11954
rect 45950 11902 46002 11954
rect 50430 11902 50482 11954
rect 4466 11734 4518 11786
rect 4570 11734 4622 11786
rect 4674 11734 4726 11786
rect 24466 11734 24518 11786
rect 24570 11734 24622 11786
rect 24674 11734 24726 11786
rect 44466 11734 44518 11786
rect 44570 11734 44622 11786
rect 44674 11734 44726 11786
rect 4622 11566 4674 11618
rect 6190 11566 6242 11618
rect 7758 11566 7810 11618
rect 10894 11566 10946 11618
rect 14030 11566 14082 11618
rect 17502 11566 17554 11618
rect 19070 11566 19122 11618
rect 25678 11566 25730 11618
rect 27582 11566 27634 11618
rect 32398 11566 32450 11618
rect 36430 11566 36482 11618
rect 37326 11566 37378 11618
rect 42590 11566 42642 11618
rect 43486 11566 43538 11618
rect 44382 11566 44434 11618
rect 46958 11566 47010 11618
rect 50318 11566 50370 11618
rect 53454 11566 53506 11618
rect 20414 11454 20466 11506
rect 21982 11454 22034 11506
rect 25118 11454 25170 11506
rect 34750 11454 34802 11506
rect 42030 11454 42082 11506
rect 44942 11454 44994 11506
rect 52110 11454 52162 11506
rect 55022 11454 55074 11506
rect 1038 11342 1090 11394
rect 3614 11342 3666 11394
rect 5182 11342 5234 11394
rect 6638 11342 6690 11394
rect 8206 11342 8258 11394
rect 9214 11342 9266 11394
rect 11454 11342 11506 11394
rect 13022 11342 13074 11394
rect 14478 11342 14530 11394
rect 16046 11342 16098 11394
rect 17838 11342 17890 11394
rect 19630 11342 19682 11394
rect 21198 11342 21250 11394
rect 22766 11342 22818 11394
rect 23550 11342 23602 11394
rect 26014 11342 26066 11394
rect 26238 11342 26290 11394
rect 31278 11342 31330 11394
rect 34414 11342 34466 11394
rect 38446 11342 38498 11394
rect 41246 11342 41298 11394
rect 41806 11342 41858 11394
rect 44046 11342 44098 11394
rect 46622 11342 46674 11394
rect 48190 11342 48242 11394
rect 49758 11342 49810 11394
rect 51326 11342 51378 11394
rect 52894 11342 52946 11394
rect 54462 11342 54514 11394
rect 1598 11230 1650 11282
rect 2606 11230 2658 11282
rect 9774 11230 9826 11282
rect 12350 11230 12402 11282
rect 15486 11230 15538 11282
rect 23998 11230 24050 11282
rect 28142 11230 28194 11282
rect 31838 11230 31890 11282
rect 32846 11230 32898 11282
rect 36878 11230 36930 11282
rect 37774 11230 37826 11282
rect 39006 11230 39058 11282
rect 43038 11230 43090 11282
rect 46062 11230 46114 11282
rect 47518 11230 47570 11282
rect 49198 11230 49250 11282
rect 26574 11118 26626 11170
rect 35982 11118 36034 11170
rect 40910 11118 40962 11170
rect 3806 10950 3858 11002
rect 3910 10950 3962 11002
rect 4014 10950 4066 11002
rect 23806 10950 23858 11002
rect 23910 10950 23962 11002
rect 24014 10950 24066 11002
rect 43806 10950 43858 11002
rect 43910 10950 43962 11002
rect 44014 10950 44066 11002
rect 3390 10782 3442 10834
rect 6414 10782 6466 10834
rect 7982 10782 8034 10834
rect 14814 10782 14866 10834
rect 41582 10782 41634 10834
rect 49646 10782 49698 10834
rect 50878 10782 50930 10834
rect 52558 10782 52610 10834
rect 2046 10670 2098 10722
rect 5518 10670 5570 10722
rect 16494 10670 16546 10722
rect 18286 10670 18338 10722
rect 19518 10670 19570 10722
rect 21870 10670 21922 10722
rect 23774 10670 23826 10722
rect 25566 10670 25618 10722
rect 26238 10670 26290 10722
rect 34974 10670 35026 10722
rect 54574 10670 54626 10722
rect 56142 10670 56194 10722
rect 2830 10558 2882 10610
rect 4398 10558 4450 10610
rect 5070 10558 5122 10610
rect 7422 10558 7474 10610
rect 8990 10558 9042 10610
rect 9550 10558 9602 10610
rect 13470 10558 13522 10610
rect 20078 10558 20130 10610
rect 24670 10558 24722 10610
rect 25230 10558 25282 10610
rect 29934 10558 29986 10610
rect 42254 10558 42306 10610
rect 47294 10558 47346 10610
rect 48750 10558 48802 10610
rect 52110 10558 52162 10610
rect 55134 10558 55186 10610
rect 9886 10446 9938 10498
rect 12126 10446 12178 10498
rect 13918 10446 13970 10498
rect 14254 10446 14306 10498
rect 15822 10446 15874 10498
rect 17726 10446 17778 10498
rect 17950 10446 18002 10498
rect 21086 10446 21138 10498
rect 24222 10446 24274 10498
rect 26686 10446 26738 10498
rect 30382 10446 30434 10498
rect 40686 10446 40738 10498
rect 40798 10446 40850 10498
rect 41246 10446 41298 10498
rect 42142 10446 42194 10498
rect 46846 10446 46898 10498
rect 47742 10446 47794 10498
rect 48302 10446 48354 10498
rect 51438 10446 51490 10498
rect 53566 10446 53618 10498
rect 11118 10334 11170 10386
rect 11566 10334 11618 10386
rect 18622 10334 18674 10386
rect 23326 10334 23378 10386
rect 27806 10334 27858 10386
rect 31614 10334 31666 10386
rect 34414 10334 34466 10386
rect 40462 10334 40514 10386
rect 4466 10166 4518 10218
rect 4570 10166 4622 10218
rect 4674 10166 4726 10218
rect 24466 10166 24518 10218
rect 24570 10166 24622 10218
rect 24674 10166 24726 10218
rect 44466 10166 44518 10218
rect 44570 10166 44622 10218
rect 44674 10166 44726 10218
rect 17950 9998 18002 10050
rect 21086 9998 21138 10050
rect 23998 9998 24050 10050
rect 25118 9998 25170 10050
rect 30046 9998 30098 10050
rect 46398 9998 46450 10050
rect 2270 9886 2322 9938
rect 5294 9886 5346 9938
rect 17390 9886 17442 9938
rect 18846 9886 18898 9938
rect 21534 9886 21586 9938
rect 27582 9886 27634 9938
rect 46958 9886 47010 9938
rect 49086 9886 49138 9938
rect 50206 9886 50258 9938
rect 3054 9774 3106 9826
rect 7534 9774 7586 9826
rect 10446 9774 10498 9826
rect 12014 9774 12066 9826
rect 12910 9774 12962 9826
rect 15150 9774 15202 9826
rect 18286 9774 18338 9826
rect 20974 9774 21026 9826
rect 21982 9774 22034 9826
rect 27806 9774 27858 9826
rect 42590 9774 42642 9826
rect 48526 9774 48578 9826
rect 49422 9774 49474 9826
rect 50990 9774 51042 9826
rect 52558 9774 52610 9826
rect 54126 9774 54178 9826
rect 4286 9662 4338 9714
rect 6862 9662 6914 9714
rect 9438 9662 9490 9714
rect 11006 9662 11058 9714
rect 13358 9662 13410 9714
rect 14142 9662 14194 9714
rect 20638 9662 20690 9714
rect 23550 9662 23602 9714
rect 25678 9662 25730 9714
rect 30606 9662 30658 9714
rect 51998 9662 52050 9714
rect 53566 9662 53618 9714
rect 26686 9550 26738 9602
rect 27022 9550 27074 9602
rect 42478 9550 42530 9602
rect 55134 9550 55186 9602
rect 3806 9382 3858 9434
rect 3910 9382 3962 9434
rect 4014 9382 4066 9434
rect 23806 9382 23858 9434
rect 23910 9382 23962 9434
rect 24014 9382 24066 9434
rect 43806 9382 43858 9434
rect 43910 9382 43962 9434
rect 44014 9382 44066 9434
rect 2046 9214 2098 9266
rect 53006 9214 53058 9266
rect 18062 9102 18114 9154
rect 20974 9102 21026 9154
rect 36318 9102 36370 9154
rect 41358 9102 41410 9154
rect 46062 9102 46114 9154
rect 51102 9102 51154 9154
rect 3838 8990 3890 9042
rect 5070 8990 5122 9042
rect 5854 8990 5906 9042
rect 9998 8990 10050 9042
rect 11342 8990 11394 9042
rect 12126 8990 12178 9042
rect 13358 8990 13410 9042
rect 18622 8990 18674 9042
rect 21310 8990 21362 9042
rect 21870 8990 21922 9042
rect 22654 8990 22706 9042
rect 23214 8990 23266 9042
rect 24110 8990 24162 9042
rect 26686 8990 26738 9042
rect 31726 8990 31778 9042
rect 33294 8990 33346 9042
rect 34974 8990 35026 9042
rect 36766 8990 36818 9042
rect 38558 8990 38610 9042
rect 39902 8990 39954 9042
rect 40014 8990 40066 9042
rect 40686 8990 40738 9042
rect 41806 8990 41858 9042
rect 42254 8990 42306 9042
rect 43150 8990 43202 9042
rect 45614 8990 45666 9042
rect 48414 8990 48466 9042
rect 48974 8990 49026 9042
rect 49310 8990 49362 9042
rect 51998 8990 52050 9042
rect 2606 8878 2658 8930
rect 3502 8878 3554 8930
rect 4398 8878 4450 8930
rect 5518 8878 5570 8930
rect 6414 8878 6466 8930
rect 10446 8878 10498 8930
rect 12014 8878 12066 8930
rect 12910 8878 12962 8930
rect 27246 8878 27298 8930
rect 31950 8878 32002 8930
rect 32510 8878 32562 8930
rect 38110 8878 38162 8930
rect 39566 8878 39618 8930
rect 41470 8878 41522 8930
rect 42478 8878 42530 8930
rect 47742 8878 47794 8930
rect 49870 8878 49922 8930
rect 50206 8878 50258 8930
rect 53566 8878 53618 8930
rect 54350 8878 54402 8930
rect 55134 8878 55186 8930
rect 55918 8878 55970 8930
rect 2942 8766 2994 8818
rect 11006 8766 11058 8818
rect 21982 8766 22034 8818
rect 31390 8766 31442 8818
rect 33854 8766 33906 8818
rect 39790 8766 39842 8818
rect 40798 8766 40850 8818
rect 48078 8766 48130 8818
rect 4466 8598 4518 8650
rect 4570 8598 4622 8650
rect 4674 8598 4726 8650
rect 24466 8598 24518 8650
rect 24570 8598 24622 8650
rect 24674 8598 24726 8650
rect 44466 8598 44518 8650
rect 44570 8598 44622 8650
rect 44674 8598 44726 8650
rect 2270 8318 2322 8370
rect 4062 8318 4114 8370
rect 13806 8318 13858 8370
rect 14926 8318 14978 8370
rect 18398 8318 18450 8370
rect 18510 8318 18562 8370
rect 28030 8318 28082 8370
rect 28926 8318 28978 8370
rect 31166 8318 31218 8370
rect 34078 8318 34130 8370
rect 35758 8318 35810 8370
rect 36094 8318 36146 8370
rect 36654 8318 36706 8370
rect 37998 8318 38050 8370
rect 39006 8318 39058 8370
rect 41134 8318 41186 8370
rect 41582 8318 41634 8370
rect 41918 8318 41970 8370
rect 42142 8318 42194 8370
rect 42254 8318 42306 8370
rect 50318 8318 50370 8370
rect 51774 8318 51826 8370
rect 53342 8318 53394 8370
rect 2606 8206 2658 8258
rect 3166 8206 3218 8258
rect 4398 8206 4450 8258
rect 7758 8206 7810 8258
rect 13582 8206 13634 8258
rect 14478 8206 14530 8258
rect 18734 8206 18786 8258
rect 19070 8206 19122 8258
rect 28478 8206 28530 8258
rect 29486 8206 29538 8258
rect 31614 8206 31666 8258
rect 33630 8206 33682 8258
rect 35086 8206 35138 8258
rect 37886 8206 37938 8258
rect 38670 8206 38722 8258
rect 40798 8206 40850 8258
rect 41022 8206 41074 8258
rect 41358 8206 41410 8258
rect 49758 8206 49810 8258
rect 50990 8206 51042 8258
rect 52558 8206 52610 8258
rect 54126 8206 54178 8258
rect 1262 8094 1314 8146
rect 3502 8094 3554 8146
rect 4958 8094 5010 8146
rect 8206 8094 8258 8146
rect 34638 8094 34690 8146
rect 55134 8094 55186 8146
rect 12798 7982 12850 8034
rect 13134 7982 13186 8034
rect 18958 7982 19010 8034
rect 36318 7982 36370 8034
rect 41694 7982 41746 8034
rect 3806 7814 3858 7866
rect 3910 7814 3962 7866
rect 4014 7814 4066 7866
rect 23806 7814 23858 7866
rect 23910 7814 23962 7866
rect 24014 7814 24066 7866
rect 43806 7814 43858 7866
rect 43910 7814 43962 7866
rect 44014 7814 44066 7866
rect 19966 7646 20018 7698
rect 53006 7646 53058 7698
rect 56142 7646 56194 7698
rect 1598 7534 1650 7586
rect 3278 7534 3330 7586
rect 14030 7534 14082 7586
rect 16158 7534 16210 7586
rect 19630 7534 19682 7586
rect 36318 7534 36370 7586
rect 42590 7534 42642 7586
rect 50542 7534 50594 7586
rect 54574 7534 54626 7586
rect 1038 7422 1090 7474
rect 2830 7422 2882 7474
rect 3726 7422 3778 7474
rect 8318 7422 8370 7474
rect 12238 7422 12290 7474
rect 18622 7422 18674 7474
rect 18958 7422 19010 7474
rect 19294 7422 19346 7474
rect 28926 7422 28978 7474
rect 36766 7422 36818 7474
rect 37102 7422 37154 7474
rect 37998 7422 38050 7474
rect 38446 7422 38498 7474
rect 39342 7422 39394 7474
rect 43038 7422 43090 7474
rect 49982 7422 50034 7474
rect 50878 7422 50930 7474
rect 52110 7422 52162 7474
rect 55246 7422 55298 7474
rect 2494 7310 2546 7362
rect 4286 7310 4338 7362
rect 8654 7310 8706 7362
rect 17726 7310 17778 7362
rect 18286 7310 18338 7362
rect 19742 7310 19794 7362
rect 29150 7310 29202 7362
rect 29486 7310 29538 7362
rect 51438 7310 51490 7362
rect 53566 7310 53618 7362
rect 1934 7198 1986 7250
rect 9886 7198 9938 7250
rect 11902 7198 11954 7250
rect 12126 7198 12178 7250
rect 13470 7198 13522 7250
rect 16606 7198 16658 7250
rect 18398 7198 18450 7250
rect 18846 7198 18898 7250
rect 28590 7198 28642 7250
rect 37326 7198 37378 7250
rect 4466 7030 4518 7082
rect 4570 7030 4622 7082
rect 4674 7030 4726 7082
rect 24466 7030 24518 7082
rect 24570 7030 24622 7082
rect 24674 7030 24726 7082
rect 44466 7030 44518 7082
rect 44570 7030 44622 7082
rect 44674 7030 44726 7082
rect 1038 6862 1090 6914
rect 2830 6862 2882 6914
rect 18622 6862 18674 6914
rect 22878 6862 22930 6914
rect 45838 6862 45890 6914
rect 16718 6750 16770 6802
rect 17278 6750 17330 6802
rect 18734 6750 18786 6802
rect 21646 6750 21698 6802
rect 25118 6750 25170 6802
rect 41134 6750 41186 6802
rect 42030 6750 42082 6802
rect 43374 6750 43426 6802
rect 43710 6750 43762 6802
rect 1934 6638 1986 6690
rect 10558 6638 10610 6690
rect 11006 6638 11058 6690
rect 11118 6638 11170 6690
rect 11230 6638 11282 6690
rect 11566 6638 11618 6690
rect 11790 6638 11842 6690
rect 12126 6638 12178 6690
rect 12350 6638 12402 6690
rect 18286 6638 18338 6690
rect 18846 6638 18898 6690
rect 21310 6638 21362 6690
rect 24782 6638 24834 6690
rect 26350 6638 26402 6690
rect 31278 6638 31330 6690
rect 31838 6638 31890 6690
rect 42254 6638 42306 6690
rect 42814 6638 42866 6690
rect 50542 6638 50594 6690
rect 51102 6638 51154 6690
rect 51438 6638 51490 6690
rect 52558 6638 52610 6690
rect 54126 6638 54178 6690
rect 1486 6526 1538 6578
rect 2382 6526 2434 6578
rect 3390 6526 3442 6578
rect 12014 6526 12066 6578
rect 46286 6526 46338 6578
rect 51886 6526 51938 6578
rect 53566 6526 53618 6578
rect 10670 6414 10722 6466
rect 41470 6414 41522 6466
rect 43150 6414 43202 6466
rect 55134 6414 55186 6466
rect 3806 6246 3858 6298
rect 3910 6246 3962 6298
rect 4014 6246 4066 6298
rect 23806 6246 23858 6298
rect 23910 6246 23962 6298
rect 24014 6246 24066 6298
rect 43806 6246 43858 6298
rect 43910 6246 43962 6298
rect 44014 6246 44066 6298
rect 9438 6078 9490 6130
rect 11566 6078 11618 6130
rect 27022 6078 27074 6130
rect 32622 6078 32674 6130
rect 32958 6078 33010 6130
rect 37326 6078 37378 6130
rect 53006 6078 53058 6130
rect 56142 6078 56194 6130
rect 1598 5966 1650 6018
rect 7310 5966 7362 6018
rect 7870 5966 7922 6018
rect 22206 5966 22258 6018
rect 25118 5966 25170 6018
rect 25678 5966 25730 6018
rect 28478 5966 28530 6018
rect 30494 5966 30546 6018
rect 37214 5966 37266 6018
rect 38558 5966 38610 6018
rect 41806 5966 41858 6018
rect 49422 5966 49474 6018
rect 54574 5966 54626 6018
rect 1038 5854 1090 5906
rect 1934 5854 1986 5906
rect 6750 5854 6802 5906
rect 11678 5854 11730 5906
rect 21646 5854 21698 5906
rect 26238 5854 26290 5906
rect 27694 5854 27746 5906
rect 29038 5854 29090 5906
rect 38446 5854 38498 5906
rect 38782 5854 38834 5906
rect 39566 5854 39618 5906
rect 42254 5854 42306 5906
rect 48974 5854 49026 5906
rect 52110 5854 52162 5906
rect 53678 5854 53730 5906
rect 2494 5742 2546 5794
rect 8206 5742 8258 5794
rect 27806 5742 27858 5794
rect 30830 5742 30882 5794
rect 32062 5742 32114 5794
rect 33182 5742 33234 5794
rect 33630 5742 33682 5794
rect 38110 5742 38162 5794
rect 55134 5742 55186 5794
rect 24670 5630 24722 5682
rect 26686 5630 26738 5682
rect 37102 5630 37154 5682
rect 39230 5630 39282 5682
rect 39454 5630 39506 5682
rect 4466 5462 4518 5514
rect 4570 5462 4622 5514
rect 4674 5462 4726 5514
rect 24466 5462 24518 5514
rect 24570 5462 24622 5514
rect 24674 5462 24726 5514
rect 44466 5462 44518 5514
rect 44570 5462 44622 5514
rect 44674 5462 44726 5514
rect 30942 5294 30994 5346
rect 39454 5294 39506 5346
rect 53230 5294 53282 5346
rect 11902 5182 11954 5234
rect 12462 5182 12514 5234
rect 13470 5182 13522 5234
rect 21310 5182 21362 5234
rect 22990 5182 23042 5234
rect 23214 5182 23266 5234
rect 31502 5182 31554 5234
rect 34526 5182 34578 5234
rect 1150 5070 1202 5122
rect 1598 5070 1650 5122
rect 2046 5070 2098 5122
rect 12910 5070 12962 5122
rect 13358 5070 13410 5122
rect 14142 5070 14194 5122
rect 14702 5070 14754 5122
rect 15598 5070 15650 5122
rect 21870 5070 21922 5122
rect 22318 5070 22370 5122
rect 38670 5070 38722 5122
rect 38782 5070 38834 5122
rect 39118 5070 39170 5122
rect 39454 5070 39506 5122
rect 39790 5070 39842 5122
rect 51998 5070 52050 5122
rect 54126 5070 54178 5122
rect 54910 5070 54962 5122
rect 2494 4958 2546 5010
rect 11902 4958 11954 5010
rect 12126 4958 12178 5010
rect 22654 4958 22706 5010
rect 34190 4958 34242 5010
rect 52446 4958 52498 5010
rect 53678 4958 53730 5010
rect 35758 4846 35810 4898
rect 3806 4678 3858 4730
rect 3910 4678 3962 4730
rect 4014 4678 4066 4730
rect 23806 4678 23858 4730
rect 23910 4678 23962 4730
rect 24014 4678 24066 4730
rect 43806 4678 43858 4730
rect 43910 4678 43962 4730
rect 44014 4678 44066 4730
rect 10894 4510 10946 4562
rect 17950 4510 18002 4562
rect 22990 4510 23042 4562
rect 39454 4510 39506 4562
rect 54574 4510 54626 4562
rect 56142 4510 56194 4562
rect 9326 4398 9378 4450
rect 11790 4398 11842 4450
rect 13470 4398 13522 4450
rect 15150 4398 15202 4450
rect 34974 4398 35026 4450
rect 53118 4398 53170 4450
rect 1038 4286 1090 4338
rect 12238 4286 12290 4338
rect 14030 4286 14082 4338
rect 18286 4286 18338 4338
rect 21310 4286 21362 4338
rect 27582 4286 27634 4338
rect 28478 4286 28530 4338
rect 34526 4286 34578 4338
rect 39566 4286 39618 4338
rect 44494 4286 44546 4338
rect 45054 4286 45106 4338
rect 49870 4286 49922 4338
rect 53566 4286 53618 4338
rect 1598 4174 1650 4226
rect 9662 4174 9714 4226
rect 18510 4174 18562 4226
rect 19070 4174 19122 4226
rect 21758 4174 21810 4226
rect 27022 4174 27074 4226
rect 27246 4174 27298 4226
rect 50430 4174 50482 4226
rect 52670 4174 52722 4226
rect 55134 4174 55186 4226
rect 15710 4062 15762 4114
rect 27470 4062 27522 4114
rect 28590 4062 28642 4114
rect 28814 4062 28866 4114
rect 34414 4062 34466 4114
rect 4466 3894 4518 3946
rect 4570 3894 4622 3946
rect 4674 3894 4726 3946
rect 24466 3894 24518 3946
rect 24570 3894 24622 3946
rect 24674 3894 24726 3946
rect 44466 3894 44518 3946
rect 44570 3894 44622 3946
rect 44674 3894 44726 3946
rect 19630 3726 19682 3778
rect 26910 3726 26962 3778
rect 27246 3726 27298 3778
rect 29710 3726 29762 3778
rect 36206 3726 36258 3778
rect 37326 3726 37378 3778
rect 51662 3726 51714 3778
rect 17950 3614 18002 3666
rect 26798 3614 26850 3666
rect 27358 3614 27410 3666
rect 52558 3614 52610 3666
rect 54126 3614 54178 3666
rect 54910 3614 54962 3666
rect 9438 3502 9490 3554
rect 18398 3502 18450 3554
rect 28590 3502 28642 3554
rect 28926 3502 28978 3554
rect 29262 3502 29314 3554
rect 35758 3502 35810 3554
rect 52222 3502 52274 3554
rect 9886 3390 9938 3442
rect 19182 3390 19234 3442
rect 28814 3390 28866 3442
rect 29598 3390 29650 3442
rect 53566 3390 53618 3442
rect 29934 3278 29986 3330
rect 3806 3110 3858 3162
rect 3910 3110 3962 3162
rect 4014 3110 4066 3162
rect 23806 3110 23858 3162
rect 23910 3110 23962 3162
rect 24014 3110 24066 3162
rect 43806 3110 43858 3162
rect 43910 3110 43962 3162
rect 44014 3110 44066 3162
rect 26910 2942 26962 2994
rect 38222 2942 38274 2994
rect 54574 2942 54626 2994
rect 56142 2942 56194 2994
rect 25342 2830 25394 2882
rect 28926 2830 28978 2882
rect 41582 2830 41634 2882
rect 48414 2830 48466 2882
rect 21646 2718 21698 2770
rect 29262 2718 29314 2770
rect 29822 2718 29874 2770
rect 30382 2718 30434 2770
rect 30942 2718 30994 2770
rect 31950 2718 32002 2770
rect 35310 2718 35362 2770
rect 36542 2718 36594 2770
rect 40574 2718 40626 2770
rect 47854 2718 47906 2770
rect 50878 2718 50930 2770
rect 51998 2718 52050 2770
rect 53566 2718 53618 2770
rect 55358 2718 55410 2770
rect 22094 2606 22146 2658
rect 25678 2606 25730 2658
rect 29934 2606 29986 2658
rect 33070 2606 33122 2658
rect 35758 2606 35810 2658
rect 36990 2606 37042 2658
rect 51438 2606 51490 2658
rect 52782 2606 52834 2658
rect 32510 2494 32562 2546
rect 40014 2494 40066 2546
rect 42142 2494 42194 2546
rect 4466 2326 4518 2378
rect 4570 2326 4622 2378
rect 4674 2326 4726 2378
rect 24466 2326 24518 2378
rect 24570 2326 24622 2378
rect 24674 2326 24726 2378
rect 44466 2326 44518 2378
rect 44570 2326 44622 2378
rect 44674 2326 44726 2378
rect 26350 2158 26402 2210
rect 28702 2158 28754 2210
rect 30158 2158 30210 2210
rect 36654 2158 36706 2210
rect 41134 2158 41186 2210
rect 49086 2158 49138 2210
rect 49870 2158 49922 2210
rect 50766 2158 50818 2210
rect 12910 2046 12962 2098
rect 23998 2046 24050 2098
rect 25118 2046 25170 2098
rect 28142 2046 28194 2098
rect 29598 2046 29650 2098
rect 37214 2046 37266 2098
rect 37886 2046 37938 2098
rect 41694 2046 41746 2098
rect 51326 2046 51378 2098
rect 51662 2046 51714 2098
rect 52222 2046 52274 2098
rect 52558 2046 52610 2098
rect 54910 2046 54962 2098
rect 23550 1934 23602 1986
rect 24782 1934 24834 1986
rect 38446 1934 38498 1986
rect 47070 1934 47122 1986
rect 49310 1934 49362 1986
rect 54126 1934 54178 1986
rect 47406 1822 47458 1874
rect 50318 1822 50370 1874
rect 53566 1822 53618 1874
rect 11902 1710 11954 1762
rect 3806 1542 3858 1594
rect 3910 1542 3962 1594
rect 4014 1542 4066 1594
rect 23806 1542 23858 1594
rect 23910 1542 23962 1594
rect 24014 1542 24066 1594
rect 43806 1542 43858 1594
rect 43910 1542 43962 1594
rect 44014 1542 44066 1594
rect 53566 1374 53618 1426
rect 56142 1374 56194 1426
rect 4174 1262 4226 1314
rect 5518 1262 5570 1314
rect 7422 1262 7474 1314
rect 51998 1262 52050 1314
rect 6526 1150 6578 1202
rect 10894 1150 10946 1202
rect 14926 1150 14978 1202
rect 25678 1150 25730 1202
rect 50990 1150 51042 1202
rect 52558 1150 52610 1202
rect 55134 1150 55186 1202
rect 2158 1038 2210 1090
rect 8094 1038 8146 1090
rect 10110 1038 10162 1090
rect 14142 1038 14194 1090
rect 26126 1038 26178 1090
rect 1598 926 1650 978
rect 3614 926 3666 978
rect 4466 758 4518 810
rect 4570 758 4622 810
rect 4674 758 4726 810
rect 24466 758 24518 810
rect 24570 758 24622 810
rect 24674 758 24726 810
rect 44466 758 44518 810
rect 44570 758 44622 810
rect 44674 758 44726 810
<< metal2 >>
rect 672 14112 784 14224
rect 1120 14112 1232 14224
rect 1568 14112 1680 14224
rect 2016 14112 2128 14224
rect 2464 14112 2576 14224
rect 2912 14112 3024 14224
rect 3360 14112 3472 14224
rect 3808 14112 3920 14224
rect 4256 14112 4368 14224
rect 4704 14112 4816 14224
rect 5152 14112 5264 14224
rect 5600 14112 5712 14224
rect 6048 14112 6160 14224
rect 6496 14112 6608 14224
rect 6944 14112 7056 14224
rect 7392 14112 7504 14224
rect 7840 14112 7952 14224
rect 8288 14112 8400 14224
rect 8736 14112 8848 14224
rect 9184 14112 9296 14224
rect 9632 14112 9744 14224
rect 10080 14112 10192 14224
rect 10528 14112 10640 14224
rect 10976 14112 11088 14224
rect 11424 14112 11536 14224
rect 11872 14112 11984 14224
rect 12320 14112 12432 14224
rect 12768 14112 12880 14224
rect 13216 14112 13328 14224
rect 13664 14112 13776 14224
rect 14112 14112 14224 14224
rect 14560 14112 14672 14224
rect 15008 14112 15120 14224
rect 15456 14112 15568 14224
rect 15904 14112 16016 14224
rect 16352 14112 16464 14224
rect 16800 14112 16912 14224
rect 17248 14112 17360 14224
rect 17696 14112 17808 14224
rect 18144 14112 18256 14224
rect 18592 14112 18704 14224
rect 19040 14112 19152 14224
rect 19488 14112 19600 14224
rect 19936 14112 20048 14224
rect 20384 14112 20496 14224
rect 20832 14112 20944 14224
rect 21084 14196 21140 14206
rect 588 13076 644 13086
rect 252 12180 308 12190
rect 252 8036 308 12124
rect 588 10836 644 13020
rect 700 11620 756 14112
rect 1148 11844 1204 14112
rect 1148 11778 1204 11788
rect 1484 13524 1540 13534
rect 700 11564 1316 11620
rect 1036 11394 1092 11406
rect 1036 11342 1038 11394
rect 1090 11342 1092 11394
rect 588 10780 980 10836
rect 252 7970 308 7980
rect 812 9268 868 9278
rect 812 4116 868 9212
rect 924 4340 980 10780
rect 1036 9044 1092 11342
rect 1036 8978 1092 8988
rect 1148 10836 1204 10846
rect 1036 7700 1092 7710
rect 1036 7474 1092 7644
rect 1036 7422 1038 7474
rect 1090 7422 1092 7474
rect 1036 7410 1092 7422
rect 1036 7252 1092 7262
rect 1036 6914 1092 7196
rect 1036 6862 1038 6914
rect 1090 6862 1092 6914
rect 1036 6850 1092 6862
rect 1036 6356 1092 6366
rect 1036 5906 1092 6300
rect 1036 5854 1038 5906
rect 1090 5854 1092 5906
rect 1036 5842 1092 5854
rect 1148 5122 1204 10780
rect 1260 8146 1316 11564
rect 1484 10836 1540 13468
rect 1596 11956 1652 14112
rect 1596 11890 1652 11900
rect 1932 11732 1988 11742
rect 1484 10770 1540 10780
rect 1596 11282 1652 11294
rect 1596 11230 1598 11282
rect 1650 11230 1652 11282
rect 1484 10164 1540 10174
rect 1484 8428 1540 10108
rect 1596 9828 1652 11230
rect 1596 9762 1652 9772
rect 1820 11284 1876 11294
rect 1820 8428 1876 11228
rect 1932 10500 1988 11676
rect 2044 10722 2100 14112
rect 2380 13972 2436 13982
rect 2156 13412 2212 13422
rect 2156 13186 2212 13356
rect 2156 13134 2158 13186
rect 2210 13134 2212 13186
rect 2156 13122 2212 13134
rect 2268 12404 2324 12414
rect 2268 12310 2324 12348
rect 2268 11956 2324 11966
rect 2044 10670 2046 10722
rect 2098 10670 2100 10722
rect 2044 10658 2100 10670
rect 2156 11844 2212 11854
rect 1932 10434 1988 10444
rect 1484 8372 1652 8428
rect 1260 8094 1262 8146
rect 1314 8094 1316 8146
rect 1260 8082 1316 8094
rect 1596 7586 1652 8372
rect 1596 7534 1598 7586
rect 1650 7534 1652 7586
rect 1596 7522 1652 7534
rect 1708 8372 1876 8428
rect 1932 9380 1988 9390
rect 1932 8428 1988 9324
rect 2044 9268 2100 9278
rect 2156 9268 2212 11788
rect 2268 9938 2324 11900
rect 2268 9886 2270 9938
rect 2322 9886 2324 9938
rect 2268 9874 2324 9886
rect 2044 9266 2212 9268
rect 2044 9214 2046 9266
rect 2098 9214 2212 9266
rect 2044 9212 2212 9214
rect 2268 9604 2324 9614
rect 2044 9202 2100 9212
rect 1932 8372 2100 8428
rect 1596 7252 1652 7262
rect 1148 5070 1150 5122
rect 1202 5070 1204 5122
rect 1148 5058 1204 5070
rect 1372 6580 1428 6590
rect 1036 4340 1092 4350
rect 924 4338 1092 4340
rect 924 4286 1038 4338
rect 1090 4286 1092 4338
rect 924 4284 1092 4286
rect 1036 4274 1092 4284
rect 812 4050 868 4060
rect 1372 3220 1428 6524
rect 1484 6578 1540 6590
rect 1484 6526 1486 6578
rect 1538 6526 1540 6578
rect 1484 4116 1540 6526
rect 1596 6018 1652 7196
rect 1596 5966 1598 6018
rect 1650 5966 1652 6018
rect 1596 5954 1652 5966
rect 1708 5908 1764 8372
rect 1932 7252 1988 7262
rect 1820 7250 1988 7252
rect 1820 7198 1934 7250
rect 1986 7198 1988 7250
rect 1820 7196 1988 7198
rect 1820 6804 1876 7196
rect 1932 7186 1988 7196
rect 1820 6738 1876 6748
rect 1932 6690 1988 6702
rect 1932 6638 1934 6690
rect 1986 6638 1988 6690
rect 1932 6132 1988 6638
rect 1932 6066 1988 6076
rect 1932 5908 1988 5918
rect 1708 5906 1988 5908
rect 1708 5854 1934 5906
rect 1986 5854 1988 5906
rect 1708 5852 1988 5854
rect 1932 5842 1988 5852
rect 1596 5124 1652 5134
rect 1596 5122 1764 5124
rect 1596 5070 1598 5122
rect 1650 5070 1764 5122
rect 1596 5068 1764 5070
rect 1596 5058 1652 5068
rect 1708 4900 1764 5068
rect 2044 5122 2100 8372
rect 2268 8370 2324 9548
rect 2380 9380 2436 13916
rect 2492 11284 2548 14112
rect 2716 12962 2772 12974
rect 2716 12910 2718 12962
rect 2770 12910 2772 12962
rect 2604 11284 2660 11294
rect 2492 11282 2660 11284
rect 2492 11230 2606 11282
rect 2658 11230 2660 11282
rect 2492 11228 2660 11230
rect 2604 11218 2660 11228
rect 2716 10724 2772 12910
rect 2828 12740 2884 12750
rect 2828 12178 2884 12684
rect 2828 12126 2830 12178
rect 2882 12126 2884 12178
rect 2828 12114 2884 12126
rect 2940 12180 2996 14112
rect 3388 12404 3444 14112
rect 3612 13524 3668 13534
rect 3388 12338 3444 12348
rect 3500 12628 3556 12638
rect 2940 12114 2996 12124
rect 3388 12180 3444 12190
rect 3388 10834 3444 12124
rect 3388 10782 3390 10834
rect 3442 10782 3444 10834
rect 3388 10770 3444 10782
rect 2716 10658 2772 10668
rect 2828 10612 2884 10622
rect 2828 10518 2884 10556
rect 2380 9314 2436 9324
rect 2716 10500 2772 10510
rect 2604 8930 2660 8942
rect 2604 8878 2606 8930
rect 2658 8878 2660 8930
rect 2604 8708 2660 8878
rect 2268 8318 2270 8370
rect 2322 8318 2324 8370
rect 2268 8306 2324 8318
rect 2492 8652 2660 8708
rect 2380 7588 2436 7598
rect 2492 7588 2548 8652
rect 2604 8258 2660 8270
rect 2604 8206 2606 8258
rect 2658 8206 2660 8258
rect 2604 8148 2660 8206
rect 2604 8082 2660 8092
rect 2492 7532 2660 7588
rect 2380 6578 2436 7532
rect 2492 7362 2548 7374
rect 2492 7310 2494 7362
rect 2546 7310 2548 7362
rect 2492 6692 2548 7310
rect 2492 6626 2548 6636
rect 2380 6526 2382 6578
rect 2434 6526 2436 6578
rect 2380 6514 2436 6526
rect 2492 5794 2548 5806
rect 2492 5742 2494 5794
rect 2546 5742 2548 5794
rect 2492 5348 2548 5742
rect 2492 5282 2548 5292
rect 2044 5070 2046 5122
rect 2098 5070 2100 5122
rect 2044 5058 2100 5070
rect 1708 4834 1764 4844
rect 2492 5010 2548 5022
rect 2492 4958 2494 5010
rect 2546 4958 2548 5010
rect 2268 4564 2324 4574
rect 1484 4050 1540 4060
rect 1596 4226 1652 4238
rect 1596 4174 1598 4226
rect 1650 4174 1652 4226
rect 1596 3780 1652 4174
rect 1596 3714 1652 3724
rect 1372 3154 1428 3164
rect 1260 2884 1316 2894
rect 1260 980 1316 2828
rect 2268 1428 2324 4508
rect 2492 4564 2548 4958
rect 2492 4498 2548 4508
rect 2604 4340 2660 7532
rect 2716 6916 2772 10444
rect 2828 10388 2884 10398
rect 2828 7474 2884 10332
rect 3052 9826 3108 9838
rect 3052 9774 3054 9826
rect 3106 9774 3108 9826
rect 2940 8818 2996 8830
rect 2940 8766 2942 8818
rect 2994 8766 2996 8818
rect 2940 8596 2996 8766
rect 2940 8530 2996 8540
rect 2828 7422 2830 7474
rect 2882 7422 2884 7474
rect 2828 7410 2884 7422
rect 2828 6916 2884 6926
rect 2716 6914 2884 6916
rect 2716 6862 2830 6914
rect 2882 6862 2884 6914
rect 2716 6860 2884 6862
rect 2828 6850 2884 6860
rect 3052 5796 3108 9774
rect 3500 9156 3556 12572
rect 3612 12290 3668 13468
rect 3724 13188 3780 13198
rect 3724 13094 3780 13132
rect 3836 12740 3892 14112
rect 4284 13412 4340 14112
rect 4732 13524 4788 14112
rect 4732 13458 4788 13468
rect 4284 13346 4340 13356
rect 4464 13356 4728 13366
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4464 13290 4728 13300
rect 4284 12964 4340 12974
rect 4284 12870 4340 12908
rect 3836 12684 4340 12740
rect 3804 12572 4068 12582
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 3804 12506 4068 12516
rect 3612 12238 3614 12290
rect 3666 12238 3668 12290
rect 3612 12226 3668 12238
rect 3612 11394 3668 11406
rect 3612 11342 3614 11394
rect 3666 11342 3668 11394
rect 3612 10500 3668 11342
rect 3804 11004 4068 11014
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 3804 10938 4068 10948
rect 3612 10434 3668 10444
rect 4172 10724 4228 10734
rect 3804 9436 4068 9446
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 3804 9370 4068 9380
rect 3836 9268 3892 9278
rect 3500 9100 3668 9156
rect 3500 8932 3556 8942
rect 3500 8838 3556 8876
rect 3164 8260 3220 8270
rect 3164 8166 3220 8204
rect 3500 8148 3556 8158
rect 3500 8054 3556 8092
rect 3052 5730 3108 5740
rect 3164 7700 3220 7710
rect 3164 5460 3220 7644
rect 3276 7586 3332 7598
rect 3276 7534 3278 7586
rect 3330 7534 3332 7586
rect 3276 5908 3332 7534
rect 3612 7476 3668 9100
rect 3836 9042 3892 9212
rect 3836 8990 3838 9042
rect 3890 8990 3892 9042
rect 3836 8978 3892 8990
rect 4060 8372 4116 8382
rect 4060 8278 4116 8316
rect 3804 7868 4068 7878
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 3804 7802 4068 7812
rect 3724 7476 3780 7486
rect 3612 7474 3780 7476
rect 3612 7422 3726 7474
rect 3778 7422 3780 7474
rect 3612 7420 3780 7422
rect 3724 7410 3780 7420
rect 4172 7476 4228 10668
rect 4284 9714 4340 12684
rect 5068 12292 5124 12302
rect 5068 12198 5124 12236
rect 4396 12180 4452 12190
rect 4396 12086 4452 12124
rect 4956 12068 5012 12078
rect 4464 11788 4728 11798
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4464 11722 4728 11732
rect 4620 11620 4676 11630
rect 4620 11526 4676 11564
rect 4396 10724 4452 10734
rect 4396 10610 4452 10668
rect 4396 10558 4398 10610
rect 4450 10558 4452 10610
rect 4396 10546 4452 10558
rect 4956 10612 5012 12012
rect 5180 11620 5236 14112
rect 5628 13188 5684 14112
rect 5628 13122 5684 13132
rect 5964 13188 6020 13198
rect 5964 13094 6020 13132
rect 5964 12964 6020 12974
rect 5180 11554 5236 11564
rect 5404 12178 5460 12190
rect 5404 12126 5406 12178
rect 5458 12126 5460 12178
rect 5180 11394 5236 11406
rect 5180 11342 5182 11394
rect 5234 11342 5236 11394
rect 5180 10948 5236 11342
rect 5180 10882 5236 10892
rect 5292 11396 5348 11406
rect 4956 10546 5012 10556
rect 5068 10610 5124 10622
rect 5068 10558 5070 10610
rect 5122 10558 5124 10610
rect 4464 10220 4728 10230
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4464 10154 4728 10164
rect 5068 9940 5124 10558
rect 5068 9874 5124 9884
rect 5180 10500 5236 10510
rect 4284 9662 4286 9714
rect 4338 9662 4340 9714
rect 4284 9650 4340 9662
rect 5068 9042 5124 9054
rect 5068 8990 5070 9042
rect 5122 8990 5124 9042
rect 4396 8930 4452 8942
rect 4396 8878 4398 8930
rect 4450 8878 4452 8930
rect 4396 8820 4452 8878
rect 4396 8754 4452 8764
rect 4464 8652 4728 8662
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4464 8586 4728 8596
rect 4396 8258 4452 8270
rect 4396 8206 4398 8258
rect 4450 8206 4452 8258
rect 4396 8036 4452 8206
rect 4396 7970 4452 7980
rect 4956 8146 5012 8158
rect 4956 8094 4958 8146
rect 5010 8094 5012 8146
rect 4172 7410 4228 7420
rect 4284 7362 4340 7374
rect 4284 7310 4286 7362
rect 4338 7310 4340 7362
rect 3276 5842 3332 5852
rect 3388 6578 3444 6590
rect 3388 6526 3390 6578
rect 3442 6526 3444 6578
rect 3388 5684 3444 6526
rect 3804 6300 4068 6310
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 3804 6234 4068 6244
rect 3388 5618 3444 5628
rect 3164 5394 3220 5404
rect 3804 4732 4068 4742
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 3804 4666 4068 4676
rect 2604 4274 2660 4284
rect 3804 3164 4068 3174
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 3804 3098 4068 3108
rect 4284 2100 4340 7310
rect 4464 7084 4728 7094
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4464 7018 4728 7028
rect 4464 5516 4728 5526
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4464 5450 4728 5460
rect 4464 3948 4728 3958
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4464 3882 4728 3892
rect 4464 2380 4728 2390
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4464 2314 4728 2324
rect 4284 2034 4340 2044
rect 4956 1652 5012 8094
rect 5068 3556 5124 8990
rect 5180 5572 5236 10444
rect 5292 9938 5348 11340
rect 5292 9886 5294 9938
rect 5346 9886 5348 9938
rect 5292 9874 5348 9886
rect 5404 8708 5460 12126
rect 5516 11060 5572 11070
rect 5516 10722 5572 11004
rect 5516 10670 5518 10722
rect 5570 10670 5572 10722
rect 5516 10658 5572 10670
rect 5628 10948 5684 10958
rect 5628 9156 5684 10892
rect 5628 9090 5684 9100
rect 5852 10836 5908 10846
rect 5852 9042 5908 10780
rect 5852 8990 5854 9042
rect 5906 8990 5908 9042
rect 5852 8978 5908 8990
rect 5516 8932 5572 8942
rect 5516 8930 5796 8932
rect 5516 8878 5518 8930
rect 5570 8878 5796 8930
rect 5516 8876 5796 8878
rect 5516 8866 5572 8876
rect 5404 8652 5684 8708
rect 5180 5506 5236 5516
rect 5404 8484 5460 8494
rect 5068 3490 5124 3500
rect 5180 5012 5236 5022
rect 3804 1596 4068 1606
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 4956 1586 5012 1596
rect 5068 3332 5124 3342
rect 3804 1530 4068 1540
rect 2268 1362 2324 1372
rect 4172 1316 4228 1326
rect 4172 1222 4228 1260
rect 5068 1204 5124 3276
rect 5180 2996 5236 4956
rect 5180 2930 5236 2940
rect 5292 4228 5348 4238
rect 5292 2212 5348 4172
rect 5404 2772 5460 8428
rect 5628 6132 5684 8652
rect 5740 6244 5796 8876
rect 5964 6356 6020 12908
rect 6076 11956 6132 14112
rect 6524 13188 6580 14112
rect 6076 11890 6132 11900
rect 6412 13132 6580 13188
rect 6188 11620 6244 11630
rect 6188 11526 6244 11564
rect 6412 10834 6468 13132
rect 6412 10782 6414 10834
rect 6466 10782 6468 10834
rect 6412 10770 6468 10782
rect 6524 12962 6580 12974
rect 6524 12910 6526 12962
rect 6578 12910 6580 12962
rect 6188 9716 6244 9726
rect 6188 7252 6244 9660
rect 6412 8930 6468 8942
rect 6412 8878 6414 8930
rect 6466 8878 6468 8930
rect 6188 7186 6244 7196
rect 6300 8820 6356 8830
rect 5964 6300 6244 6356
rect 5740 6188 6020 6244
rect 5628 6076 5908 6132
rect 5740 5572 5796 5582
rect 5404 2706 5460 2716
rect 5628 3444 5684 3454
rect 5292 2146 5348 2156
rect 5516 1316 5572 1326
rect 5068 1138 5124 1148
rect 5404 1314 5572 1316
rect 5404 1262 5518 1314
rect 5570 1262 5572 1314
rect 5404 1260 5572 1262
rect 2156 1090 2212 1102
rect 2156 1038 2158 1090
rect 2210 1038 2212 1090
rect 1596 980 1652 990
rect 1260 914 1316 924
rect 1372 978 1652 980
rect 1372 926 1598 978
rect 1650 926 1652 978
rect 1372 924 1652 926
rect 1372 112 1428 924
rect 1596 914 1652 924
rect 2156 308 2212 1038
rect 3612 980 3668 990
rect 2156 242 2212 252
rect 3388 978 3668 980
rect 3388 926 3614 978
rect 3666 926 3668 978
rect 3388 924 3668 926
rect 3388 112 3444 924
rect 3612 914 3668 924
rect 4464 812 4728 822
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4464 746 4728 756
rect 5404 112 5460 1260
rect 5516 1250 5572 1260
rect 5628 532 5684 3388
rect 5740 3108 5796 5516
rect 5740 3042 5796 3052
rect 5852 2884 5908 6076
rect 5852 2818 5908 2828
rect 5964 756 6020 6188
rect 6188 5124 6244 6300
rect 6188 5058 6244 5068
rect 6188 4900 6244 4910
rect 6076 4340 6132 4350
rect 6076 2436 6132 4284
rect 6076 2370 6132 2380
rect 6188 1764 6244 4844
rect 6300 4452 6356 8764
rect 6412 8708 6468 8878
rect 6412 8642 6468 8652
rect 6524 8260 6580 12910
rect 6972 12180 7028 14112
rect 6748 12124 7028 12180
rect 7308 13748 7364 13758
rect 7308 12178 7364 13692
rect 7420 13188 7476 14112
rect 7420 13122 7476 13132
rect 7532 13412 7588 13422
rect 7532 13186 7588 13356
rect 7532 13134 7534 13186
rect 7586 13134 7588 13186
rect 7532 13122 7588 13134
rect 7308 12126 7310 12178
rect 7362 12126 7364 12178
rect 6748 11620 6804 12124
rect 7308 12114 7364 12126
rect 6748 11554 6804 11564
rect 6860 11956 6916 11966
rect 6412 8204 6580 8260
rect 6636 11394 6692 11406
rect 6636 11342 6638 11394
rect 6690 11342 6692 11394
rect 6412 4676 6468 8204
rect 6412 4610 6468 4620
rect 6524 8036 6580 8046
rect 6524 4564 6580 7980
rect 6636 7924 6692 11342
rect 6860 9714 6916 11900
rect 6972 11954 7028 11966
rect 6972 11902 6974 11954
rect 7026 11902 7028 11954
rect 6972 11844 7028 11902
rect 6972 11778 7028 11788
rect 7756 11620 7812 11630
rect 7756 11526 7812 11564
rect 7868 10836 7924 14112
rect 8204 13300 8260 13310
rect 8092 12962 8148 12974
rect 8092 12910 8094 12962
rect 8146 12910 8148 12962
rect 7980 10836 8036 10846
rect 7868 10834 8036 10836
rect 7868 10782 7982 10834
rect 8034 10782 8036 10834
rect 7868 10780 8036 10782
rect 7980 10770 8036 10780
rect 7420 10612 7476 10622
rect 7420 10518 7476 10556
rect 6860 9662 6862 9714
rect 6914 9662 6916 9714
rect 6860 9650 6916 9662
rect 7532 9826 7588 9838
rect 7532 9774 7534 9826
rect 7586 9774 7588 9826
rect 7532 8820 7588 9774
rect 7532 8754 7588 8764
rect 7980 9828 8036 9838
rect 7756 8260 7812 8270
rect 7756 8166 7812 8204
rect 6636 7858 6692 7868
rect 7868 7364 7924 7374
rect 6636 7140 6692 7150
rect 6636 5012 6692 7084
rect 7308 6020 7364 6030
rect 7308 5926 7364 5964
rect 7868 6018 7924 7308
rect 7868 5966 7870 6018
rect 7922 5966 7924 6018
rect 7868 5954 7924 5966
rect 6748 5908 6804 5918
rect 6748 5814 6804 5852
rect 6636 4946 6692 4956
rect 6524 4498 6580 4508
rect 6300 4386 6356 4396
rect 7980 3892 8036 9772
rect 7980 3826 8036 3836
rect 6188 1698 6244 1708
rect 6524 2660 6580 2670
rect 6524 1202 6580 2604
rect 8092 1988 8148 12910
rect 8204 12290 8260 13244
rect 8204 12238 8206 12290
rect 8258 12238 8260 12290
rect 8204 12226 8260 12238
rect 8204 12068 8260 12078
rect 8204 11394 8260 12012
rect 8316 11844 8372 14112
rect 8316 11778 8372 11788
rect 8764 11620 8820 14112
rect 9212 12964 9268 14112
rect 9660 13412 9716 14112
rect 9660 13346 9716 13356
rect 10108 13300 10164 14112
rect 10108 13234 10164 13244
rect 9772 13188 9828 13198
rect 9772 13094 9828 13132
rect 10108 13076 10164 13086
rect 9212 12908 9492 12964
rect 8764 11554 8820 11564
rect 9100 12066 9156 12078
rect 9100 12014 9102 12066
rect 9154 12014 9156 12066
rect 8204 11342 8206 11394
rect 8258 11342 8260 11394
rect 8204 11330 8260 11342
rect 8428 11172 8484 11182
rect 8428 8372 8484 11116
rect 8988 10836 9044 10846
rect 8988 10610 9044 10780
rect 8988 10558 8990 10610
rect 9042 10558 9044 10610
rect 8988 10546 9044 10558
rect 8428 8306 8484 8316
rect 8652 8260 8708 8270
rect 8204 8146 8260 8158
rect 8204 8094 8206 8146
rect 8258 8094 8260 8146
rect 8204 6132 8260 8094
rect 8316 7474 8372 7486
rect 8316 7422 8318 7474
rect 8370 7422 8372 7474
rect 8316 7364 8372 7422
rect 8316 7298 8372 7308
rect 8652 7362 8708 8204
rect 8652 7310 8654 7362
rect 8706 7310 8708 7362
rect 8652 7298 8708 7310
rect 8204 6066 8260 6076
rect 8204 5908 8260 5918
rect 8204 5794 8260 5852
rect 8204 5742 8206 5794
rect 8258 5742 8260 5794
rect 8204 5730 8260 5742
rect 9100 3220 9156 12014
rect 9212 11394 9268 11406
rect 9212 11342 9214 11394
rect 9266 11342 9268 11394
rect 9212 10164 9268 11342
rect 9212 10098 9268 10108
rect 9436 9714 9492 12908
rect 10108 12402 10164 13020
rect 10108 12350 10110 12402
rect 10162 12350 10164 12402
rect 10108 12338 10164 12350
rect 10220 12962 10276 12974
rect 10220 12910 10222 12962
rect 10274 12910 10276 12962
rect 10108 11844 10164 11854
rect 9772 11282 9828 11294
rect 9772 11230 9774 11282
rect 9826 11230 9828 11282
rect 9436 9662 9438 9714
rect 9490 9662 9492 9714
rect 9436 9650 9492 9662
rect 9548 10610 9604 10622
rect 9548 10558 9550 10610
rect 9602 10558 9604 10610
rect 9324 7364 9380 7374
rect 9324 4450 9380 7308
rect 9548 7364 9604 10558
rect 9548 7298 9604 7308
rect 9660 8932 9716 8942
rect 9436 6692 9492 6702
rect 9436 6130 9492 6636
rect 9436 6078 9438 6130
rect 9490 6078 9492 6130
rect 9436 6066 9492 6078
rect 9324 4398 9326 4450
rect 9378 4398 9380 4450
rect 9324 4386 9380 4398
rect 9660 4228 9716 8876
rect 9772 8596 9828 11230
rect 9884 10498 9940 10510
rect 9884 10446 9886 10498
rect 9938 10446 9940 10498
rect 9884 10164 9940 10446
rect 9884 10098 9940 10108
rect 10108 9716 10164 11788
rect 10108 9650 10164 9660
rect 9772 8530 9828 8540
rect 9996 9042 10052 9054
rect 9996 8990 9998 9042
rect 10050 8990 10052 9042
rect 9436 4226 9716 4228
rect 9436 4174 9662 4226
rect 9714 4174 9716 4226
rect 9436 4172 9716 4174
rect 9436 3554 9492 4172
rect 9660 4162 9716 4172
rect 9772 8372 9828 8382
rect 9772 4228 9828 8316
rect 9884 7250 9940 7262
rect 9884 7198 9886 7250
rect 9938 7198 9940 7250
rect 9884 6804 9940 7198
rect 9884 6738 9940 6748
rect 9772 4162 9828 4172
rect 9996 3892 10052 8990
rect 10108 8148 10164 8158
rect 10108 6356 10164 8092
rect 10108 6290 10164 6300
rect 9436 3502 9438 3554
rect 9490 3502 9492 3554
rect 9436 3490 9492 3502
rect 9772 3836 10052 3892
rect 9100 3154 9156 3164
rect 9548 3444 9604 3454
rect 8092 1922 8148 1932
rect 9100 2884 9156 2894
rect 6524 1150 6526 1202
rect 6578 1150 6580 1202
rect 6524 1138 6580 1150
rect 7420 1314 7476 1326
rect 7420 1262 7422 1314
rect 7474 1262 7476 1314
rect 5964 690 6020 700
rect 5628 466 5684 476
rect 7420 112 7476 1262
rect 9100 1316 9156 2828
rect 9548 1428 9604 3388
rect 9548 1362 9604 1372
rect 9660 2996 9716 3006
rect 9100 1250 9156 1260
rect 8092 1090 8148 1102
rect 8092 1038 8094 1090
rect 8146 1038 8148 1090
rect 8092 868 8148 1038
rect 8092 802 8148 812
rect 9660 868 9716 2940
rect 9772 1876 9828 3836
rect 9884 3442 9940 3454
rect 9884 3390 9886 3442
rect 9938 3390 9940 3442
rect 9884 3388 9940 3390
rect 9884 3332 10052 3388
rect 9772 1810 9828 1820
rect 9884 3108 9940 3118
rect 9660 802 9716 812
rect 9884 644 9940 3052
rect 9996 1652 10052 3332
rect 9996 1586 10052 1596
rect 9884 578 9940 588
rect 10108 1090 10164 1102
rect 10108 1038 10110 1090
rect 10162 1038 10164 1090
rect 9436 196 9492 206
rect 9436 112 9492 140
rect 10108 196 10164 1038
rect 10220 420 10276 12910
rect 10444 12180 10500 12190
rect 10332 12178 10500 12180
rect 10332 12126 10446 12178
rect 10498 12126 10500 12178
rect 10332 12124 10500 12126
rect 10332 7700 10388 12124
rect 10444 12114 10500 12124
rect 10444 9828 10500 9838
rect 10444 9734 10500 9772
rect 10556 9716 10612 14112
rect 10780 13860 10836 13870
rect 10780 10612 10836 13804
rect 11004 13076 11060 14112
rect 11340 13300 11396 13310
rect 11340 13186 11396 13244
rect 11340 13134 11342 13186
rect 11394 13134 11396 13186
rect 11340 13122 11396 13134
rect 11004 13010 11060 13020
rect 11452 12516 11508 14112
rect 10892 12460 11508 12516
rect 11788 13412 11844 13422
rect 10892 11618 10948 12460
rect 11004 12292 11060 12302
rect 11004 12178 11060 12236
rect 11004 12126 11006 12178
rect 11058 12126 11060 12178
rect 11004 12114 11060 12126
rect 11788 12180 11844 13356
rect 11900 13188 11956 14112
rect 11900 13122 11956 13132
rect 11900 12964 11956 12974
rect 11900 12962 12292 12964
rect 11900 12910 11902 12962
rect 11954 12910 12292 12962
rect 11900 12908 12292 12910
rect 11900 12898 11956 12908
rect 12012 12404 12068 12414
rect 12012 12310 12068 12348
rect 11788 12114 11844 12124
rect 12012 12180 12068 12190
rect 10892 11566 10894 11618
rect 10946 11566 10948 11618
rect 10892 11554 10948 11566
rect 11228 11956 11284 11966
rect 10780 10546 10836 10556
rect 11116 10386 11172 10398
rect 11116 10334 11118 10386
rect 11170 10334 11172 10386
rect 11116 10164 11172 10334
rect 11116 10098 11172 10108
rect 11004 9716 11060 9726
rect 10556 9714 11060 9716
rect 10556 9662 11006 9714
rect 11058 9662 11060 9714
rect 10556 9660 11060 9662
rect 11004 9650 11060 9660
rect 10892 9380 10948 9390
rect 10332 7634 10388 7644
rect 10444 8930 10500 8942
rect 10444 8878 10446 8930
rect 10498 8878 10500 8930
rect 10332 7476 10388 7486
rect 10332 4228 10388 7420
rect 10444 7028 10500 8878
rect 10444 6962 10500 6972
rect 10556 6804 10612 6814
rect 10556 6690 10612 6748
rect 10556 6638 10558 6690
rect 10610 6638 10612 6690
rect 10556 6626 10612 6638
rect 10892 6692 10948 9324
rect 10892 6626 10948 6636
rect 11004 8818 11060 8830
rect 11004 8766 11006 8818
rect 11058 8766 11060 8818
rect 11004 6690 11060 8766
rect 11228 6916 11284 11900
rect 12012 11844 12068 12124
rect 12012 11778 12068 11788
rect 11452 11396 11508 11406
rect 11452 11394 11732 11396
rect 11452 11342 11454 11394
rect 11506 11342 11732 11394
rect 11452 11340 11732 11342
rect 11452 11330 11508 11340
rect 11564 10388 11620 10398
rect 11452 10386 11620 10388
rect 11452 10334 11566 10386
rect 11618 10334 11620 10386
rect 11452 10332 11620 10334
rect 11228 6850 11284 6860
rect 11340 9044 11396 9054
rect 11452 9044 11508 10332
rect 11564 10322 11620 10332
rect 11340 9042 11508 9044
rect 11340 8990 11342 9042
rect 11394 8990 11508 9042
rect 11340 8988 11508 8990
rect 11004 6638 11006 6690
rect 11058 6638 11060 6690
rect 11004 6626 11060 6638
rect 11116 6692 11172 6702
rect 11116 6598 11172 6636
rect 11228 6690 11284 6702
rect 11228 6638 11230 6690
rect 11282 6638 11284 6690
rect 10668 6468 10724 6478
rect 11228 6468 11284 6638
rect 10668 6466 11284 6468
rect 10668 6414 10670 6466
rect 10722 6414 11284 6466
rect 10668 6412 11284 6414
rect 10668 6402 10724 6412
rect 11340 6356 11396 8988
rect 11676 7364 11732 11340
rect 11900 10724 11956 10734
rect 11676 7298 11732 7308
rect 11788 9828 11844 9838
rect 10332 4162 10388 4172
rect 10780 6300 11396 6356
rect 11452 7252 11508 7262
rect 10780 2436 10836 6300
rect 10892 5908 10948 5918
rect 10892 5236 10948 5852
rect 10892 4562 10948 5180
rect 10892 4510 10894 4562
rect 10946 4510 10948 4562
rect 10892 4498 10948 4510
rect 11452 3388 11508 7196
rect 11788 6916 11844 9772
rect 11900 9156 11956 10668
rect 12124 10500 12180 10510
rect 12124 10406 12180 10444
rect 12124 10164 12180 10174
rect 12012 9826 12068 9838
rect 12012 9774 12014 9826
rect 12066 9774 12068 9826
rect 12012 9716 12068 9774
rect 12012 9650 12068 9660
rect 11900 9090 11956 9100
rect 12012 9492 12068 9502
rect 12012 8930 12068 9436
rect 12012 8878 12014 8930
rect 12066 8878 12068 8930
rect 12012 7476 12068 8878
rect 12124 9042 12180 10108
rect 12236 9604 12292 12908
rect 12348 11282 12404 14112
rect 12572 13972 12628 13982
rect 12348 11230 12350 11282
rect 12402 11230 12404 11282
rect 12348 11218 12404 11230
rect 12460 13636 12516 13646
rect 12460 11060 12516 13580
rect 12460 10994 12516 11004
rect 12236 9538 12292 9548
rect 12572 9268 12628 13916
rect 12796 12404 12852 14112
rect 13244 13300 13300 14112
rect 13244 13234 13300 13244
rect 13356 13188 13412 13198
rect 13356 13074 13412 13132
rect 13356 13022 13358 13074
rect 13410 13022 13412 13074
rect 13356 13010 13412 13022
rect 12796 12338 12852 12348
rect 13692 12292 13748 14112
rect 14140 13188 14196 14112
rect 14028 13132 14196 13188
rect 14476 13412 14532 13422
rect 13692 12236 13972 12292
rect 13804 12066 13860 12078
rect 13804 12014 13806 12066
rect 13858 12014 13860 12066
rect 13244 11956 13300 11966
rect 13244 11862 13300 11900
rect 13020 11394 13076 11406
rect 13020 11342 13022 11394
rect 13074 11342 13076 11394
rect 12908 9826 12964 9838
rect 12908 9774 12910 9826
rect 12962 9774 12964 9826
rect 12908 9492 12964 9774
rect 12908 9426 12964 9436
rect 12572 9202 12628 9212
rect 12124 8990 12126 9042
rect 12178 8990 12180 9042
rect 12124 8260 12180 8990
rect 12908 8930 12964 8942
rect 12908 8878 12910 8930
rect 12962 8878 12964 8930
rect 12124 8194 12180 8204
rect 12684 8596 12740 8606
rect 12012 7410 12068 7420
rect 12236 8036 12292 8046
rect 12236 7474 12292 7980
rect 12236 7422 12238 7474
rect 12290 7422 12292 7474
rect 12236 7410 12292 7422
rect 12460 7588 12516 7598
rect 11900 7252 11956 7262
rect 12124 7252 12180 7262
rect 11900 7250 12068 7252
rect 11900 7198 11902 7250
rect 11954 7198 12068 7250
rect 11900 7196 12068 7198
rect 11900 7186 11956 7196
rect 11788 6860 11956 6916
rect 11564 6690 11620 6702
rect 11564 6638 11566 6690
rect 11618 6638 11620 6690
rect 11564 6130 11620 6638
rect 11788 6692 11844 6702
rect 11788 6598 11844 6636
rect 11900 6468 11956 6860
rect 12012 6804 12068 7196
rect 12124 7250 12292 7252
rect 12124 7198 12126 7250
rect 12178 7198 12292 7250
rect 12124 7196 12292 7198
rect 12124 7186 12180 7196
rect 12236 6804 12292 7196
rect 12012 6748 12180 6804
rect 12124 6690 12180 6748
rect 12124 6638 12126 6690
rect 12178 6638 12180 6690
rect 12124 6626 12180 6638
rect 11564 6078 11566 6130
rect 11618 6078 11620 6130
rect 11564 6066 11620 6078
rect 11788 6412 11956 6468
rect 12012 6578 12068 6590
rect 12012 6526 12014 6578
rect 12066 6526 12068 6578
rect 11676 5908 11732 5918
rect 11676 5814 11732 5852
rect 10780 2370 10836 2380
rect 10892 3332 11508 3388
rect 11564 5796 11620 5806
rect 10892 1202 10948 3332
rect 11564 1428 11620 5740
rect 11788 4450 11844 6412
rect 11900 5236 11956 5246
rect 11900 5142 11956 5180
rect 11900 5012 11956 5022
rect 11900 4918 11956 4956
rect 11788 4398 11790 4450
rect 11842 4398 11844 4450
rect 11788 4386 11844 4398
rect 12012 3388 12068 6526
rect 12124 5236 12180 5246
rect 12124 5010 12180 5180
rect 12236 5124 12292 6748
rect 12236 5058 12292 5068
rect 12348 6690 12404 6702
rect 12348 6638 12350 6690
rect 12402 6638 12404 6690
rect 12124 4958 12126 5010
rect 12178 4958 12180 5010
rect 12124 4946 12180 4958
rect 12348 5012 12404 6638
rect 12460 6020 12516 7532
rect 12460 5954 12516 5964
rect 12572 7476 12628 7486
rect 12348 4946 12404 4956
rect 12460 5572 12516 5582
rect 12460 5234 12516 5516
rect 12460 5182 12462 5234
rect 12514 5182 12516 5234
rect 12460 4788 12516 5182
rect 12236 4732 12516 4788
rect 12572 4788 12628 7420
rect 12684 6468 12740 8540
rect 12796 8036 12852 8046
rect 12796 7942 12852 7980
rect 12684 6402 12740 6412
rect 12796 7700 12852 7710
rect 12236 4338 12292 4732
rect 12572 4722 12628 4732
rect 12236 4286 12238 4338
rect 12290 4286 12292 4338
rect 12236 4274 12292 4286
rect 12012 3332 12180 3388
rect 12124 2660 12180 3332
rect 12124 2594 12180 2604
rect 12348 2660 12404 2670
rect 12236 2100 12292 2110
rect 12348 2100 12404 2604
rect 12292 2044 12404 2100
rect 12236 2034 12292 2044
rect 11564 1362 11620 1372
rect 11900 1762 11956 1774
rect 11900 1710 11902 1762
rect 11954 1710 11956 1762
rect 10892 1150 10894 1202
rect 10946 1150 10948 1202
rect 10892 1138 10948 1150
rect 10220 354 10276 364
rect 10108 130 10164 140
rect 11452 196 11508 206
rect 11452 112 11508 140
rect 11900 196 11956 1710
rect 12796 532 12852 7644
rect 12908 5460 12964 8878
rect 13020 8596 13076 11342
rect 13244 11060 13300 11070
rect 13020 8530 13076 8540
rect 13132 10276 13188 10286
rect 13132 8372 13188 10220
rect 13132 8306 13188 8316
rect 12908 5394 12964 5404
rect 13020 8260 13076 8270
rect 12908 5124 12964 5134
rect 13020 5124 13076 8204
rect 13132 8034 13188 8046
rect 13132 7982 13134 8034
rect 13186 7982 13188 8034
rect 13132 7252 13188 7982
rect 13132 7186 13188 7196
rect 13244 5572 13300 11004
rect 13468 10610 13524 10622
rect 13468 10558 13470 10610
rect 13522 10558 13524 10610
rect 13356 10164 13412 10174
rect 13356 9714 13412 10108
rect 13356 9662 13358 9714
rect 13410 9662 13412 9714
rect 13356 9650 13412 9662
rect 13356 9042 13412 9054
rect 13356 8990 13358 9042
rect 13410 8990 13412 9042
rect 13356 8484 13412 8990
rect 13356 8418 13412 8428
rect 13468 7812 13524 10558
rect 13804 8932 13860 12014
rect 13916 11396 13972 12236
rect 14028 11618 14084 13132
rect 14028 11566 14030 11618
rect 14082 11566 14084 11618
rect 14028 11554 14084 11566
rect 14140 12962 14196 12974
rect 14140 12910 14142 12962
rect 14194 12910 14196 12962
rect 14140 11508 14196 12910
rect 14140 11442 14196 11452
rect 14364 12964 14420 12974
rect 13916 11340 14084 11396
rect 13804 8866 13860 8876
rect 13916 10498 13972 10510
rect 13916 10446 13918 10498
rect 13970 10446 13972 10498
rect 13692 8820 13748 8830
rect 13580 8260 13636 8270
rect 13580 8166 13636 8204
rect 13468 7746 13524 7756
rect 13468 7252 13524 7262
rect 13468 7158 13524 7196
rect 13244 5506 13300 5516
rect 13356 6132 13412 6142
rect 12908 5122 13076 5124
rect 12908 5070 12910 5122
rect 12962 5070 13076 5122
rect 12908 5068 13076 5070
rect 13356 5122 13412 6076
rect 13468 5236 13524 5246
rect 13468 5142 13524 5180
rect 13356 5070 13358 5122
rect 13410 5070 13412 5122
rect 12908 5058 12964 5068
rect 13356 5058 13412 5070
rect 13468 4676 13524 4686
rect 13468 4450 13524 4620
rect 13692 4676 13748 8764
rect 13804 8370 13860 8382
rect 13804 8318 13806 8370
rect 13858 8318 13860 8370
rect 13804 8260 13860 8318
rect 13804 8194 13860 8204
rect 13692 4610 13748 4620
rect 13468 4398 13470 4450
rect 13522 4398 13524 4450
rect 13468 4386 13524 4398
rect 13356 3668 13412 3678
rect 13356 3388 13412 3612
rect 13244 3332 13412 3388
rect 13244 3266 13300 3276
rect 12908 2996 12964 3006
rect 12908 2098 12964 2940
rect 12908 2046 12910 2098
rect 12962 2046 12964 2098
rect 12908 2034 12964 2046
rect 12796 466 12852 476
rect 13804 1876 13860 1886
rect 13804 308 13860 1820
rect 13916 1092 13972 10446
rect 14028 9716 14084 11340
rect 14252 10500 14308 10510
rect 14252 10406 14308 10444
rect 14140 9716 14196 9726
rect 14028 9714 14196 9716
rect 14028 9662 14142 9714
rect 14194 9662 14196 9714
rect 14028 9660 14196 9662
rect 14140 9650 14196 9660
rect 14364 9380 14420 12908
rect 14476 11394 14532 13356
rect 14588 12292 14644 14112
rect 14812 14084 14868 14094
rect 14812 12852 14868 14028
rect 15036 13188 15092 14112
rect 15036 13122 15092 13132
rect 14924 13076 14980 13086
rect 14924 12982 14980 13020
rect 14812 12796 14980 12852
rect 14812 12404 14868 12414
rect 14812 12310 14868 12348
rect 14588 12236 14756 12292
rect 14476 11342 14478 11394
rect 14530 11342 14532 11394
rect 14476 11330 14532 11342
rect 14588 11620 14644 11630
rect 14476 10500 14532 10510
rect 14476 10276 14532 10444
rect 14476 10210 14532 10220
rect 14028 9324 14420 9380
rect 14028 7586 14084 9324
rect 14028 7534 14030 7586
rect 14082 7534 14084 7586
rect 14028 7522 14084 7534
rect 14252 8596 14308 8606
rect 14028 6132 14084 6142
rect 14028 4338 14084 6076
rect 14140 5124 14196 5134
rect 14140 5030 14196 5068
rect 14028 4286 14030 4338
rect 14082 4286 14084 4338
rect 14028 4274 14084 4286
rect 14252 3556 14308 8540
rect 14476 8258 14532 8270
rect 14476 8206 14478 8258
rect 14530 8206 14532 8258
rect 14476 8148 14532 8206
rect 14476 8082 14532 8092
rect 14252 3490 14308 3500
rect 14588 3388 14644 11564
rect 14700 10836 14756 12236
rect 14812 10836 14868 10846
rect 14700 10834 14868 10836
rect 14700 10782 14814 10834
rect 14866 10782 14868 10834
rect 14700 10780 14868 10782
rect 14812 10770 14868 10780
rect 14924 8370 14980 12796
rect 15372 12066 15428 12078
rect 15372 12014 15374 12066
rect 15426 12014 15428 12066
rect 15148 9828 15204 9838
rect 15148 9826 15316 9828
rect 15148 9774 15150 9826
rect 15202 9774 15316 9826
rect 15148 9772 15316 9774
rect 15148 9762 15204 9772
rect 14924 8318 14926 8370
rect 14978 8318 14980 8370
rect 14924 8306 14980 8318
rect 14700 5122 14756 5134
rect 14700 5070 14702 5122
rect 14754 5070 14756 5122
rect 14700 5012 14756 5070
rect 14700 4946 14756 4956
rect 15148 4564 15204 4574
rect 15148 4450 15204 4508
rect 15148 4398 15150 4450
rect 15202 4398 15204 4450
rect 15148 4386 15204 4398
rect 15260 3668 15316 9772
rect 15372 8484 15428 12014
rect 15484 11282 15540 14112
rect 15484 11230 15486 11282
rect 15538 11230 15540 11282
rect 15484 11218 15540 11230
rect 15708 12962 15764 12974
rect 15708 12910 15710 12962
rect 15762 12910 15764 12962
rect 15708 10276 15764 12910
rect 15932 12404 15988 14112
rect 16380 13748 16436 14112
rect 16380 13692 16548 13748
rect 15932 12338 15988 12348
rect 16380 12404 16436 12414
rect 16380 12310 16436 12348
rect 16044 11394 16100 11406
rect 16044 11342 16046 11394
rect 16098 11342 16100 11394
rect 15708 10210 15764 10220
rect 15820 10498 15876 10510
rect 15820 10446 15822 10498
rect 15874 10446 15876 10498
rect 15820 10164 15876 10446
rect 15820 10098 15876 10108
rect 15372 8418 15428 8428
rect 15596 5572 15652 5582
rect 15596 5122 15652 5516
rect 15596 5070 15598 5122
rect 15650 5070 15652 5122
rect 15596 5058 15652 5070
rect 15260 3602 15316 3612
rect 15708 5012 15764 5022
rect 15708 4114 15764 4956
rect 15708 4062 15710 4114
rect 15762 4062 15764 4114
rect 14140 3332 14644 3388
rect 15708 3444 15764 4062
rect 15820 4340 15876 4350
rect 15820 3892 15876 4284
rect 15820 3826 15876 3836
rect 16044 3892 16100 11342
rect 16492 10722 16548 13692
rect 16716 13524 16772 13534
rect 16492 10670 16494 10722
rect 16546 10670 16548 10722
rect 16492 10658 16548 10670
rect 16604 11956 16660 11966
rect 16604 9492 16660 11900
rect 16716 11620 16772 13468
rect 16828 13076 16884 14112
rect 16828 13010 16884 13020
rect 17276 12404 17332 14112
rect 17388 13188 17444 13198
rect 17388 13094 17444 13132
rect 17724 12628 17780 14112
rect 17276 12338 17332 12348
rect 17500 12572 17780 12628
rect 17836 12962 17892 12974
rect 17836 12910 17838 12962
rect 17890 12910 17892 12962
rect 16716 11554 16772 11564
rect 16940 12066 16996 12078
rect 16940 12014 16942 12066
rect 16994 12014 16996 12066
rect 16940 11620 16996 12014
rect 16940 11554 16996 11564
rect 17164 11844 17220 11854
rect 17164 10500 17220 11788
rect 17500 11618 17556 12572
rect 17500 11566 17502 11618
rect 17554 11566 17556 11618
rect 17500 11554 17556 11566
rect 17836 11620 17892 12910
rect 17948 12404 18004 12414
rect 18172 12404 18228 14112
rect 18620 13188 18676 14112
rect 18620 13122 18676 13132
rect 18956 13188 19012 13198
rect 18956 13094 19012 13132
rect 17948 12402 18228 12404
rect 17948 12350 17950 12402
rect 18002 12350 18228 12402
rect 17948 12348 18228 12350
rect 18284 12404 18340 12414
rect 17948 12338 18004 12348
rect 18284 11732 18340 12348
rect 18396 12180 18452 12190
rect 18396 12086 18452 12124
rect 18284 11666 18340 11676
rect 17836 11564 18004 11620
rect 17836 11394 17892 11406
rect 17836 11342 17838 11394
rect 17890 11342 17892 11394
rect 17164 10434 17220 10444
rect 17388 10500 17444 10510
rect 17388 9938 17444 10444
rect 17388 9886 17390 9938
rect 17442 9886 17444 9938
rect 17388 9874 17444 9886
rect 17724 10498 17780 10510
rect 17724 10446 17726 10498
rect 17778 10446 17780 10498
rect 17724 9828 17780 10446
rect 17836 9940 17892 11342
rect 17948 10948 18004 11564
rect 19068 11618 19124 14112
rect 19516 13188 19572 14112
rect 19404 13132 19572 13188
rect 19964 13188 20020 14112
rect 19068 11566 19070 11618
rect 19122 11566 19124 11618
rect 19068 11554 19124 11566
rect 19292 12962 19348 12974
rect 19292 12910 19294 12962
rect 19346 12910 19348 12962
rect 17948 10882 18004 10892
rect 18284 10724 18340 10734
rect 18060 10668 18284 10724
rect 17948 10498 18004 10510
rect 17948 10446 17950 10498
rect 18002 10446 18004 10498
rect 17948 10276 18004 10446
rect 17948 10210 18004 10220
rect 17948 10052 18004 10062
rect 18060 10052 18116 10668
rect 18284 10630 18340 10668
rect 18620 10388 18676 10398
rect 18396 10386 18676 10388
rect 18396 10334 18622 10386
rect 18674 10334 18676 10386
rect 18396 10332 18676 10334
rect 17948 10050 18116 10052
rect 17948 9998 17950 10050
rect 18002 9998 18116 10050
rect 17948 9996 18116 9998
rect 18172 10276 18228 10286
rect 17948 9986 18004 9996
rect 17836 9874 17892 9884
rect 17724 9762 17780 9772
rect 18172 9604 18228 10220
rect 18284 9828 18340 9838
rect 18284 9734 18340 9772
rect 18172 9548 18340 9604
rect 16604 9426 16660 9436
rect 17948 9492 18004 9502
rect 17948 9044 18004 9436
rect 18284 9380 18340 9548
rect 18060 9156 18116 9166
rect 18060 9062 18116 9100
rect 17948 8978 18004 8988
rect 18284 9044 18340 9324
rect 16492 8820 16548 8830
rect 16156 8148 16212 8158
rect 16156 7586 16212 8092
rect 16156 7534 16158 7586
rect 16210 7534 16212 7586
rect 16156 6916 16212 7534
rect 16156 6850 16212 6860
rect 16044 3826 16100 3836
rect 16156 5012 16212 5022
rect 15708 3378 15764 3388
rect 14140 2884 14196 3332
rect 14140 2818 14196 2828
rect 14924 1316 14980 1326
rect 14924 1202 14980 1260
rect 14924 1150 14926 1202
rect 14978 1150 14980 1202
rect 14924 1138 14980 1150
rect 13916 1026 13972 1036
rect 14140 1090 14196 1102
rect 14140 1038 14142 1090
rect 14194 1038 14196 1090
rect 13804 242 13860 252
rect 11900 130 11956 140
rect 13468 196 13524 206
rect 13468 112 13524 140
rect 14140 196 14196 1038
rect 14140 130 14196 140
rect 15484 196 15540 206
rect 15484 112 15540 140
rect 15820 196 15876 206
rect 1344 0 1456 112
rect 3360 0 3472 112
rect 5376 0 5488 112
rect 7392 0 7504 112
rect 9408 0 9520 112
rect 11424 0 11536 112
rect 13440 0 13552 112
rect 15456 0 15568 112
rect 15820 84 15876 140
rect 16156 84 16212 4956
rect 16492 1652 16548 8764
rect 17500 8708 17556 8718
rect 17052 7812 17108 7822
rect 16604 7250 16660 7262
rect 16604 7198 16606 7250
rect 16658 7198 16660 7250
rect 16604 6804 16660 7198
rect 17052 7028 17108 7756
rect 17052 6962 17108 6972
rect 17276 7028 17332 7038
rect 16828 6916 16884 6926
rect 16716 6804 16772 6814
rect 16604 6802 16772 6804
rect 16604 6750 16718 6802
rect 16770 6750 16772 6802
rect 16604 6748 16772 6750
rect 16604 5348 16660 6748
rect 16716 6738 16772 6748
rect 16716 6356 16772 6366
rect 16828 6356 16884 6860
rect 17276 6802 17332 6972
rect 17276 6750 17278 6802
rect 17330 6750 17332 6802
rect 17276 6738 17332 6750
rect 16772 6300 16884 6356
rect 17388 6468 17444 6478
rect 16716 6290 16772 6300
rect 16604 5282 16660 5292
rect 17388 4900 17444 6412
rect 17500 6020 17556 8652
rect 18284 8148 18340 8988
rect 18396 8370 18452 10332
rect 18620 10322 18676 10332
rect 18844 10052 18900 10062
rect 18844 9938 18900 9996
rect 18844 9886 18846 9938
rect 18898 9886 18900 9938
rect 18844 9874 18900 9886
rect 19292 9380 19348 12910
rect 19404 12290 19460 13132
rect 19964 13122 20020 13132
rect 20188 13636 20244 13646
rect 19404 12238 19406 12290
rect 19458 12238 19460 12290
rect 19404 12226 19460 12238
rect 20076 12066 20132 12078
rect 20076 12014 20078 12066
rect 20130 12014 20132 12066
rect 20076 11732 20132 12014
rect 20076 11666 20132 11676
rect 20188 11508 20244 13580
rect 20076 11452 20244 11508
rect 20300 12180 20356 12190
rect 19516 11396 19572 11406
rect 19516 10722 19572 11340
rect 19628 11396 19684 11406
rect 19628 11394 19908 11396
rect 19628 11342 19630 11394
rect 19682 11342 19908 11394
rect 19628 11340 19908 11342
rect 19628 11330 19684 11340
rect 19516 10670 19518 10722
rect 19570 10670 19572 10722
rect 19516 10658 19572 10670
rect 19292 9314 19348 9324
rect 19404 10612 19460 10622
rect 19404 9268 19460 10556
rect 19404 9202 19460 9212
rect 18620 9156 18676 9166
rect 18620 9042 18676 9100
rect 18620 8990 18622 9042
rect 18674 8990 18676 9042
rect 18620 8978 18676 8990
rect 18620 8428 18900 8484
rect 18396 8318 18398 8370
rect 18450 8318 18452 8370
rect 18396 8306 18452 8318
rect 18508 8372 18564 8382
rect 18620 8372 18676 8428
rect 18508 8370 18676 8372
rect 18508 8318 18510 8370
rect 18562 8318 18676 8370
rect 18508 8316 18676 8318
rect 18844 8372 18900 8428
rect 18844 8316 19012 8372
rect 18508 8306 18564 8316
rect 18732 8260 18788 8270
rect 18956 8260 19012 8316
rect 19068 8260 19124 8270
rect 18732 8258 18900 8260
rect 18732 8206 18734 8258
rect 18786 8206 18900 8258
rect 18732 8204 18900 8206
rect 18956 8258 19236 8260
rect 18956 8206 19070 8258
rect 19122 8206 19236 8258
rect 18956 8204 19236 8206
rect 18732 8194 18788 8204
rect 18284 8092 18564 8148
rect 17612 7364 17668 7374
rect 17612 6468 17668 7308
rect 17724 7364 17780 7374
rect 18284 7364 18340 7374
rect 17724 7362 18284 7364
rect 17724 7310 17726 7362
rect 17778 7310 18284 7362
rect 17724 7308 18284 7310
rect 17724 7298 17780 7308
rect 18284 7270 18340 7308
rect 18396 7250 18452 7262
rect 18396 7198 18398 7250
rect 18450 7198 18452 7250
rect 18396 6804 18452 7198
rect 18396 6738 18452 6748
rect 18284 6692 18340 6702
rect 17612 6402 17668 6412
rect 17948 6690 18340 6692
rect 17948 6638 18286 6690
rect 18338 6638 18340 6690
rect 17948 6636 18340 6638
rect 17500 5954 17556 5964
rect 17388 4834 17444 4844
rect 16828 4676 16884 4686
rect 16828 2436 16884 4620
rect 17948 4562 18004 6636
rect 18284 6626 18340 6636
rect 17948 4510 17950 4562
rect 18002 4510 18004 4562
rect 17948 4498 18004 4510
rect 18284 4338 18340 4350
rect 18284 4286 18286 4338
rect 18338 4286 18340 4338
rect 17948 3668 18004 3678
rect 17948 3574 18004 3612
rect 18172 3556 18228 3566
rect 18172 2884 18228 3500
rect 18284 3556 18340 4286
rect 18508 4226 18564 8092
rect 18620 7474 18676 7486
rect 18620 7422 18622 7474
rect 18674 7422 18676 7474
rect 18620 6914 18676 7422
rect 18732 7476 18788 7486
rect 18844 7476 18900 8204
rect 19068 8194 19124 8204
rect 18956 8036 19012 8046
rect 18956 8034 19124 8036
rect 18956 7982 18958 8034
rect 19010 7982 19124 8034
rect 18956 7980 19124 7982
rect 18956 7970 19012 7980
rect 18956 7476 19012 7486
rect 18844 7474 19012 7476
rect 18844 7422 18958 7474
rect 19010 7422 19012 7474
rect 18844 7420 19012 7422
rect 18732 7252 18788 7420
rect 18956 7410 19012 7420
rect 18844 7252 18900 7262
rect 18732 7250 18900 7252
rect 18732 7198 18846 7250
rect 18898 7198 18900 7250
rect 18732 7196 18900 7198
rect 18844 7186 18900 7196
rect 19068 7028 19124 7980
rect 18620 6862 18622 6914
rect 18674 6862 18676 6914
rect 18620 6850 18676 6862
rect 18732 6972 19124 7028
rect 18732 6802 18788 6972
rect 18732 6750 18734 6802
rect 18786 6750 18788 6802
rect 18732 6738 18788 6750
rect 18844 6804 18900 6814
rect 18844 6690 18900 6748
rect 18844 6638 18846 6690
rect 18898 6638 18900 6690
rect 18844 6626 18900 6638
rect 18508 4174 18510 4226
rect 18562 4174 18564 4226
rect 18508 4162 18564 4174
rect 18620 6580 18676 6590
rect 18396 3556 18452 3566
rect 18284 3554 18452 3556
rect 18284 3502 18398 3554
rect 18450 3502 18452 3554
rect 18284 3500 18452 3502
rect 18284 3444 18340 3500
rect 18396 3490 18452 3500
rect 18284 3378 18340 3388
rect 18172 2818 18228 2828
rect 17164 2660 17220 2670
rect 16828 2370 16884 2380
rect 16940 2548 16996 2558
rect 16828 1764 16884 1774
rect 16492 1586 16548 1596
rect 16716 1652 16772 1662
rect 16716 532 16772 1596
rect 16716 466 16772 476
rect 16828 420 16884 1708
rect 16940 1204 16996 2492
rect 17052 1764 17108 1774
rect 17052 1428 17108 1708
rect 17052 1362 17108 1372
rect 16940 1138 16996 1148
rect 17164 868 17220 2604
rect 17164 802 17220 812
rect 16828 354 16884 364
rect 17500 196 17556 206
rect 17500 112 17556 140
rect 18620 196 18676 6524
rect 19180 6356 19236 8204
rect 19628 7586 19684 7598
rect 19628 7534 19630 7586
rect 19682 7534 19684 7586
rect 19292 7476 19348 7486
rect 19628 7476 19684 7534
rect 19292 7474 19684 7476
rect 19292 7422 19294 7474
rect 19346 7422 19684 7474
rect 19292 7420 19684 7422
rect 19292 7410 19348 7420
rect 19740 7364 19796 7374
rect 19740 7270 19796 7308
rect 19852 6580 19908 11340
rect 20076 10610 20132 11452
rect 20076 10558 20078 10610
rect 20130 10558 20132 10610
rect 20076 10546 20132 10558
rect 20188 11284 20244 11294
rect 20076 10164 20132 10174
rect 19964 8820 20020 8830
rect 19964 7698 20020 8764
rect 19964 7646 19966 7698
rect 20018 7646 20020 7698
rect 19964 7634 20020 7646
rect 19852 6514 19908 6524
rect 20076 6356 20132 10108
rect 20188 9828 20244 11228
rect 20300 10388 20356 12124
rect 20412 11506 20468 14112
rect 20636 13748 20692 13758
rect 20524 12964 20580 12974
rect 20524 12870 20580 12908
rect 20412 11454 20414 11506
rect 20466 11454 20468 11506
rect 20412 11442 20468 11454
rect 20300 10322 20356 10332
rect 20188 9762 20244 9772
rect 20300 9716 20356 9726
rect 20300 8260 20356 9660
rect 20300 8194 20356 8204
rect 20524 9716 20580 9726
rect 20412 8036 20468 8046
rect 20524 8036 20580 9660
rect 20636 9714 20692 13692
rect 20748 13300 20804 13310
rect 20748 9828 20804 13244
rect 20860 12516 20916 14112
rect 20860 12450 20916 12460
rect 20860 12292 20916 12302
rect 20860 12198 20916 12236
rect 21084 11060 21140 14140
rect 21280 14112 21392 14224
rect 21728 14112 21840 14224
rect 22176 14112 22288 14224
rect 22624 14112 22736 14224
rect 23072 14112 23184 14224
rect 23520 14112 23632 14224
rect 23968 14112 24080 14224
rect 24416 14112 24528 14224
rect 24864 14112 24976 14224
rect 25312 14112 25424 14224
rect 25760 14112 25872 14224
rect 26208 14112 26320 14224
rect 26656 14112 26768 14224
rect 27104 14112 27216 14224
rect 27552 14112 27664 14224
rect 28000 14112 28112 14224
rect 28448 14112 28560 14224
rect 28896 14112 29008 14224
rect 29344 14112 29456 14224
rect 29792 14112 29904 14224
rect 30240 14112 30352 14224
rect 30688 14112 30800 14224
rect 31136 14112 31248 14224
rect 31584 14112 31696 14224
rect 32032 14112 32144 14224
rect 32480 14112 32592 14224
rect 32928 14112 33040 14224
rect 33376 14112 33488 14224
rect 33824 14112 33936 14224
rect 34272 14112 34384 14224
rect 34524 14196 34580 14206
rect 21196 13300 21252 13310
rect 21196 11620 21252 13244
rect 21308 12740 21364 14112
rect 21308 12674 21364 12684
rect 21420 13860 21476 13870
rect 21420 12628 21476 13804
rect 21532 12852 21588 12862
rect 21756 12852 21812 14112
rect 21532 12850 21812 12852
rect 21532 12798 21534 12850
rect 21586 12798 21812 12850
rect 21532 12796 21812 12798
rect 22092 12962 22148 12974
rect 22092 12910 22094 12962
rect 22146 12910 22148 12962
rect 21532 12786 21588 12796
rect 21980 12740 22036 12750
rect 21644 12628 21700 12638
rect 21420 12572 21588 12628
rect 21308 12404 21364 12414
rect 21308 11844 21364 12348
rect 21420 12180 21476 12190
rect 21420 12086 21476 12124
rect 21308 11788 21476 11844
rect 21196 11564 21364 11620
rect 21196 11396 21252 11406
rect 21196 11302 21252 11340
rect 20748 9762 20804 9772
rect 20860 11004 21140 11060
rect 20636 9662 20638 9714
rect 20690 9662 20692 9714
rect 20636 9650 20692 9662
rect 20860 9156 20916 11004
rect 21084 10500 21140 10510
rect 21084 10406 21140 10444
rect 21084 10276 21140 10286
rect 21084 10050 21140 10220
rect 21084 9998 21086 10050
rect 21138 9998 21140 10050
rect 21084 9986 21140 9998
rect 20860 9090 20916 9100
rect 20972 9826 21028 9838
rect 20972 9774 20974 9826
rect 21026 9774 21028 9826
rect 20972 9154 21028 9774
rect 21308 9268 21364 11564
rect 20972 9102 20974 9154
rect 21026 9102 21028 9154
rect 20972 9090 21028 9102
rect 21196 9212 21364 9268
rect 20468 7980 20580 8036
rect 20636 8036 20692 8046
rect 20412 7970 20468 7980
rect 19180 6290 19236 6300
rect 19852 6300 20132 6356
rect 19068 4226 19124 4238
rect 19068 4174 19070 4226
rect 19122 4174 19124 4226
rect 19068 3780 19124 4174
rect 19068 3714 19124 3724
rect 19180 3892 19236 3902
rect 19180 3442 19236 3836
rect 19628 3780 19684 3790
rect 19628 3686 19684 3724
rect 19180 3390 19182 3442
rect 19234 3390 19236 3442
rect 19180 3378 19236 3390
rect 19852 2660 19908 6300
rect 20524 5908 20580 5918
rect 20300 5796 20356 5806
rect 20188 4564 20244 4574
rect 19852 2594 19908 2604
rect 20076 3556 20132 3566
rect 20076 2548 20132 3500
rect 20076 2482 20132 2492
rect 20188 1764 20244 4508
rect 18620 130 18676 140
rect 19516 1708 20244 1764
rect 19516 112 19572 1708
rect 15820 28 16212 84
rect 17472 0 17584 112
rect 19488 0 19600 112
rect 20300 84 20356 5740
rect 20412 5236 20468 5246
rect 20412 1428 20468 5180
rect 20412 1362 20468 1372
rect 20524 532 20580 5852
rect 20636 2996 20692 7980
rect 21196 7924 21252 9212
rect 21308 9044 21364 9054
rect 21308 8950 21364 8988
rect 21196 7858 21252 7868
rect 21308 8148 21364 8158
rect 21308 7364 21364 8092
rect 21196 7252 21252 7262
rect 20636 2930 20692 2940
rect 20748 6580 20804 6590
rect 20748 2772 20804 6524
rect 21196 6468 21252 7196
rect 21196 6402 21252 6412
rect 21308 6690 21364 7308
rect 21308 6638 21310 6690
rect 21362 6638 21364 6690
rect 21308 5460 21364 6638
rect 21196 5404 21364 5460
rect 21196 5012 21252 5404
rect 21308 5236 21364 5246
rect 21420 5236 21476 11788
rect 21532 9938 21588 12572
rect 21532 9886 21534 9938
rect 21586 9886 21588 9938
rect 21532 9874 21588 9886
rect 21644 9044 21700 12572
rect 21868 12516 21924 12526
rect 21868 10722 21924 12460
rect 21980 11506 22036 12684
rect 21980 11454 21982 11506
rect 22034 11454 22036 11506
rect 21980 11442 22036 11454
rect 21868 10670 21870 10722
rect 21922 10670 21924 10722
rect 21868 10658 21924 10670
rect 21980 10612 22036 10622
rect 21980 9828 22036 10556
rect 22092 10052 22148 12910
rect 22204 12290 22260 14112
rect 22652 13186 22708 14112
rect 23100 13636 23156 14112
rect 23100 13580 23492 13636
rect 22652 13134 22654 13186
rect 22706 13134 22708 13186
rect 22652 13122 22708 13134
rect 22876 13412 22932 13422
rect 22204 12238 22206 12290
rect 22258 12238 22260 12290
rect 22204 12226 22260 12238
rect 22428 13076 22484 13086
rect 22204 12068 22260 12078
rect 22204 11060 22260 12012
rect 22204 10994 22260 11004
rect 22092 9986 22148 9996
rect 21868 9826 22036 9828
rect 21868 9774 21982 9826
rect 22034 9774 22036 9826
rect 21868 9772 22036 9774
rect 21644 8978 21700 8988
rect 21756 9268 21812 9278
rect 21532 8484 21588 8494
rect 21532 5460 21588 8428
rect 21756 8148 21812 9212
rect 21868 9042 21924 9772
rect 21980 9762 22036 9772
rect 21868 8990 21870 9042
rect 21922 8990 21924 9042
rect 21868 8978 21924 8990
rect 21980 8820 22036 8830
rect 21980 8726 22036 8764
rect 21756 8082 21812 8092
rect 22204 8372 22260 8382
rect 21644 7924 21700 7934
rect 21644 7364 21700 7868
rect 21644 7298 21700 7308
rect 21980 7364 22036 7374
rect 21644 7140 21700 7150
rect 21644 6802 21700 7084
rect 21644 6750 21646 6802
rect 21698 6750 21700 6802
rect 21644 5906 21700 6750
rect 21644 5854 21646 5906
rect 21698 5854 21700 5906
rect 21644 5842 21700 5854
rect 21532 5394 21588 5404
rect 21308 5234 21476 5236
rect 21308 5182 21310 5234
rect 21362 5182 21476 5234
rect 21308 5180 21476 5182
rect 21308 5170 21364 5180
rect 21868 5124 21924 5134
rect 21868 5030 21924 5068
rect 21196 4956 21364 5012
rect 20972 4452 21028 4462
rect 20972 4228 21028 4396
rect 21308 4338 21364 4956
rect 21308 4286 21310 4338
rect 21362 4286 21364 4338
rect 21308 4274 21364 4286
rect 21532 4676 21588 4686
rect 20972 4162 21028 4172
rect 21196 4228 21252 4238
rect 21196 3556 21252 4172
rect 21196 3490 21252 3500
rect 20748 2706 20804 2716
rect 21532 2660 21588 4620
rect 21756 4226 21812 4238
rect 21756 4174 21758 4226
rect 21810 4174 21812 4226
rect 21756 4004 21812 4174
rect 21644 2772 21700 2782
rect 21756 2772 21812 3948
rect 21980 3556 22036 7308
rect 22204 6018 22260 8316
rect 22204 5966 22206 6018
rect 22258 5966 22260 6018
rect 22204 5954 22260 5966
rect 22316 8260 22372 8270
rect 22316 5796 22372 8204
rect 22428 6692 22484 13020
rect 22652 12516 22708 12526
rect 22428 6626 22484 6636
rect 22540 10500 22596 10510
rect 22204 5740 22372 5796
rect 22428 6020 22484 6030
rect 22540 6020 22596 10444
rect 22652 9716 22708 12460
rect 22764 11394 22820 11406
rect 22764 11342 22766 11394
rect 22818 11342 22820 11394
rect 22764 10500 22820 11342
rect 22764 10434 22820 10444
rect 22652 9650 22708 9660
rect 22652 9042 22708 9054
rect 22652 8990 22654 9042
rect 22706 8990 22708 9042
rect 22652 6916 22708 8990
rect 22764 8708 22820 8718
rect 22764 8372 22820 8652
rect 22764 8306 22820 8316
rect 22876 7140 22932 13356
rect 23212 13412 23268 13422
rect 22988 12964 23044 12974
rect 22988 12178 23044 12908
rect 23212 12516 23268 13356
rect 23436 12964 23492 13580
rect 23548 13188 23604 14112
rect 23772 14084 23828 14094
rect 23548 13122 23604 13132
rect 23660 13748 23716 13758
rect 23436 12908 23604 12964
rect 23436 12516 23492 12526
rect 23212 12450 23268 12460
rect 23324 12460 23436 12516
rect 22988 12126 22990 12178
rect 23042 12126 23044 12178
rect 22988 12114 23044 12126
rect 23100 11396 23156 11406
rect 22988 10388 23044 10398
rect 22988 10052 23044 10332
rect 22988 9986 23044 9996
rect 23100 9716 23156 11340
rect 23324 10612 23380 12460
rect 23436 12450 23492 12460
rect 23548 12402 23604 12908
rect 23548 12350 23550 12402
rect 23602 12350 23604 12402
rect 23548 12338 23604 12350
rect 23548 11844 23604 11854
rect 23548 11394 23604 11788
rect 23548 11342 23550 11394
rect 23602 11342 23604 11394
rect 23548 11330 23604 11342
rect 23660 10724 23716 13692
rect 23772 13076 23828 14028
rect 23884 13076 23940 13086
rect 23772 13074 23940 13076
rect 23772 13022 23886 13074
rect 23938 13022 23940 13074
rect 23772 13020 23940 13022
rect 23884 13010 23940 13020
rect 23996 13076 24052 14112
rect 24444 13524 24500 14112
rect 24892 13748 24948 14112
rect 24892 13692 25172 13748
rect 24332 13468 24500 13524
rect 24332 13078 24388 13468
rect 24464 13356 24728 13366
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 25116 13300 25172 13692
rect 24464 13290 24728 13300
rect 24892 13244 25172 13300
rect 24332 13022 24612 13078
rect 23996 13010 24052 13020
rect 23772 12852 23828 12862
rect 24444 12852 24500 12862
rect 23828 12850 24500 12852
rect 23828 12798 24446 12850
rect 24498 12798 24500 12850
rect 23828 12796 24500 12798
rect 23772 12786 23828 12796
rect 24444 12786 24500 12796
rect 24556 12628 24612 13022
rect 24780 13076 24836 13086
rect 23804 12572 24068 12582
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 23804 12506 24068 12516
rect 24220 12572 24612 12628
rect 24668 12628 24724 12638
rect 24220 11508 24276 12572
rect 24556 12180 24612 12190
rect 24668 12180 24724 12572
rect 24556 12178 24724 12180
rect 24556 12126 24558 12178
rect 24610 12126 24724 12178
rect 24556 12124 24724 12126
rect 24556 12114 24612 12124
rect 24780 11956 24836 13020
rect 24892 12292 24948 13244
rect 25116 12292 25172 12302
rect 25340 12292 25396 14112
rect 25676 12852 25732 12862
rect 24892 12236 25060 12292
rect 24892 11956 24948 11966
rect 24780 11954 24948 11956
rect 24780 11902 24894 11954
rect 24946 11902 24948 11954
rect 24780 11900 24948 11902
rect 24892 11890 24948 11900
rect 24464 11788 24728 11798
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24464 11722 24728 11732
rect 24220 11452 24724 11508
rect 23996 11284 24052 11294
rect 23996 11190 24052 11228
rect 24444 11172 24500 11182
rect 24332 11116 24444 11172
rect 23804 11004 24068 11014
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 23804 10938 24068 10948
rect 23772 10724 23828 10734
rect 24332 10724 24388 11116
rect 24444 11106 24500 11116
rect 23660 10722 23828 10724
rect 23660 10670 23774 10722
rect 23826 10670 23828 10722
rect 23660 10668 23828 10670
rect 23772 10658 23828 10668
rect 24108 10668 24388 10724
rect 23212 10556 23380 10612
rect 23212 10276 23268 10556
rect 23212 10210 23268 10220
rect 23324 10386 23380 10398
rect 23324 10334 23326 10386
rect 23378 10334 23380 10386
rect 23324 10164 23380 10334
rect 23324 10098 23380 10108
rect 23436 10276 23492 10286
rect 23100 9650 23156 9660
rect 23212 10052 23268 10062
rect 23212 9042 23268 9996
rect 23436 9940 23492 10220
rect 23996 10052 24052 10062
rect 23996 9958 24052 9996
rect 23212 8990 23214 9042
rect 23266 8990 23268 9042
rect 23212 8978 23268 8990
rect 23324 9884 23492 9940
rect 23100 8820 23156 8830
rect 22876 7084 23044 7140
rect 22876 6916 22932 6926
rect 22652 6914 22932 6916
rect 22652 6862 22878 6914
rect 22930 6862 22932 6914
rect 22652 6860 22932 6862
rect 22652 6356 22708 6860
rect 22876 6850 22932 6860
rect 22652 6290 22708 6300
rect 22988 6356 23044 7084
rect 22988 6290 23044 6300
rect 22540 5964 22932 6020
rect 22092 5684 22148 5694
rect 22092 4340 22148 5628
rect 22092 4274 22148 4284
rect 21980 3490 22036 3500
rect 22204 3388 22260 5740
rect 22316 5124 22372 5134
rect 22316 5030 22372 5068
rect 22428 4564 22484 5964
rect 22652 5796 22708 5806
rect 22540 5124 22596 5134
rect 22540 4788 22596 5068
rect 22652 5012 22708 5740
rect 22652 5010 22820 5012
rect 22652 4958 22654 5010
rect 22706 4958 22820 5010
rect 22652 4956 22820 4958
rect 22652 4946 22708 4956
rect 22540 4722 22596 4732
rect 22428 4508 22596 4564
rect 21644 2770 21812 2772
rect 21644 2718 21646 2770
rect 21698 2718 21812 2770
rect 21644 2716 21812 2718
rect 21868 3332 21924 3342
rect 21644 2706 21700 2716
rect 21532 2594 21588 2604
rect 21756 2436 21812 2446
rect 21644 1876 21700 1886
rect 21644 1652 21700 1820
rect 21644 1586 21700 1596
rect 20524 466 20580 476
rect 21532 1204 21588 1214
rect 21532 112 21588 1148
rect 20300 18 20356 28
rect 21504 0 21616 112
rect 21756 84 21812 2380
rect 21868 1316 21924 3276
rect 21980 3332 22260 3388
rect 22428 4340 22484 4350
rect 21980 2996 22036 3332
rect 21980 2930 22036 2940
rect 21868 1250 21924 1260
rect 22092 2658 22148 2670
rect 22092 2606 22094 2658
rect 22146 2606 22148 2658
rect 22092 1316 22148 2606
rect 22428 1988 22484 4284
rect 22540 2436 22596 4508
rect 22540 2370 22596 2380
rect 22652 3444 22708 3454
rect 22428 1922 22484 1932
rect 22092 1250 22148 1260
rect 22652 868 22708 3388
rect 22764 2548 22820 4956
rect 22876 4340 22932 5964
rect 22988 5234 23044 5246
rect 22988 5182 22990 5234
rect 23042 5182 23044 5234
rect 22988 4562 23044 5182
rect 22988 4510 22990 4562
rect 23042 4510 23044 4562
rect 22988 4498 23044 4510
rect 22876 4284 23044 4340
rect 22764 2482 22820 2492
rect 22876 3444 22932 3454
rect 22876 980 22932 3388
rect 22876 914 22932 924
rect 22652 802 22708 812
rect 22988 308 23044 4284
rect 23100 3220 23156 8764
rect 23212 5572 23268 5582
rect 23324 5572 23380 9884
rect 23548 9828 23604 9838
rect 23548 9714 23604 9772
rect 23548 9662 23550 9714
rect 23602 9662 23604 9714
rect 23548 9650 23604 9662
rect 24108 9604 24164 10668
rect 24668 10610 24724 11452
rect 24668 10558 24670 10610
rect 24722 10558 24724 10610
rect 24668 10546 24724 10558
rect 24220 10498 24276 10510
rect 24220 10446 24222 10498
rect 24274 10446 24276 10498
rect 24220 10276 24276 10446
rect 24892 10500 24948 10510
rect 24220 10210 24276 10220
rect 24464 10220 24728 10230
rect 24332 10164 24388 10174
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24464 10154 24728 10164
rect 24332 10052 24388 10108
rect 24332 9996 24612 10052
rect 24556 9940 24612 9996
rect 24556 9874 24612 9884
rect 23660 9548 24164 9604
rect 23548 9380 23604 9390
rect 23548 6916 23604 9324
rect 23660 7812 23716 9548
rect 24220 9492 24276 9502
rect 23804 9436 24068 9446
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 23804 9370 24068 9380
rect 24108 9044 24164 9054
rect 24108 8950 24164 8988
rect 24220 8484 24276 9436
rect 24444 9268 24500 9278
rect 24332 9212 24444 9268
rect 24332 8596 24388 9212
rect 24444 9202 24500 9212
rect 24464 8652 24728 8662
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24464 8586 24728 8596
rect 24332 8530 24388 8540
rect 23996 8428 24276 8484
rect 24892 8484 24948 10444
rect 25004 10052 25060 12236
rect 25116 11506 25172 12236
rect 25116 11454 25118 11506
rect 25170 11454 25172 11506
rect 25116 11442 25172 11454
rect 25228 12236 25396 12292
rect 25452 12850 25732 12852
rect 25452 12798 25678 12850
rect 25730 12798 25732 12850
rect 25452 12796 25732 12798
rect 25228 10610 25284 12236
rect 25340 11956 25396 11966
rect 25340 11862 25396 11900
rect 25228 10558 25230 10610
rect 25282 10558 25284 10610
rect 25228 10546 25284 10558
rect 25228 10164 25284 10174
rect 25116 10052 25172 10062
rect 25004 10050 25172 10052
rect 25004 9998 25118 10050
rect 25170 9998 25172 10050
rect 25004 9996 25172 9998
rect 25116 9986 25172 9996
rect 25228 9604 25284 10108
rect 25228 9538 25284 9548
rect 25452 9268 25508 12796
rect 25676 12786 25732 12796
rect 25564 12404 25620 12414
rect 25564 11956 25620 12348
rect 25564 11890 25620 11900
rect 25676 11620 25732 11630
rect 25788 11620 25844 14112
rect 26012 13860 26068 13870
rect 25900 12066 25956 12078
rect 25900 12014 25902 12066
rect 25954 12014 25956 12066
rect 25900 11844 25956 12014
rect 25900 11778 25956 11788
rect 25676 11618 25844 11620
rect 25676 11566 25678 11618
rect 25730 11566 25844 11618
rect 25676 11564 25844 11566
rect 26012 11620 26068 13804
rect 26236 13636 26292 14112
rect 26236 13570 26292 13580
rect 26236 13188 26292 13198
rect 26684 13188 26740 14112
rect 26908 14084 26964 14094
rect 26236 13186 26740 13188
rect 26236 13134 26238 13186
rect 26290 13134 26740 13186
rect 26236 13132 26740 13134
rect 26796 13188 26852 13198
rect 26236 13122 26292 13132
rect 26572 12852 26628 12862
rect 25676 11554 25732 11564
rect 26012 11554 26068 11564
rect 26124 12850 26628 12852
rect 26124 12798 26574 12850
rect 26626 12798 26628 12850
rect 26124 12796 26628 12798
rect 26012 11394 26068 11406
rect 26012 11342 26014 11394
rect 26066 11342 26068 11394
rect 25452 9202 25508 9212
rect 25564 10722 25620 10734
rect 25564 10670 25566 10722
rect 25618 10670 25620 10722
rect 25564 9940 25620 10670
rect 25564 9044 25620 9884
rect 25564 8978 25620 8988
rect 25676 9714 25732 9726
rect 25676 9662 25678 9714
rect 25730 9662 25732 9714
rect 25228 8932 25284 8942
rect 25284 8876 25396 8932
rect 25228 8866 25284 8876
rect 24892 8428 25284 8484
rect 23996 8036 24052 8428
rect 25228 8372 25284 8428
rect 25340 8372 25396 8876
rect 25340 8316 25620 8372
rect 25228 8306 25284 8316
rect 24220 8260 24276 8270
rect 24220 8148 24276 8204
rect 24220 8092 24388 8148
rect 24332 8036 24388 8092
rect 24780 8036 24836 8046
rect 23996 7980 24276 8036
rect 24332 7980 24780 8036
rect 23804 7868 24068 7878
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 23804 7802 24068 7812
rect 23660 7746 23716 7756
rect 24220 7140 24276 7980
rect 24780 7970 24836 7980
rect 24444 7700 24500 7710
rect 24220 7074 24276 7084
rect 24332 7644 24444 7700
rect 24108 6916 24164 6926
rect 23548 6860 23716 6916
rect 23548 6692 23604 6702
rect 23548 6244 23604 6636
rect 23548 6178 23604 6188
rect 23268 5516 23380 5572
rect 23212 5234 23268 5516
rect 23212 5182 23214 5234
rect 23266 5182 23268 5234
rect 23212 5170 23268 5182
rect 23660 4340 23716 6860
rect 24164 6860 24276 6916
rect 24108 6850 24164 6860
rect 24220 6356 24276 6860
rect 24332 6692 24388 7644
rect 24444 7634 24500 7644
rect 25228 7700 25284 7710
rect 24464 7084 24728 7094
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 24464 7018 24728 7028
rect 25116 6804 25172 6814
rect 25004 6802 25172 6804
rect 25004 6750 25118 6802
rect 25170 6750 25172 6802
rect 25004 6748 25172 6750
rect 24332 6626 24388 6636
rect 24780 6692 24836 6702
rect 24836 6636 24948 6692
rect 24780 6598 24836 6636
rect 23804 6300 24068 6310
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 24220 6290 24276 6300
rect 23804 6234 24068 6244
rect 24668 5684 24724 5722
rect 24668 5618 24724 5628
rect 24464 5516 24728 5526
rect 24332 5460 24388 5470
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24464 5450 24728 5460
rect 23804 4732 24068 4742
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 23804 4666 24068 4676
rect 24332 4676 24388 5404
rect 24332 4610 24388 4620
rect 23660 4274 23716 4284
rect 24892 4004 24948 6636
rect 25004 5684 25060 6748
rect 25116 6738 25172 6748
rect 25116 6018 25172 6030
rect 25116 5966 25118 6018
rect 25170 5966 25172 6018
rect 25116 5908 25172 5966
rect 25116 5842 25172 5852
rect 25228 5684 25284 7644
rect 25340 7252 25396 7262
rect 25340 6916 25396 7196
rect 25340 6850 25396 6860
rect 25564 6468 25620 8316
rect 25676 7252 25732 9662
rect 25676 7186 25732 7196
rect 25788 9492 25844 9502
rect 25788 6692 25844 9436
rect 25788 6626 25844 6636
rect 25900 9044 25956 9054
rect 25564 6412 25844 6468
rect 25452 6356 25508 6366
rect 25508 6300 25732 6356
rect 25452 6290 25508 6300
rect 25676 6018 25732 6300
rect 25676 5966 25678 6018
rect 25730 5966 25732 6018
rect 25676 5954 25732 5966
rect 25004 5618 25060 5628
rect 25116 5628 25284 5684
rect 25116 4228 25172 5628
rect 25116 4162 25172 4172
rect 25228 5460 25284 5470
rect 24464 3948 24728 3958
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24892 3938 24948 3948
rect 24464 3882 24728 3892
rect 23100 3154 23156 3164
rect 23324 3556 23380 3566
rect 23212 2996 23268 3006
rect 23212 980 23268 2940
rect 23324 1764 23380 3500
rect 24332 3220 24388 3230
rect 23804 3164 24068 3174
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 23804 3098 24068 3108
rect 24220 3108 24276 3118
rect 23436 2884 23492 2894
rect 23436 2548 23492 2828
rect 23436 2482 23492 2492
rect 23996 2884 24052 2894
rect 23996 2098 24052 2828
rect 24108 2212 24164 2222
rect 24220 2212 24276 3052
rect 24332 2436 24388 3164
rect 25228 3108 25284 5404
rect 25340 4564 25396 4574
rect 25340 3780 25396 4508
rect 25340 3714 25396 3724
rect 25452 4004 25508 4014
rect 25452 3556 25508 3948
rect 25228 3042 25284 3052
rect 25340 3500 25508 3556
rect 25340 2884 25396 3500
rect 25788 3388 25844 6412
rect 25452 3332 25844 3388
rect 25452 3108 25508 3332
rect 25452 3042 25508 3052
rect 24892 2882 25396 2884
rect 24892 2830 25342 2882
rect 25394 2830 25396 2882
rect 24892 2828 25396 2830
rect 24332 2370 24388 2380
rect 24464 2380 24728 2390
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24464 2314 24728 2324
rect 24164 2156 24276 2212
rect 24108 2146 24164 2156
rect 23996 2046 23998 2098
rect 24050 2046 24052 2098
rect 23996 2034 24052 2046
rect 23548 1988 23604 1998
rect 23548 1894 23604 1932
rect 24780 1988 24836 1998
rect 24892 1988 24948 2828
rect 25340 2818 25396 2828
rect 25676 2660 25732 2670
rect 25564 2548 25620 2558
rect 24780 1986 24948 1988
rect 24780 1934 24782 1986
rect 24834 1934 24948 1986
rect 24780 1932 24948 1934
rect 25116 2098 25172 2110
rect 25116 2046 25118 2098
rect 25170 2046 25172 2098
rect 25116 1988 25172 2046
rect 24780 1922 24836 1932
rect 25116 1922 25172 1932
rect 23324 1698 23380 1708
rect 24332 1652 24388 1662
rect 23804 1596 24068 1606
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 23804 1530 24068 1540
rect 23212 914 23268 924
rect 23548 1428 23604 1438
rect 22988 242 23044 252
rect 23548 112 23604 1372
rect 24332 868 24388 1596
rect 24332 802 24388 812
rect 24464 812 24728 822
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24464 746 24728 756
rect 25564 112 25620 2492
rect 25676 1202 25732 2604
rect 25900 1428 25956 8988
rect 26012 6244 26068 11342
rect 26124 10052 26180 12796
rect 26572 12786 26628 12796
rect 26236 12066 26292 12078
rect 26236 12014 26238 12066
rect 26290 12014 26292 12066
rect 26236 11394 26292 12014
rect 26236 11342 26238 11394
rect 26290 11342 26292 11394
rect 26236 11330 26292 11342
rect 26684 11620 26740 11630
rect 26572 11172 26628 11182
rect 26124 9986 26180 9996
rect 26236 11170 26628 11172
rect 26236 11118 26574 11170
rect 26626 11118 26628 11170
rect 26236 11116 26628 11118
rect 26236 10722 26292 11116
rect 26572 11106 26628 11116
rect 26236 10670 26238 10722
rect 26290 10670 26292 10722
rect 26012 6178 26068 6188
rect 26124 9828 26180 9838
rect 26012 4788 26068 4798
rect 26012 3332 26068 4732
rect 26012 3266 26068 3276
rect 26124 1540 26180 9772
rect 26236 8148 26292 10670
rect 26684 10498 26740 11564
rect 26684 10446 26686 10498
rect 26738 10446 26740 10498
rect 26684 10434 26740 10446
rect 26796 10276 26852 13132
rect 26908 11396 26964 14028
rect 27132 13186 27188 14112
rect 27132 13134 27134 13186
rect 27186 13134 27188 13186
rect 27132 13122 27188 13134
rect 27468 13412 27524 13422
rect 26908 11330 26964 11340
rect 27020 12852 27076 12862
rect 26796 10210 26852 10220
rect 26908 10948 26964 10958
rect 26908 10052 26964 10892
rect 26908 9986 26964 9996
rect 27020 9828 27076 12796
rect 27244 12290 27300 12302
rect 27244 12238 27246 12290
rect 27298 12238 27300 12290
rect 26908 9772 27076 9828
rect 27132 10388 27188 10398
rect 26684 9602 26740 9614
rect 26684 9550 26686 9602
rect 26738 9550 26740 9602
rect 26684 9042 26740 9550
rect 26684 8990 26686 9042
rect 26738 8990 26740 9042
rect 26684 8978 26740 8990
rect 26236 8082 26292 8092
rect 26348 8932 26404 8942
rect 26348 7364 26404 8876
rect 26908 8820 26964 9772
rect 26908 8754 26964 8764
rect 27020 9602 27076 9614
rect 27020 9550 27022 9602
rect 27074 9550 27076 9602
rect 26348 7298 26404 7308
rect 27020 7812 27076 9550
rect 27132 8820 27188 10332
rect 27244 10052 27300 12238
rect 27468 10612 27524 13356
rect 27580 13188 27636 14112
rect 28028 13524 28084 14112
rect 28028 13458 28084 13468
rect 27804 13188 27860 13198
rect 27580 13186 27860 13188
rect 27580 13134 27806 13186
rect 27858 13134 27860 13186
rect 27580 13132 27860 13134
rect 27804 13122 27860 13132
rect 27916 13076 27972 13086
rect 27580 11620 27636 11630
rect 27580 11526 27636 11564
rect 27916 10948 27972 13020
rect 28252 12964 28308 12974
rect 28140 11282 28196 11294
rect 28140 11230 28142 11282
rect 28194 11230 28196 11282
rect 27468 10546 27524 10556
rect 27580 10892 27972 10948
rect 28028 11060 28084 11070
rect 27580 10164 27636 10892
rect 27244 9492 27300 9996
rect 27244 9426 27300 9436
rect 27468 10108 27636 10164
rect 27692 10724 27748 10734
rect 27132 8754 27188 8764
rect 27244 8930 27300 8942
rect 27244 8878 27246 8930
rect 27298 8878 27300 8930
rect 27132 7812 27188 7822
rect 27020 7756 27132 7812
rect 26460 7252 26516 7262
rect 26348 6692 26404 6702
rect 26348 6598 26404 6636
rect 26236 6580 26292 6590
rect 26236 5906 26292 6524
rect 26460 6356 26516 7196
rect 27020 6804 27076 7756
rect 27132 7746 27188 7756
rect 26460 6290 26516 6300
rect 26908 6748 27076 6804
rect 26236 5854 26238 5906
rect 26290 5854 26292 5906
rect 26236 5842 26292 5854
rect 26348 6244 26404 6254
rect 26348 4676 26404 6188
rect 26908 5908 26964 6748
rect 27020 6580 27076 6590
rect 27020 6130 27076 6524
rect 27020 6078 27022 6130
rect 27074 6078 27076 6130
rect 27020 6066 27076 6078
rect 26796 5852 26964 5908
rect 26796 5796 26852 5852
rect 26796 5730 26852 5740
rect 26684 5682 26740 5694
rect 26684 5630 26686 5682
rect 26738 5630 26740 5682
rect 26348 4610 26404 4620
rect 26572 5236 26628 5246
rect 26572 4676 26628 5180
rect 26572 4610 26628 4620
rect 26684 4340 26740 5630
rect 27244 5460 27300 8878
rect 27468 8708 27524 10108
rect 27580 9940 27636 9950
rect 27580 9846 27636 9884
rect 27468 8642 27524 8652
rect 27692 8708 27748 10668
rect 27804 10386 27860 10398
rect 27804 10334 27806 10386
rect 27858 10334 27860 10386
rect 27804 9826 27860 10334
rect 28028 9940 28084 11004
rect 28140 10276 28196 11230
rect 28140 10210 28196 10220
rect 28252 10164 28308 12908
rect 28364 12850 28420 12862
rect 28364 12798 28366 12850
rect 28418 12798 28420 12850
rect 28364 11060 28420 12798
rect 28476 12180 28532 14112
rect 28924 13972 28980 14112
rect 28924 13906 28980 13916
rect 28812 13748 28868 13758
rect 28700 13636 28756 13646
rect 28476 12114 28532 12124
rect 28588 13524 28644 13534
rect 28588 11508 28644 13468
rect 28700 13186 28756 13580
rect 28700 13134 28702 13186
rect 28754 13134 28756 13186
rect 28700 13122 28756 13134
rect 28588 11442 28644 11452
rect 28700 12404 28756 12414
rect 28364 10994 28420 11004
rect 28588 10724 28644 10734
rect 28476 10388 28532 10398
rect 28588 10388 28644 10668
rect 28532 10332 28644 10388
rect 28700 10388 28756 12348
rect 28812 11620 28868 13692
rect 29036 13188 29092 13198
rect 28812 11554 28868 11564
rect 28924 12404 28980 12414
rect 28476 10322 28532 10332
rect 28700 10322 28756 10332
rect 28252 10098 28308 10108
rect 28028 9884 28420 9940
rect 27804 9774 27806 9826
rect 27858 9774 27860 9826
rect 27804 9762 27860 9774
rect 27692 8642 27748 8652
rect 27916 9492 27972 9502
rect 27916 8148 27972 9436
rect 28252 9268 28308 9278
rect 28028 8372 28084 8382
rect 28028 8278 28084 8316
rect 27916 8092 28084 8148
rect 27244 5394 27300 5404
rect 27692 6692 27748 6702
rect 27692 5906 27748 6636
rect 27692 5854 27694 5906
rect 27746 5854 27748 5906
rect 26684 4274 26740 4284
rect 26796 5236 26852 5246
rect 26796 3666 26852 5180
rect 27580 4340 27636 4350
rect 27580 4246 27636 4284
rect 27020 4226 27076 4238
rect 27020 4174 27022 4226
rect 27074 4174 27076 4226
rect 26908 3780 26964 3790
rect 27020 3780 27076 4174
rect 26908 3778 27076 3780
rect 26908 3726 26910 3778
rect 26962 3726 27076 3778
rect 26908 3724 27076 3726
rect 27244 4226 27300 4238
rect 27244 4174 27246 4226
rect 27298 4174 27300 4226
rect 27244 3778 27300 4174
rect 27244 3726 27246 3778
rect 27298 3726 27300 3778
rect 26908 3714 26964 3724
rect 27244 3714 27300 3726
rect 27356 4116 27412 4126
rect 26796 3614 26798 3666
rect 26850 3614 26852 3666
rect 26796 3388 26852 3614
rect 27356 3666 27412 4060
rect 27356 3614 27358 3666
rect 27410 3614 27412 3666
rect 27356 3388 27412 3614
rect 26348 3332 26852 3388
rect 26908 3332 27412 3388
rect 27468 4114 27524 4126
rect 27468 4062 27470 4114
rect 27522 4062 27524 4114
rect 27468 3332 27524 4062
rect 26348 2210 26404 3332
rect 26908 2994 26964 3332
rect 27468 3266 27524 3276
rect 26908 2942 26910 2994
rect 26962 2942 26964 2994
rect 26908 2930 26964 2942
rect 27580 3220 27636 3230
rect 26348 2158 26350 2210
rect 26402 2158 26404 2210
rect 26348 2146 26404 2158
rect 26796 2324 26852 2334
rect 26348 1540 26404 1550
rect 26124 1484 26348 1540
rect 26348 1474 26404 1484
rect 25900 1362 25956 1372
rect 25676 1150 25678 1202
rect 25730 1150 25732 1202
rect 25676 1138 25732 1150
rect 26796 1204 26852 2268
rect 26796 1138 26852 1148
rect 26124 1092 26180 1102
rect 26124 998 26180 1036
rect 27580 112 27636 3164
rect 27692 2772 27748 5854
rect 27804 5796 27860 5806
rect 27804 5702 27860 5740
rect 28028 3668 28084 8092
rect 28028 3602 28084 3612
rect 27692 2706 27748 2716
rect 28140 3108 28196 3118
rect 28140 2098 28196 3052
rect 28140 2046 28142 2098
rect 28194 2046 28196 2098
rect 28140 2034 28196 2046
rect 28252 1652 28308 9212
rect 28364 5572 28420 9884
rect 28812 9604 28868 9614
rect 28700 8372 28756 8382
rect 28476 8258 28532 8270
rect 28476 8206 28478 8258
rect 28530 8206 28532 8258
rect 28476 7364 28532 8206
rect 28700 8036 28756 8316
rect 28700 7970 28756 7980
rect 28476 7298 28532 7308
rect 28588 7250 28644 7262
rect 28588 7198 28590 7250
rect 28642 7198 28644 7250
rect 28476 6244 28532 6254
rect 28476 6018 28532 6188
rect 28476 5966 28478 6018
rect 28530 5966 28532 6018
rect 28476 5954 28532 5966
rect 28364 5506 28420 5516
rect 28476 4340 28532 4350
rect 28588 4340 28644 7198
rect 28812 6468 28868 9548
rect 28924 9044 28980 12348
rect 29036 11620 29092 13132
rect 29148 12852 29204 12862
rect 29148 12758 29204 12796
rect 29372 12180 29428 14112
rect 29820 13188 29876 14112
rect 30044 13188 30100 13198
rect 29820 13186 30100 13188
rect 29820 13134 30046 13186
rect 30098 13134 30100 13186
rect 29820 13132 30100 13134
rect 30044 13122 30100 13132
rect 29372 12114 29428 12124
rect 29484 12852 29540 12862
rect 29036 11554 29092 11564
rect 28924 8978 28980 8988
rect 29036 11396 29092 11406
rect 28924 8596 28980 8606
rect 28924 8370 28980 8540
rect 28924 8318 28926 8370
rect 28978 8318 28980 8370
rect 28924 8306 28980 8318
rect 29036 7812 29092 11340
rect 29484 10724 29540 12796
rect 30268 12740 30324 14112
rect 30716 13188 30772 14112
rect 30716 13122 30772 13132
rect 30828 13300 30884 13310
rect 30604 12850 30660 12862
rect 30604 12798 30606 12850
rect 30658 12798 30660 12850
rect 30268 12684 30548 12740
rect 30492 12178 30548 12684
rect 30492 12126 30494 12178
rect 30546 12126 30548 12178
rect 30492 12114 30548 12126
rect 30604 12068 30660 12798
rect 30604 12002 30660 12012
rect 30716 12292 30772 12302
rect 30044 11956 30100 11966
rect 29484 10658 29540 10668
rect 29820 10724 29876 10734
rect 28924 7756 29092 7812
rect 29148 10612 29204 10622
rect 28924 7700 28980 7756
rect 29148 7700 29204 10556
rect 29820 9492 29876 10668
rect 29820 9426 29876 9436
rect 29932 10610 29988 10622
rect 29932 10558 29934 10610
rect 29986 10558 29988 10610
rect 29708 8708 29764 8718
rect 28924 7634 28980 7644
rect 29036 7644 29204 7700
rect 29484 8260 29540 8270
rect 28924 7474 28980 7486
rect 28924 7422 28926 7474
rect 28978 7422 28980 7474
rect 28924 7364 28980 7422
rect 29036 7476 29092 7644
rect 29036 7410 29092 7420
rect 28924 7298 28980 7308
rect 29148 7362 29204 7374
rect 29148 7310 29150 7362
rect 29202 7310 29204 7362
rect 29148 6692 29204 7310
rect 29484 7362 29540 8204
rect 29484 7310 29486 7362
rect 29538 7310 29540 7362
rect 29484 7298 29540 7310
rect 29596 7476 29652 7486
rect 29148 6626 29204 6636
rect 29260 7252 29316 7262
rect 28812 6402 28868 6412
rect 29036 6468 29092 6478
rect 29036 5906 29092 6412
rect 29036 5854 29038 5906
rect 29090 5854 29092 5906
rect 29036 5796 29092 5854
rect 29036 5730 29092 5740
rect 29260 5796 29316 7196
rect 29260 5730 29316 5740
rect 28476 4338 28644 4340
rect 28476 4286 28478 4338
rect 28530 4286 28644 4338
rect 28476 4284 28644 4286
rect 28700 5460 28756 5470
rect 28476 4274 28532 4284
rect 28588 4116 28644 4126
rect 28588 4022 28644 4060
rect 28700 3780 28756 5404
rect 29036 4228 29092 4238
rect 28812 4116 28868 4126
rect 28812 4114 28980 4116
rect 28812 4062 28814 4114
rect 28866 4062 28980 4114
rect 28812 4060 28980 4062
rect 28812 4050 28868 4060
rect 28476 3724 28756 3780
rect 28476 2548 28532 3724
rect 28588 3554 28644 3566
rect 28588 3502 28590 3554
rect 28642 3502 28644 3554
rect 28588 3332 28644 3502
rect 28924 3554 28980 4060
rect 28924 3502 28926 3554
rect 28978 3502 28980 3554
rect 28924 3490 28980 3502
rect 28812 3444 28868 3454
rect 28812 3350 28868 3388
rect 28588 3266 28644 3276
rect 28924 2996 28980 3006
rect 28924 2884 28980 2940
rect 28476 2482 28532 2492
rect 28700 2882 28980 2884
rect 28700 2830 28926 2882
rect 28978 2830 28980 2882
rect 28700 2828 28980 2830
rect 28700 2210 28756 2828
rect 28924 2818 28980 2828
rect 28700 2158 28702 2210
rect 28754 2158 28756 2210
rect 28700 2146 28756 2158
rect 28812 2548 28868 2558
rect 28812 1764 28868 2492
rect 28252 1586 28308 1596
rect 28476 1708 28868 1764
rect 28476 644 28532 1708
rect 29036 1316 29092 4172
rect 29596 3780 29652 7420
rect 29708 7140 29764 8652
rect 29932 8428 29988 10558
rect 30044 10500 30100 11900
rect 30380 10500 30436 10510
rect 30044 10498 30436 10500
rect 30044 10446 30382 10498
rect 30434 10446 30436 10498
rect 30044 10444 30436 10446
rect 30044 10050 30100 10444
rect 30380 10434 30436 10444
rect 30044 9998 30046 10050
rect 30098 9998 30100 10050
rect 30044 9986 30100 9998
rect 30156 10164 30212 10174
rect 30156 9492 30212 10108
rect 30604 9716 30660 9726
rect 30604 9622 30660 9660
rect 30268 9492 30324 9502
rect 30156 9436 30268 9492
rect 30268 9426 30324 9436
rect 30716 8932 30772 12236
rect 30828 10724 30884 13244
rect 30828 10658 30884 10668
rect 30940 12740 30996 12750
rect 30828 10388 30884 10398
rect 30828 9044 30884 10332
rect 30828 8978 30884 8988
rect 30716 8866 30772 8876
rect 30940 8596 30996 12684
rect 30940 8530 30996 8540
rect 31052 12066 31108 12078
rect 31052 12014 31054 12066
rect 31106 12014 31108 12066
rect 29932 8372 30548 8428
rect 30044 8148 30100 8372
rect 30044 8082 30100 8092
rect 29708 7074 29764 7084
rect 30156 7028 30212 7038
rect 29820 6692 29876 6702
rect 29596 3714 29652 3724
rect 29708 5236 29764 5246
rect 29708 3778 29764 5180
rect 29708 3726 29710 3778
rect 29762 3726 29764 3778
rect 29708 3714 29764 3726
rect 29260 3554 29316 3566
rect 29260 3502 29262 3554
rect 29314 3502 29316 3554
rect 29036 1250 29092 1260
rect 29148 3444 29204 3454
rect 29260 3444 29316 3502
rect 29820 3556 29876 6636
rect 30156 6132 30212 6972
rect 30156 6066 30212 6076
rect 30380 6356 30436 6366
rect 30156 5572 30212 5582
rect 30212 5516 30324 5572
rect 30156 5506 30212 5516
rect 29932 4564 29988 4574
rect 30156 4564 30212 4574
rect 29988 4508 30100 4564
rect 29932 4498 29988 4508
rect 29820 3490 29876 3500
rect 29596 3444 29652 3454
rect 29260 3442 29652 3444
rect 29260 3390 29598 3442
rect 29650 3390 29652 3442
rect 29260 3388 29652 3390
rect 28476 578 28532 588
rect 29148 420 29204 3388
rect 29596 3378 29652 3388
rect 29932 3330 29988 3342
rect 29932 3278 29934 3330
rect 29986 3278 29988 3330
rect 29260 2772 29316 2782
rect 29260 2678 29316 2716
rect 29820 2772 29876 2782
rect 29820 2678 29876 2716
rect 29932 2658 29988 3278
rect 30044 3108 30100 4508
rect 30156 3220 30212 4508
rect 30268 3556 30324 5516
rect 30380 5236 30436 6300
rect 30492 6018 30548 8372
rect 30828 6804 30884 6814
rect 30492 5966 30494 6018
rect 30546 5966 30548 6018
rect 30492 5954 30548 5966
rect 30604 6356 30660 6366
rect 30492 5684 30548 5694
rect 30492 5348 30548 5628
rect 30492 5282 30548 5292
rect 30380 5170 30436 5180
rect 30492 4676 30548 4686
rect 30268 3490 30324 3500
rect 30380 4116 30436 4126
rect 30156 3154 30212 3164
rect 30044 3042 30100 3052
rect 29932 2606 29934 2658
rect 29986 2606 29988 2658
rect 29932 2594 29988 2606
rect 30156 2772 30212 2782
rect 30156 2210 30212 2716
rect 30380 2770 30436 4060
rect 30380 2718 30382 2770
rect 30434 2718 30436 2770
rect 30380 2706 30436 2718
rect 30156 2158 30158 2210
rect 30210 2158 30212 2210
rect 30156 2146 30212 2158
rect 30268 2660 30324 2670
rect 29596 2100 29652 2110
rect 29596 2006 29652 2044
rect 30268 1540 30324 2604
rect 30492 2324 30548 4620
rect 30604 3892 30660 6300
rect 30828 5794 30884 6748
rect 30828 5742 30830 5794
rect 30882 5742 30884 5794
rect 30828 5348 30884 5742
rect 30940 5348 30996 5358
rect 30828 5346 30996 5348
rect 30828 5294 30942 5346
rect 30994 5294 30996 5346
rect 30828 5292 30996 5294
rect 30940 5282 30996 5292
rect 30604 3826 30660 3836
rect 30604 3220 30660 3230
rect 30604 2548 30660 3164
rect 31052 2996 31108 12014
rect 31164 12068 31220 14112
rect 31500 13188 31556 13198
rect 31500 13094 31556 13132
rect 31612 13076 31668 14112
rect 31612 13010 31668 13020
rect 31724 13188 31780 13198
rect 31500 12404 31556 12414
rect 31500 12290 31556 12348
rect 31500 12238 31502 12290
rect 31554 12238 31556 12290
rect 31500 12226 31556 12238
rect 31164 12002 31220 12012
rect 31724 11508 31780 13132
rect 31948 12850 32004 12862
rect 31948 12798 31950 12850
rect 32002 12798 32004 12850
rect 31948 12516 32004 12798
rect 31948 12450 32004 12460
rect 31948 11954 32004 11966
rect 31948 11902 31950 11954
rect 32002 11902 32004 11954
rect 31948 11732 32004 11902
rect 31948 11666 32004 11676
rect 32060 11620 32116 14112
rect 32396 12962 32452 12974
rect 32396 12910 32398 12962
rect 32450 12910 32452 12962
rect 32284 12180 32340 12190
rect 32284 12086 32340 12124
rect 32396 12068 32452 12910
rect 32508 12180 32564 14112
rect 32732 13860 32788 13870
rect 32508 12114 32564 12124
rect 32620 12292 32676 12302
rect 32396 12002 32452 12012
rect 32396 11620 32452 11630
rect 32060 11618 32452 11620
rect 32060 11566 32398 11618
rect 32450 11566 32452 11618
rect 32060 11564 32452 11566
rect 32396 11554 32452 11564
rect 31724 11442 31780 11452
rect 31276 11396 31332 11406
rect 31276 11302 31332 11340
rect 31500 11396 31556 11406
rect 31500 10836 31556 11340
rect 31836 11284 31892 11294
rect 31836 11190 31892 11228
rect 31500 10770 31556 10780
rect 32620 10724 32676 12236
rect 32732 11060 32788 13804
rect 32956 13188 33012 14112
rect 32956 13122 33012 13132
rect 33292 13076 33348 13086
rect 33292 12982 33348 13020
rect 32956 12850 33012 12862
rect 32956 12798 32958 12850
rect 33010 12798 33012 12850
rect 32956 12292 33012 12798
rect 32956 12226 33012 12236
rect 33180 12180 33236 12190
rect 33180 12086 33236 12124
rect 33404 12180 33460 14112
rect 33740 13860 33796 13870
rect 33628 13412 33684 13422
rect 33404 12114 33460 12124
rect 33516 12852 33572 12862
rect 32844 12068 32900 12078
rect 32844 12066 33124 12068
rect 32844 12014 32846 12066
rect 32898 12014 33124 12066
rect 32844 12012 33124 12014
rect 32844 12002 32900 12012
rect 32732 10994 32788 11004
rect 32844 11282 32900 11294
rect 32844 11230 32846 11282
rect 32898 11230 32900 11282
rect 32620 10658 32676 10668
rect 32396 10500 32452 10510
rect 31612 10388 31668 10398
rect 31612 10386 32004 10388
rect 31612 10334 31614 10386
rect 31666 10334 32004 10386
rect 31612 10332 32004 10334
rect 31612 10322 31668 10332
rect 31724 9042 31780 9054
rect 31724 8990 31726 9042
rect 31778 8990 31780 9042
rect 31388 8818 31444 8830
rect 31388 8766 31390 8818
rect 31442 8766 31444 8818
rect 31276 8484 31332 8494
rect 31164 8372 31332 8428
rect 31388 8428 31444 8766
rect 31388 8372 31668 8428
rect 31164 8370 31220 8372
rect 31164 8318 31166 8370
rect 31218 8318 31220 8370
rect 31164 8306 31220 8318
rect 31612 8258 31668 8372
rect 31612 8206 31614 8258
rect 31666 8206 31668 8258
rect 31612 8194 31668 8206
rect 31724 7812 31780 8990
rect 31948 8930 32004 10332
rect 31948 8878 31950 8930
rect 32002 8878 32004 8930
rect 31948 8866 32004 8878
rect 32060 8820 32116 8830
rect 32060 7924 32116 8764
rect 32060 7858 32116 7868
rect 32172 8596 32228 8606
rect 31724 7746 31780 7756
rect 31164 7252 31220 7262
rect 31164 5460 31220 7196
rect 31612 6804 31668 6814
rect 31276 6692 31332 6702
rect 31276 6598 31332 6636
rect 31164 5394 31220 5404
rect 31500 5460 31556 5470
rect 31500 5234 31556 5404
rect 31500 5182 31502 5234
rect 31554 5182 31556 5234
rect 31500 5170 31556 5182
rect 31052 2930 31108 2940
rect 30604 2482 30660 2492
rect 30940 2770 30996 2782
rect 30940 2718 30942 2770
rect 30994 2718 30996 2770
rect 30940 2548 30996 2718
rect 30492 2258 30548 2268
rect 30940 1652 30996 2492
rect 30940 1586 30996 1596
rect 31164 1988 31220 1998
rect 30268 1474 30324 1484
rect 31164 1204 31220 1932
rect 31164 1138 31220 1148
rect 31388 1988 31444 1998
rect 31388 532 31444 1932
rect 31388 466 31444 476
rect 29148 354 29204 364
rect 29596 196 29652 206
rect 29596 112 29652 140
rect 31612 112 31668 6748
rect 31836 6690 31892 6702
rect 31836 6638 31838 6690
rect 31890 6638 31892 6690
rect 31836 6132 31892 6638
rect 31836 6066 31892 6076
rect 31948 6244 32004 6254
rect 31948 2770 32004 6188
rect 32060 5796 32116 5806
rect 32060 5702 32116 5740
rect 32060 5348 32116 5358
rect 32060 4788 32116 5292
rect 32172 5124 32228 8540
rect 32396 8148 32452 10444
rect 32620 9044 32676 9054
rect 32508 8932 32564 8942
rect 32508 8838 32564 8876
rect 32396 8082 32452 8092
rect 32620 6804 32676 8988
rect 32620 6738 32676 6748
rect 32620 6132 32676 6142
rect 32620 6038 32676 6076
rect 32172 5058 32228 5068
rect 32060 4722 32116 4732
rect 32284 5012 32340 5022
rect 32060 4452 32116 4462
rect 32060 3108 32116 4396
rect 32060 3042 32116 3052
rect 31948 2718 31950 2770
rect 32002 2718 32004 2770
rect 31948 2706 32004 2718
rect 32284 2436 32340 4956
rect 32844 2772 32900 11230
rect 32956 7812 33012 7822
rect 32956 6130 33012 7756
rect 32956 6078 32958 6130
rect 33010 6078 33012 6130
rect 32956 6066 33012 6078
rect 33068 3220 33124 12012
rect 33516 11620 33572 12796
rect 33628 12290 33684 13356
rect 33628 12238 33630 12290
rect 33682 12238 33684 12290
rect 33628 12226 33684 12238
rect 33516 11554 33572 11564
rect 33516 11172 33572 11182
rect 33180 10164 33236 10174
rect 33180 8820 33236 10108
rect 33292 9940 33348 9950
rect 33292 9042 33348 9884
rect 33516 9604 33572 11116
rect 33516 9538 33572 9548
rect 33740 9380 33796 13804
rect 33852 13636 33908 14112
rect 33852 13570 33908 13580
rect 34188 13188 34244 13198
rect 34188 13094 34244 13132
rect 33292 8990 33294 9042
rect 33346 8990 33348 9042
rect 33292 8978 33348 8990
rect 33404 9324 33796 9380
rect 33852 12850 33908 12862
rect 33852 12798 33854 12850
rect 33906 12798 33908 12850
rect 33404 9044 33460 9324
rect 33852 9044 33908 12798
rect 34188 12404 34244 12414
rect 34076 12180 34132 12190
rect 34076 12086 34132 12124
rect 33404 8978 33460 8988
rect 33740 8988 33908 9044
rect 33964 11956 34020 11966
rect 34188 11956 34244 12348
rect 34300 12180 34356 14112
rect 34524 12516 34580 14140
rect 34720 14112 34832 14224
rect 35168 14112 35280 14224
rect 35616 14112 35728 14224
rect 36064 14112 36176 14224
rect 36512 14112 36624 14224
rect 36960 14112 37072 14224
rect 37408 14112 37520 14224
rect 37856 14112 37968 14224
rect 38304 14112 38416 14224
rect 38752 14112 38864 14224
rect 39200 14112 39312 14224
rect 39648 14112 39760 14224
rect 40096 14112 40208 14224
rect 40544 14112 40656 14224
rect 40992 14112 41104 14224
rect 41440 14112 41552 14224
rect 41888 14112 42000 14224
rect 42336 14112 42448 14224
rect 42784 14112 42896 14224
rect 43232 14112 43344 14224
rect 43680 14112 43792 14224
rect 44128 14112 44240 14224
rect 44576 14112 44688 14224
rect 45024 14112 45136 14224
rect 45472 14112 45584 14224
rect 45920 14112 46032 14224
rect 46368 14112 46480 14224
rect 46816 14112 46928 14224
rect 47264 14112 47376 14224
rect 47712 14112 47824 14224
rect 48160 14112 48272 14224
rect 48608 14112 48720 14224
rect 49056 14112 49168 14224
rect 49504 14112 49616 14224
rect 49952 14112 50064 14224
rect 50400 14112 50512 14224
rect 50848 14112 50960 14224
rect 51296 14112 51408 14224
rect 51744 14112 51856 14224
rect 52192 14112 52304 14224
rect 52640 14112 52752 14224
rect 53088 14112 53200 14224
rect 53536 14112 53648 14224
rect 53984 14112 54096 14224
rect 54432 14112 54544 14224
rect 54880 14112 54992 14224
rect 55328 14112 55440 14224
rect 55776 14112 55888 14224
rect 56224 14112 56336 14224
rect 56672 14112 56784 14224
rect 34748 13188 34804 14112
rect 35196 13524 35252 14112
rect 35196 13458 35252 13468
rect 35308 13636 35364 13646
rect 34748 13122 34804 13132
rect 35308 13186 35364 13580
rect 35644 13636 35700 14112
rect 35644 13570 35700 13580
rect 35308 13134 35310 13186
rect 35362 13134 35364 13186
rect 35308 13122 35364 13134
rect 35868 13076 35924 13086
rect 34748 12852 34804 12862
rect 34748 12850 35140 12852
rect 34748 12798 34750 12850
rect 34802 12798 35140 12850
rect 34748 12796 35140 12798
rect 34748 12786 34804 12796
rect 34524 12460 34804 12516
rect 34300 12114 34356 12124
rect 34524 12290 34580 12302
rect 34524 12238 34526 12290
rect 34578 12238 34580 12290
rect 34412 12068 34468 12078
rect 34188 11900 34356 11956
rect 33180 8754 33236 8764
rect 33516 8932 33572 8942
rect 33516 8484 33572 8876
rect 33516 8418 33572 8428
rect 33628 8820 33684 8830
rect 33628 8258 33684 8764
rect 33740 8428 33796 8988
rect 33852 8820 33908 8830
rect 33852 8726 33908 8764
rect 33740 8372 33908 8428
rect 33628 8206 33630 8258
rect 33682 8206 33684 8258
rect 33628 8194 33684 8206
rect 33852 7028 33908 8372
rect 33964 7252 34020 11900
rect 34188 10276 34244 10286
rect 34076 9940 34132 9950
rect 34076 9156 34132 9884
rect 34188 9380 34244 10220
rect 34188 9314 34244 9324
rect 34076 9100 34244 9156
rect 34076 8820 34132 8830
rect 34076 8370 34132 8764
rect 34076 8318 34078 8370
rect 34130 8318 34132 8370
rect 34076 8306 34132 8318
rect 33964 7186 34020 7196
rect 33852 6962 33908 6972
rect 33404 6804 33460 6814
rect 33180 5796 33236 5806
rect 33180 5702 33236 5740
rect 33068 3154 33124 3164
rect 32844 2706 32900 2716
rect 33068 2660 33124 2670
rect 33068 2566 33124 2604
rect 32508 2548 32564 2558
rect 32508 2454 32564 2492
rect 32284 2370 32340 2380
rect 32284 1764 32340 1774
rect 32060 1540 32116 1550
rect 31948 1484 32060 1540
rect 31724 1428 31780 1438
rect 31948 1428 32004 1484
rect 32060 1474 32116 1484
rect 31780 1372 32004 1428
rect 31724 1362 31780 1372
rect 31948 756 32004 766
rect 31948 196 32004 700
rect 31948 130 32004 140
rect 21756 18 21812 28
rect 23520 0 23632 112
rect 25536 0 25648 112
rect 27552 0 27664 112
rect 29568 0 29680 112
rect 31584 0 31696 112
rect 32284 84 32340 1708
rect 33404 1540 33460 6748
rect 33628 6244 33684 6254
rect 33628 5794 33684 6188
rect 33628 5742 33630 5794
rect 33682 5742 33684 5794
rect 33628 5730 33684 5742
rect 34188 5010 34244 9100
rect 34300 7476 34356 11900
rect 34412 11394 34468 12012
rect 34524 11508 34580 12238
rect 34524 11442 34580 11452
rect 34748 11506 34804 12460
rect 34972 12180 35028 12190
rect 34972 12086 35028 12124
rect 34748 11454 34750 11506
rect 34802 11454 34804 11506
rect 34412 11342 34414 11394
rect 34466 11342 34468 11394
rect 34412 11330 34468 11342
rect 34412 10386 34468 10398
rect 34412 10334 34414 10386
rect 34466 10334 34468 10386
rect 34412 10276 34468 10334
rect 34412 10210 34468 10220
rect 34748 10276 34804 11454
rect 34972 11844 35028 11854
rect 34972 10948 35028 11788
rect 34748 10210 34804 10220
rect 34860 10892 35028 10948
rect 34300 7410 34356 7420
rect 34636 8146 34692 8158
rect 34636 8094 34638 8146
rect 34690 8094 34692 8146
rect 34188 4958 34190 5010
rect 34242 4958 34244 5010
rect 34188 4946 34244 4958
rect 34524 5234 34580 5246
rect 34524 5182 34526 5234
rect 34578 5182 34580 5234
rect 34524 4338 34580 5182
rect 34524 4286 34526 4338
rect 34578 4286 34580 4338
rect 34524 4274 34580 4286
rect 34412 4114 34468 4126
rect 34412 4062 34414 4114
rect 34466 4062 34468 4114
rect 34412 4004 34468 4062
rect 34412 3938 34468 3948
rect 34524 4116 34580 4126
rect 34524 2324 34580 4060
rect 34524 2258 34580 2268
rect 34636 1764 34692 8094
rect 34748 7028 34804 7038
rect 34748 1988 34804 6972
rect 34860 6468 34916 10892
rect 34972 10724 35028 10734
rect 34972 10630 35028 10668
rect 34972 9044 35028 9054
rect 34972 8950 35028 8988
rect 34972 8708 35028 8718
rect 34972 7924 35028 8652
rect 35084 8258 35140 12796
rect 35756 12850 35812 12862
rect 35756 12798 35758 12850
rect 35810 12798 35812 12850
rect 35196 12516 35252 12526
rect 35196 10276 35252 12460
rect 35196 10210 35252 10220
rect 35308 12404 35364 12414
rect 35308 8428 35364 12348
rect 35420 12068 35476 12078
rect 35420 9940 35476 12012
rect 35532 12068 35588 12078
rect 35532 12066 35700 12068
rect 35532 12014 35534 12066
rect 35586 12014 35700 12066
rect 35532 12012 35700 12014
rect 35532 12002 35588 12012
rect 35532 11284 35588 11294
rect 35532 10388 35588 11228
rect 35532 10322 35588 10332
rect 35420 9874 35476 9884
rect 35532 10052 35588 10062
rect 35308 8372 35476 8428
rect 35084 8206 35086 8258
rect 35138 8206 35140 8258
rect 35084 8036 35140 8206
rect 35308 8260 35364 8270
rect 35420 8260 35476 8372
rect 35364 8204 35476 8260
rect 35308 8194 35364 8204
rect 35084 7970 35140 7980
rect 34972 7858 35028 7868
rect 35308 7140 35364 7150
rect 35196 6692 35252 6702
rect 34860 6402 34916 6412
rect 35084 6468 35140 6478
rect 34972 5012 35028 5022
rect 34972 4450 35028 4956
rect 34972 4398 34974 4450
rect 35026 4398 35028 4450
rect 34972 4386 35028 4398
rect 35084 4116 35140 6412
rect 35196 5796 35252 6636
rect 35308 6020 35364 7084
rect 35532 6244 35588 9996
rect 35644 6356 35700 12012
rect 35756 11844 35812 12798
rect 35756 11778 35812 11788
rect 35756 9940 35812 9950
rect 35756 9268 35812 9884
rect 35868 9380 35924 13020
rect 36092 11620 36148 14112
rect 36204 13188 36260 13198
rect 36204 13094 36260 13132
rect 36316 12068 36372 12078
rect 36316 11974 36372 12012
rect 36428 11620 36484 11630
rect 36092 11618 36484 11620
rect 36092 11566 36430 11618
rect 36482 11566 36484 11618
rect 36092 11564 36484 11566
rect 36428 11554 36484 11564
rect 36540 11620 36596 14112
rect 36876 12964 36932 12974
rect 36764 12850 36820 12862
rect 36764 12798 36766 12850
rect 36818 12798 36820 12850
rect 36764 12628 36820 12798
rect 36764 12562 36820 12572
rect 36876 12404 36932 12908
rect 36988 12852 37044 14112
rect 37436 13860 37492 14112
rect 37436 13794 37492 13804
rect 37100 13524 37156 13534
rect 37100 13186 37156 13468
rect 37100 13134 37102 13186
rect 37154 13134 37156 13186
rect 37100 13122 37156 13134
rect 37884 12964 37940 14112
rect 37996 13636 38052 13646
rect 37996 13186 38052 13580
rect 37996 13134 37998 13186
rect 38050 13134 38052 13186
rect 37996 13122 38052 13134
rect 37884 12908 38052 12964
rect 36988 12786 37044 12796
rect 37212 12852 37268 12862
rect 36764 12348 36932 12404
rect 36540 11554 36596 11564
rect 36652 12292 36708 12302
rect 35980 11508 36036 11518
rect 35980 11170 36036 11452
rect 35980 11118 35982 11170
rect 36034 11118 36036 11170
rect 35980 9604 36036 11118
rect 35980 9538 36036 9548
rect 36316 11396 36372 11406
rect 35868 9324 36260 9380
rect 35756 9212 35924 9268
rect 35756 8372 35812 8382
rect 35756 8278 35812 8316
rect 35644 6290 35700 6300
rect 35308 5954 35364 5964
rect 35420 6188 35588 6244
rect 35196 5740 35364 5796
rect 34972 4060 35140 4116
rect 34748 1922 34804 1932
rect 34860 3892 34916 3902
rect 34636 1698 34692 1708
rect 33404 1474 33460 1484
rect 33628 1652 33684 1662
rect 33628 112 33684 1596
rect 33740 1428 33796 1438
rect 33740 868 33796 1372
rect 33740 802 33796 812
rect 34860 868 34916 3836
rect 34860 802 34916 812
rect 34972 644 35028 4060
rect 35308 4004 35364 5740
rect 35308 3938 35364 3948
rect 35084 3892 35140 3902
rect 35084 1428 35140 3836
rect 35196 3668 35252 3678
rect 35196 1764 35252 3612
rect 35308 3332 35364 3342
rect 35308 2770 35364 3276
rect 35308 2718 35310 2770
rect 35362 2718 35364 2770
rect 35308 2706 35364 2718
rect 35196 1698 35252 1708
rect 35084 1362 35140 1372
rect 35420 1204 35476 6188
rect 35532 6020 35588 6030
rect 35532 3444 35588 5964
rect 35756 4900 35812 4910
rect 35756 4806 35812 4844
rect 35756 3556 35812 3566
rect 35868 3556 35924 9212
rect 36092 8370 36148 8382
rect 36092 8318 36094 8370
rect 36146 8318 36148 8370
rect 36092 7700 36148 8318
rect 36092 7634 36148 7644
rect 36204 3778 36260 9324
rect 36316 9154 36372 11340
rect 36652 10612 36708 12236
rect 36540 10556 36708 10612
rect 36540 10164 36596 10556
rect 36764 10276 36820 12348
rect 36988 12292 37044 12302
rect 36876 12180 36932 12190
rect 36876 12086 36932 12124
rect 36876 11284 36932 11294
rect 36876 11190 36932 11228
rect 36764 10220 36932 10276
rect 36540 10108 36820 10164
rect 36316 9102 36318 9154
rect 36370 9102 36372 9154
rect 36316 9090 36372 9102
rect 36540 9940 36596 9950
rect 36428 8372 36484 8382
rect 36316 8036 36372 8046
rect 36316 7942 36372 7980
rect 36316 7588 36372 7598
rect 36428 7588 36484 8316
rect 36316 7586 36484 7588
rect 36316 7534 36318 7586
rect 36370 7534 36484 7586
rect 36316 7532 36484 7534
rect 36540 7588 36596 9884
rect 36764 9042 36820 10108
rect 36876 9828 36932 10220
rect 36988 10164 37044 12236
rect 36988 10098 37044 10108
rect 36876 9772 37044 9828
rect 36764 8990 36766 9042
rect 36818 8990 36820 9042
rect 36652 8932 36708 8942
rect 36652 8370 36708 8876
rect 36652 8318 36654 8370
rect 36706 8318 36708 8370
rect 36652 8306 36708 8318
rect 36764 8372 36820 8990
rect 36764 8306 36820 8316
rect 36876 9604 36932 9614
rect 36988 9604 37044 9772
rect 37100 9604 37156 9614
rect 36988 9548 37100 9604
rect 36316 7522 36372 7532
rect 36540 7522 36596 7532
rect 36652 7476 36708 7486
rect 36652 5796 36708 7420
rect 36764 7476 36820 7486
rect 36876 7476 36932 9548
rect 37100 9538 37156 9548
rect 36764 7474 36932 7476
rect 36764 7422 36766 7474
rect 36818 7422 36932 7474
rect 36764 7420 36932 7422
rect 37100 8036 37156 8046
rect 37100 7474 37156 7980
rect 37100 7422 37102 7474
rect 37154 7422 37156 7474
rect 36764 7410 36820 7420
rect 37100 7410 37156 7422
rect 36652 5730 36708 5740
rect 36988 6692 37044 6702
rect 36988 5348 37044 6636
rect 37212 6580 37268 12796
rect 37660 12850 37716 12862
rect 37660 12798 37662 12850
rect 37714 12798 37716 12850
rect 37324 11620 37380 11630
rect 37324 11526 37380 11564
rect 37324 10276 37380 10286
rect 37324 9156 37380 10220
rect 37324 9090 37380 9100
rect 37548 8484 37604 8494
rect 37548 8036 37604 8428
rect 37548 7970 37604 7980
rect 37436 7700 37492 7710
rect 37212 6514 37268 6524
rect 37324 7250 37380 7262
rect 37324 7198 37326 7250
rect 37378 7198 37380 7250
rect 37212 6244 37268 6254
rect 37212 6018 37268 6188
rect 37324 6130 37380 7198
rect 37324 6078 37326 6130
rect 37378 6078 37380 6130
rect 37324 6066 37380 6078
rect 37212 5966 37214 6018
rect 37266 5966 37268 6018
rect 37212 5954 37268 5966
rect 37436 5908 37492 7644
rect 37324 5852 37492 5908
rect 36988 5282 37044 5292
rect 37100 5682 37156 5694
rect 37100 5630 37102 5682
rect 37154 5630 37156 5682
rect 37100 5012 37156 5630
rect 37100 4946 37156 4956
rect 37212 5348 37268 5358
rect 37212 4788 37268 5292
rect 36204 3726 36206 3778
rect 36258 3726 36260 3778
rect 35756 3554 36148 3556
rect 35756 3502 35758 3554
rect 35810 3502 36148 3554
rect 35756 3500 36148 3502
rect 35756 3490 35812 3500
rect 35532 3378 35588 3388
rect 36092 3108 36148 3500
rect 36204 3332 36260 3726
rect 36204 3266 36260 3276
rect 36764 4732 37268 4788
rect 36092 3052 36596 3108
rect 36540 2770 36596 3052
rect 36540 2718 36542 2770
rect 36594 2718 36596 2770
rect 36540 2706 36596 2718
rect 35756 2658 35812 2670
rect 35756 2606 35758 2658
rect 35810 2606 35812 2658
rect 35420 1138 35476 1148
rect 35644 2548 35700 2558
rect 34972 578 35028 588
rect 35644 112 35700 2492
rect 35756 1540 35812 2606
rect 36652 2212 36708 2222
rect 36652 2118 36708 2156
rect 36764 1652 36820 4732
rect 36876 4564 36932 4574
rect 36876 1988 36932 4508
rect 37212 3892 37268 3902
rect 36988 2658 37044 2670
rect 36988 2606 36990 2658
rect 37042 2606 37044 2658
rect 36988 2212 37044 2606
rect 36988 2146 37044 2156
rect 37212 2098 37268 3836
rect 37324 3778 37380 5852
rect 37660 5796 37716 12798
rect 37884 12740 37940 12750
rect 37772 12178 37828 12190
rect 37772 12126 37774 12178
rect 37826 12126 37828 12178
rect 37772 12068 37828 12126
rect 37772 12002 37828 12012
rect 37772 11282 37828 11294
rect 37772 11230 37774 11282
rect 37826 11230 37828 11282
rect 37772 6580 37828 11230
rect 37884 8428 37940 12684
rect 37996 11620 38052 12908
rect 37996 11554 38052 11564
rect 38108 12740 38164 12750
rect 38108 9940 38164 12684
rect 38332 12180 38388 14112
rect 38444 12852 38500 12862
rect 38444 12758 38500 12796
rect 38220 12124 38388 12180
rect 38220 10164 38276 12124
rect 38332 11956 38388 11966
rect 38780 11956 38836 14112
rect 39228 13300 39284 14112
rect 39228 13234 39284 13244
rect 39676 13076 39732 14112
rect 39676 13010 39732 13020
rect 40124 12964 40180 14112
rect 40572 13188 40628 14112
rect 40796 13188 40852 13198
rect 40572 13186 40852 13188
rect 40572 13134 40798 13186
rect 40850 13134 40852 13186
rect 40572 13132 40852 13134
rect 40796 13122 40852 13132
rect 41020 13188 41076 14112
rect 41020 13122 41076 13132
rect 41356 13748 41412 13758
rect 41356 13074 41412 13692
rect 41468 13636 41524 14112
rect 41468 13570 41524 13580
rect 41692 13188 41748 13198
rect 41692 13094 41748 13132
rect 41916 13188 41972 14112
rect 41916 13122 41972 13132
rect 41356 13022 41358 13074
rect 41410 13022 41412 13074
rect 41356 13010 41412 13022
rect 40124 12898 40180 12908
rect 42140 12850 42196 12862
rect 42140 12798 42142 12850
rect 42194 12798 42196 12850
rect 40124 12516 40180 12526
rect 38332 11954 38500 11956
rect 38332 11902 38334 11954
rect 38386 11902 38500 11954
rect 38332 11900 38500 11902
rect 38332 11890 38388 11900
rect 38220 10098 38276 10108
rect 38444 11394 38500 11900
rect 38780 11890 38836 11900
rect 39452 11954 39508 11966
rect 39452 11902 39454 11954
rect 39506 11902 39508 11954
rect 38444 11342 38446 11394
rect 38498 11342 38500 11394
rect 38444 10052 38500 11342
rect 39004 11282 39060 11294
rect 39004 11230 39006 11282
rect 39058 11230 39060 11282
rect 38444 9986 38500 9996
rect 38556 10948 38612 10958
rect 38108 9884 38276 9940
rect 38108 8930 38164 8942
rect 38108 8878 38110 8930
rect 38162 8878 38164 8930
rect 37884 8362 37940 8372
rect 37996 8370 38052 8382
rect 37996 8318 37998 8370
rect 38050 8318 38052 8370
rect 37884 8258 37940 8270
rect 37884 8206 37886 8258
rect 37938 8206 37940 8258
rect 37884 7700 37940 8206
rect 37996 8260 38052 8318
rect 37996 8194 38052 8204
rect 37884 7140 37940 7644
rect 37884 7074 37940 7084
rect 37996 7474 38052 7486
rect 37996 7422 37998 7474
rect 38050 7422 38052 7474
rect 37772 6514 37828 6524
rect 37884 6244 37940 6254
rect 37884 5908 37940 6188
rect 37996 6020 38052 7422
rect 38108 6132 38164 8878
rect 38220 7364 38276 9884
rect 38220 7298 38276 7308
rect 38332 9156 38388 9166
rect 38332 6692 38388 9100
rect 38556 9044 38612 10892
rect 38444 9042 38612 9044
rect 38444 8990 38558 9042
rect 38610 8990 38612 9042
rect 38444 8988 38612 8990
rect 38444 8596 38500 8988
rect 38556 8978 38612 8988
rect 38780 9604 38836 9614
rect 38444 8540 38724 8596
rect 38444 7474 38500 8540
rect 38444 7422 38446 7474
rect 38498 7422 38500 7474
rect 38444 7410 38500 7422
rect 38556 8428 38612 8438
rect 38332 6626 38388 6636
rect 38108 6076 38388 6132
rect 37996 5964 38276 6020
rect 37884 5852 38164 5908
rect 37436 5740 37716 5796
rect 38108 5794 38164 5852
rect 38108 5742 38110 5794
rect 38162 5742 38164 5794
rect 37436 4116 37492 5740
rect 38108 5730 38164 5742
rect 38220 5572 38276 5964
rect 38108 5516 38276 5572
rect 38108 4900 38164 5516
rect 38108 4834 38164 4844
rect 38220 5012 38276 5022
rect 37996 4788 38052 4798
rect 37436 4050 37492 4060
rect 37884 4452 37940 4462
rect 37324 3726 37326 3778
rect 37378 3726 37380 3778
rect 37324 3714 37380 3726
rect 37212 2046 37214 2098
rect 37266 2046 37268 2098
rect 37212 2034 37268 2046
rect 37660 3556 37716 3566
rect 36876 1932 37044 1988
rect 36764 1586 36820 1596
rect 35756 1474 35812 1484
rect 36988 980 37044 1932
rect 36988 914 37044 924
rect 37660 112 37716 3500
rect 37884 2098 37940 4396
rect 37996 4228 38052 4732
rect 37996 4162 38052 4172
rect 38220 2994 38276 4956
rect 38332 3108 38388 6076
rect 38556 6018 38612 8372
rect 38668 8258 38724 8540
rect 38668 8206 38670 8258
rect 38722 8206 38724 8258
rect 38668 8194 38724 8206
rect 38780 7588 38836 9548
rect 39004 9604 39060 11230
rect 39004 9538 39060 9548
rect 39116 11284 39172 11294
rect 39004 8372 39060 8382
rect 39004 8278 39060 8316
rect 38780 7522 38836 7532
rect 39116 7252 39172 11228
rect 39452 10500 39508 11902
rect 40124 11844 40180 12460
rect 42140 12404 42196 12798
rect 42140 12338 42196 12348
rect 41356 12292 41412 12302
rect 41356 12198 41412 12236
rect 40124 11778 40180 11788
rect 40348 12068 40404 12078
rect 40236 10612 40292 10622
rect 39452 10434 39508 10444
rect 39900 10500 39956 10510
rect 39676 10388 39732 10398
rect 39564 8932 39620 8942
rect 39564 8838 39620 8876
rect 39340 8260 39396 8270
rect 39340 7474 39396 8204
rect 39340 7422 39342 7474
rect 39394 7422 39396 7474
rect 39340 7410 39396 7422
rect 39452 7476 39508 7486
rect 39116 7186 39172 7196
rect 39452 7140 39508 7420
rect 39452 7074 39508 7084
rect 39676 7140 39732 10332
rect 39900 9042 39956 10444
rect 40236 10052 40292 10556
rect 40236 9986 40292 9996
rect 40348 9492 40404 12012
rect 42252 12068 42308 12078
rect 42252 11974 42308 12012
rect 41692 11956 41748 11966
rect 41244 11508 41300 11518
rect 41244 11394 41300 11452
rect 41244 11342 41246 11394
rect 41298 11342 41300 11394
rect 41244 11330 41300 11342
rect 41580 11508 41636 11518
rect 40908 11172 40964 11182
rect 40572 11170 40964 11172
rect 40572 11118 40910 11170
rect 40962 11118 40964 11170
rect 40572 11116 40964 11118
rect 40460 10388 40516 10398
rect 40460 10294 40516 10332
rect 40348 9426 40404 9436
rect 40124 9380 40180 9390
rect 39900 8990 39902 9042
rect 39954 8990 39956 9042
rect 39900 8978 39956 8990
rect 40012 9044 40068 9054
rect 40012 8950 40068 8988
rect 39788 8820 39844 8830
rect 40124 8820 40180 9324
rect 39788 8726 39844 8764
rect 40012 8764 40180 8820
rect 39676 7074 39732 7084
rect 39788 7364 39844 7374
rect 39788 6916 39844 7308
rect 38556 5966 38558 6018
rect 38610 5966 38612 6018
rect 38556 5954 38612 5966
rect 39564 6860 39844 6916
rect 38444 5906 38500 5918
rect 38444 5854 38446 5906
rect 38498 5854 38500 5906
rect 38444 5572 38500 5854
rect 38780 5908 38836 5918
rect 38780 5906 39396 5908
rect 38780 5854 38782 5906
rect 38834 5854 39396 5906
rect 38780 5852 39396 5854
rect 38780 5842 38836 5852
rect 39228 5684 39284 5694
rect 38780 5682 39284 5684
rect 38780 5630 39230 5682
rect 39282 5630 39284 5682
rect 38780 5628 39284 5630
rect 38780 5572 38836 5628
rect 39228 5618 39284 5628
rect 38444 5516 38836 5572
rect 39340 5348 39396 5852
rect 39564 5906 39620 6860
rect 39900 6804 39956 6814
rect 39564 5854 39566 5906
rect 39618 5854 39620 5906
rect 39564 5842 39620 5854
rect 39788 6748 39900 6804
rect 39452 5684 39508 5694
rect 39452 5682 39620 5684
rect 39452 5630 39454 5682
rect 39506 5630 39620 5682
rect 39452 5628 39620 5630
rect 39452 5618 39508 5628
rect 39452 5348 39508 5358
rect 39340 5346 39508 5348
rect 39340 5294 39454 5346
rect 39506 5294 39508 5346
rect 39340 5292 39508 5294
rect 39452 5282 39508 5292
rect 38668 5122 38724 5134
rect 38668 5070 38670 5122
rect 38722 5070 38724 5122
rect 38668 5012 38724 5070
rect 38780 5124 38836 5134
rect 39116 5124 39172 5134
rect 38780 5122 39172 5124
rect 38780 5070 38782 5122
rect 38834 5070 39118 5122
rect 39170 5070 39172 5122
rect 38780 5068 39172 5070
rect 38780 5058 38836 5068
rect 39116 5058 39172 5068
rect 39452 5122 39508 5134
rect 39452 5070 39454 5122
rect 39506 5070 39508 5122
rect 38668 4946 38724 4956
rect 39452 4562 39508 5070
rect 39452 4510 39454 4562
rect 39506 4510 39508 4562
rect 39452 4498 39508 4510
rect 39564 4900 39620 5628
rect 39788 5122 39844 6748
rect 39900 6738 39956 6748
rect 40012 5684 40068 8764
rect 40236 8484 40292 8494
rect 40236 8148 40292 8428
rect 40236 8082 40292 8092
rect 40572 7364 40628 11116
rect 40908 11106 40964 11116
rect 41580 10834 41636 11452
rect 41580 10782 41582 10834
rect 41634 10782 41636 10834
rect 41580 10770 41636 10782
rect 40684 10500 40740 10510
rect 40684 10406 40740 10444
rect 40796 10500 40852 10510
rect 41244 10500 41300 10510
rect 40796 10498 41300 10500
rect 40796 10446 40798 10498
rect 40850 10446 41246 10498
rect 41298 10446 41300 10498
rect 40796 10444 41300 10446
rect 40796 10434 40852 10444
rect 41244 10434 41300 10444
rect 41580 10500 41636 10510
rect 40908 10276 40964 10286
rect 40684 9044 40740 9054
rect 40684 8950 40740 8988
rect 40796 8818 40852 8830
rect 40796 8766 40798 8818
rect 40850 8766 40852 8818
rect 40796 8258 40852 8766
rect 40796 8206 40798 8258
rect 40850 8206 40852 8258
rect 40796 8194 40852 8206
rect 40908 7924 40964 10220
rect 41244 10164 41300 10174
rect 41132 9044 41188 9054
rect 41132 8370 41188 8988
rect 41132 8318 41134 8370
rect 41186 8318 41188 8370
rect 41132 8306 41188 8318
rect 41020 8260 41076 8270
rect 41020 8166 41076 8204
rect 40908 7858 40964 7868
rect 40572 7298 40628 7308
rect 40012 5618 40068 5628
rect 40124 7252 40180 7262
rect 40124 5572 40180 7196
rect 40460 7028 40516 7038
rect 40124 5506 40180 5516
rect 40236 6916 40292 6926
rect 39788 5070 39790 5122
rect 39842 5070 39844 5122
rect 39788 5058 39844 5070
rect 39564 4338 39620 4844
rect 40236 4900 40292 6860
rect 40460 6692 40516 6972
rect 41244 6916 41300 10108
rect 41356 9156 41412 9166
rect 41356 9062 41412 9100
rect 41468 8930 41524 8942
rect 41468 8878 41470 8930
rect 41522 8878 41524 8930
rect 41468 8820 41524 8878
rect 41468 8754 41524 8764
rect 41580 8370 41636 10444
rect 41580 8318 41582 8370
rect 41634 8318 41636 8370
rect 41580 8306 41636 8318
rect 41244 6850 41300 6860
rect 41356 8258 41412 8270
rect 41356 8206 41358 8258
rect 41410 8206 41412 8258
rect 41132 6804 41188 6814
rect 41132 6710 41188 6748
rect 40460 6626 40516 6636
rect 41356 6692 41412 8206
rect 41468 8260 41524 8270
rect 41692 8260 41748 11900
rect 41916 11954 41972 11966
rect 41916 11902 41918 11954
rect 41970 11902 41972 11954
rect 41916 11508 41972 11902
rect 41916 11442 41972 11452
rect 42028 11732 42084 11742
rect 42028 11508 42084 11676
rect 42364 11620 42420 14112
rect 42700 12852 42756 12862
rect 42700 12178 42756 12796
rect 42700 12126 42702 12178
rect 42754 12126 42756 12178
rect 42700 11732 42756 12126
rect 42812 12180 42868 14112
rect 42924 13636 42980 13646
rect 42924 13186 42980 13580
rect 42924 13134 42926 13186
rect 42978 13134 42980 13186
rect 42924 13122 42980 13134
rect 43036 12964 43092 12974
rect 42812 12114 42868 12124
rect 42924 12628 42980 12638
rect 42700 11666 42756 11676
rect 42812 11956 42868 11966
rect 42588 11620 42644 11630
rect 42364 11618 42644 11620
rect 42364 11566 42590 11618
rect 42642 11566 42644 11618
rect 42364 11564 42644 11566
rect 42588 11554 42644 11564
rect 42028 11506 42196 11508
rect 42028 11454 42030 11506
rect 42082 11454 42196 11506
rect 42028 11452 42196 11454
rect 42028 11442 42084 11452
rect 41804 11396 41860 11406
rect 41804 11302 41860 11340
rect 42140 10498 42196 11452
rect 42364 11396 42420 11406
rect 42252 10612 42308 10650
rect 42252 10546 42308 10556
rect 42140 10446 42142 10498
rect 42194 10446 42196 10498
rect 42140 10434 42196 10446
rect 42252 10388 42308 10398
rect 41804 9042 41860 9054
rect 41804 8990 41806 9042
rect 41858 8990 41860 9042
rect 41804 8428 41860 8990
rect 42252 9042 42308 10332
rect 42252 8990 42254 9042
rect 42306 8990 42308 9042
rect 42252 8978 42308 8990
rect 41916 8596 41972 8606
rect 41972 8540 42084 8596
rect 41916 8530 41972 8540
rect 41804 8372 41972 8428
rect 41916 8370 41972 8372
rect 41916 8318 41918 8370
rect 41970 8318 41972 8370
rect 41916 8306 41972 8318
rect 41692 8204 41860 8260
rect 41468 8036 41524 8204
rect 41692 8036 41748 8046
rect 41468 8034 41748 8036
rect 41468 7982 41694 8034
rect 41746 7982 41748 8034
rect 41468 7980 41748 7982
rect 41692 7970 41748 7980
rect 41804 7364 41860 8204
rect 42028 7700 42084 8540
rect 42140 8370 42196 8382
rect 42140 8318 42142 8370
rect 42194 8318 42196 8370
rect 42140 8260 42196 8318
rect 42252 8372 42308 8382
rect 42252 8278 42308 8316
rect 42140 8194 42196 8204
rect 42364 8148 42420 11340
rect 42588 9826 42644 9838
rect 42588 9774 42590 9826
rect 42642 9774 42644 9826
rect 42476 9602 42532 9614
rect 42476 9550 42478 9602
rect 42530 9550 42532 9602
rect 42476 8930 42532 9550
rect 42476 8878 42478 8930
rect 42530 8878 42532 8930
rect 42476 8866 42532 8878
rect 42252 8092 42420 8148
rect 42588 8148 42644 9774
rect 42812 8148 42868 11900
rect 42924 8428 42980 12572
rect 43036 11732 43092 12908
rect 43036 11666 43092 11676
rect 43260 11620 43316 14112
rect 43484 14084 43540 14094
rect 43484 13074 43540 14028
rect 43484 13022 43486 13074
rect 43538 13022 43540 13074
rect 43484 13010 43540 13022
rect 43708 12740 43764 14112
rect 43820 13188 43876 13198
rect 43820 13094 43876 13132
rect 44156 12964 44212 14112
rect 44604 13636 44660 14112
rect 44604 13570 44660 13580
rect 44940 13524 44996 13534
rect 44464 13356 44728 13366
rect 44520 13300 44568 13356
rect 44624 13300 44672 13356
rect 44464 13290 44728 13300
rect 44940 13074 44996 13468
rect 44940 13022 44942 13074
rect 44994 13022 44996 13074
rect 44940 13010 44996 13022
rect 44156 12898 44212 12908
rect 44380 12852 44436 12862
rect 44380 12758 44436 12796
rect 44604 12740 44660 12750
rect 43708 12684 44324 12740
rect 43804 12572 44068 12582
rect 43596 12516 43652 12526
rect 43860 12516 43908 12572
rect 43964 12516 44012 12572
rect 43804 12506 44068 12516
rect 43484 11620 43540 11630
rect 43260 11618 43540 11620
rect 43260 11566 43486 11618
rect 43538 11566 43540 11618
rect 43260 11564 43540 11566
rect 43484 11554 43540 11564
rect 43036 11282 43092 11294
rect 43036 11230 43038 11282
rect 43090 11230 43092 11282
rect 43036 9940 43092 11230
rect 43036 9874 43092 9884
rect 43260 11284 43316 11294
rect 43148 9044 43204 9054
rect 43148 8950 43204 8988
rect 42924 8372 43092 8428
rect 42028 7644 42196 7700
rect 41804 7308 41972 7364
rect 41356 6626 41412 6636
rect 41804 7140 41860 7150
rect 41468 6468 41524 6478
rect 41468 6374 41524 6412
rect 41804 6018 41860 7084
rect 41804 5966 41806 6018
rect 41858 5966 41860 6018
rect 41804 5954 41860 5966
rect 40236 4834 40292 4844
rect 40460 5236 40516 5246
rect 39564 4286 39566 4338
rect 39618 4286 39620 4338
rect 39564 4274 39620 4286
rect 39004 4228 39060 4238
rect 39004 3388 39060 4172
rect 38332 3042 38388 3052
rect 38780 3332 39060 3388
rect 39116 4004 39172 4014
rect 38780 2996 38836 3332
rect 38220 2942 38222 2994
rect 38274 2942 38276 2994
rect 38220 2930 38276 2942
rect 38556 2940 38836 2996
rect 37884 2046 37886 2098
rect 37938 2046 37940 2098
rect 37884 2034 37940 2046
rect 38444 1986 38500 1998
rect 38444 1934 38446 1986
rect 38498 1934 38500 1986
rect 38444 644 38500 1934
rect 38444 578 38500 588
rect 38556 308 38612 2940
rect 38668 2772 38724 2782
rect 38668 532 38724 2716
rect 39116 2100 39172 3948
rect 39116 2034 39172 2044
rect 39676 4004 39732 4014
rect 38780 1988 38836 1998
rect 38780 868 38836 1932
rect 38780 802 38836 812
rect 38668 466 38724 476
rect 38556 242 38612 252
rect 39676 112 39732 3948
rect 40348 3780 40404 3790
rect 40348 3108 40404 3724
rect 40348 3042 40404 3052
rect 40460 2660 40516 5180
rect 41916 5236 41972 7308
rect 42028 7140 42084 7150
rect 42028 6802 42084 7084
rect 42028 6750 42030 6802
rect 42082 6750 42084 6802
rect 42028 6738 42084 6750
rect 41916 5170 41972 5180
rect 42140 5012 42196 7644
rect 42252 6690 42308 8092
rect 42588 8082 42644 8092
rect 42700 8092 42868 8148
rect 42924 8260 42980 8270
rect 42588 7588 42644 7598
rect 42588 7494 42644 7532
rect 42252 6638 42254 6690
rect 42306 6638 42308 6690
rect 42252 6626 42308 6638
rect 42364 6804 42420 6814
rect 42252 6468 42308 6478
rect 42252 5906 42308 6412
rect 42252 5854 42254 5906
rect 42306 5854 42308 5906
rect 42252 5842 42308 5854
rect 42364 5348 42420 6748
rect 42364 5282 42420 5292
rect 42140 4946 42196 4956
rect 41132 4788 41188 4798
rect 40572 2772 40628 2782
rect 40572 2678 40628 2716
rect 40460 2594 40516 2604
rect 40012 2548 40068 2558
rect 40012 2454 40068 2492
rect 41132 2210 41188 4732
rect 42252 4676 42308 4686
rect 41692 4452 41748 4462
rect 41580 3108 41636 3118
rect 41580 2882 41636 3052
rect 41580 2830 41582 2882
rect 41634 2830 41636 2882
rect 41580 2818 41636 2830
rect 41132 2158 41134 2210
rect 41186 2158 41188 2210
rect 41132 2146 41188 2158
rect 41692 2098 41748 4396
rect 42028 3556 42084 3566
rect 42028 3220 42084 3500
rect 41692 2046 41694 2098
rect 41746 2046 41748 2098
rect 41692 2034 41748 2046
rect 41804 3164 42084 3220
rect 41804 1876 41860 3164
rect 41692 1820 41860 1876
rect 42028 2996 42084 3006
rect 41692 112 41748 1820
rect 42028 1540 42084 2940
rect 42028 1474 42084 1484
rect 42140 2546 42196 2558
rect 42140 2494 42142 2546
rect 42194 2494 42196 2546
rect 42140 196 42196 2494
rect 42252 2548 42308 4620
rect 42700 3108 42756 8092
rect 42812 6692 42868 6702
rect 42812 6598 42868 6636
rect 42700 3042 42756 3052
rect 42252 2482 42308 2492
rect 42924 1988 42980 8204
rect 43036 7474 43092 8372
rect 43260 7812 43316 11228
rect 43260 7746 43316 7756
rect 43372 10612 43428 10622
rect 43036 7422 43038 7474
rect 43090 7422 43092 7474
rect 43036 7140 43092 7422
rect 43036 7074 43092 7084
rect 43260 7588 43316 7598
rect 43148 6468 43204 6478
rect 43148 6374 43204 6412
rect 43260 3892 43316 7532
rect 43372 7476 43428 10556
rect 43596 9268 43652 12460
rect 44156 12180 44212 12190
rect 44156 12086 44212 12124
rect 44156 11620 44212 11630
rect 44268 11620 44324 12684
rect 44604 12290 44660 12684
rect 44604 12238 44606 12290
rect 44658 12238 44660 12290
rect 44604 12226 44660 12238
rect 45052 12180 45108 14112
rect 45500 13300 45556 14112
rect 45948 13412 46004 14112
rect 45948 13346 46004 13356
rect 45500 13244 45892 13300
rect 45052 12114 45108 12124
rect 45500 13076 45556 13086
rect 45388 12068 45444 12078
rect 45052 11954 45108 11966
rect 45052 11902 45054 11954
rect 45106 11902 45108 11954
rect 44464 11788 44728 11798
rect 44520 11732 44568 11788
rect 44624 11732 44672 11788
rect 44464 11722 44728 11732
rect 44380 11620 44436 11630
rect 44268 11618 44436 11620
rect 44268 11566 44382 11618
rect 44434 11566 44436 11618
rect 44268 11564 44436 11566
rect 44044 11396 44100 11406
rect 44044 11302 44100 11340
rect 43804 11004 44068 11014
rect 43860 10948 43908 11004
rect 43964 10948 44012 11004
rect 43804 10938 44068 10948
rect 44156 10948 44212 11564
rect 44380 11554 44436 11564
rect 44940 11508 44996 11518
rect 44940 11414 44996 11452
rect 44156 10882 44212 10892
rect 44268 10612 44324 10622
rect 44268 10164 44324 10556
rect 44828 10388 44884 10398
rect 44464 10220 44728 10230
rect 44520 10164 44568 10220
rect 44624 10164 44672 10220
rect 44464 10154 44728 10164
rect 44268 10098 44324 10108
rect 43804 9436 44068 9446
rect 43860 9380 43908 9436
rect 43964 9380 44012 9436
rect 43804 9370 44068 9380
rect 43596 9202 43652 9212
rect 44464 8652 44728 8662
rect 44520 8596 44568 8652
rect 44624 8596 44672 8652
rect 44464 8586 44728 8596
rect 43804 7868 44068 7878
rect 43860 7812 43908 7868
rect 43964 7812 44012 7868
rect 43804 7802 44068 7812
rect 43372 6802 43428 7420
rect 43372 6750 43374 6802
rect 43426 6750 43428 6802
rect 43372 6738 43428 6750
rect 43484 7252 43540 7262
rect 43372 5908 43428 5918
rect 43372 4116 43428 5852
rect 43484 5124 43540 7196
rect 43708 7140 43764 7150
rect 43708 6802 43764 7084
rect 44464 7084 44728 7094
rect 43708 6750 43710 6802
rect 43762 6750 43764 6802
rect 43708 6738 43764 6750
rect 44268 7028 44324 7038
rect 44520 7028 44568 7084
rect 44624 7028 44672 7084
rect 44464 7018 44728 7028
rect 44268 6356 44324 6972
rect 44380 6356 44436 6366
rect 43804 6300 44068 6310
rect 44268 6300 44380 6356
rect 43596 6244 43652 6254
rect 43860 6244 43908 6300
rect 43964 6244 44012 6300
rect 44380 6290 44436 6300
rect 43804 6234 44068 6244
rect 43596 6132 43652 6188
rect 44380 6132 44436 6142
rect 43596 6076 44380 6132
rect 44380 6066 44436 6076
rect 44268 5796 44324 5806
rect 44268 5684 44324 5740
rect 44716 5684 44772 5694
rect 44268 5628 44716 5684
rect 44716 5618 44772 5628
rect 44464 5516 44728 5526
rect 44520 5460 44568 5516
rect 44624 5460 44672 5516
rect 44464 5450 44728 5460
rect 44492 5236 44548 5246
rect 43484 5058 43540 5068
rect 43708 5124 43764 5134
rect 43708 4900 43764 5068
rect 43484 4844 43764 4900
rect 43484 4788 43540 4844
rect 44156 4788 44212 4798
rect 43484 4722 43540 4732
rect 43804 4732 44068 4742
rect 43860 4676 43908 4732
rect 43964 4676 44012 4732
rect 43804 4666 44068 4676
rect 43372 4050 43428 4060
rect 44044 4004 44100 4014
rect 44156 4004 44212 4732
rect 44492 4338 44548 5180
rect 44492 4286 44494 4338
rect 44546 4286 44548 4338
rect 44492 4274 44548 4286
rect 44100 3948 44212 4004
rect 44464 3948 44728 3958
rect 44044 3938 44100 3948
rect 44520 3892 44568 3948
rect 44624 3892 44672 3948
rect 44464 3882 44728 3892
rect 43260 3826 43316 3836
rect 43804 3164 44068 3174
rect 43860 3108 43908 3164
rect 43964 3108 44012 3164
rect 43804 3098 44068 3108
rect 44828 3108 44884 10332
rect 45052 6020 45108 11902
rect 45388 10388 45444 12012
rect 45500 11396 45556 13020
rect 45612 12068 45668 12078
rect 45612 12066 45780 12068
rect 45612 12014 45614 12066
rect 45666 12014 45780 12066
rect 45612 12012 45780 12014
rect 45612 12002 45668 12012
rect 45500 11330 45556 11340
rect 45388 10322 45444 10332
rect 45612 9042 45668 9054
rect 45612 8990 45614 9042
rect 45666 8990 45668 9042
rect 45052 5954 45108 5964
rect 45500 8372 45556 8382
rect 45164 5236 45220 5246
rect 45052 4340 45108 4350
rect 45052 4246 45108 4284
rect 45164 3332 45220 5180
rect 45164 3266 45220 3276
rect 45276 5012 45332 5022
rect 44828 3042 44884 3052
rect 42924 1922 42980 1932
rect 44268 2436 44324 2446
rect 43804 1596 44068 1606
rect 43860 1540 43908 1596
rect 43964 1540 44012 1596
rect 43804 1530 44068 1540
rect 44044 1428 44100 1438
rect 42140 130 42196 140
rect 43708 644 43764 654
rect 43708 112 43764 588
rect 44044 420 44100 1372
rect 44268 1428 44324 2380
rect 44464 2380 44728 2390
rect 44520 2324 44568 2380
rect 44624 2324 44672 2380
rect 44464 2314 44728 2324
rect 45276 1652 45332 4956
rect 45500 4452 45556 8316
rect 45500 4386 45556 4396
rect 45612 3388 45668 8990
rect 45724 7140 45780 12012
rect 45836 11172 45892 13244
rect 45948 12852 46004 12862
rect 45948 12758 46004 12796
rect 46396 12180 46452 14112
rect 46844 13188 46900 14112
rect 46732 13132 46900 13188
rect 46956 13972 47012 13982
rect 46172 12124 46452 12180
rect 46620 12964 46676 12974
rect 45948 11954 46004 11966
rect 45948 11902 45950 11954
rect 46002 11902 46004 11954
rect 45948 11844 46004 11902
rect 45948 11778 46004 11788
rect 46060 11284 46116 11294
rect 46172 11284 46228 12124
rect 46508 12066 46564 12078
rect 46508 12014 46510 12066
rect 46562 12014 46564 12066
rect 46508 11508 46564 12014
rect 46620 11620 46676 12908
rect 46732 11732 46788 13132
rect 46844 12962 46900 12974
rect 46844 12910 46846 12962
rect 46898 12910 46900 12962
rect 46844 11956 46900 12910
rect 46844 11890 46900 11900
rect 46844 11732 46900 11742
rect 46732 11676 46844 11732
rect 46844 11666 46900 11676
rect 46620 11554 46676 11564
rect 46956 11618 47012 13916
rect 47180 13188 47236 13198
rect 46956 11566 46958 11618
rect 47010 11566 47012 11618
rect 46956 11554 47012 11566
rect 47068 11956 47124 11966
rect 46508 11442 46564 11452
rect 46620 11394 46676 11406
rect 46620 11342 46622 11394
rect 46674 11342 46676 11394
rect 46620 11284 46676 11342
rect 46172 11228 46676 11284
rect 46060 11190 46116 11228
rect 45836 11116 46004 11172
rect 45724 7074 45780 7084
rect 45836 6916 45892 6926
rect 45836 6822 45892 6860
rect 45948 6244 46004 11116
rect 46172 11060 46228 11070
rect 46060 10276 46116 10286
rect 46060 9154 46116 10220
rect 46060 9102 46062 9154
rect 46114 9102 46116 9154
rect 46060 9090 46116 9102
rect 45948 6178 46004 6188
rect 46172 4340 46228 11004
rect 47068 10612 47124 11900
rect 47068 10546 47124 10556
rect 46844 10498 46900 10510
rect 46844 10446 46846 10498
rect 46898 10446 46900 10498
rect 46396 10052 46452 10062
rect 46396 9958 46452 9996
rect 46844 8148 46900 10446
rect 47180 10388 47236 13132
rect 47292 10610 47348 14112
rect 47628 13636 47684 13646
rect 47292 10558 47294 10610
rect 47346 10558 47348 10610
rect 47292 10546 47348 10558
rect 47516 11282 47572 11294
rect 47516 11230 47518 11282
rect 47570 11230 47572 11282
rect 47516 10612 47572 11230
rect 47516 10546 47572 10556
rect 47628 10500 47684 13580
rect 47740 10724 47796 14112
rect 47852 13748 47908 13758
rect 47852 12850 47908 13692
rect 48188 13188 48244 14112
rect 48188 13122 48244 13132
rect 47852 12798 47854 12850
rect 47906 12798 47908 12850
rect 47852 12786 47908 12798
rect 47964 12964 48020 12974
rect 47964 12402 48020 12908
rect 47964 12350 47966 12402
rect 48018 12350 48020 12402
rect 47964 12338 48020 12350
rect 48412 12962 48468 12974
rect 48412 12910 48414 12962
rect 48466 12910 48468 12962
rect 48412 12292 48468 12910
rect 48636 12964 48692 14112
rect 49084 13524 49140 14112
rect 49084 13458 49140 13468
rect 49308 13860 49364 13870
rect 48972 13188 49028 13198
rect 48972 13094 49028 13132
rect 48636 12908 49140 12964
rect 49084 12402 49140 12908
rect 49084 12350 49086 12402
rect 49138 12350 49140 12402
rect 49084 12338 49140 12350
rect 48412 12226 48468 12236
rect 48412 12068 48468 12078
rect 48188 11394 48244 11406
rect 48188 11342 48190 11394
rect 48242 11342 48244 11394
rect 48188 10724 48244 11342
rect 47740 10668 47908 10724
rect 47740 10500 47796 10510
rect 47628 10498 47796 10500
rect 47628 10446 47742 10498
rect 47794 10446 47796 10498
rect 47628 10444 47796 10446
rect 47740 10434 47796 10444
rect 47180 10332 47348 10388
rect 46956 10164 47012 10174
rect 46956 9938 47012 10108
rect 46956 9886 46958 9938
rect 47010 9886 47012 9938
rect 46956 9874 47012 9886
rect 46844 8082 46900 8092
rect 47180 9156 47236 9166
rect 47068 7700 47124 7710
rect 46284 6578 46340 6590
rect 46284 6526 46286 6578
rect 46338 6526 46340 6578
rect 46284 4900 46340 6526
rect 47068 6580 47124 7644
rect 47068 6514 47124 6524
rect 47180 5012 47236 9100
rect 47180 4946 47236 4956
rect 46284 4834 46340 4844
rect 46172 4274 46228 4284
rect 47292 3388 47348 10332
rect 47740 8932 47796 8942
rect 47852 8932 47908 10668
rect 48188 10658 48244 10668
rect 48300 10500 48356 10510
rect 48300 10406 48356 10444
rect 48412 9042 48468 12012
rect 48524 12066 48580 12078
rect 48524 12014 48526 12066
rect 48578 12014 48580 12066
rect 48524 11508 48580 12014
rect 49196 11732 49252 11742
rect 48524 11442 48580 11452
rect 49084 11620 49140 11630
rect 48860 11172 48916 11182
rect 48748 10610 48804 10622
rect 48748 10558 48750 10610
rect 48802 10558 48804 10610
rect 48412 8990 48414 9042
rect 48466 8990 48468 9042
rect 48412 8978 48468 8990
rect 48524 9826 48580 9838
rect 48524 9774 48526 9826
rect 48578 9774 48580 9826
rect 47740 8930 47908 8932
rect 47740 8878 47742 8930
rect 47794 8878 47908 8930
rect 47740 8876 47908 8878
rect 47740 8866 47796 8876
rect 48076 8820 48132 8830
rect 48076 8726 48132 8764
rect 48412 8708 48468 8718
rect 48076 7812 48132 7822
rect 47404 5572 47460 5582
rect 47404 5012 47460 5516
rect 47404 4946 47460 4956
rect 45612 3332 45780 3388
rect 45724 1764 45780 3332
rect 47180 3332 47348 3388
rect 47852 3556 47908 3566
rect 47068 1988 47124 1998
rect 47180 1988 47236 3332
rect 47852 2770 47908 3500
rect 48076 3220 48132 7756
rect 48300 7476 48356 7486
rect 48300 6020 48356 7420
rect 48300 5954 48356 5964
rect 48076 3154 48132 3164
rect 48412 2882 48468 8652
rect 48524 4788 48580 9774
rect 48524 4722 48580 4732
rect 48636 6356 48692 6366
rect 48636 2884 48692 6300
rect 48748 2996 48804 10558
rect 48860 9492 48916 11116
rect 49084 11060 49140 11564
rect 49196 11282 49252 11676
rect 49196 11230 49198 11282
rect 49250 11230 49252 11282
rect 49196 11218 49252 11230
rect 49084 11004 49252 11060
rect 49084 10052 49140 10062
rect 49084 9938 49140 9996
rect 49084 9886 49086 9938
rect 49138 9886 49140 9938
rect 49084 9874 49140 9886
rect 48860 9426 48916 9436
rect 48972 9044 49028 9054
rect 48972 8950 49028 8988
rect 49084 8820 49140 8830
rect 48972 5908 49028 5918
rect 48972 5814 49028 5852
rect 48748 2930 48804 2940
rect 48412 2830 48414 2882
rect 48466 2830 48468 2882
rect 48412 2818 48468 2830
rect 48524 2828 48692 2884
rect 47852 2718 47854 2770
rect 47906 2718 47908 2770
rect 47852 2706 47908 2718
rect 47068 1986 47236 1988
rect 47068 1934 47070 1986
rect 47122 1934 47236 1986
rect 47068 1932 47236 1934
rect 47068 1922 47124 1932
rect 45276 1586 45332 1596
rect 45612 1708 45780 1764
rect 47404 1874 47460 1886
rect 47404 1822 47406 1874
rect 47458 1822 47460 1874
rect 44268 1362 44324 1372
rect 44464 812 44728 822
rect 44520 756 44568 812
rect 44624 756 44672 812
rect 44464 746 44728 756
rect 45612 644 45668 1708
rect 45612 578 45668 588
rect 45724 1540 45780 1550
rect 44044 354 44100 364
rect 45724 112 45780 1484
rect 47404 532 47460 1822
rect 48524 868 48580 2828
rect 48636 2660 48692 2670
rect 48636 1092 48692 2604
rect 49084 2210 49140 8764
rect 49196 7476 49252 11004
rect 49308 9042 49364 13804
rect 49532 11620 49588 14112
rect 49980 13076 50036 14112
rect 49980 13010 50036 13020
rect 50428 12404 50484 14112
rect 50428 12338 50484 12348
rect 50652 12962 50708 12974
rect 50652 12910 50654 12962
rect 50706 12910 50708 12962
rect 49532 11554 49588 11564
rect 50092 12066 50148 12078
rect 50092 12014 50094 12066
rect 50146 12014 50148 12066
rect 49756 11394 49812 11406
rect 49756 11342 49758 11394
rect 49810 11342 49812 11394
rect 49644 11060 49700 11070
rect 49644 10834 49700 11004
rect 49644 10782 49646 10834
rect 49698 10782 49700 10834
rect 49644 10770 49700 10782
rect 49756 10164 49812 11342
rect 49756 10098 49812 10108
rect 49420 9826 49476 9838
rect 49420 9774 49422 9826
rect 49474 9774 49476 9826
rect 49420 9604 49476 9774
rect 49420 9538 49476 9548
rect 49308 8990 49310 9042
rect 49362 8990 49364 9042
rect 49308 8978 49364 8990
rect 49980 9268 50036 9278
rect 49868 8930 49924 8942
rect 49868 8878 49870 8930
rect 49922 8878 49924 8930
rect 49196 7410 49252 7420
rect 49644 8820 49700 8830
rect 49420 6020 49476 6030
rect 49420 5926 49476 5964
rect 49084 2158 49086 2210
rect 49138 2158 49140 2210
rect 49084 2146 49140 2158
rect 49308 1986 49364 1998
rect 49308 1934 49310 1986
rect 49362 1934 49364 1986
rect 49308 1652 49364 1934
rect 49308 1586 49364 1596
rect 48636 1026 48692 1036
rect 48524 802 48580 812
rect 47404 466 47460 476
rect 49644 420 49700 8764
rect 49868 8484 49924 8878
rect 49868 8418 49924 8428
rect 49756 8258 49812 8270
rect 49756 8206 49758 8258
rect 49810 8206 49812 8258
rect 49756 980 49812 8206
rect 49980 7474 50036 9212
rect 49980 7422 49982 7474
rect 50034 7422 50036 7474
rect 49980 7410 50036 7422
rect 49868 6916 49924 6926
rect 49868 4338 49924 6860
rect 50092 5124 50148 12014
rect 50428 11956 50484 11966
rect 50428 11862 50484 11900
rect 50316 11620 50372 11630
rect 50316 11526 50372 11564
rect 50204 9940 50260 9950
rect 50204 9846 50260 9884
rect 50204 8932 50260 8942
rect 50204 8838 50260 8876
rect 50316 8372 50372 8382
rect 50316 8278 50372 8316
rect 50540 7588 50596 7598
rect 50540 7494 50596 7532
rect 50540 6692 50596 6702
rect 50540 6598 50596 6636
rect 50092 5058 50148 5068
rect 50652 5012 50708 12910
rect 50876 12740 50932 14112
rect 51100 13524 51156 13534
rect 51100 13186 51156 13468
rect 51100 13134 51102 13186
rect 51154 13134 51156 13186
rect 51100 13122 51156 13134
rect 50876 12674 50932 12684
rect 50988 12068 51044 12078
rect 50988 12066 51268 12068
rect 50988 12014 50990 12066
rect 51042 12014 51268 12066
rect 50988 12012 51268 12014
rect 50988 12002 51044 12012
rect 50876 11396 50932 11406
rect 49868 4286 49870 4338
rect 49922 4286 49924 4338
rect 49868 4274 49924 4286
rect 50316 4956 50708 5012
rect 50764 11172 50820 11182
rect 49868 2548 49924 2558
rect 49868 2210 49924 2492
rect 49868 2158 49870 2210
rect 49922 2158 49924 2210
rect 49868 2146 49924 2158
rect 50316 1874 50372 4956
rect 50428 4226 50484 4238
rect 50428 4174 50430 4226
rect 50482 4174 50484 4226
rect 50428 3668 50484 4174
rect 50428 3602 50484 3612
rect 50652 3332 50708 3342
rect 50652 2212 50708 3276
rect 50764 2772 50820 11116
rect 50876 10834 50932 11340
rect 50876 10782 50878 10834
rect 50930 10782 50932 10834
rect 50876 10770 50932 10782
rect 50988 9828 51044 9838
rect 50988 9734 51044 9772
rect 51100 9156 51156 9166
rect 51100 9062 51156 9100
rect 50988 8258 51044 8270
rect 50988 8206 50990 8258
rect 51042 8206 51044 8258
rect 50876 7476 50932 7486
rect 50876 7382 50932 7420
rect 50988 6916 51044 8206
rect 50988 6850 51044 6860
rect 51100 6692 51156 6702
rect 51100 6598 51156 6636
rect 50876 2772 50932 2782
rect 50764 2770 50932 2772
rect 50764 2718 50878 2770
rect 50930 2718 50932 2770
rect 50764 2716 50932 2718
rect 50876 2706 50932 2716
rect 51212 2772 51268 12012
rect 51324 11620 51380 14112
rect 51324 11554 51380 11564
rect 51660 13412 51716 13422
rect 51324 11394 51380 11406
rect 51324 11342 51326 11394
rect 51378 11342 51380 11394
rect 51324 10276 51380 11342
rect 51436 10500 51492 10510
rect 51436 10406 51492 10444
rect 51324 10210 51380 10220
rect 51548 10276 51604 10286
rect 51436 7364 51492 7374
rect 51436 7270 51492 7308
rect 51436 6690 51492 6702
rect 51436 6638 51438 6690
rect 51490 6638 51492 6690
rect 51212 2706 51268 2716
rect 51324 3332 51380 3342
rect 50764 2212 50820 2222
rect 50652 2210 50820 2212
rect 50652 2158 50766 2210
rect 50818 2158 50820 2210
rect 50652 2156 50820 2158
rect 50764 2146 50820 2156
rect 51324 2098 51380 3276
rect 51436 2884 51492 6638
rect 51548 3556 51604 10220
rect 51660 3778 51716 13356
rect 51772 13300 51828 14112
rect 51772 13234 51828 13244
rect 52220 13188 52276 14112
rect 52220 13122 52276 13132
rect 52332 12964 52388 12974
rect 52668 12964 52724 14112
rect 53116 13412 53172 14112
rect 53116 13346 53172 13356
rect 52892 13076 52948 13086
rect 52892 12982 52948 13020
rect 52332 12962 52500 12964
rect 52332 12910 52334 12962
rect 52386 12910 52500 12962
rect 52332 12908 52500 12910
rect 52668 12908 52836 12964
rect 52332 12898 52388 12908
rect 52108 12740 52164 12750
rect 52108 11506 52164 12684
rect 52108 11454 52110 11506
rect 52162 11454 52164 11506
rect 52108 11442 52164 11454
rect 52220 12178 52276 12190
rect 52220 12126 52222 12178
rect 52274 12126 52276 12178
rect 51996 10724 52052 10734
rect 51884 10500 51940 10510
rect 51772 10276 51828 10286
rect 51772 8370 51828 10220
rect 51772 8318 51774 8370
rect 51826 8318 51828 8370
rect 51772 8306 51828 8318
rect 51884 6578 51940 10444
rect 51996 9714 52052 10668
rect 52108 10612 52164 10622
rect 52108 10518 52164 10556
rect 51996 9662 51998 9714
rect 52050 9662 52052 9714
rect 51996 9650 52052 9662
rect 51996 9044 52052 9054
rect 51996 8950 52052 8988
rect 52108 8932 52164 8942
rect 52108 7700 52164 8876
rect 52220 8372 52276 12126
rect 52220 8306 52276 8316
rect 52332 9492 52388 9502
rect 52108 7634 52164 7644
rect 52108 7474 52164 7486
rect 52108 7422 52110 7474
rect 52162 7422 52164 7474
rect 52108 7252 52164 7422
rect 52108 7186 52164 7196
rect 51884 6526 51886 6578
rect 51938 6526 51940 6578
rect 51884 6514 51940 6526
rect 52108 5906 52164 5918
rect 52108 5854 52110 5906
rect 52162 5854 52164 5906
rect 52108 5236 52164 5854
rect 52108 5170 52164 5180
rect 51660 3726 51662 3778
rect 51714 3726 51716 3778
rect 51660 3714 51716 3726
rect 51884 5124 51940 5134
rect 51548 3500 51828 3556
rect 51436 2828 51604 2884
rect 51324 2046 51326 2098
rect 51378 2046 51380 2098
rect 51324 2034 51380 2046
rect 51436 2658 51492 2670
rect 51436 2606 51438 2658
rect 51490 2606 51492 2658
rect 50316 1822 50318 1874
rect 50370 1822 50372 1874
rect 50316 1810 50372 1822
rect 51436 1876 51492 2606
rect 51436 1810 51492 1820
rect 51548 1540 51604 2828
rect 51660 2100 51716 2110
rect 51660 2006 51716 2044
rect 51548 1474 51604 1484
rect 50988 1316 51044 1326
rect 50988 1202 51044 1260
rect 50988 1150 50990 1202
rect 51042 1150 51044 1202
rect 50988 1138 51044 1150
rect 49756 914 49812 924
rect 49644 354 49700 364
rect 49756 756 49812 766
rect 47740 196 47796 206
rect 47740 112 47796 140
rect 49756 112 49812 700
rect 51772 112 51828 3500
rect 51884 2100 51940 5068
rect 51996 5122 52052 5134
rect 51996 5070 51998 5122
rect 52050 5070 52052 5122
rect 51996 5012 52052 5070
rect 51996 4956 52164 5012
rect 51996 2772 52052 2782
rect 51996 2678 52052 2716
rect 51884 2034 51940 2044
rect 52108 1428 52164 4956
rect 52332 4900 52388 9436
rect 52444 7588 52500 12908
rect 52556 12404 52612 12414
rect 52556 12310 52612 12348
rect 52556 11620 52612 11630
rect 52780 11620 52836 12908
rect 53564 12292 53620 14112
rect 53788 13524 53844 13534
rect 53564 12236 53732 12292
rect 53564 12066 53620 12078
rect 53564 12014 53566 12066
rect 53618 12014 53620 12066
rect 53452 11620 53508 11630
rect 52780 11618 53508 11620
rect 52780 11566 53454 11618
rect 53506 11566 53508 11618
rect 52780 11564 53508 11566
rect 52556 10834 52612 11564
rect 53452 11554 53508 11564
rect 52892 11396 52948 11406
rect 52556 10782 52558 10834
rect 52610 10782 52612 10834
rect 52556 10770 52612 10782
rect 52780 11394 52948 11396
rect 52780 11342 52894 11394
rect 52946 11342 52948 11394
rect 52780 11340 52948 11342
rect 52556 9826 52612 9838
rect 52556 9774 52558 9826
rect 52610 9774 52612 9826
rect 52556 8484 52612 9774
rect 52556 8418 52612 8428
rect 52556 8260 52612 8270
rect 52556 8166 52612 8204
rect 52444 7522 52500 7532
rect 52556 6690 52612 6702
rect 52556 6638 52558 6690
rect 52610 6638 52612 6690
rect 52556 5684 52612 6638
rect 52556 5618 52612 5628
rect 52332 4834 52388 4844
rect 52444 5010 52500 5022
rect 52444 4958 52446 5010
rect 52498 4958 52500 5010
rect 52332 4340 52388 4350
rect 52220 3556 52276 3566
rect 52220 3462 52276 3500
rect 52332 2660 52388 4284
rect 52332 2594 52388 2604
rect 52220 2100 52276 2110
rect 52220 2006 52276 2044
rect 52108 1362 52164 1372
rect 51996 1314 52052 1326
rect 51996 1262 51998 1314
rect 52050 1262 52052 1314
rect 51996 980 52052 1262
rect 52444 1204 52500 4958
rect 52556 4676 52612 4686
rect 52556 3666 52612 4620
rect 52668 4228 52724 4238
rect 52668 4134 52724 4172
rect 52556 3614 52558 3666
rect 52610 3614 52612 3666
rect 52556 3602 52612 3614
rect 52780 3332 52836 11340
rect 52892 11330 52948 11340
rect 53564 10724 53620 12014
rect 52892 10668 53620 10724
rect 52892 6692 52948 10668
rect 53564 10500 53620 10510
rect 53452 10498 53620 10500
rect 53452 10446 53566 10498
rect 53618 10446 53620 10498
rect 53452 10444 53620 10446
rect 53004 9268 53060 9278
rect 53004 9174 53060 9212
rect 53340 8372 53396 8382
rect 53340 8278 53396 8316
rect 53004 7924 53060 7934
rect 53004 7698 53060 7868
rect 53004 7646 53006 7698
rect 53058 7646 53060 7698
rect 53004 7634 53060 7646
rect 53452 7476 53508 10444
rect 53564 10434 53620 10444
rect 53564 9716 53620 9726
rect 53676 9716 53732 12236
rect 53788 9940 53844 13468
rect 53788 9874 53844 9884
rect 53900 10500 53956 10510
rect 53564 9714 53732 9716
rect 53564 9662 53566 9714
rect 53618 9662 53732 9714
rect 53564 9660 53732 9662
rect 53564 9650 53620 9660
rect 53676 9492 53732 9502
rect 53564 8930 53620 8942
rect 53564 8878 53566 8930
rect 53618 8878 53620 8930
rect 53564 8596 53620 8878
rect 53564 8530 53620 8540
rect 52892 6626 52948 6636
rect 53340 7420 53508 7476
rect 53228 6580 53284 6590
rect 53004 6244 53060 6254
rect 53004 6130 53060 6188
rect 53004 6078 53006 6130
rect 53058 6078 53060 6130
rect 53004 6066 53060 6078
rect 53228 5346 53284 6524
rect 53228 5294 53230 5346
rect 53282 5294 53284 5346
rect 53228 5282 53284 5294
rect 53116 4452 53172 4462
rect 53116 4358 53172 4396
rect 52780 3266 52836 3276
rect 52556 3220 52612 3230
rect 52556 2098 52612 3164
rect 53340 2884 53396 7420
rect 53564 7364 53620 7374
rect 53452 7362 53620 7364
rect 53452 7310 53566 7362
rect 53618 7310 53620 7362
rect 53452 7308 53620 7310
rect 53452 6132 53508 7308
rect 53564 7298 53620 7308
rect 53564 6580 53620 6590
rect 53564 6486 53620 6524
rect 53452 6066 53508 6076
rect 53676 5906 53732 9436
rect 53900 6580 53956 10444
rect 54012 9268 54068 14112
rect 54124 13300 54180 13310
rect 54124 12402 54180 13244
rect 54348 12964 54404 12974
rect 54124 12350 54126 12402
rect 54178 12350 54180 12402
rect 54124 12338 54180 12350
rect 54236 12962 54404 12964
rect 54236 12910 54350 12962
rect 54402 12910 54404 12962
rect 54236 12908 54404 12910
rect 54012 9202 54068 9212
rect 54124 9826 54180 9838
rect 54124 9774 54126 9826
rect 54178 9774 54180 9826
rect 54124 8428 54180 9774
rect 53900 6514 53956 6524
rect 54012 8372 54180 8428
rect 53676 5854 53678 5906
rect 53730 5854 53732 5906
rect 53676 5842 53732 5854
rect 53676 5012 53732 5022
rect 53676 4918 53732 4956
rect 53564 4564 53620 4574
rect 53564 4338 53620 4508
rect 53564 4286 53566 4338
rect 53618 4286 53620 4338
rect 53564 4274 53620 4286
rect 53564 3444 53620 3454
rect 53564 3350 53620 3388
rect 53340 2818 53396 2828
rect 53564 3108 53620 3118
rect 54012 3108 54068 8372
rect 54124 8258 54180 8270
rect 54124 8206 54126 8258
rect 54178 8206 54180 8258
rect 54124 8036 54180 8206
rect 54124 7970 54180 7980
rect 54124 6690 54180 6702
rect 54124 6638 54126 6690
rect 54178 6638 54180 6690
rect 54124 5796 54180 6638
rect 54124 5730 54180 5740
rect 54124 5122 54180 5134
rect 54124 5070 54126 5122
rect 54178 5070 54180 5122
rect 54124 4900 54180 5070
rect 54124 4834 54180 4844
rect 54236 4340 54292 12908
rect 54348 12898 54404 12908
rect 54460 12292 54516 14112
rect 54908 13748 54964 14112
rect 54908 13682 54964 13692
rect 54908 13188 54964 13198
rect 54908 13094 54964 13132
rect 55356 12964 55412 14112
rect 55356 12898 55412 12908
rect 55692 13412 55748 13422
rect 54348 12236 54516 12292
rect 54684 12628 54740 12638
rect 54348 11396 54404 12236
rect 54348 11330 54404 11340
rect 54460 11394 54516 11406
rect 54460 11342 54462 11394
rect 54514 11342 54516 11394
rect 54348 8930 54404 8942
rect 54348 8878 54350 8930
rect 54402 8878 54404 8930
rect 54348 8596 54404 8878
rect 54348 8530 54404 8540
rect 54236 4274 54292 4284
rect 54124 3780 54180 3790
rect 54124 3666 54180 3724
rect 54124 3614 54126 3666
rect 54178 3614 54180 3666
rect 54124 3602 54180 3614
rect 53564 2770 53620 3052
rect 53564 2718 53566 2770
rect 53618 2718 53620 2770
rect 53564 2706 53620 2718
rect 53676 3052 54068 3108
rect 52780 2660 52836 2670
rect 52780 2566 52836 2604
rect 52556 2046 52558 2098
rect 52610 2046 52612 2098
rect 52556 2034 52612 2046
rect 53564 1876 53620 1886
rect 53564 1782 53620 1820
rect 53564 1428 53620 1438
rect 53564 1334 53620 1372
rect 52556 1204 52612 1214
rect 52444 1202 52612 1204
rect 52444 1150 52558 1202
rect 52610 1150 52612 1202
rect 52444 1148 52612 1150
rect 52556 1138 52612 1148
rect 51996 914 52052 924
rect 53676 644 53732 3052
rect 54124 1986 54180 1998
rect 54124 1934 54126 1986
rect 54178 1934 54180 1986
rect 54124 1764 54180 1934
rect 54124 1698 54180 1708
rect 53676 578 53732 588
rect 53788 868 53844 878
rect 53788 112 53844 812
rect 54460 756 54516 11342
rect 54572 10722 54628 10734
rect 54572 10670 54574 10722
rect 54626 10670 54628 10722
rect 54572 10164 54628 10670
rect 54684 10276 54740 12572
rect 55692 12402 55748 13356
rect 55692 12350 55694 12402
rect 55746 12350 55748 12402
rect 55692 12338 55748 12350
rect 55244 12178 55300 12190
rect 55244 12126 55246 12178
rect 55298 12126 55300 12178
rect 55020 11508 55076 11518
rect 55020 11414 55076 11452
rect 55132 10836 55188 10846
rect 55132 10610 55188 10780
rect 55132 10558 55134 10610
rect 55186 10558 55188 10610
rect 55132 10546 55188 10558
rect 54684 10210 54740 10220
rect 54572 10098 54628 10108
rect 55244 10052 55300 12126
rect 55580 11284 55636 11294
rect 55244 9986 55300 9996
rect 55468 10388 55524 10398
rect 55132 9602 55188 9614
rect 55132 9550 55134 9602
rect 55186 9550 55188 9602
rect 55132 9492 55188 9550
rect 55132 9426 55188 9436
rect 55132 8932 55188 8942
rect 55132 8838 55188 8876
rect 55468 8372 55524 10332
rect 55132 8316 55524 8372
rect 55580 8372 55636 11228
rect 55804 10500 55860 14112
rect 56252 12852 56308 14112
rect 56252 12786 56308 12796
rect 56364 13972 56420 13982
rect 55804 10434 55860 10444
rect 56140 10722 56196 10734
rect 56140 10670 56142 10722
rect 56194 10670 56196 10722
rect 56140 9044 56196 10670
rect 56364 9156 56420 13916
rect 56364 9090 56420 9100
rect 56140 8978 56196 8988
rect 55132 8146 55188 8316
rect 55580 8306 55636 8316
rect 55916 8930 55972 8942
rect 55916 8878 55918 8930
rect 55970 8878 55972 8930
rect 55132 8094 55134 8146
rect 55186 8094 55188 8146
rect 55132 8082 55188 8094
rect 55916 8148 55972 8878
rect 55916 8082 55972 8092
rect 56140 7700 56196 7710
rect 56140 7606 56196 7644
rect 54572 7586 54628 7598
rect 54572 7534 54574 7586
rect 54626 7534 54628 7586
rect 54572 7252 54628 7534
rect 54572 7186 54628 7196
rect 55244 7474 55300 7486
rect 55244 7422 55246 7474
rect 55298 7422 55300 7474
rect 55132 6466 55188 6478
rect 55132 6414 55134 6466
rect 55186 6414 55188 6466
rect 55132 6356 55188 6414
rect 55244 6468 55300 7422
rect 55244 6402 55300 6412
rect 55356 7140 55412 7150
rect 55132 6290 55188 6300
rect 54572 6018 54628 6030
rect 54572 5966 54574 6018
rect 54626 5966 54628 6018
rect 54572 5908 54628 5966
rect 54572 5842 54628 5852
rect 55132 5794 55188 5806
rect 55132 5742 55134 5794
rect 55186 5742 55188 5794
rect 55132 5348 55188 5742
rect 55132 5282 55188 5292
rect 54908 5124 54964 5134
rect 54908 5030 54964 5068
rect 54572 4564 54628 4574
rect 54572 4470 54628 4508
rect 55132 4226 55188 4238
rect 55132 4174 55134 4226
rect 55186 4174 55188 4226
rect 55132 4116 55188 4174
rect 55132 4050 55188 4060
rect 54908 3668 54964 3678
rect 54908 3574 54964 3612
rect 54572 3220 54628 3230
rect 54572 2994 54628 3164
rect 54572 2942 54574 2994
rect 54626 2942 54628 2994
rect 54572 2930 54628 2942
rect 55356 2770 55412 7084
rect 56140 6804 56196 6814
rect 56140 6130 56196 6748
rect 56700 6244 56756 14112
rect 57036 13076 57092 13086
rect 57036 11060 57092 13020
rect 57036 10994 57092 11004
rect 57260 12180 57316 12190
rect 57260 7924 57316 12124
rect 57260 7858 57316 7868
rect 56700 6178 56756 6188
rect 56140 6078 56142 6130
rect 56194 6078 56196 6130
rect 56140 6066 56196 6078
rect 56140 5460 56196 5470
rect 56140 4562 56196 5404
rect 56140 4510 56142 4562
rect 56194 4510 56196 4562
rect 56140 4498 56196 4510
rect 56140 4116 56196 4126
rect 56140 2994 56196 4060
rect 56140 2942 56142 2994
rect 56194 2942 56196 2994
rect 56140 2930 56196 2942
rect 57036 3444 57092 3454
rect 55356 2718 55358 2770
rect 55410 2718 55412 2770
rect 55356 2706 55412 2718
rect 56140 2772 56196 2782
rect 54908 2324 54964 2334
rect 54908 2098 54964 2268
rect 54908 2046 54910 2098
rect 54962 2046 54964 2098
rect 54908 2034 54964 2046
rect 56140 1426 56196 2716
rect 56140 1374 56142 1426
rect 56194 1374 56196 1426
rect 56140 1362 56196 1374
rect 56924 2660 56980 2670
rect 55132 1204 55188 1214
rect 55132 1110 55188 1148
rect 54460 690 54516 700
rect 55804 1092 55860 1102
rect 55804 112 55860 1036
rect 32284 18 32340 28
rect 33600 0 33712 112
rect 35616 0 35728 112
rect 37632 0 37744 112
rect 39648 0 39760 112
rect 41664 0 41776 112
rect 43680 0 43792 112
rect 45696 0 45808 112
rect 47712 0 47824 112
rect 49728 0 49840 112
rect 51744 0 51856 112
rect 53760 0 53872 112
rect 55776 0 55888 112
rect 56924 84 56980 2604
rect 57036 532 57092 3388
rect 57036 466 57092 476
rect 56924 18 56980 28
<< via2 >>
rect 21084 14140 21140 14196
rect 588 13020 644 13076
rect 252 12124 308 12180
rect 1148 11788 1204 11844
rect 1484 13468 1540 13524
rect 252 7980 308 8036
rect 812 9212 868 9268
rect 1036 8988 1092 9044
rect 1148 10780 1204 10836
rect 1036 7644 1092 7700
rect 1036 7196 1092 7252
rect 1036 6300 1092 6356
rect 1596 11900 1652 11956
rect 1932 11676 1988 11732
rect 1484 10780 1540 10836
rect 1484 10108 1540 10164
rect 1596 9772 1652 9828
rect 1820 11228 1876 11284
rect 2380 13916 2436 13972
rect 2156 13356 2212 13412
rect 2268 12402 2324 12404
rect 2268 12350 2270 12402
rect 2270 12350 2322 12402
rect 2322 12350 2324 12402
rect 2268 12348 2324 12350
rect 2268 11900 2324 11956
rect 2156 11788 2212 11844
rect 1932 10444 1988 10500
rect 1932 9324 1988 9380
rect 2268 9548 2324 9604
rect 1596 7196 1652 7252
rect 1372 6524 1428 6580
rect 812 4060 868 4116
rect 1820 6748 1876 6804
rect 1932 6076 1988 6132
rect 2828 12684 2884 12740
rect 3612 13468 3668 13524
rect 3388 12348 3444 12404
rect 3500 12572 3556 12628
rect 2940 12124 2996 12180
rect 3388 12124 3444 12180
rect 2716 10668 2772 10724
rect 2828 10610 2884 10612
rect 2828 10558 2830 10610
rect 2830 10558 2882 10610
rect 2882 10558 2884 10610
rect 2828 10556 2884 10558
rect 2380 9324 2436 9380
rect 2716 10444 2772 10500
rect 2380 7532 2436 7588
rect 2604 8092 2660 8148
rect 2492 6636 2548 6692
rect 2492 5292 2548 5348
rect 1708 4844 1764 4900
rect 2268 4508 2324 4564
rect 1484 4060 1540 4116
rect 1596 3724 1652 3780
rect 1372 3164 1428 3220
rect 1260 2828 1316 2884
rect 2492 4508 2548 4564
rect 2828 10332 2884 10388
rect 2940 8540 2996 8596
rect 3724 13186 3780 13188
rect 3724 13134 3726 13186
rect 3726 13134 3778 13186
rect 3778 13134 3780 13186
rect 3724 13132 3780 13134
rect 4732 13468 4788 13524
rect 4284 13356 4340 13412
rect 4464 13354 4520 13356
rect 4464 13302 4466 13354
rect 4466 13302 4518 13354
rect 4518 13302 4520 13354
rect 4464 13300 4520 13302
rect 4568 13354 4624 13356
rect 4568 13302 4570 13354
rect 4570 13302 4622 13354
rect 4622 13302 4624 13354
rect 4568 13300 4624 13302
rect 4672 13354 4728 13356
rect 4672 13302 4674 13354
rect 4674 13302 4726 13354
rect 4726 13302 4728 13354
rect 4672 13300 4728 13302
rect 4284 12962 4340 12964
rect 4284 12910 4286 12962
rect 4286 12910 4338 12962
rect 4338 12910 4340 12962
rect 4284 12908 4340 12910
rect 3804 12570 3860 12572
rect 3804 12518 3806 12570
rect 3806 12518 3858 12570
rect 3858 12518 3860 12570
rect 3804 12516 3860 12518
rect 3908 12570 3964 12572
rect 3908 12518 3910 12570
rect 3910 12518 3962 12570
rect 3962 12518 3964 12570
rect 3908 12516 3964 12518
rect 4012 12570 4068 12572
rect 4012 12518 4014 12570
rect 4014 12518 4066 12570
rect 4066 12518 4068 12570
rect 4012 12516 4068 12518
rect 3804 11002 3860 11004
rect 3804 10950 3806 11002
rect 3806 10950 3858 11002
rect 3858 10950 3860 11002
rect 3804 10948 3860 10950
rect 3908 11002 3964 11004
rect 3908 10950 3910 11002
rect 3910 10950 3962 11002
rect 3962 10950 3964 11002
rect 3908 10948 3964 10950
rect 4012 11002 4068 11004
rect 4012 10950 4014 11002
rect 4014 10950 4066 11002
rect 4066 10950 4068 11002
rect 4012 10948 4068 10950
rect 3612 10444 3668 10500
rect 4172 10668 4228 10724
rect 3804 9434 3860 9436
rect 3804 9382 3806 9434
rect 3806 9382 3858 9434
rect 3858 9382 3860 9434
rect 3804 9380 3860 9382
rect 3908 9434 3964 9436
rect 3908 9382 3910 9434
rect 3910 9382 3962 9434
rect 3962 9382 3964 9434
rect 3908 9380 3964 9382
rect 4012 9434 4068 9436
rect 4012 9382 4014 9434
rect 4014 9382 4066 9434
rect 4066 9382 4068 9434
rect 4012 9380 4068 9382
rect 3836 9212 3892 9268
rect 3500 8930 3556 8932
rect 3500 8878 3502 8930
rect 3502 8878 3554 8930
rect 3554 8878 3556 8930
rect 3500 8876 3556 8878
rect 3164 8258 3220 8260
rect 3164 8206 3166 8258
rect 3166 8206 3218 8258
rect 3218 8206 3220 8258
rect 3164 8204 3220 8206
rect 3500 8146 3556 8148
rect 3500 8094 3502 8146
rect 3502 8094 3554 8146
rect 3554 8094 3556 8146
rect 3500 8092 3556 8094
rect 3052 5740 3108 5796
rect 3164 7644 3220 7700
rect 4060 8370 4116 8372
rect 4060 8318 4062 8370
rect 4062 8318 4114 8370
rect 4114 8318 4116 8370
rect 4060 8316 4116 8318
rect 3804 7866 3860 7868
rect 3804 7814 3806 7866
rect 3806 7814 3858 7866
rect 3858 7814 3860 7866
rect 3804 7812 3860 7814
rect 3908 7866 3964 7868
rect 3908 7814 3910 7866
rect 3910 7814 3962 7866
rect 3962 7814 3964 7866
rect 3908 7812 3964 7814
rect 4012 7866 4068 7868
rect 4012 7814 4014 7866
rect 4014 7814 4066 7866
rect 4066 7814 4068 7866
rect 4012 7812 4068 7814
rect 5068 12290 5124 12292
rect 5068 12238 5070 12290
rect 5070 12238 5122 12290
rect 5122 12238 5124 12290
rect 5068 12236 5124 12238
rect 4396 12178 4452 12180
rect 4396 12126 4398 12178
rect 4398 12126 4450 12178
rect 4450 12126 4452 12178
rect 4396 12124 4452 12126
rect 4956 12012 5012 12068
rect 4464 11786 4520 11788
rect 4464 11734 4466 11786
rect 4466 11734 4518 11786
rect 4518 11734 4520 11786
rect 4464 11732 4520 11734
rect 4568 11786 4624 11788
rect 4568 11734 4570 11786
rect 4570 11734 4622 11786
rect 4622 11734 4624 11786
rect 4568 11732 4624 11734
rect 4672 11786 4728 11788
rect 4672 11734 4674 11786
rect 4674 11734 4726 11786
rect 4726 11734 4728 11786
rect 4672 11732 4728 11734
rect 4620 11618 4676 11620
rect 4620 11566 4622 11618
rect 4622 11566 4674 11618
rect 4674 11566 4676 11618
rect 4620 11564 4676 11566
rect 4396 10668 4452 10724
rect 5628 13132 5684 13188
rect 5964 13186 6020 13188
rect 5964 13134 5966 13186
rect 5966 13134 6018 13186
rect 6018 13134 6020 13186
rect 5964 13132 6020 13134
rect 5964 12908 6020 12964
rect 5180 11564 5236 11620
rect 5180 10892 5236 10948
rect 5292 11340 5348 11396
rect 4956 10556 5012 10612
rect 4464 10218 4520 10220
rect 4464 10166 4466 10218
rect 4466 10166 4518 10218
rect 4518 10166 4520 10218
rect 4464 10164 4520 10166
rect 4568 10218 4624 10220
rect 4568 10166 4570 10218
rect 4570 10166 4622 10218
rect 4622 10166 4624 10218
rect 4568 10164 4624 10166
rect 4672 10218 4728 10220
rect 4672 10166 4674 10218
rect 4674 10166 4726 10218
rect 4726 10166 4728 10218
rect 4672 10164 4728 10166
rect 5068 9884 5124 9940
rect 5180 10444 5236 10500
rect 4396 8764 4452 8820
rect 4464 8650 4520 8652
rect 4464 8598 4466 8650
rect 4466 8598 4518 8650
rect 4518 8598 4520 8650
rect 4464 8596 4520 8598
rect 4568 8650 4624 8652
rect 4568 8598 4570 8650
rect 4570 8598 4622 8650
rect 4622 8598 4624 8650
rect 4568 8596 4624 8598
rect 4672 8650 4728 8652
rect 4672 8598 4674 8650
rect 4674 8598 4726 8650
rect 4726 8598 4728 8650
rect 4672 8596 4728 8598
rect 4396 7980 4452 8036
rect 4172 7420 4228 7476
rect 3276 5852 3332 5908
rect 3804 6298 3860 6300
rect 3804 6246 3806 6298
rect 3806 6246 3858 6298
rect 3858 6246 3860 6298
rect 3804 6244 3860 6246
rect 3908 6298 3964 6300
rect 3908 6246 3910 6298
rect 3910 6246 3962 6298
rect 3962 6246 3964 6298
rect 3908 6244 3964 6246
rect 4012 6298 4068 6300
rect 4012 6246 4014 6298
rect 4014 6246 4066 6298
rect 4066 6246 4068 6298
rect 4012 6244 4068 6246
rect 3388 5628 3444 5684
rect 3164 5404 3220 5460
rect 3804 4730 3860 4732
rect 3804 4678 3806 4730
rect 3806 4678 3858 4730
rect 3858 4678 3860 4730
rect 3804 4676 3860 4678
rect 3908 4730 3964 4732
rect 3908 4678 3910 4730
rect 3910 4678 3962 4730
rect 3962 4678 3964 4730
rect 3908 4676 3964 4678
rect 4012 4730 4068 4732
rect 4012 4678 4014 4730
rect 4014 4678 4066 4730
rect 4066 4678 4068 4730
rect 4012 4676 4068 4678
rect 2604 4284 2660 4340
rect 3804 3162 3860 3164
rect 3804 3110 3806 3162
rect 3806 3110 3858 3162
rect 3858 3110 3860 3162
rect 3804 3108 3860 3110
rect 3908 3162 3964 3164
rect 3908 3110 3910 3162
rect 3910 3110 3962 3162
rect 3962 3110 3964 3162
rect 3908 3108 3964 3110
rect 4012 3162 4068 3164
rect 4012 3110 4014 3162
rect 4014 3110 4066 3162
rect 4066 3110 4068 3162
rect 4012 3108 4068 3110
rect 4464 7082 4520 7084
rect 4464 7030 4466 7082
rect 4466 7030 4518 7082
rect 4518 7030 4520 7082
rect 4464 7028 4520 7030
rect 4568 7082 4624 7084
rect 4568 7030 4570 7082
rect 4570 7030 4622 7082
rect 4622 7030 4624 7082
rect 4568 7028 4624 7030
rect 4672 7082 4728 7084
rect 4672 7030 4674 7082
rect 4674 7030 4726 7082
rect 4726 7030 4728 7082
rect 4672 7028 4728 7030
rect 4464 5514 4520 5516
rect 4464 5462 4466 5514
rect 4466 5462 4518 5514
rect 4518 5462 4520 5514
rect 4464 5460 4520 5462
rect 4568 5514 4624 5516
rect 4568 5462 4570 5514
rect 4570 5462 4622 5514
rect 4622 5462 4624 5514
rect 4568 5460 4624 5462
rect 4672 5514 4728 5516
rect 4672 5462 4674 5514
rect 4674 5462 4726 5514
rect 4726 5462 4728 5514
rect 4672 5460 4728 5462
rect 4464 3946 4520 3948
rect 4464 3894 4466 3946
rect 4466 3894 4518 3946
rect 4518 3894 4520 3946
rect 4464 3892 4520 3894
rect 4568 3946 4624 3948
rect 4568 3894 4570 3946
rect 4570 3894 4622 3946
rect 4622 3894 4624 3946
rect 4568 3892 4624 3894
rect 4672 3946 4728 3948
rect 4672 3894 4674 3946
rect 4674 3894 4726 3946
rect 4726 3894 4728 3946
rect 4672 3892 4728 3894
rect 4464 2378 4520 2380
rect 4464 2326 4466 2378
rect 4466 2326 4518 2378
rect 4518 2326 4520 2378
rect 4464 2324 4520 2326
rect 4568 2378 4624 2380
rect 4568 2326 4570 2378
rect 4570 2326 4622 2378
rect 4622 2326 4624 2378
rect 4568 2324 4624 2326
rect 4672 2378 4728 2380
rect 4672 2326 4674 2378
rect 4674 2326 4726 2378
rect 4726 2326 4728 2378
rect 4672 2324 4728 2326
rect 4284 2044 4340 2100
rect 5516 11004 5572 11060
rect 5628 10892 5684 10948
rect 5628 9100 5684 9156
rect 5852 10780 5908 10836
rect 5180 5516 5236 5572
rect 5404 8428 5460 8484
rect 5068 3500 5124 3556
rect 5180 4956 5236 5012
rect 3804 1594 3860 1596
rect 3804 1542 3806 1594
rect 3806 1542 3858 1594
rect 3858 1542 3860 1594
rect 3804 1540 3860 1542
rect 3908 1594 3964 1596
rect 3908 1542 3910 1594
rect 3910 1542 3962 1594
rect 3962 1542 3964 1594
rect 3908 1540 3964 1542
rect 4012 1594 4068 1596
rect 4012 1542 4014 1594
rect 4014 1542 4066 1594
rect 4066 1542 4068 1594
rect 4956 1596 5012 1652
rect 5068 3276 5124 3332
rect 4012 1540 4068 1542
rect 2268 1372 2324 1428
rect 4172 1314 4228 1316
rect 4172 1262 4174 1314
rect 4174 1262 4226 1314
rect 4226 1262 4228 1314
rect 4172 1260 4228 1262
rect 5180 2940 5236 2996
rect 5292 4172 5348 4228
rect 6076 11900 6132 11956
rect 6188 11618 6244 11620
rect 6188 11566 6190 11618
rect 6190 11566 6242 11618
rect 6242 11566 6244 11618
rect 6188 11564 6244 11566
rect 6188 9660 6244 9716
rect 6188 7196 6244 7252
rect 6300 8764 6356 8820
rect 5740 5516 5796 5572
rect 5404 2716 5460 2772
rect 5628 3388 5684 3444
rect 5292 2156 5348 2212
rect 5068 1148 5124 1204
rect 1260 924 1316 980
rect 2156 252 2212 308
rect 4464 810 4520 812
rect 4464 758 4466 810
rect 4466 758 4518 810
rect 4518 758 4520 810
rect 4464 756 4520 758
rect 4568 810 4624 812
rect 4568 758 4570 810
rect 4570 758 4622 810
rect 4622 758 4624 810
rect 4568 756 4624 758
rect 4672 810 4728 812
rect 4672 758 4674 810
rect 4674 758 4726 810
rect 4726 758 4728 810
rect 4672 756 4728 758
rect 5740 3052 5796 3108
rect 5852 2828 5908 2884
rect 6188 5068 6244 5124
rect 6188 4844 6244 4900
rect 6076 4284 6132 4340
rect 6076 2380 6132 2436
rect 6412 8652 6468 8708
rect 7308 13692 7364 13748
rect 7420 13132 7476 13188
rect 7532 13356 7588 13412
rect 6748 11564 6804 11620
rect 6860 11900 6916 11956
rect 6412 4620 6468 4676
rect 6524 7980 6580 8036
rect 6972 11788 7028 11844
rect 7756 11618 7812 11620
rect 7756 11566 7758 11618
rect 7758 11566 7810 11618
rect 7810 11566 7812 11618
rect 7756 11564 7812 11566
rect 8204 13244 8260 13300
rect 7420 10610 7476 10612
rect 7420 10558 7422 10610
rect 7422 10558 7474 10610
rect 7474 10558 7476 10610
rect 7420 10556 7476 10558
rect 7532 8764 7588 8820
rect 7980 9772 8036 9828
rect 7756 8258 7812 8260
rect 7756 8206 7758 8258
rect 7758 8206 7810 8258
rect 7810 8206 7812 8258
rect 7756 8204 7812 8206
rect 6636 7868 6692 7924
rect 7868 7308 7924 7364
rect 6636 7084 6692 7140
rect 7308 6018 7364 6020
rect 7308 5966 7310 6018
rect 7310 5966 7362 6018
rect 7362 5966 7364 6018
rect 7308 5964 7364 5966
rect 6748 5906 6804 5908
rect 6748 5854 6750 5906
rect 6750 5854 6802 5906
rect 6802 5854 6804 5906
rect 6748 5852 6804 5854
rect 6636 4956 6692 5012
rect 6524 4508 6580 4564
rect 6300 4396 6356 4452
rect 7980 3836 8036 3892
rect 6188 1708 6244 1764
rect 6524 2604 6580 2660
rect 8204 12012 8260 12068
rect 8316 11788 8372 11844
rect 9660 13356 9716 13412
rect 10108 13244 10164 13300
rect 9772 13186 9828 13188
rect 9772 13134 9774 13186
rect 9774 13134 9826 13186
rect 9826 13134 9828 13186
rect 9772 13132 9828 13134
rect 10108 13020 10164 13076
rect 8764 11564 8820 11620
rect 8428 11116 8484 11172
rect 8988 10780 9044 10836
rect 8428 8316 8484 8372
rect 8652 8204 8708 8260
rect 8316 7308 8372 7364
rect 8204 6076 8260 6132
rect 8204 5852 8260 5908
rect 9212 10108 9268 10164
rect 10108 11788 10164 11844
rect 9324 7308 9380 7364
rect 9548 7308 9604 7364
rect 9660 8876 9716 8932
rect 9436 6636 9492 6692
rect 9884 10108 9940 10164
rect 10108 9660 10164 9716
rect 9772 8540 9828 8596
rect 9772 8316 9828 8372
rect 9884 6748 9940 6804
rect 9772 4172 9828 4228
rect 10108 8092 10164 8148
rect 10108 6300 10164 6356
rect 9100 3164 9156 3220
rect 9548 3388 9604 3444
rect 8092 1932 8148 1988
rect 9100 2828 9156 2884
rect 5964 700 6020 756
rect 5628 476 5684 532
rect 9548 1372 9604 1428
rect 9660 2940 9716 2996
rect 9100 1260 9156 1316
rect 8092 812 8148 868
rect 9772 1820 9828 1876
rect 9884 3052 9940 3108
rect 9660 812 9716 868
rect 9996 1596 10052 1652
rect 9884 588 9940 644
rect 9436 140 9492 196
rect 10444 9826 10500 9828
rect 10444 9774 10446 9826
rect 10446 9774 10498 9826
rect 10498 9774 10500 9826
rect 10444 9772 10500 9774
rect 10780 13804 10836 13860
rect 11340 13244 11396 13300
rect 11004 13020 11060 13076
rect 11788 13356 11844 13412
rect 11004 12236 11060 12292
rect 11900 13132 11956 13188
rect 12012 12402 12068 12404
rect 12012 12350 12014 12402
rect 12014 12350 12066 12402
rect 12066 12350 12068 12402
rect 12012 12348 12068 12350
rect 11788 12124 11844 12180
rect 12012 12124 12068 12180
rect 11228 11900 11284 11956
rect 10780 10556 10836 10612
rect 11116 10108 11172 10164
rect 10892 9324 10948 9380
rect 10332 7644 10388 7700
rect 10332 7420 10388 7476
rect 10444 6972 10500 7028
rect 10556 6748 10612 6804
rect 10892 6636 10948 6692
rect 12012 11788 12068 11844
rect 11228 6860 11284 6916
rect 11116 6690 11172 6692
rect 11116 6638 11118 6690
rect 11118 6638 11170 6690
rect 11170 6638 11172 6690
rect 11116 6636 11172 6638
rect 11900 10668 11956 10724
rect 11676 7308 11732 7364
rect 11788 9772 11844 9828
rect 10332 4172 10388 4228
rect 11452 7196 11508 7252
rect 10892 5852 10948 5908
rect 10892 5180 10948 5236
rect 12124 10498 12180 10500
rect 12124 10446 12126 10498
rect 12126 10446 12178 10498
rect 12178 10446 12180 10498
rect 12124 10444 12180 10446
rect 12124 10108 12180 10164
rect 12012 9660 12068 9716
rect 11900 9100 11956 9156
rect 12012 9436 12068 9492
rect 12572 13916 12628 13972
rect 12460 13580 12516 13636
rect 12460 11004 12516 11060
rect 12236 9548 12292 9604
rect 13244 13244 13300 13300
rect 13356 13132 13412 13188
rect 12796 12348 12852 12404
rect 14476 13356 14532 13412
rect 13244 11954 13300 11956
rect 13244 11902 13246 11954
rect 13246 11902 13298 11954
rect 13298 11902 13300 11954
rect 13244 11900 13300 11902
rect 12908 9436 12964 9492
rect 12572 9212 12628 9268
rect 12124 8204 12180 8260
rect 12684 8540 12740 8596
rect 12012 7420 12068 7476
rect 12236 7980 12292 8036
rect 12460 7532 12516 7588
rect 11788 6690 11844 6692
rect 11788 6638 11790 6690
rect 11790 6638 11842 6690
rect 11842 6638 11844 6690
rect 11788 6636 11844 6638
rect 12236 6748 12292 6804
rect 11676 5906 11732 5908
rect 11676 5854 11678 5906
rect 11678 5854 11730 5906
rect 11730 5854 11732 5906
rect 11676 5852 11732 5854
rect 10780 2380 10836 2436
rect 11564 5740 11620 5796
rect 11900 5234 11956 5236
rect 11900 5182 11902 5234
rect 11902 5182 11954 5234
rect 11954 5182 11956 5234
rect 11900 5180 11956 5182
rect 11900 5010 11956 5012
rect 11900 4958 11902 5010
rect 11902 4958 11954 5010
rect 11954 4958 11956 5010
rect 11900 4956 11956 4958
rect 12124 5180 12180 5236
rect 12236 5068 12292 5124
rect 12460 5964 12516 6020
rect 12572 7420 12628 7476
rect 12348 4956 12404 5012
rect 12460 5516 12516 5572
rect 12796 8034 12852 8036
rect 12796 7982 12798 8034
rect 12798 7982 12850 8034
rect 12850 7982 12852 8034
rect 12796 7980 12852 7982
rect 12684 6412 12740 6468
rect 12796 7644 12852 7700
rect 12572 4732 12628 4788
rect 12124 2604 12180 2660
rect 12348 2604 12404 2660
rect 12236 2044 12292 2100
rect 11564 1372 11620 1428
rect 10220 364 10276 420
rect 10108 140 10164 196
rect 11452 140 11508 196
rect 13244 11004 13300 11060
rect 13020 8540 13076 8596
rect 13132 10220 13188 10276
rect 13132 8316 13188 8372
rect 12908 5404 12964 5460
rect 13020 8204 13076 8260
rect 13132 7196 13188 7252
rect 13356 10108 13412 10164
rect 13356 8428 13412 8484
rect 14140 11452 14196 11508
rect 14364 12908 14420 12964
rect 13804 8876 13860 8932
rect 13692 8764 13748 8820
rect 13580 8258 13636 8260
rect 13580 8206 13582 8258
rect 13582 8206 13634 8258
rect 13634 8206 13636 8258
rect 13580 8204 13636 8206
rect 13468 7756 13524 7812
rect 13468 7250 13524 7252
rect 13468 7198 13470 7250
rect 13470 7198 13522 7250
rect 13522 7198 13524 7250
rect 13468 7196 13524 7198
rect 13244 5516 13300 5572
rect 13356 6076 13412 6132
rect 13468 5234 13524 5236
rect 13468 5182 13470 5234
rect 13470 5182 13522 5234
rect 13522 5182 13524 5234
rect 13468 5180 13524 5182
rect 13468 4620 13524 4676
rect 13804 8204 13860 8260
rect 13692 4620 13748 4676
rect 13356 3612 13412 3668
rect 13244 3276 13300 3332
rect 12908 2940 12964 2996
rect 12796 476 12852 532
rect 13804 1820 13860 1876
rect 14252 10498 14308 10500
rect 14252 10446 14254 10498
rect 14254 10446 14306 10498
rect 14306 10446 14308 10498
rect 14252 10444 14308 10446
rect 14812 14028 14868 14084
rect 15036 13132 15092 13188
rect 14924 13074 14980 13076
rect 14924 13022 14926 13074
rect 14926 13022 14978 13074
rect 14978 13022 14980 13074
rect 14924 13020 14980 13022
rect 14812 12402 14868 12404
rect 14812 12350 14814 12402
rect 14814 12350 14866 12402
rect 14866 12350 14868 12402
rect 14812 12348 14868 12350
rect 14588 11564 14644 11620
rect 14476 10444 14532 10500
rect 14476 10220 14532 10276
rect 14252 8540 14308 8596
rect 14028 6076 14084 6132
rect 14140 5122 14196 5124
rect 14140 5070 14142 5122
rect 14142 5070 14194 5122
rect 14194 5070 14196 5122
rect 14140 5068 14196 5070
rect 14476 8092 14532 8148
rect 14252 3500 14308 3556
rect 14700 4956 14756 5012
rect 15148 4508 15204 4564
rect 15932 12348 15988 12404
rect 16380 12402 16436 12404
rect 16380 12350 16382 12402
rect 16382 12350 16434 12402
rect 16434 12350 16436 12402
rect 16380 12348 16436 12350
rect 15708 10220 15764 10276
rect 15820 10108 15876 10164
rect 15372 8428 15428 8484
rect 15596 5516 15652 5572
rect 15260 3612 15316 3668
rect 15708 4956 15764 5012
rect 15820 4284 15876 4340
rect 15820 3836 15876 3892
rect 16716 13468 16772 13524
rect 16604 11900 16660 11956
rect 16828 13020 16884 13076
rect 17388 13186 17444 13188
rect 17388 13134 17390 13186
rect 17390 13134 17442 13186
rect 17442 13134 17444 13186
rect 17388 13132 17444 13134
rect 17276 12348 17332 12404
rect 16716 11564 16772 11620
rect 16940 11564 16996 11620
rect 17164 11788 17220 11844
rect 18620 13132 18676 13188
rect 18956 13186 19012 13188
rect 18956 13134 18958 13186
rect 18958 13134 19010 13186
rect 19010 13134 19012 13186
rect 18956 13132 19012 13134
rect 18284 12348 18340 12404
rect 18396 12178 18452 12180
rect 18396 12126 18398 12178
rect 18398 12126 18450 12178
rect 18450 12126 18452 12178
rect 18396 12124 18452 12126
rect 18284 11676 18340 11732
rect 17164 10444 17220 10500
rect 17388 10444 17444 10500
rect 19964 13132 20020 13188
rect 17948 10892 18004 10948
rect 18284 10722 18340 10724
rect 18284 10670 18286 10722
rect 18286 10670 18338 10722
rect 18338 10670 18340 10722
rect 18284 10668 18340 10670
rect 17948 10220 18004 10276
rect 18172 10220 18228 10276
rect 17836 9884 17892 9940
rect 17724 9772 17780 9828
rect 18284 9826 18340 9828
rect 18284 9774 18286 9826
rect 18286 9774 18338 9826
rect 18338 9774 18340 9826
rect 18284 9772 18340 9774
rect 16604 9436 16660 9492
rect 17948 9436 18004 9492
rect 18284 9324 18340 9380
rect 18060 9154 18116 9156
rect 18060 9102 18062 9154
rect 18062 9102 18114 9154
rect 18114 9102 18116 9154
rect 18060 9100 18116 9102
rect 17948 8988 18004 9044
rect 18284 8988 18340 9044
rect 16492 8764 16548 8820
rect 16156 8092 16212 8148
rect 16156 6860 16212 6916
rect 16044 3836 16100 3892
rect 16156 4956 16212 5012
rect 15708 3388 15764 3444
rect 14140 2828 14196 2884
rect 14924 1260 14980 1316
rect 13916 1036 13972 1092
rect 13804 252 13860 308
rect 11900 140 11956 196
rect 13468 140 13524 196
rect 14140 140 14196 196
rect 15484 140 15540 196
rect 15820 140 15876 196
rect 17500 8652 17556 8708
rect 17052 7756 17108 7812
rect 17052 6972 17108 7028
rect 17276 6972 17332 7028
rect 16828 6860 16884 6916
rect 16716 6300 16772 6356
rect 17388 6412 17444 6468
rect 16604 5292 16660 5348
rect 18844 9996 18900 10052
rect 20188 13580 20244 13636
rect 20076 11676 20132 11732
rect 20300 12124 20356 12180
rect 19516 11340 19572 11396
rect 19292 9324 19348 9380
rect 19404 10556 19460 10612
rect 19404 9212 19460 9268
rect 18620 9100 18676 9156
rect 17612 7308 17668 7364
rect 18284 7362 18340 7364
rect 18284 7310 18286 7362
rect 18286 7310 18338 7362
rect 18338 7310 18340 7362
rect 18284 7308 18340 7310
rect 18396 6748 18452 6804
rect 17612 6412 17668 6468
rect 17500 5964 17556 6020
rect 17388 4844 17444 4900
rect 16828 4620 16884 4676
rect 17948 3666 18004 3668
rect 17948 3614 17950 3666
rect 17950 3614 18002 3666
rect 18002 3614 18004 3666
rect 17948 3612 18004 3614
rect 18172 3500 18228 3556
rect 18732 7420 18788 7476
rect 18844 6748 18900 6804
rect 18620 6524 18676 6580
rect 18284 3388 18340 3444
rect 18172 2828 18228 2884
rect 17164 2604 17220 2660
rect 16828 2380 16884 2436
rect 16940 2492 16996 2548
rect 16828 1708 16884 1764
rect 16492 1596 16548 1652
rect 16716 1596 16772 1652
rect 16716 476 16772 532
rect 17052 1708 17108 1764
rect 17052 1372 17108 1428
rect 16940 1148 16996 1204
rect 17164 812 17220 868
rect 16828 364 16884 420
rect 17500 140 17556 196
rect 19740 7362 19796 7364
rect 19740 7310 19742 7362
rect 19742 7310 19794 7362
rect 19794 7310 19796 7362
rect 19740 7308 19796 7310
rect 20188 11228 20244 11284
rect 20076 10108 20132 10164
rect 19964 8764 20020 8820
rect 19852 6524 19908 6580
rect 20636 13692 20692 13748
rect 20524 12962 20580 12964
rect 20524 12910 20526 12962
rect 20526 12910 20578 12962
rect 20578 12910 20580 12962
rect 20524 12908 20580 12910
rect 20300 10332 20356 10388
rect 20188 9772 20244 9828
rect 20300 9660 20356 9716
rect 20300 8204 20356 8260
rect 20524 9660 20580 9716
rect 20748 13244 20804 13300
rect 20860 12460 20916 12516
rect 20860 12290 20916 12292
rect 20860 12238 20862 12290
rect 20862 12238 20914 12290
rect 20914 12238 20916 12290
rect 20860 12236 20916 12238
rect 34524 14140 34580 14196
rect 21196 13244 21252 13300
rect 21308 12684 21364 12740
rect 21420 13804 21476 13860
rect 21980 12684 22036 12740
rect 21308 12348 21364 12404
rect 21420 12178 21476 12180
rect 21420 12126 21422 12178
rect 21422 12126 21474 12178
rect 21474 12126 21476 12178
rect 21420 12124 21476 12126
rect 21196 11394 21252 11396
rect 21196 11342 21198 11394
rect 21198 11342 21250 11394
rect 21250 11342 21252 11394
rect 21196 11340 21252 11342
rect 20748 9772 20804 9828
rect 21084 10498 21140 10500
rect 21084 10446 21086 10498
rect 21086 10446 21138 10498
rect 21138 10446 21140 10498
rect 21084 10444 21140 10446
rect 21084 10220 21140 10276
rect 20860 9100 20916 9156
rect 20412 7980 20468 8036
rect 20636 7980 20692 8036
rect 19180 6300 19236 6356
rect 19068 3724 19124 3780
rect 19180 3836 19236 3892
rect 19628 3778 19684 3780
rect 19628 3726 19630 3778
rect 19630 3726 19682 3778
rect 19682 3726 19684 3778
rect 19628 3724 19684 3726
rect 20524 5852 20580 5908
rect 20300 5740 20356 5796
rect 20188 4508 20244 4564
rect 19852 2604 19908 2660
rect 20076 3500 20132 3556
rect 20076 2492 20132 2548
rect 18620 140 18676 196
rect 20412 5180 20468 5236
rect 20412 1372 20468 1428
rect 21308 9042 21364 9044
rect 21308 8990 21310 9042
rect 21310 8990 21362 9042
rect 21362 8990 21364 9042
rect 21308 8988 21364 8990
rect 21196 7868 21252 7924
rect 21308 8092 21364 8148
rect 21308 7308 21364 7364
rect 21196 7196 21252 7252
rect 20636 2940 20692 2996
rect 20748 6524 20804 6580
rect 21196 6412 21252 6468
rect 21644 12572 21700 12628
rect 21868 12460 21924 12516
rect 21980 10556 22036 10612
rect 22876 13356 22932 13412
rect 22428 13020 22484 13076
rect 22204 12012 22260 12068
rect 22204 11004 22260 11060
rect 22092 9996 22148 10052
rect 21644 8988 21700 9044
rect 21756 9212 21812 9268
rect 21532 8428 21588 8484
rect 21980 8818 22036 8820
rect 21980 8766 21982 8818
rect 21982 8766 22034 8818
rect 22034 8766 22036 8818
rect 21980 8764 22036 8766
rect 21756 8092 21812 8148
rect 22204 8316 22260 8372
rect 21644 7868 21700 7924
rect 21644 7308 21700 7364
rect 21980 7308 22036 7364
rect 21644 7084 21700 7140
rect 21532 5404 21588 5460
rect 21868 5122 21924 5124
rect 21868 5070 21870 5122
rect 21870 5070 21922 5122
rect 21922 5070 21924 5122
rect 21868 5068 21924 5070
rect 20972 4396 21028 4452
rect 21532 4620 21588 4676
rect 20972 4172 21028 4228
rect 21196 4172 21252 4228
rect 21196 3500 21252 3556
rect 20748 2716 20804 2772
rect 21756 3948 21812 4004
rect 22316 8204 22372 8260
rect 22652 12460 22708 12516
rect 22428 6636 22484 6692
rect 22540 10444 22596 10500
rect 22428 5964 22484 6020
rect 22764 10444 22820 10500
rect 22652 9660 22708 9716
rect 22764 8652 22820 8708
rect 22764 8316 22820 8372
rect 23212 13356 23268 13412
rect 22988 12908 23044 12964
rect 23772 14028 23828 14084
rect 23548 13132 23604 13188
rect 23660 13692 23716 13748
rect 23212 12460 23268 12516
rect 23436 12460 23492 12516
rect 23100 11340 23156 11396
rect 22988 10332 23044 10388
rect 22988 9996 23044 10052
rect 23548 11788 23604 11844
rect 23996 13020 24052 13076
rect 24464 13354 24520 13356
rect 24464 13302 24466 13354
rect 24466 13302 24518 13354
rect 24518 13302 24520 13354
rect 24464 13300 24520 13302
rect 24568 13354 24624 13356
rect 24568 13302 24570 13354
rect 24570 13302 24622 13354
rect 24622 13302 24624 13354
rect 24568 13300 24624 13302
rect 24672 13354 24728 13356
rect 24672 13302 24674 13354
rect 24674 13302 24726 13354
rect 24726 13302 24728 13354
rect 24672 13300 24728 13302
rect 23772 12796 23828 12852
rect 24780 13020 24836 13076
rect 23804 12570 23860 12572
rect 23804 12518 23806 12570
rect 23806 12518 23858 12570
rect 23858 12518 23860 12570
rect 23804 12516 23860 12518
rect 23908 12570 23964 12572
rect 23908 12518 23910 12570
rect 23910 12518 23962 12570
rect 23962 12518 23964 12570
rect 23908 12516 23964 12518
rect 24012 12570 24068 12572
rect 24012 12518 24014 12570
rect 24014 12518 24066 12570
rect 24066 12518 24068 12570
rect 24012 12516 24068 12518
rect 24668 12572 24724 12628
rect 24464 11786 24520 11788
rect 24464 11734 24466 11786
rect 24466 11734 24518 11786
rect 24518 11734 24520 11786
rect 24464 11732 24520 11734
rect 24568 11786 24624 11788
rect 24568 11734 24570 11786
rect 24570 11734 24622 11786
rect 24622 11734 24624 11786
rect 24568 11732 24624 11734
rect 24672 11786 24728 11788
rect 24672 11734 24674 11786
rect 24674 11734 24726 11786
rect 24726 11734 24728 11786
rect 24672 11732 24728 11734
rect 23996 11282 24052 11284
rect 23996 11230 23998 11282
rect 23998 11230 24050 11282
rect 24050 11230 24052 11282
rect 23996 11228 24052 11230
rect 24444 11116 24500 11172
rect 23804 11002 23860 11004
rect 23804 10950 23806 11002
rect 23806 10950 23858 11002
rect 23858 10950 23860 11002
rect 23804 10948 23860 10950
rect 23908 11002 23964 11004
rect 23908 10950 23910 11002
rect 23910 10950 23962 11002
rect 23962 10950 23964 11002
rect 23908 10948 23964 10950
rect 24012 11002 24068 11004
rect 24012 10950 24014 11002
rect 24014 10950 24066 11002
rect 24066 10950 24068 11002
rect 24012 10948 24068 10950
rect 23212 10220 23268 10276
rect 23324 10108 23380 10164
rect 23436 10220 23492 10276
rect 23100 9660 23156 9716
rect 23212 9996 23268 10052
rect 23996 10050 24052 10052
rect 23996 9998 23998 10050
rect 23998 9998 24050 10050
rect 24050 9998 24052 10050
rect 23996 9996 24052 9998
rect 23100 8764 23156 8820
rect 22652 6300 22708 6356
rect 22988 6300 23044 6356
rect 22092 5628 22148 5684
rect 22092 4284 22148 4340
rect 21980 3500 22036 3556
rect 22316 5122 22372 5124
rect 22316 5070 22318 5122
rect 22318 5070 22370 5122
rect 22370 5070 22372 5122
rect 22316 5068 22372 5070
rect 22652 5740 22708 5796
rect 22540 5068 22596 5124
rect 22540 4732 22596 4788
rect 21868 3276 21924 3332
rect 21532 2604 21588 2660
rect 21756 2380 21812 2436
rect 21644 1820 21700 1876
rect 21644 1596 21700 1652
rect 20524 476 20580 532
rect 21532 1148 21588 1204
rect 20300 28 20356 84
rect 22428 4284 22484 4340
rect 21980 2940 22036 2996
rect 21868 1260 21924 1316
rect 22540 2380 22596 2436
rect 22652 3388 22708 3444
rect 22428 1932 22484 1988
rect 22092 1260 22148 1316
rect 22764 2492 22820 2548
rect 22876 3388 22932 3444
rect 22876 924 22932 980
rect 22652 812 22708 868
rect 23548 9772 23604 9828
rect 24220 10220 24276 10276
rect 24892 10444 24948 10500
rect 24464 10218 24520 10220
rect 24332 10108 24388 10164
rect 24464 10166 24466 10218
rect 24466 10166 24518 10218
rect 24518 10166 24520 10218
rect 24464 10164 24520 10166
rect 24568 10218 24624 10220
rect 24568 10166 24570 10218
rect 24570 10166 24622 10218
rect 24622 10166 24624 10218
rect 24568 10164 24624 10166
rect 24672 10218 24728 10220
rect 24672 10166 24674 10218
rect 24674 10166 24726 10218
rect 24726 10166 24728 10218
rect 24672 10164 24728 10166
rect 24556 9884 24612 9940
rect 23548 9324 23604 9380
rect 23804 9434 23860 9436
rect 23804 9382 23806 9434
rect 23806 9382 23858 9434
rect 23858 9382 23860 9434
rect 23804 9380 23860 9382
rect 23908 9434 23964 9436
rect 23908 9382 23910 9434
rect 23910 9382 23962 9434
rect 23962 9382 23964 9434
rect 23908 9380 23964 9382
rect 24012 9434 24068 9436
rect 24012 9382 24014 9434
rect 24014 9382 24066 9434
rect 24066 9382 24068 9434
rect 24012 9380 24068 9382
rect 24220 9436 24276 9492
rect 24108 9042 24164 9044
rect 24108 8990 24110 9042
rect 24110 8990 24162 9042
rect 24162 8990 24164 9042
rect 24108 8988 24164 8990
rect 24444 9212 24500 9268
rect 24332 8540 24388 8596
rect 24464 8650 24520 8652
rect 24464 8598 24466 8650
rect 24466 8598 24518 8650
rect 24518 8598 24520 8650
rect 24464 8596 24520 8598
rect 24568 8650 24624 8652
rect 24568 8598 24570 8650
rect 24570 8598 24622 8650
rect 24622 8598 24624 8650
rect 24568 8596 24624 8598
rect 24672 8650 24728 8652
rect 24672 8598 24674 8650
rect 24674 8598 24726 8650
rect 24726 8598 24728 8650
rect 24672 8596 24728 8598
rect 25116 12236 25172 12292
rect 25340 11954 25396 11956
rect 25340 11902 25342 11954
rect 25342 11902 25394 11954
rect 25394 11902 25396 11954
rect 25340 11900 25396 11902
rect 25228 10108 25284 10164
rect 25228 9548 25284 9604
rect 25564 12348 25620 12404
rect 25564 11900 25620 11956
rect 26012 13804 26068 13860
rect 25900 11788 25956 11844
rect 26236 13580 26292 13636
rect 26908 14028 26964 14084
rect 26796 13132 26852 13188
rect 26012 11564 26068 11620
rect 25452 9212 25508 9268
rect 25564 9884 25620 9940
rect 25564 8988 25620 9044
rect 25228 8876 25284 8932
rect 25228 8316 25284 8372
rect 24220 8204 24276 8260
rect 24780 7980 24836 8036
rect 23660 7756 23716 7812
rect 23804 7866 23860 7868
rect 23804 7814 23806 7866
rect 23806 7814 23858 7866
rect 23858 7814 23860 7866
rect 23804 7812 23860 7814
rect 23908 7866 23964 7868
rect 23908 7814 23910 7866
rect 23910 7814 23962 7866
rect 23962 7814 23964 7866
rect 23908 7812 23964 7814
rect 24012 7866 24068 7868
rect 24012 7814 24014 7866
rect 24014 7814 24066 7866
rect 24066 7814 24068 7866
rect 24012 7812 24068 7814
rect 24220 7084 24276 7140
rect 24444 7644 24500 7700
rect 23548 6636 23604 6692
rect 23548 6188 23604 6244
rect 23212 5516 23268 5572
rect 24108 6860 24164 6916
rect 25228 7644 25284 7700
rect 24464 7082 24520 7084
rect 24464 7030 24466 7082
rect 24466 7030 24518 7082
rect 24518 7030 24520 7082
rect 24464 7028 24520 7030
rect 24568 7082 24624 7084
rect 24568 7030 24570 7082
rect 24570 7030 24622 7082
rect 24622 7030 24624 7082
rect 24568 7028 24624 7030
rect 24672 7082 24728 7084
rect 24672 7030 24674 7082
rect 24674 7030 24726 7082
rect 24726 7030 24728 7082
rect 24672 7028 24728 7030
rect 24332 6636 24388 6692
rect 24780 6690 24836 6692
rect 24780 6638 24782 6690
rect 24782 6638 24834 6690
rect 24834 6638 24836 6690
rect 24780 6636 24836 6638
rect 23804 6298 23860 6300
rect 23804 6246 23806 6298
rect 23806 6246 23858 6298
rect 23858 6246 23860 6298
rect 23804 6244 23860 6246
rect 23908 6298 23964 6300
rect 23908 6246 23910 6298
rect 23910 6246 23962 6298
rect 23962 6246 23964 6298
rect 23908 6244 23964 6246
rect 24012 6298 24068 6300
rect 24012 6246 24014 6298
rect 24014 6246 24066 6298
rect 24066 6246 24068 6298
rect 24220 6300 24276 6356
rect 24012 6244 24068 6246
rect 24668 5682 24724 5684
rect 24668 5630 24670 5682
rect 24670 5630 24722 5682
rect 24722 5630 24724 5682
rect 24668 5628 24724 5630
rect 24464 5514 24520 5516
rect 24332 5404 24388 5460
rect 24464 5462 24466 5514
rect 24466 5462 24518 5514
rect 24518 5462 24520 5514
rect 24464 5460 24520 5462
rect 24568 5514 24624 5516
rect 24568 5462 24570 5514
rect 24570 5462 24622 5514
rect 24622 5462 24624 5514
rect 24568 5460 24624 5462
rect 24672 5514 24728 5516
rect 24672 5462 24674 5514
rect 24674 5462 24726 5514
rect 24726 5462 24728 5514
rect 24672 5460 24728 5462
rect 23804 4730 23860 4732
rect 23804 4678 23806 4730
rect 23806 4678 23858 4730
rect 23858 4678 23860 4730
rect 23804 4676 23860 4678
rect 23908 4730 23964 4732
rect 23908 4678 23910 4730
rect 23910 4678 23962 4730
rect 23962 4678 23964 4730
rect 23908 4676 23964 4678
rect 24012 4730 24068 4732
rect 24012 4678 24014 4730
rect 24014 4678 24066 4730
rect 24066 4678 24068 4730
rect 24012 4676 24068 4678
rect 24332 4620 24388 4676
rect 23660 4284 23716 4340
rect 25116 5852 25172 5908
rect 25340 7196 25396 7252
rect 25340 6860 25396 6916
rect 25676 7196 25732 7252
rect 25788 9436 25844 9492
rect 25788 6636 25844 6692
rect 25900 8988 25956 9044
rect 25452 6300 25508 6356
rect 25004 5628 25060 5684
rect 25116 4172 25172 4228
rect 25228 5404 25284 5460
rect 24464 3946 24520 3948
rect 24464 3894 24466 3946
rect 24466 3894 24518 3946
rect 24518 3894 24520 3946
rect 24464 3892 24520 3894
rect 24568 3946 24624 3948
rect 24568 3894 24570 3946
rect 24570 3894 24622 3946
rect 24622 3894 24624 3946
rect 24568 3892 24624 3894
rect 24672 3946 24728 3948
rect 24672 3894 24674 3946
rect 24674 3894 24726 3946
rect 24726 3894 24728 3946
rect 24892 3948 24948 4004
rect 24672 3892 24728 3894
rect 23100 3164 23156 3220
rect 23324 3500 23380 3556
rect 23212 2940 23268 2996
rect 23804 3162 23860 3164
rect 23804 3110 23806 3162
rect 23806 3110 23858 3162
rect 23858 3110 23860 3162
rect 23804 3108 23860 3110
rect 23908 3162 23964 3164
rect 23908 3110 23910 3162
rect 23910 3110 23962 3162
rect 23962 3110 23964 3162
rect 23908 3108 23964 3110
rect 24012 3162 24068 3164
rect 24012 3110 24014 3162
rect 24014 3110 24066 3162
rect 24066 3110 24068 3162
rect 24332 3164 24388 3220
rect 24012 3108 24068 3110
rect 24220 3052 24276 3108
rect 23436 2828 23492 2884
rect 23436 2492 23492 2548
rect 23996 2828 24052 2884
rect 25340 4508 25396 4564
rect 25340 3724 25396 3780
rect 25452 3948 25508 4004
rect 25228 3052 25284 3108
rect 25452 3052 25508 3108
rect 24332 2380 24388 2436
rect 24464 2378 24520 2380
rect 24464 2326 24466 2378
rect 24466 2326 24518 2378
rect 24518 2326 24520 2378
rect 24464 2324 24520 2326
rect 24568 2378 24624 2380
rect 24568 2326 24570 2378
rect 24570 2326 24622 2378
rect 24622 2326 24624 2378
rect 24568 2324 24624 2326
rect 24672 2378 24728 2380
rect 24672 2326 24674 2378
rect 24674 2326 24726 2378
rect 24726 2326 24728 2378
rect 24672 2324 24728 2326
rect 24108 2156 24164 2212
rect 23548 1986 23604 1988
rect 23548 1934 23550 1986
rect 23550 1934 23602 1986
rect 23602 1934 23604 1986
rect 23548 1932 23604 1934
rect 25676 2658 25732 2660
rect 25676 2606 25678 2658
rect 25678 2606 25730 2658
rect 25730 2606 25732 2658
rect 25676 2604 25732 2606
rect 25564 2492 25620 2548
rect 25116 1932 25172 1988
rect 23324 1708 23380 1764
rect 23804 1594 23860 1596
rect 23804 1542 23806 1594
rect 23806 1542 23858 1594
rect 23858 1542 23860 1594
rect 23804 1540 23860 1542
rect 23908 1594 23964 1596
rect 23908 1542 23910 1594
rect 23910 1542 23962 1594
rect 23962 1542 23964 1594
rect 23908 1540 23964 1542
rect 24012 1594 24068 1596
rect 24012 1542 24014 1594
rect 24014 1542 24066 1594
rect 24066 1542 24068 1594
rect 24012 1540 24068 1542
rect 24332 1596 24388 1652
rect 23212 924 23268 980
rect 23548 1372 23604 1428
rect 22988 252 23044 308
rect 24332 812 24388 868
rect 24464 810 24520 812
rect 24464 758 24466 810
rect 24466 758 24518 810
rect 24518 758 24520 810
rect 24464 756 24520 758
rect 24568 810 24624 812
rect 24568 758 24570 810
rect 24570 758 24622 810
rect 24622 758 24624 810
rect 24568 756 24624 758
rect 24672 810 24728 812
rect 24672 758 24674 810
rect 24674 758 24726 810
rect 24726 758 24728 810
rect 24672 756 24728 758
rect 26684 11564 26740 11620
rect 26124 9996 26180 10052
rect 26012 6188 26068 6244
rect 26124 9772 26180 9828
rect 26012 4732 26068 4788
rect 26012 3276 26068 3332
rect 27468 13356 27524 13412
rect 26908 11340 26964 11396
rect 27020 12796 27076 12852
rect 26796 10220 26852 10276
rect 26908 10892 26964 10948
rect 26908 9996 26964 10052
rect 27132 10332 27188 10388
rect 26236 8092 26292 8148
rect 26348 8876 26404 8932
rect 26908 8764 26964 8820
rect 26348 7308 26404 7364
rect 28028 13468 28084 13524
rect 27916 13020 27972 13076
rect 27580 11618 27636 11620
rect 27580 11566 27582 11618
rect 27582 11566 27634 11618
rect 27634 11566 27636 11618
rect 27580 11564 27636 11566
rect 28252 12908 28308 12964
rect 27468 10556 27524 10612
rect 28028 11004 28084 11060
rect 27244 9996 27300 10052
rect 27244 9436 27300 9492
rect 27692 10668 27748 10724
rect 27132 8764 27188 8820
rect 27132 7756 27188 7812
rect 26460 7196 26516 7252
rect 26348 6690 26404 6692
rect 26348 6638 26350 6690
rect 26350 6638 26402 6690
rect 26402 6638 26404 6690
rect 26348 6636 26404 6638
rect 26236 6524 26292 6580
rect 26460 6300 26516 6356
rect 26348 6188 26404 6244
rect 27020 6524 27076 6580
rect 26796 5740 26852 5796
rect 26348 4620 26404 4676
rect 26572 5180 26628 5236
rect 26572 4620 26628 4676
rect 27580 9938 27636 9940
rect 27580 9886 27582 9938
rect 27582 9886 27634 9938
rect 27634 9886 27636 9938
rect 27580 9884 27636 9886
rect 27468 8652 27524 8708
rect 28140 10220 28196 10276
rect 28924 13916 28980 13972
rect 28812 13692 28868 13748
rect 28700 13580 28756 13636
rect 28476 12124 28532 12180
rect 28588 13468 28644 13524
rect 28588 11452 28644 11508
rect 28700 12348 28756 12404
rect 28364 11004 28420 11060
rect 28588 10668 28644 10724
rect 28476 10332 28532 10388
rect 29036 13132 29092 13188
rect 28812 11564 28868 11620
rect 28924 12348 28980 12404
rect 28700 10332 28756 10388
rect 28252 10108 28308 10164
rect 27692 8652 27748 8708
rect 27916 9436 27972 9492
rect 28252 9212 28308 9268
rect 28028 8370 28084 8372
rect 28028 8318 28030 8370
rect 28030 8318 28082 8370
rect 28082 8318 28084 8370
rect 28028 8316 28084 8318
rect 27244 5404 27300 5460
rect 27692 6636 27748 6692
rect 26684 4284 26740 4340
rect 26796 5180 26852 5236
rect 27580 4338 27636 4340
rect 27580 4286 27582 4338
rect 27582 4286 27634 4338
rect 27634 4286 27636 4338
rect 27580 4284 27636 4286
rect 27356 4060 27412 4116
rect 27468 3276 27524 3332
rect 27580 3164 27636 3220
rect 26796 2268 26852 2324
rect 26348 1484 26404 1540
rect 25900 1372 25956 1428
rect 26796 1148 26852 1204
rect 26124 1090 26180 1092
rect 26124 1038 26126 1090
rect 26126 1038 26178 1090
rect 26178 1038 26180 1090
rect 26124 1036 26180 1038
rect 27804 5794 27860 5796
rect 27804 5742 27806 5794
rect 27806 5742 27858 5794
rect 27858 5742 27860 5794
rect 27804 5740 27860 5742
rect 28028 3612 28084 3668
rect 27692 2716 27748 2772
rect 28140 3052 28196 3108
rect 28812 9548 28868 9604
rect 28700 8316 28756 8372
rect 28700 7980 28756 8036
rect 28476 7308 28532 7364
rect 28476 6188 28532 6244
rect 28364 5516 28420 5572
rect 29148 12850 29204 12852
rect 29148 12798 29150 12850
rect 29150 12798 29202 12850
rect 29202 12798 29204 12850
rect 29148 12796 29204 12798
rect 29372 12124 29428 12180
rect 29484 12796 29540 12852
rect 29036 11564 29092 11620
rect 28924 8988 28980 9044
rect 29036 11340 29092 11396
rect 28924 8540 28980 8596
rect 30716 13132 30772 13188
rect 30828 13244 30884 13300
rect 30604 12012 30660 12068
rect 30716 12236 30772 12292
rect 30044 11900 30100 11956
rect 29484 10668 29540 10724
rect 29820 10668 29876 10724
rect 29148 10556 29204 10612
rect 29820 9436 29876 9492
rect 29708 8652 29764 8708
rect 28924 7644 28980 7700
rect 29484 8258 29540 8260
rect 29484 8206 29486 8258
rect 29486 8206 29538 8258
rect 29538 8206 29540 8258
rect 29484 8204 29540 8206
rect 29036 7420 29092 7476
rect 28924 7308 28980 7364
rect 29596 7420 29652 7476
rect 29148 6636 29204 6692
rect 29260 7196 29316 7252
rect 28812 6412 28868 6468
rect 29036 6412 29092 6468
rect 29036 5740 29092 5796
rect 29260 5740 29316 5796
rect 28700 5404 28756 5460
rect 28588 4114 28644 4116
rect 28588 4062 28590 4114
rect 28590 4062 28642 4114
rect 28642 4062 28644 4114
rect 28588 4060 28644 4062
rect 29036 4172 29092 4228
rect 28812 3442 28868 3444
rect 28812 3390 28814 3442
rect 28814 3390 28866 3442
rect 28866 3390 28868 3442
rect 28812 3388 28868 3390
rect 28588 3276 28644 3332
rect 28924 2940 28980 2996
rect 28476 2492 28532 2548
rect 28812 2492 28868 2548
rect 28252 1596 28308 1652
rect 30156 10108 30212 10164
rect 30604 9714 30660 9716
rect 30604 9662 30606 9714
rect 30606 9662 30658 9714
rect 30658 9662 30660 9714
rect 30604 9660 30660 9662
rect 30268 9436 30324 9492
rect 30828 10668 30884 10724
rect 30940 12684 30996 12740
rect 30828 10332 30884 10388
rect 30828 8988 30884 9044
rect 30716 8876 30772 8932
rect 30940 8540 30996 8596
rect 30044 8092 30100 8148
rect 29708 7084 29764 7140
rect 30156 6972 30212 7028
rect 29820 6636 29876 6692
rect 29596 3724 29652 3780
rect 29708 5180 29764 5236
rect 29036 1260 29092 1316
rect 29148 3388 29204 3444
rect 30156 6076 30212 6132
rect 30380 6300 30436 6356
rect 30156 5516 30212 5572
rect 29932 4508 29988 4564
rect 29820 3500 29876 3556
rect 28476 588 28532 644
rect 29260 2770 29316 2772
rect 29260 2718 29262 2770
rect 29262 2718 29314 2770
rect 29314 2718 29316 2770
rect 29260 2716 29316 2718
rect 29820 2770 29876 2772
rect 29820 2718 29822 2770
rect 29822 2718 29874 2770
rect 29874 2718 29876 2770
rect 29820 2716 29876 2718
rect 30156 4508 30212 4564
rect 30828 6748 30884 6804
rect 30604 6300 30660 6356
rect 30492 5628 30548 5684
rect 30492 5292 30548 5348
rect 30380 5180 30436 5236
rect 30492 4620 30548 4676
rect 30268 3500 30324 3556
rect 30380 4060 30436 4116
rect 30156 3164 30212 3220
rect 30044 3052 30100 3108
rect 30156 2716 30212 2772
rect 30268 2604 30324 2660
rect 29596 2098 29652 2100
rect 29596 2046 29598 2098
rect 29598 2046 29650 2098
rect 29650 2046 29652 2098
rect 29596 2044 29652 2046
rect 30604 3836 30660 3892
rect 30604 3164 30660 3220
rect 31500 13186 31556 13188
rect 31500 13134 31502 13186
rect 31502 13134 31554 13186
rect 31554 13134 31556 13186
rect 31500 13132 31556 13134
rect 31612 13020 31668 13076
rect 31724 13132 31780 13188
rect 31500 12348 31556 12404
rect 31164 12012 31220 12068
rect 31948 12460 32004 12516
rect 31948 11676 32004 11732
rect 32284 12178 32340 12180
rect 32284 12126 32286 12178
rect 32286 12126 32338 12178
rect 32338 12126 32340 12178
rect 32284 12124 32340 12126
rect 32732 13804 32788 13860
rect 32508 12124 32564 12180
rect 32620 12236 32676 12292
rect 32396 12012 32452 12068
rect 31724 11452 31780 11508
rect 31276 11394 31332 11396
rect 31276 11342 31278 11394
rect 31278 11342 31330 11394
rect 31330 11342 31332 11394
rect 31276 11340 31332 11342
rect 31500 11340 31556 11396
rect 31836 11282 31892 11284
rect 31836 11230 31838 11282
rect 31838 11230 31890 11282
rect 31890 11230 31892 11282
rect 31836 11228 31892 11230
rect 31500 10780 31556 10836
rect 32956 13132 33012 13188
rect 33292 13074 33348 13076
rect 33292 13022 33294 13074
rect 33294 13022 33346 13074
rect 33346 13022 33348 13074
rect 33292 13020 33348 13022
rect 32956 12236 33012 12292
rect 33180 12178 33236 12180
rect 33180 12126 33182 12178
rect 33182 12126 33234 12178
rect 33234 12126 33236 12178
rect 33180 12124 33236 12126
rect 33740 13804 33796 13860
rect 33628 13356 33684 13412
rect 33404 12124 33460 12180
rect 33516 12796 33572 12852
rect 32732 11004 32788 11060
rect 32620 10668 32676 10724
rect 32396 10444 32452 10500
rect 31276 8428 31332 8484
rect 32060 8764 32116 8820
rect 32060 7868 32116 7924
rect 32172 8540 32228 8596
rect 31724 7756 31780 7812
rect 31164 7196 31220 7252
rect 31612 6748 31668 6804
rect 31276 6690 31332 6692
rect 31276 6638 31278 6690
rect 31278 6638 31330 6690
rect 31330 6638 31332 6690
rect 31276 6636 31332 6638
rect 31164 5404 31220 5460
rect 31500 5404 31556 5460
rect 31052 2940 31108 2996
rect 30604 2492 30660 2548
rect 30940 2492 30996 2548
rect 30492 2268 30548 2324
rect 30940 1596 30996 1652
rect 31164 1932 31220 1988
rect 30268 1484 30324 1540
rect 31164 1148 31220 1204
rect 31388 1932 31444 1988
rect 31388 476 31444 532
rect 29148 364 29204 420
rect 29596 140 29652 196
rect 31836 6076 31892 6132
rect 31948 6188 32004 6244
rect 32060 5794 32116 5796
rect 32060 5742 32062 5794
rect 32062 5742 32114 5794
rect 32114 5742 32116 5794
rect 32060 5740 32116 5742
rect 32060 5292 32116 5348
rect 32620 8988 32676 9044
rect 32508 8930 32564 8932
rect 32508 8878 32510 8930
rect 32510 8878 32562 8930
rect 32562 8878 32564 8930
rect 32508 8876 32564 8878
rect 32396 8092 32452 8148
rect 32620 6748 32676 6804
rect 32620 6130 32676 6132
rect 32620 6078 32622 6130
rect 32622 6078 32674 6130
rect 32674 6078 32676 6130
rect 32620 6076 32676 6078
rect 32172 5068 32228 5124
rect 32060 4732 32116 4788
rect 32284 4956 32340 5012
rect 32060 4396 32116 4452
rect 32060 3052 32116 3108
rect 32956 7756 33012 7812
rect 33516 11564 33572 11620
rect 33516 11116 33572 11172
rect 33180 10108 33236 10164
rect 33292 9884 33348 9940
rect 33516 9548 33572 9604
rect 33852 13580 33908 13636
rect 34188 13186 34244 13188
rect 34188 13134 34190 13186
rect 34190 13134 34242 13186
rect 34242 13134 34244 13186
rect 34188 13132 34244 13134
rect 34188 12348 34244 12404
rect 34076 12178 34132 12180
rect 34076 12126 34078 12178
rect 34078 12126 34130 12178
rect 34130 12126 34132 12178
rect 34076 12124 34132 12126
rect 33404 8988 33460 9044
rect 33964 11900 34020 11956
rect 35196 13468 35252 13524
rect 35308 13580 35364 13636
rect 34748 13132 34804 13188
rect 35644 13580 35700 13636
rect 35868 13020 35924 13076
rect 34300 12124 34356 12180
rect 34412 12012 34468 12068
rect 33180 8764 33236 8820
rect 33516 8876 33572 8932
rect 33516 8428 33572 8484
rect 33628 8764 33684 8820
rect 33852 8818 33908 8820
rect 33852 8766 33854 8818
rect 33854 8766 33906 8818
rect 33906 8766 33908 8818
rect 33852 8764 33908 8766
rect 34188 10220 34244 10276
rect 34076 9884 34132 9940
rect 34188 9324 34244 9380
rect 34076 8764 34132 8820
rect 33964 7196 34020 7252
rect 33852 6972 33908 7028
rect 33404 6748 33460 6804
rect 33180 5794 33236 5796
rect 33180 5742 33182 5794
rect 33182 5742 33234 5794
rect 33234 5742 33236 5794
rect 33180 5740 33236 5742
rect 33068 3164 33124 3220
rect 32844 2716 32900 2772
rect 33068 2658 33124 2660
rect 33068 2606 33070 2658
rect 33070 2606 33122 2658
rect 33122 2606 33124 2658
rect 33068 2604 33124 2606
rect 32508 2546 32564 2548
rect 32508 2494 32510 2546
rect 32510 2494 32562 2546
rect 32562 2494 32564 2546
rect 32508 2492 32564 2494
rect 32284 2380 32340 2436
rect 32284 1708 32340 1764
rect 32060 1484 32116 1540
rect 31724 1372 31780 1428
rect 31948 700 32004 756
rect 31948 140 32004 196
rect 21756 28 21812 84
rect 33628 6188 33684 6244
rect 34524 11452 34580 11508
rect 34972 12178 35028 12180
rect 34972 12126 34974 12178
rect 34974 12126 35026 12178
rect 35026 12126 35028 12178
rect 34972 12124 35028 12126
rect 34412 10220 34468 10276
rect 34972 11788 35028 11844
rect 34748 10220 34804 10276
rect 34300 7420 34356 7476
rect 34412 3948 34468 4004
rect 34524 4060 34580 4116
rect 34524 2268 34580 2324
rect 34748 6972 34804 7028
rect 34972 10722 35028 10724
rect 34972 10670 34974 10722
rect 34974 10670 35026 10722
rect 35026 10670 35028 10722
rect 34972 10668 35028 10670
rect 34972 9042 35028 9044
rect 34972 8990 34974 9042
rect 34974 8990 35026 9042
rect 35026 8990 35028 9042
rect 34972 8988 35028 8990
rect 34972 8652 35028 8708
rect 35196 12460 35252 12516
rect 35196 10220 35252 10276
rect 35308 12348 35364 12404
rect 35420 12012 35476 12068
rect 35532 11228 35588 11284
rect 35532 10332 35588 10388
rect 35420 9884 35476 9940
rect 35532 9996 35588 10052
rect 35308 8204 35364 8260
rect 35084 7980 35140 8036
rect 34972 7868 35028 7924
rect 35308 7084 35364 7140
rect 35196 6636 35252 6692
rect 34860 6412 34916 6468
rect 35084 6412 35140 6468
rect 34972 4956 35028 5012
rect 35756 11788 35812 11844
rect 35756 9884 35812 9940
rect 36204 13186 36260 13188
rect 36204 13134 36206 13186
rect 36206 13134 36258 13186
rect 36258 13134 36260 13186
rect 36204 13132 36260 13134
rect 36316 12066 36372 12068
rect 36316 12014 36318 12066
rect 36318 12014 36370 12066
rect 36370 12014 36372 12066
rect 36316 12012 36372 12014
rect 36876 12908 36932 12964
rect 36764 12572 36820 12628
rect 37436 13804 37492 13860
rect 37100 13468 37156 13524
rect 37996 13580 38052 13636
rect 36988 12796 37044 12852
rect 37212 12796 37268 12852
rect 36540 11564 36596 11620
rect 36652 12236 36708 12292
rect 35980 11452 36036 11508
rect 35980 9548 36036 9604
rect 36316 11340 36372 11396
rect 35756 8370 35812 8372
rect 35756 8318 35758 8370
rect 35758 8318 35810 8370
rect 35810 8318 35812 8370
rect 35756 8316 35812 8318
rect 35644 6300 35700 6356
rect 35308 5964 35364 6020
rect 34748 1932 34804 1988
rect 34860 3836 34916 3892
rect 34636 1708 34692 1764
rect 33404 1484 33460 1540
rect 33628 1596 33684 1652
rect 33740 1372 33796 1428
rect 33740 812 33796 868
rect 34860 812 34916 868
rect 35308 3948 35364 4004
rect 35084 3836 35140 3892
rect 35196 3612 35252 3668
rect 35308 3276 35364 3332
rect 35196 1708 35252 1764
rect 35084 1372 35140 1428
rect 35532 5964 35588 6020
rect 35756 4898 35812 4900
rect 35756 4846 35758 4898
rect 35758 4846 35810 4898
rect 35810 4846 35812 4898
rect 35756 4844 35812 4846
rect 36092 7644 36148 7700
rect 36988 12236 37044 12292
rect 36876 12178 36932 12180
rect 36876 12126 36878 12178
rect 36878 12126 36930 12178
rect 36930 12126 36932 12178
rect 36876 12124 36932 12126
rect 36876 11282 36932 11284
rect 36876 11230 36878 11282
rect 36878 11230 36930 11282
rect 36930 11230 36932 11282
rect 36876 11228 36932 11230
rect 36540 9884 36596 9940
rect 36428 8316 36484 8372
rect 36316 8034 36372 8036
rect 36316 7982 36318 8034
rect 36318 7982 36370 8034
rect 36370 7982 36372 8034
rect 36316 7980 36372 7982
rect 36988 10108 37044 10164
rect 36652 8876 36708 8932
rect 36764 8316 36820 8372
rect 36876 9548 36932 9604
rect 37100 9548 37156 9604
rect 36540 7532 36596 7588
rect 36652 7420 36708 7476
rect 37100 7980 37156 8036
rect 36652 5740 36708 5796
rect 36988 6636 37044 6692
rect 37324 11618 37380 11620
rect 37324 11566 37326 11618
rect 37326 11566 37378 11618
rect 37378 11566 37380 11618
rect 37324 11564 37380 11566
rect 37324 10220 37380 10276
rect 37324 9100 37380 9156
rect 37548 8428 37604 8484
rect 37548 7980 37604 8036
rect 37436 7644 37492 7700
rect 37212 6524 37268 6580
rect 37212 6188 37268 6244
rect 36988 5292 37044 5348
rect 37100 4956 37156 5012
rect 37212 5292 37268 5348
rect 35532 3388 35588 3444
rect 36204 3276 36260 3332
rect 35420 1148 35476 1204
rect 35644 2492 35700 2548
rect 34972 588 35028 644
rect 36652 2210 36708 2212
rect 36652 2158 36654 2210
rect 36654 2158 36706 2210
rect 36706 2158 36708 2210
rect 36652 2156 36708 2158
rect 36876 4508 36932 4564
rect 37212 3836 37268 3892
rect 36988 2156 37044 2212
rect 37884 12684 37940 12740
rect 37772 12012 37828 12068
rect 37996 11564 38052 11620
rect 38108 12684 38164 12740
rect 38444 12850 38500 12852
rect 38444 12798 38446 12850
rect 38446 12798 38498 12850
rect 38498 12798 38500 12850
rect 38444 12796 38500 12798
rect 39228 13244 39284 13300
rect 39676 13020 39732 13076
rect 41020 13132 41076 13188
rect 41356 13692 41412 13748
rect 41468 13580 41524 13636
rect 41692 13186 41748 13188
rect 41692 13134 41694 13186
rect 41694 13134 41746 13186
rect 41746 13134 41748 13186
rect 41692 13132 41748 13134
rect 41916 13132 41972 13188
rect 40124 12908 40180 12964
rect 40124 12460 40180 12516
rect 38220 10108 38276 10164
rect 38780 11900 38836 11956
rect 38444 9996 38500 10052
rect 38556 10892 38612 10948
rect 37884 8372 37940 8428
rect 37996 8204 38052 8260
rect 37884 7644 37940 7700
rect 37884 7084 37940 7140
rect 37772 6524 37828 6580
rect 37884 6188 37940 6244
rect 38220 7308 38276 7364
rect 38332 9100 38388 9156
rect 38780 9548 38836 9604
rect 38556 8372 38612 8428
rect 38332 6636 38388 6692
rect 38108 4844 38164 4900
rect 38220 4956 38276 5012
rect 37996 4732 38052 4788
rect 37436 4060 37492 4116
rect 37884 4396 37940 4452
rect 37660 3500 37716 3556
rect 36764 1596 36820 1652
rect 35756 1484 35812 1540
rect 36988 924 37044 980
rect 37996 4172 38052 4228
rect 39004 9548 39060 9604
rect 39116 11228 39172 11284
rect 39004 8370 39060 8372
rect 39004 8318 39006 8370
rect 39006 8318 39058 8370
rect 39058 8318 39060 8370
rect 39004 8316 39060 8318
rect 38780 7532 38836 7588
rect 42140 12348 42196 12404
rect 41356 12290 41412 12292
rect 41356 12238 41358 12290
rect 41358 12238 41410 12290
rect 41410 12238 41412 12290
rect 41356 12236 41412 12238
rect 40124 11788 40180 11844
rect 40348 12012 40404 12068
rect 40236 10556 40292 10612
rect 39452 10444 39508 10500
rect 39900 10444 39956 10500
rect 39676 10332 39732 10388
rect 39564 8930 39620 8932
rect 39564 8878 39566 8930
rect 39566 8878 39618 8930
rect 39618 8878 39620 8930
rect 39564 8876 39620 8878
rect 39340 8204 39396 8260
rect 39452 7420 39508 7476
rect 39116 7196 39172 7252
rect 39452 7084 39508 7140
rect 40236 9996 40292 10052
rect 42252 12066 42308 12068
rect 42252 12014 42254 12066
rect 42254 12014 42306 12066
rect 42306 12014 42308 12066
rect 42252 12012 42308 12014
rect 41692 11900 41748 11956
rect 41244 11452 41300 11508
rect 41580 11452 41636 11508
rect 40460 10386 40516 10388
rect 40460 10334 40462 10386
rect 40462 10334 40514 10386
rect 40514 10334 40516 10386
rect 40460 10332 40516 10334
rect 40348 9436 40404 9492
rect 40124 9324 40180 9380
rect 40012 9042 40068 9044
rect 40012 8990 40014 9042
rect 40014 8990 40066 9042
rect 40066 8990 40068 9042
rect 40012 8988 40068 8990
rect 39788 8818 39844 8820
rect 39788 8766 39790 8818
rect 39790 8766 39842 8818
rect 39842 8766 39844 8818
rect 39788 8764 39844 8766
rect 39676 7084 39732 7140
rect 39788 7308 39844 7364
rect 39900 6748 39956 6804
rect 38668 4956 38724 5012
rect 40236 8428 40292 8484
rect 40236 8092 40292 8148
rect 40684 10498 40740 10500
rect 40684 10446 40686 10498
rect 40686 10446 40738 10498
rect 40738 10446 40740 10498
rect 40684 10444 40740 10446
rect 41580 10444 41636 10500
rect 40908 10220 40964 10276
rect 40684 9042 40740 9044
rect 40684 8990 40686 9042
rect 40686 8990 40738 9042
rect 40738 8990 40740 9042
rect 40684 8988 40740 8990
rect 41244 10108 41300 10164
rect 41132 8988 41188 9044
rect 41020 8258 41076 8260
rect 41020 8206 41022 8258
rect 41022 8206 41074 8258
rect 41074 8206 41076 8258
rect 41020 8204 41076 8206
rect 40908 7868 40964 7924
rect 40572 7308 40628 7364
rect 40012 5628 40068 5684
rect 40124 7196 40180 7252
rect 40460 6972 40516 7028
rect 40124 5516 40180 5572
rect 40236 6860 40292 6916
rect 39564 4844 39620 4900
rect 41356 9154 41412 9156
rect 41356 9102 41358 9154
rect 41358 9102 41410 9154
rect 41410 9102 41412 9154
rect 41356 9100 41412 9102
rect 41468 8764 41524 8820
rect 41244 6860 41300 6916
rect 41132 6802 41188 6804
rect 41132 6750 41134 6802
rect 41134 6750 41186 6802
rect 41186 6750 41188 6802
rect 41132 6748 41188 6750
rect 40460 6636 40516 6692
rect 41468 8204 41524 8260
rect 41916 11452 41972 11508
rect 42028 11676 42084 11732
rect 42700 12796 42756 12852
rect 42924 13580 42980 13636
rect 43036 12908 43092 12964
rect 42812 12124 42868 12180
rect 42924 12572 42980 12628
rect 42700 11676 42756 11732
rect 42812 11900 42868 11956
rect 41804 11394 41860 11396
rect 41804 11342 41806 11394
rect 41806 11342 41858 11394
rect 41858 11342 41860 11394
rect 41804 11340 41860 11342
rect 42364 11340 42420 11396
rect 42252 10610 42308 10612
rect 42252 10558 42254 10610
rect 42254 10558 42306 10610
rect 42306 10558 42308 10610
rect 42252 10556 42308 10558
rect 42252 10332 42308 10388
rect 41916 8540 41972 8596
rect 42252 8370 42308 8372
rect 42252 8318 42254 8370
rect 42254 8318 42306 8370
rect 42306 8318 42308 8370
rect 42252 8316 42308 8318
rect 42140 8204 42196 8260
rect 43036 11676 43092 11732
rect 43484 14028 43540 14084
rect 43820 13186 43876 13188
rect 43820 13134 43822 13186
rect 43822 13134 43874 13186
rect 43874 13134 43876 13186
rect 43820 13132 43876 13134
rect 44604 13580 44660 13636
rect 44940 13468 44996 13524
rect 44464 13354 44520 13356
rect 44464 13302 44466 13354
rect 44466 13302 44518 13354
rect 44518 13302 44520 13354
rect 44464 13300 44520 13302
rect 44568 13354 44624 13356
rect 44568 13302 44570 13354
rect 44570 13302 44622 13354
rect 44622 13302 44624 13354
rect 44568 13300 44624 13302
rect 44672 13354 44728 13356
rect 44672 13302 44674 13354
rect 44674 13302 44726 13354
rect 44726 13302 44728 13354
rect 44672 13300 44728 13302
rect 44156 12908 44212 12964
rect 44380 12850 44436 12852
rect 44380 12798 44382 12850
rect 44382 12798 44434 12850
rect 44434 12798 44436 12850
rect 44380 12796 44436 12798
rect 43804 12570 43860 12572
rect 43596 12460 43652 12516
rect 43804 12518 43806 12570
rect 43806 12518 43858 12570
rect 43858 12518 43860 12570
rect 43804 12516 43860 12518
rect 43908 12570 43964 12572
rect 43908 12518 43910 12570
rect 43910 12518 43962 12570
rect 43962 12518 43964 12570
rect 43908 12516 43964 12518
rect 44012 12570 44068 12572
rect 44012 12518 44014 12570
rect 44014 12518 44066 12570
rect 44066 12518 44068 12570
rect 44012 12516 44068 12518
rect 43036 9884 43092 9940
rect 43260 11228 43316 11284
rect 43148 9042 43204 9044
rect 43148 8990 43150 9042
rect 43150 8990 43202 9042
rect 43202 8990 43204 9042
rect 43148 8988 43204 8990
rect 42588 8092 42644 8148
rect 41356 6636 41412 6692
rect 41804 7084 41860 7140
rect 41468 6466 41524 6468
rect 41468 6414 41470 6466
rect 41470 6414 41522 6466
rect 41522 6414 41524 6466
rect 41468 6412 41524 6414
rect 40236 4844 40292 4900
rect 40460 5180 40516 5236
rect 39004 4172 39060 4228
rect 38332 3052 38388 3108
rect 39116 3948 39172 4004
rect 38444 588 38500 644
rect 38668 2716 38724 2772
rect 39116 2044 39172 2100
rect 39676 3948 39732 4004
rect 38780 1932 38836 1988
rect 38780 812 38836 868
rect 38668 476 38724 532
rect 38556 252 38612 308
rect 40348 3724 40404 3780
rect 40348 3052 40404 3108
rect 42028 7084 42084 7140
rect 41916 5180 41972 5236
rect 42924 8204 42980 8260
rect 42588 7586 42644 7588
rect 42588 7534 42590 7586
rect 42590 7534 42642 7586
rect 42642 7534 42644 7586
rect 42588 7532 42644 7534
rect 42364 6748 42420 6804
rect 42252 6412 42308 6468
rect 42364 5292 42420 5348
rect 42140 4956 42196 5012
rect 41132 4732 41188 4788
rect 40572 2770 40628 2772
rect 40572 2718 40574 2770
rect 40574 2718 40626 2770
rect 40626 2718 40628 2770
rect 40572 2716 40628 2718
rect 40460 2604 40516 2660
rect 40012 2546 40068 2548
rect 40012 2494 40014 2546
rect 40014 2494 40066 2546
rect 40066 2494 40068 2546
rect 40012 2492 40068 2494
rect 42252 4620 42308 4676
rect 41692 4396 41748 4452
rect 41580 3052 41636 3108
rect 42028 3500 42084 3556
rect 42028 2940 42084 2996
rect 42028 1484 42084 1540
rect 42812 6690 42868 6692
rect 42812 6638 42814 6690
rect 42814 6638 42866 6690
rect 42866 6638 42868 6690
rect 42812 6636 42868 6638
rect 42700 3052 42756 3108
rect 42252 2492 42308 2548
rect 43260 7756 43316 7812
rect 43372 10556 43428 10612
rect 43036 7084 43092 7140
rect 43260 7532 43316 7588
rect 43148 6466 43204 6468
rect 43148 6414 43150 6466
rect 43150 6414 43202 6466
rect 43202 6414 43204 6466
rect 43148 6412 43204 6414
rect 44156 12178 44212 12180
rect 44156 12126 44158 12178
rect 44158 12126 44210 12178
rect 44210 12126 44212 12178
rect 44156 12124 44212 12126
rect 44156 11564 44212 11620
rect 44604 12684 44660 12740
rect 45948 13356 46004 13412
rect 45052 12124 45108 12180
rect 45500 13020 45556 13076
rect 45388 12012 45444 12068
rect 44464 11786 44520 11788
rect 44464 11734 44466 11786
rect 44466 11734 44518 11786
rect 44518 11734 44520 11786
rect 44464 11732 44520 11734
rect 44568 11786 44624 11788
rect 44568 11734 44570 11786
rect 44570 11734 44622 11786
rect 44622 11734 44624 11786
rect 44568 11732 44624 11734
rect 44672 11786 44728 11788
rect 44672 11734 44674 11786
rect 44674 11734 44726 11786
rect 44726 11734 44728 11786
rect 44672 11732 44728 11734
rect 44044 11394 44100 11396
rect 44044 11342 44046 11394
rect 44046 11342 44098 11394
rect 44098 11342 44100 11394
rect 44044 11340 44100 11342
rect 43804 11002 43860 11004
rect 43804 10950 43806 11002
rect 43806 10950 43858 11002
rect 43858 10950 43860 11002
rect 43804 10948 43860 10950
rect 43908 11002 43964 11004
rect 43908 10950 43910 11002
rect 43910 10950 43962 11002
rect 43962 10950 43964 11002
rect 43908 10948 43964 10950
rect 44012 11002 44068 11004
rect 44012 10950 44014 11002
rect 44014 10950 44066 11002
rect 44066 10950 44068 11002
rect 44012 10948 44068 10950
rect 44940 11506 44996 11508
rect 44940 11454 44942 11506
rect 44942 11454 44994 11506
rect 44994 11454 44996 11506
rect 44940 11452 44996 11454
rect 44156 10892 44212 10948
rect 44268 10556 44324 10612
rect 44828 10332 44884 10388
rect 44268 10108 44324 10164
rect 44464 10218 44520 10220
rect 44464 10166 44466 10218
rect 44466 10166 44518 10218
rect 44518 10166 44520 10218
rect 44464 10164 44520 10166
rect 44568 10218 44624 10220
rect 44568 10166 44570 10218
rect 44570 10166 44622 10218
rect 44622 10166 44624 10218
rect 44568 10164 44624 10166
rect 44672 10218 44728 10220
rect 44672 10166 44674 10218
rect 44674 10166 44726 10218
rect 44726 10166 44728 10218
rect 44672 10164 44728 10166
rect 43804 9434 43860 9436
rect 43804 9382 43806 9434
rect 43806 9382 43858 9434
rect 43858 9382 43860 9434
rect 43804 9380 43860 9382
rect 43908 9434 43964 9436
rect 43908 9382 43910 9434
rect 43910 9382 43962 9434
rect 43962 9382 43964 9434
rect 43908 9380 43964 9382
rect 44012 9434 44068 9436
rect 44012 9382 44014 9434
rect 44014 9382 44066 9434
rect 44066 9382 44068 9434
rect 44012 9380 44068 9382
rect 43596 9212 43652 9268
rect 44464 8650 44520 8652
rect 44464 8598 44466 8650
rect 44466 8598 44518 8650
rect 44518 8598 44520 8650
rect 44464 8596 44520 8598
rect 44568 8650 44624 8652
rect 44568 8598 44570 8650
rect 44570 8598 44622 8650
rect 44622 8598 44624 8650
rect 44568 8596 44624 8598
rect 44672 8650 44728 8652
rect 44672 8598 44674 8650
rect 44674 8598 44726 8650
rect 44726 8598 44728 8650
rect 44672 8596 44728 8598
rect 43804 7866 43860 7868
rect 43804 7814 43806 7866
rect 43806 7814 43858 7866
rect 43858 7814 43860 7866
rect 43804 7812 43860 7814
rect 43908 7866 43964 7868
rect 43908 7814 43910 7866
rect 43910 7814 43962 7866
rect 43962 7814 43964 7866
rect 43908 7812 43964 7814
rect 44012 7866 44068 7868
rect 44012 7814 44014 7866
rect 44014 7814 44066 7866
rect 44066 7814 44068 7866
rect 44012 7812 44068 7814
rect 43372 7420 43428 7476
rect 43484 7196 43540 7252
rect 43372 5852 43428 5908
rect 43708 7084 43764 7140
rect 44464 7082 44520 7084
rect 44268 6972 44324 7028
rect 44464 7030 44466 7082
rect 44466 7030 44518 7082
rect 44518 7030 44520 7082
rect 44464 7028 44520 7030
rect 44568 7082 44624 7084
rect 44568 7030 44570 7082
rect 44570 7030 44622 7082
rect 44622 7030 44624 7082
rect 44568 7028 44624 7030
rect 44672 7082 44728 7084
rect 44672 7030 44674 7082
rect 44674 7030 44726 7082
rect 44726 7030 44728 7082
rect 44672 7028 44728 7030
rect 44380 6300 44436 6356
rect 43804 6298 43860 6300
rect 43596 6188 43652 6244
rect 43804 6246 43806 6298
rect 43806 6246 43858 6298
rect 43858 6246 43860 6298
rect 43804 6244 43860 6246
rect 43908 6298 43964 6300
rect 43908 6246 43910 6298
rect 43910 6246 43962 6298
rect 43962 6246 43964 6298
rect 43908 6244 43964 6246
rect 44012 6298 44068 6300
rect 44012 6246 44014 6298
rect 44014 6246 44066 6298
rect 44066 6246 44068 6298
rect 44012 6244 44068 6246
rect 44380 6076 44436 6132
rect 44268 5740 44324 5796
rect 44716 5628 44772 5684
rect 44464 5514 44520 5516
rect 44464 5462 44466 5514
rect 44466 5462 44518 5514
rect 44518 5462 44520 5514
rect 44464 5460 44520 5462
rect 44568 5514 44624 5516
rect 44568 5462 44570 5514
rect 44570 5462 44622 5514
rect 44622 5462 44624 5514
rect 44568 5460 44624 5462
rect 44672 5514 44728 5516
rect 44672 5462 44674 5514
rect 44674 5462 44726 5514
rect 44726 5462 44728 5514
rect 44672 5460 44728 5462
rect 44492 5180 44548 5236
rect 43484 5068 43540 5124
rect 43708 5068 43764 5124
rect 43484 4732 43540 4788
rect 43804 4730 43860 4732
rect 43804 4678 43806 4730
rect 43806 4678 43858 4730
rect 43858 4678 43860 4730
rect 43804 4676 43860 4678
rect 43908 4730 43964 4732
rect 43908 4678 43910 4730
rect 43910 4678 43962 4730
rect 43962 4678 43964 4730
rect 43908 4676 43964 4678
rect 44012 4730 44068 4732
rect 44012 4678 44014 4730
rect 44014 4678 44066 4730
rect 44066 4678 44068 4730
rect 44012 4676 44068 4678
rect 44156 4732 44212 4788
rect 43372 4060 43428 4116
rect 44044 3948 44100 4004
rect 44464 3946 44520 3948
rect 43260 3836 43316 3892
rect 44464 3894 44466 3946
rect 44466 3894 44518 3946
rect 44518 3894 44520 3946
rect 44464 3892 44520 3894
rect 44568 3946 44624 3948
rect 44568 3894 44570 3946
rect 44570 3894 44622 3946
rect 44622 3894 44624 3946
rect 44568 3892 44624 3894
rect 44672 3946 44728 3948
rect 44672 3894 44674 3946
rect 44674 3894 44726 3946
rect 44726 3894 44728 3946
rect 44672 3892 44728 3894
rect 43804 3162 43860 3164
rect 43804 3110 43806 3162
rect 43806 3110 43858 3162
rect 43858 3110 43860 3162
rect 43804 3108 43860 3110
rect 43908 3162 43964 3164
rect 43908 3110 43910 3162
rect 43910 3110 43962 3162
rect 43962 3110 43964 3162
rect 43908 3108 43964 3110
rect 44012 3162 44068 3164
rect 44012 3110 44014 3162
rect 44014 3110 44066 3162
rect 44066 3110 44068 3162
rect 44012 3108 44068 3110
rect 45500 11340 45556 11396
rect 45388 10332 45444 10388
rect 45052 5964 45108 6020
rect 45500 8316 45556 8372
rect 45164 5180 45220 5236
rect 45052 4338 45108 4340
rect 45052 4286 45054 4338
rect 45054 4286 45106 4338
rect 45106 4286 45108 4338
rect 45052 4284 45108 4286
rect 45164 3276 45220 3332
rect 45276 4956 45332 5012
rect 44828 3052 44884 3108
rect 42924 1932 42980 1988
rect 44268 2380 44324 2436
rect 43804 1594 43860 1596
rect 43804 1542 43806 1594
rect 43806 1542 43858 1594
rect 43858 1542 43860 1594
rect 43804 1540 43860 1542
rect 43908 1594 43964 1596
rect 43908 1542 43910 1594
rect 43910 1542 43962 1594
rect 43962 1542 43964 1594
rect 43908 1540 43964 1542
rect 44012 1594 44068 1596
rect 44012 1542 44014 1594
rect 44014 1542 44066 1594
rect 44066 1542 44068 1594
rect 44012 1540 44068 1542
rect 44044 1372 44100 1428
rect 42140 140 42196 196
rect 43708 588 43764 644
rect 44464 2378 44520 2380
rect 44464 2326 44466 2378
rect 44466 2326 44518 2378
rect 44518 2326 44520 2378
rect 44464 2324 44520 2326
rect 44568 2378 44624 2380
rect 44568 2326 44570 2378
rect 44570 2326 44622 2378
rect 44622 2326 44624 2378
rect 44568 2324 44624 2326
rect 44672 2378 44728 2380
rect 44672 2326 44674 2378
rect 44674 2326 44726 2378
rect 44726 2326 44728 2378
rect 44672 2324 44728 2326
rect 45500 4396 45556 4452
rect 45948 12850 46004 12852
rect 45948 12798 45950 12850
rect 45950 12798 46002 12850
rect 46002 12798 46004 12850
rect 45948 12796 46004 12798
rect 46956 13916 47012 13972
rect 46620 12908 46676 12964
rect 45948 11788 46004 11844
rect 46060 11282 46116 11284
rect 46060 11230 46062 11282
rect 46062 11230 46114 11282
rect 46114 11230 46116 11282
rect 46060 11228 46116 11230
rect 46844 11900 46900 11956
rect 46844 11676 46900 11732
rect 46620 11564 46676 11620
rect 47180 13132 47236 13188
rect 47068 11900 47124 11956
rect 46508 11452 46564 11508
rect 45724 7084 45780 7140
rect 45836 6914 45892 6916
rect 45836 6862 45838 6914
rect 45838 6862 45890 6914
rect 45890 6862 45892 6914
rect 45836 6860 45892 6862
rect 46172 11004 46228 11060
rect 46060 10220 46116 10276
rect 45948 6188 46004 6244
rect 47068 10556 47124 10612
rect 46396 10050 46452 10052
rect 46396 9998 46398 10050
rect 46398 9998 46450 10050
rect 46450 9998 46452 10050
rect 46396 9996 46452 9998
rect 47628 13580 47684 13636
rect 47516 10556 47572 10612
rect 47852 13692 47908 13748
rect 48188 13132 48244 13188
rect 47964 12908 48020 12964
rect 49084 13468 49140 13524
rect 49308 13804 49364 13860
rect 48972 13186 49028 13188
rect 48972 13134 48974 13186
rect 48974 13134 49026 13186
rect 49026 13134 49028 13186
rect 48972 13132 49028 13134
rect 48412 12236 48468 12292
rect 48412 12012 48468 12068
rect 46956 10108 47012 10164
rect 46844 8092 46900 8148
rect 47180 9100 47236 9156
rect 47068 7644 47124 7700
rect 47068 6524 47124 6580
rect 47180 4956 47236 5012
rect 46284 4844 46340 4900
rect 46172 4284 46228 4340
rect 48188 10668 48244 10724
rect 48300 10498 48356 10500
rect 48300 10446 48302 10498
rect 48302 10446 48354 10498
rect 48354 10446 48356 10498
rect 48300 10444 48356 10446
rect 49196 11676 49252 11732
rect 48524 11452 48580 11508
rect 49084 11564 49140 11620
rect 48860 11116 48916 11172
rect 48076 8818 48132 8820
rect 48076 8766 48078 8818
rect 48078 8766 48130 8818
rect 48130 8766 48132 8818
rect 48076 8764 48132 8766
rect 48412 8652 48468 8708
rect 48076 7756 48132 7812
rect 47404 5516 47460 5572
rect 47404 4956 47460 5012
rect 47852 3500 47908 3556
rect 48300 7420 48356 7476
rect 48300 5964 48356 6020
rect 48076 3164 48132 3220
rect 48524 4732 48580 4788
rect 48636 6300 48692 6356
rect 49084 9996 49140 10052
rect 48860 9436 48916 9492
rect 48972 9042 49028 9044
rect 48972 8990 48974 9042
rect 48974 8990 49026 9042
rect 49026 8990 49028 9042
rect 48972 8988 49028 8990
rect 49084 8764 49140 8820
rect 48972 5906 49028 5908
rect 48972 5854 48974 5906
rect 48974 5854 49026 5906
rect 49026 5854 49028 5906
rect 48972 5852 49028 5854
rect 48748 2940 48804 2996
rect 45276 1596 45332 1652
rect 44268 1372 44324 1428
rect 44464 810 44520 812
rect 44464 758 44466 810
rect 44466 758 44518 810
rect 44518 758 44520 810
rect 44464 756 44520 758
rect 44568 810 44624 812
rect 44568 758 44570 810
rect 44570 758 44622 810
rect 44622 758 44624 810
rect 44568 756 44624 758
rect 44672 810 44728 812
rect 44672 758 44674 810
rect 44674 758 44726 810
rect 44726 758 44728 810
rect 44672 756 44728 758
rect 45612 588 45668 644
rect 45724 1484 45780 1540
rect 44044 364 44100 420
rect 48636 2604 48692 2660
rect 49980 13020 50036 13076
rect 50428 12348 50484 12404
rect 49532 11564 49588 11620
rect 49644 11004 49700 11060
rect 49756 10108 49812 10164
rect 49420 9548 49476 9604
rect 49980 9212 50036 9268
rect 49196 7420 49252 7476
rect 49644 8764 49700 8820
rect 49420 6018 49476 6020
rect 49420 5966 49422 6018
rect 49422 5966 49474 6018
rect 49474 5966 49476 6018
rect 49420 5964 49476 5966
rect 49308 1596 49364 1652
rect 48636 1036 48692 1092
rect 48524 812 48580 868
rect 47404 476 47460 532
rect 49868 8428 49924 8484
rect 49868 6860 49924 6916
rect 50428 11954 50484 11956
rect 50428 11902 50430 11954
rect 50430 11902 50482 11954
rect 50482 11902 50484 11954
rect 50428 11900 50484 11902
rect 50316 11618 50372 11620
rect 50316 11566 50318 11618
rect 50318 11566 50370 11618
rect 50370 11566 50372 11618
rect 50316 11564 50372 11566
rect 50204 9938 50260 9940
rect 50204 9886 50206 9938
rect 50206 9886 50258 9938
rect 50258 9886 50260 9938
rect 50204 9884 50260 9886
rect 50204 8930 50260 8932
rect 50204 8878 50206 8930
rect 50206 8878 50258 8930
rect 50258 8878 50260 8930
rect 50204 8876 50260 8878
rect 50316 8370 50372 8372
rect 50316 8318 50318 8370
rect 50318 8318 50370 8370
rect 50370 8318 50372 8370
rect 50316 8316 50372 8318
rect 50540 7586 50596 7588
rect 50540 7534 50542 7586
rect 50542 7534 50594 7586
rect 50594 7534 50596 7586
rect 50540 7532 50596 7534
rect 50540 6690 50596 6692
rect 50540 6638 50542 6690
rect 50542 6638 50594 6690
rect 50594 6638 50596 6690
rect 50540 6636 50596 6638
rect 50092 5068 50148 5124
rect 51100 13468 51156 13524
rect 50876 12684 50932 12740
rect 50876 11340 50932 11396
rect 50764 11116 50820 11172
rect 49868 2492 49924 2548
rect 50428 3612 50484 3668
rect 50652 3276 50708 3332
rect 50988 9826 51044 9828
rect 50988 9774 50990 9826
rect 50990 9774 51042 9826
rect 51042 9774 51044 9826
rect 50988 9772 51044 9774
rect 51100 9154 51156 9156
rect 51100 9102 51102 9154
rect 51102 9102 51154 9154
rect 51154 9102 51156 9154
rect 51100 9100 51156 9102
rect 50876 7474 50932 7476
rect 50876 7422 50878 7474
rect 50878 7422 50930 7474
rect 50930 7422 50932 7474
rect 50876 7420 50932 7422
rect 50988 6860 51044 6916
rect 51100 6690 51156 6692
rect 51100 6638 51102 6690
rect 51102 6638 51154 6690
rect 51154 6638 51156 6690
rect 51100 6636 51156 6638
rect 51324 11564 51380 11620
rect 51660 13356 51716 13412
rect 51436 10498 51492 10500
rect 51436 10446 51438 10498
rect 51438 10446 51490 10498
rect 51490 10446 51492 10498
rect 51436 10444 51492 10446
rect 51324 10220 51380 10276
rect 51548 10220 51604 10276
rect 51436 7362 51492 7364
rect 51436 7310 51438 7362
rect 51438 7310 51490 7362
rect 51490 7310 51492 7362
rect 51436 7308 51492 7310
rect 51212 2716 51268 2772
rect 51324 3276 51380 3332
rect 51772 13244 51828 13300
rect 52220 13132 52276 13188
rect 53116 13356 53172 13412
rect 52892 13074 52948 13076
rect 52892 13022 52894 13074
rect 52894 13022 52946 13074
rect 52946 13022 52948 13074
rect 52892 13020 52948 13022
rect 52108 12684 52164 12740
rect 51996 10668 52052 10724
rect 51884 10444 51940 10500
rect 51772 10220 51828 10276
rect 52108 10610 52164 10612
rect 52108 10558 52110 10610
rect 52110 10558 52162 10610
rect 52162 10558 52164 10610
rect 52108 10556 52164 10558
rect 51996 9042 52052 9044
rect 51996 8990 51998 9042
rect 51998 8990 52050 9042
rect 52050 8990 52052 9042
rect 51996 8988 52052 8990
rect 52108 8876 52164 8932
rect 52220 8316 52276 8372
rect 52332 9436 52388 9492
rect 52108 7644 52164 7700
rect 52108 7196 52164 7252
rect 52108 5180 52164 5236
rect 51884 5068 51940 5124
rect 51436 1820 51492 1876
rect 51660 2098 51716 2100
rect 51660 2046 51662 2098
rect 51662 2046 51714 2098
rect 51714 2046 51716 2098
rect 51660 2044 51716 2046
rect 51548 1484 51604 1540
rect 50988 1260 51044 1316
rect 49756 924 49812 980
rect 49644 364 49700 420
rect 49756 700 49812 756
rect 47740 140 47796 196
rect 51996 2770 52052 2772
rect 51996 2718 51998 2770
rect 51998 2718 52050 2770
rect 52050 2718 52052 2770
rect 51996 2716 52052 2718
rect 51884 2044 51940 2100
rect 52556 12402 52612 12404
rect 52556 12350 52558 12402
rect 52558 12350 52610 12402
rect 52610 12350 52612 12402
rect 52556 12348 52612 12350
rect 52556 11564 52612 11620
rect 53788 13468 53844 13524
rect 52556 8428 52612 8484
rect 52556 8258 52612 8260
rect 52556 8206 52558 8258
rect 52558 8206 52610 8258
rect 52610 8206 52612 8258
rect 52556 8204 52612 8206
rect 52444 7532 52500 7588
rect 52556 5628 52612 5684
rect 52332 4844 52388 4900
rect 52332 4284 52388 4340
rect 52220 3554 52276 3556
rect 52220 3502 52222 3554
rect 52222 3502 52274 3554
rect 52274 3502 52276 3554
rect 52220 3500 52276 3502
rect 52332 2604 52388 2660
rect 52220 2098 52276 2100
rect 52220 2046 52222 2098
rect 52222 2046 52274 2098
rect 52274 2046 52276 2098
rect 52220 2044 52276 2046
rect 52108 1372 52164 1428
rect 52556 4620 52612 4676
rect 52668 4226 52724 4228
rect 52668 4174 52670 4226
rect 52670 4174 52722 4226
rect 52722 4174 52724 4226
rect 52668 4172 52724 4174
rect 53004 9266 53060 9268
rect 53004 9214 53006 9266
rect 53006 9214 53058 9266
rect 53058 9214 53060 9266
rect 53004 9212 53060 9214
rect 53340 8370 53396 8372
rect 53340 8318 53342 8370
rect 53342 8318 53394 8370
rect 53394 8318 53396 8370
rect 53340 8316 53396 8318
rect 53004 7868 53060 7924
rect 53788 9884 53844 9940
rect 53900 10444 53956 10500
rect 53676 9436 53732 9492
rect 53564 8540 53620 8596
rect 52892 6636 52948 6692
rect 53228 6524 53284 6580
rect 53004 6188 53060 6244
rect 53116 4450 53172 4452
rect 53116 4398 53118 4450
rect 53118 4398 53170 4450
rect 53170 4398 53172 4450
rect 53116 4396 53172 4398
rect 52780 3276 52836 3332
rect 52556 3164 52612 3220
rect 53564 6578 53620 6580
rect 53564 6526 53566 6578
rect 53566 6526 53618 6578
rect 53618 6526 53620 6578
rect 53564 6524 53620 6526
rect 53452 6076 53508 6132
rect 54124 13244 54180 13300
rect 54012 9212 54068 9268
rect 53900 6524 53956 6580
rect 53676 5010 53732 5012
rect 53676 4958 53678 5010
rect 53678 4958 53730 5010
rect 53730 4958 53732 5010
rect 53676 4956 53732 4958
rect 53564 4508 53620 4564
rect 53564 3442 53620 3444
rect 53564 3390 53566 3442
rect 53566 3390 53618 3442
rect 53618 3390 53620 3442
rect 53564 3388 53620 3390
rect 53340 2828 53396 2884
rect 54124 7980 54180 8036
rect 54124 5740 54180 5796
rect 54124 4844 54180 4900
rect 54908 13692 54964 13748
rect 54908 13186 54964 13188
rect 54908 13134 54910 13186
rect 54910 13134 54962 13186
rect 54962 13134 54964 13186
rect 54908 13132 54964 13134
rect 55356 12908 55412 12964
rect 55692 13356 55748 13412
rect 54684 12572 54740 12628
rect 54348 11340 54404 11396
rect 54348 8540 54404 8596
rect 54236 4284 54292 4340
rect 54124 3724 54180 3780
rect 53564 3052 53620 3108
rect 52780 2658 52836 2660
rect 52780 2606 52782 2658
rect 52782 2606 52834 2658
rect 52834 2606 52836 2658
rect 52780 2604 52836 2606
rect 53564 1874 53620 1876
rect 53564 1822 53566 1874
rect 53566 1822 53618 1874
rect 53618 1822 53620 1874
rect 53564 1820 53620 1822
rect 53564 1426 53620 1428
rect 53564 1374 53566 1426
rect 53566 1374 53618 1426
rect 53618 1374 53620 1426
rect 53564 1372 53620 1374
rect 51996 924 52052 980
rect 54124 1708 54180 1764
rect 53676 588 53732 644
rect 53788 812 53844 868
rect 55020 11506 55076 11508
rect 55020 11454 55022 11506
rect 55022 11454 55074 11506
rect 55074 11454 55076 11506
rect 55020 11452 55076 11454
rect 55132 10780 55188 10836
rect 54684 10220 54740 10276
rect 54572 10108 54628 10164
rect 55580 11228 55636 11284
rect 55244 9996 55300 10052
rect 55468 10332 55524 10388
rect 55132 9436 55188 9492
rect 55132 8930 55188 8932
rect 55132 8878 55134 8930
rect 55134 8878 55186 8930
rect 55186 8878 55188 8930
rect 55132 8876 55188 8878
rect 56252 12796 56308 12852
rect 56364 13916 56420 13972
rect 55804 10444 55860 10500
rect 56364 9100 56420 9156
rect 56140 8988 56196 9044
rect 55580 8316 55636 8372
rect 55916 8092 55972 8148
rect 56140 7698 56196 7700
rect 56140 7646 56142 7698
rect 56142 7646 56194 7698
rect 56194 7646 56196 7698
rect 56140 7644 56196 7646
rect 54572 7196 54628 7252
rect 55244 6412 55300 6468
rect 55356 7084 55412 7140
rect 55132 6300 55188 6356
rect 54572 5852 54628 5908
rect 55132 5292 55188 5348
rect 54908 5122 54964 5124
rect 54908 5070 54910 5122
rect 54910 5070 54962 5122
rect 54962 5070 54964 5122
rect 54908 5068 54964 5070
rect 54572 4562 54628 4564
rect 54572 4510 54574 4562
rect 54574 4510 54626 4562
rect 54626 4510 54628 4562
rect 54572 4508 54628 4510
rect 55132 4060 55188 4116
rect 54908 3666 54964 3668
rect 54908 3614 54910 3666
rect 54910 3614 54962 3666
rect 54962 3614 54964 3666
rect 54908 3612 54964 3614
rect 54572 3164 54628 3220
rect 56140 6748 56196 6804
rect 57036 13020 57092 13076
rect 57036 11004 57092 11060
rect 57260 12124 57316 12180
rect 57260 7868 57316 7924
rect 56700 6188 56756 6244
rect 56140 5404 56196 5460
rect 56140 4060 56196 4116
rect 57036 3388 57092 3444
rect 56140 2716 56196 2772
rect 54908 2268 54964 2324
rect 56924 2604 56980 2660
rect 55132 1202 55188 1204
rect 55132 1150 55134 1202
rect 55134 1150 55186 1202
rect 55186 1150 55188 1202
rect 55132 1148 55188 1150
rect 54460 700 54516 756
rect 55804 1036 55860 1092
rect 32284 28 32340 84
rect 57036 476 57092 532
rect 56924 28 56980 84
<< metal3 >>
rect 21074 14140 21084 14196
rect 21140 14140 25340 14196
rect 25396 14140 25406 14196
rect 25564 14140 28476 14196
rect 28532 14140 28542 14196
rect 28690 14140 28700 14196
rect 28756 14140 34524 14196
rect 34580 14140 34590 14196
rect 34738 14140 34748 14196
rect 34804 14140 47012 14196
rect 25564 14084 25620 14140
rect 14802 14028 14812 14084
rect 14868 14028 23772 14084
rect 23828 14028 23838 14084
rect 24210 14028 24220 14084
rect 24276 14028 25620 14084
rect 26898 14028 26908 14084
rect 26964 14028 43484 14084
rect 43540 14028 43550 14084
rect 0 13972 112 14000
rect 46956 13972 47012 14140
rect 57344 13972 57456 14000
rect 0 13916 2380 13972
rect 2436 13916 2446 13972
rect 12562 13916 12572 13972
rect 12628 13916 25228 13972
rect 25284 13916 25294 13972
rect 25442 13916 25452 13972
rect 25508 13916 28924 13972
rect 28980 13916 28990 13972
rect 33404 13916 40236 13972
rect 40292 13916 40302 13972
rect 46946 13916 46956 13972
rect 47012 13916 47022 13972
rect 56354 13916 56364 13972
rect 56420 13916 57456 13972
rect 0 13888 112 13916
rect 10770 13804 10780 13860
rect 10836 13804 21420 13860
rect 21476 13804 21486 13860
rect 21970 13804 21980 13860
rect 22036 13804 26012 13860
rect 26068 13804 26078 13860
rect 26226 13804 26236 13860
rect 26292 13804 27244 13860
rect 27300 13804 27310 13860
rect 27468 13804 32732 13860
rect 32788 13804 32798 13860
rect 27468 13748 27524 13804
rect 33404 13748 33460 13916
rect 57344 13888 57456 13916
rect 33730 13804 33740 13860
rect 33796 13804 34748 13860
rect 34804 13804 34814 13860
rect 37426 13804 37436 13860
rect 37492 13804 49308 13860
rect 49364 13804 49374 13860
rect 7298 13692 7308 13748
rect 7364 13692 20636 13748
rect 20692 13692 20702 13748
rect 23650 13692 23660 13748
rect 23716 13692 27524 13748
rect 27682 13692 27692 13748
rect 27748 13692 28588 13748
rect 28644 13692 28654 13748
rect 28802 13692 28812 13748
rect 28868 13692 33460 13748
rect 33516 13692 41356 13748
rect 41412 13692 41422 13748
rect 47842 13692 47852 13748
rect 47908 13692 54908 13748
rect 54964 13692 54974 13748
rect 33516 13636 33572 13692
rect 12450 13580 12460 13636
rect 12516 13580 18508 13636
rect 18564 13580 18574 13636
rect 20178 13580 20188 13636
rect 20244 13580 25060 13636
rect 26226 13580 26236 13636
rect 26292 13580 28700 13636
rect 28756 13580 28766 13636
rect 28914 13580 28924 13636
rect 28980 13580 33572 13636
rect 33842 13580 33852 13636
rect 33908 13580 35308 13636
rect 35364 13580 35374 13636
rect 35634 13580 35644 13636
rect 35700 13580 37996 13636
rect 38052 13580 38062 13636
rect 41458 13580 41468 13636
rect 41524 13580 42924 13636
rect 42980 13580 42990 13636
rect 44594 13580 44604 13636
rect 44660 13580 47628 13636
rect 47684 13580 47694 13636
rect 0 13524 112 13552
rect 25004 13524 25060 13580
rect 57344 13524 57456 13552
rect 0 13468 1484 13524
rect 1540 13468 1550 13524
rect 3602 13468 3612 13524
rect 3668 13468 4732 13524
rect 4788 13468 4798 13524
rect 16706 13468 16716 13524
rect 16772 13468 24948 13524
rect 25004 13468 28028 13524
rect 28084 13468 28094 13524
rect 28578 13468 28588 13524
rect 28644 13468 33404 13524
rect 33460 13468 33470 13524
rect 35186 13468 35196 13524
rect 35252 13468 37100 13524
rect 37156 13468 37166 13524
rect 37650 13468 37660 13524
rect 37716 13468 44940 13524
rect 44996 13468 45006 13524
rect 49074 13468 49084 13524
rect 49140 13468 51100 13524
rect 51156 13468 51166 13524
rect 53778 13468 53788 13524
rect 53844 13468 57456 13524
rect 0 13440 112 13468
rect 2146 13356 2156 13412
rect 2212 13356 4284 13412
rect 4340 13356 4350 13412
rect 7522 13356 7532 13412
rect 7588 13356 9660 13412
rect 9716 13356 9726 13412
rect 11778 13356 11788 13412
rect 11844 13356 13524 13412
rect 14466 13356 14476 13412
rect 14532 13356 22876 13412
rect 22932 13356 22942 13412
rect 23202 13356 23212 13412
rect 23268 13356 24220 13412
rect 24276 13356 24286 13412
rect 4454 13300 4464 13356
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4728 13300 4738 13356
rect 13468 13300 13524 13356
rect 24454 13300 24464 13356
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24728 13300 24738 13356
rect 24892 13300 24948 13468
rect 57344 13440 57456 13468
rect 27458 13356 27468 13412
rect 27524 13356 33628 13412
rect 33684 13356 33694 13412
rect 45938 13356 45948 13412
rect 46004 13356 51660 13412
rect 51716 13356 51726 13412
rect 53106 13356 53116 13412
rect 53172 13356 55692 13412
rect 55748 13356 55758 13412
rect 44454 13300 44464 13356
rect 44520 13300 44568 13356
rect 44624 13300 44672 13356
rect 44728 13300 44738 13356
rect 8194 13244 8204 13300
rect 8260 13244 10108 13300
rect 10164 13244 10174 13300
rect 11330 13244 11340 13300
rect 11396 13244 13244 13300
rect 13300 13244 13310 13300
rect 13468 13244 20748 13300
rect 20804 13244 20814 13300
rect 21186 13244 21196 13300
rect 21252 13244 24388 13300
rect 24892 13244 29484 13300
rect 29540 13244 29550 13300
rect 30818 13244 30828 13300
rect 30884 13244 34468 13300
rect 39218 13244 39228 13300
rect 39284 13244 44100 13300
rect 51762 13244 51772 13300
rect 51828 13244 54124 13300
rect 54180 13244 54190 13300
rect 24332 13188 24388 13244
rect 3714 13132 3724 13188
rect 3780 13132 5628 13188
rect 5684 13132 5694 13188
rect 5954 13132 5964 13188
rect 6020 13132 7420 13188
rect 7476 13132 7486 13188
rect 9762 13132 9772 13188
rect 9828 13132 11900 13188
rect 11956 13132 11966 13188
rect 13346 13132 13356 13188
rect 13412 13132 15036 13188
rect 15092 13132 15102 13188
rect 17378 13132 17388 13188
rect 17444 13132 18620 13188
rect 18676 13132 18686 13188
rect 18946 13132 18956 13188
rect 19012 13132 19964 13188
rect 20020 13132 20030 13188
rect 23538 13132 23548 13188
rect 23604 13132 23642 13188
rect 24332 13132 25788 13188
rect 25844 13132 25854 13188
rect 26786 13132 26796 13188
rect 26852 13132 29036 13188
rect 29092 13132 29102 13188
rect 30706 13132 30716 13188
rect 30772 13132 31500 13188
rect 31556 13132 31566 13188
rect 31714 13132 31724 13188
rect 31780 13132 32732 13188
rect 32788 13132 32798 13188
rect 32946 13132 32956 13188
rect 33012 13132 34188 13188
rect 34244 13132 34254 13188
rect 0 13076 112 13104
rect 34412 13076 34468 13244
rect 44044 13188 44100 13244
rect 34738 13132 34748 13188
rect 34804 13132 36204 13188
rect 36260 13132 36270 13188
rect 41010 13132 41020 13188
rect 41076 13132 41692 13188
rect 41748 13132 41758 13188
rect 41906 13132 41916 13188
rect 41972 13132 43820 13188
rect 43876 13132 43886 13188
rect 44044 13132 47180 13188
rect 47236 13132 47246 13188
rect 48178 13132 48188 13188
rect 48244 13132 48972 13188
rect 49028 13132 49038 13188
rect 52210 13132 52220 13188
rect 52276 13132 54908 13188
rect 54964 13132 54974 13188
rect 57344 13076 57456 13104
rect 0 13020 588 13076
rect 644 13020 654 13076
rect 10098 13020 10108 13076
rect 10164 13020 11004 13076
rect 11060 13020 11070 13076
rect 14914 13020 14924 13076
rect 14980 13020 16828 13076
rect 16884 13020 16894 13076
rect 18498 13020 18508 13076
rect 18564 13020 22428 13076
rect 22484 13020 22494 13076
rect 23986 13020 23996 13076
rect 24052 13020 24780 13076
rect 24836 13020 24846 13076
rect 27906 13020 27916 13076
rect 27972 13020 28756 13076
rect 31602 13020 31612 13076
rect 31668 13020 33292 13076
rect 33348 13020 33358 13076
rect 33506 13020 33516 13076
rect 33572 13020 34132 13076
rect 34412 13020 35868 13076
rect 35924 13020 35934 13076
rect 39666 13020 39676 13076
rect 39732 13020 45500 13076
rect 45556 13020 45566 13076
rect 49970 13020 49980 13076
rect 50036 13020 52892 13076
rect 52948 13020 52958 13076
rect 57026 13020 57036 13076
rect 57092 13020 57456 13076
rect 0 12992 112 13020
rect 28700 12964 28756 13020
rect 34076 12964 34132 13020
rect 57344 12992 57456 13020
rect 4274 12908 4284 12964
rect 4340 12908 5964 12964
rect 6020 12908 6030 12964
rect 14354 12908 14364 12964
rect 14420 12908 20524 12964
rect 20580 12908 20590 12964
rect 22978 12908 22988 12964
rect 23044 12908 28252 12964
rect 28308 12908 28318 12964
rect 28700 12908 33852 12964
rect 33908 12908 33918 12964
rect 34076 12908 36876 12964
rect 36932 12908 36942 12964
rect 40114 12908 40124 12964
rect 40180 12908 43036 12964
rect 43092 12908 43102 12964
rect 44146 12908 44156 12964
rect 44212 12908 46620 12964
rect 46676 12908 46686 12964
rect 47954 12908 47964 12964
rect 48020 12908 55356 12964
rect 55412 12908 55422 12964
rect 23538 12796 23548 12852
rect 23604 12796 23772 12852
rect 23828 12796 23838 12852
rect 23996 12796 26236 12852
rect 26292 12796 26302 12852
rect 27010 12796 27020 12852
rect 27076 12796 29148 12852
rect 29204 12796 29214 12852
rect 29474 12796 29484 12852
rect 29540 12796 33292 12852
rect 33348 12796 33358 12852
rect 33506 12796 33516 12852
rect 33572 12796 36988 12852
rect 37044 12796 37054 12852
rect 37202 12796 37212 12852
rect 37268 12796 38444 12852
rect 38500 12796 38510 12852
rect 42690 12796 42700 12852
rect 42756 12796 44380 12852
rect 44436 12796 44446 12852
rect 45938 12796 45948 12852
rect 46004 12796 56252 12852
rect 56308 12796 56318 12852
rect 23996 12740 24052 12796
rect 2818 12684 2828 12740
rect 2884 12684 11284 12740
rect 21298 12684 21308 12740
rect 21364 12684 21980 12740
rect 22036 12684 22046 12740
rect 22204 12684 24052 12740
rect 24210 12684 24220 12740
rect 24276 12684 30940 12740
rect 30996 12684 31006 12740
rect 32722 12684 32732 12740
rect 32788 12684 37884 12740
rect 37940 12684 37950 12740
rect 38098 12684 38108 12740
rect 38164 12684 44604 12740
rect 44660 12684 44670 12740
rect 50866 12684 50876 12740
rect 50932 12684 52108 12740
rect 52164 12684 52174 12740
rect 0 12628 112 12656
rect 0 12572 3500 12628
rect 3556 12572 3566 12628
rect 0 12544 112 12572
rect 3794 12516 3804 12572
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 4068 12516 4078 12572
rect 2258 12348 2268 12404
rect 2324 12348 3388 12404
rect 3444 12348 3454 12404
rect 11228 12292 11284 12684
rect 17938 12572 17948 12628
rect 18004 12572 21644 12628
rect 21700 12572 21710 12628
rect 20850 12460 20860 12516
rect 20916 12460 21868 12516
rect 21924 12460 21934 12516
rect 22204 12404 22260 12684
rect 57344 12628 57456 12656
rect 24658 12572 24668 12628
rect 24724 12572 24892 12628
rect 24948 12572 24958 12628
rect 25218 12572 25228 12628
rect 25284 12572 33180 12628
rect 33236 12572 33246 12628
rect 36754 12572 36764 12628
rect 36820 12572 42924 12628
rect 42980 12572 42990 12628
rect 54674 12572 54684 12628
rect 54740 12572 57456 12628
rect 23794 12516 23804 12572
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 24068 12516 24078 12572
rect 43794 12516 43804 12572
rect 43860 12516 43908 12572
rect 43964 12516 44012 12572
rect 44068 12516 44078 12572
rect 57344 12544 57456 12572
rect 22642 12460 22652 12516
rect 22708 12460 23212 12516
rect 23268 12460 23278 12516
rect 23426 12460 23436 12516
rect 12002 12348 12012 12404
rect 12068 12348 12796 12404
rect 12852 12348 12862 12404
rect 14802 12348 14812 12404
rect 14868 12348 15932 12404
rect 15988 12348 15998 12404
rect 16370 12348 16380 12404
rect 16436 12348 17276 12404
rect 17332 12348 17342 12404
rect 18274 12348 18284 12404
rect 18340 12348 21308 12404
rect 21364 12348 21374 12404
rect 21522 12348 21532 12404
rect 21588 12348 22260 12404
rect 23492 12404 23548 12516
rect 24220 12460 31948 12516
rect 32004 12460 32014 12516
rect 33282 12460 33292 12516
rect 33348 12460 35196 12516
rect 35252 12460 35262 12516
rect 40114 12460 40124 12516
rect 40180 12460 43596 12516
rect 43652 12460 43662 12516
rect 24220 12404 24276 12460
rect 23492 12348 24276 12404
rect 24892 12348 25564 12404
rect 25620 12348 25630 12404
rect 25778 12348 25788 12404
rect 25844 12348 28700 12404
rect 28756 12348 28766 12404
rect 28914 12348 28924 12404
rect 28980 12348 30996 12404
rect 31490 12348 31500 12404
rect 31556 12348 34188 12404
rect 34244 12348 34254 12404
rect 35298 12348 35308 12404
rect 35364 12348 42140 12404
rect 42196 12348 42206 12404
rect 50418 12348 50428 12404
rect 50484 12348 52556 12404
rect 52612 12348 52622 12404
rect 24892 12292 24948 12348
rect 30940 12292 30996 12348
rect 5058 12236 5068 12292
rect 5124 12236 11004 12292
rect 11060 12236 11070 12292
rect 11228 12236 20860 12292
rect 20916 12236 20926 12292
rect 21084 12236 24948 12292
rect 25106 12236 25116 12292
rect 25172 12236 30716 12292
rect 30772 12236 30782 12292
rect 30940 12236 32620 12292
rect 32676 12236 32686 12292
rect 32946 12236 32956 12292
rect 33012 12236 36652 12292
rect 36708 12236 36718 12292
rect 36978 12236 36988 12292
rect 37044 12236 41356 12292
rect 41412 12236 41422 12292
rect 42588 12236 48412 12292
rect 48468 12236 48478 12292
rect 0 12180 112 12208
rect 21084 12180 21140 12236
rect 42588 12180 42644 12236
rect 57344 12180 57456 12208
rect 0 12124 252 12180
rect 308 12124 318 12180
rect 2930 12124 2940 12180
rect 2996 12124 3388 12180
rect 3444 12124 3454 12180
rect 4386 12124 4396 12180
rect 4452 12124 11788 12180
rect 11844 12124 11854 12180
rect 12002 12124 12012 12180
rect 12068 12124 18228 12180
rect 18358 12124 18396 12180
rect 18452 12124 18462 12180
rect 20290 12124 20300 12180
rect 20356 12124 21140 12180
rect 21410 12124 21420 12180
rect 21476 12124 28476 12180
rect 28532 12124 28542 12180
rect 29362 12124 29372 12180
rect 29428 12124 32284 12180
rect 32340 12124 32350 12180
rect 32498 12124 32508 12180
rect 32564 12124 33180 12180
rect 33236 12124 33246 12180
rect 33394 12124 33404 12180
rect 33460 12124 34076 12180
rect 34132 12124 34142 12180
rect 34290 12124 34300 12180
rect 34356 12124 34972 12180
rect 35028 12124 35038 12180
rect 36866 12124 36876 12180
rect 36932 12124 42644 12180
rect 42802 12124 42812 12180
rect 42868 12124 44156 12180
rect 44212 12124 44222 12180
rect 45042 12124 45052 12180
rect 45108 12124 48468 12180
rect 57250 12124 57260 12180
rect 57316 12124 57456 12180
rect 0 12096 112 12124
rect 18172 12068 18228 12124
rect 48412 12068 48468 12124
rect 57344 12096 57456 12124
rect 4946 12012 4956 12068
rect 5012 12012 7140 12068
rect 8194 12012 8204 12068
rect 8260 12012 17948 12068
rect 18004 12012 18014 12068
rect 18172 12012 21980 12068
rect 22036 12012 22046 12068
rect 22194 12012 22204 12068
rect 22260 12012 30604 12068
rect 30660 12012 30670 12068
rect 31154 12012 31164 12068
rect 31220 12012 32396 12068
rect 32452 12012 32462 12068
rect 34402 12012 34412 12068
rect 34468 12012 35420 12068
rect 35476 12012 36316 12068
rect 36372 12012 37772 12068
rect 37828 12012 37838 12068
rect 40338 12012 40348 12068
rect 40404 12012 42252 12068
rect 42308 12012 42318 12068
rect 42476 12012 45388 12068
rect 45444 12012 45454 12068
rect 48402 12012 48412 12068
rect 48468 12012 48478 12068
rect 7084 11956 7140 12012
rect 1586 11900 1596 11956
rect 1652 11900 2268 11956
rect 2324 11900 2334 11956
rect 6066 11900 6076 11956
rect 6132 11900 6860 11956
rect 6916 11900 6926 11956
rect 7084 11900 9380 11956
rect 11218 11900 11228 11956
rect 11284 11900 13244 11956
rect 13300 11900 13310 11956
rect 16594 11900 16604 11956
rect 16660 11900 25340 11956
rect 25396 11900 25406 11956
rect 25554 11900 25564 11956
rect 25620 11900 30044 11956
rect 30100 11900 30110 11956
rect 33954 11900 33964 11956
rect 34020 11900 36036 11956
rect 38770 11900 38780 11956
rect 38836 11900 41692 11956
rect 41748 11900 41758 11956
rect 1138 11788 1148 11844
rect 1204 11788 2156 11844
rect 2212 11788 2222 11844
rect 6962 11788 6972 11844
rect 7028 11788 8316 11844
rect 8372 11788 8382 11844
rect 0 11732 112 11760
rect 4454 11732 4464 11788
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4728 11732 4738 11788
rect 9324 11732 9380 11900
rect 35980 11844 36036 11900
rect 42476 11844 42532 12012
rect 42802 11900 42812 11956
rect 42868 11900 46844 11956
rect 46900 11900 46910 11956
rect 47058 11900 47068 11956
rect 47124 11900 50428 11956
rect 50484 11900 50494 11956
rect 10098 11788 10108 11844
rect 10164 11788 12012 11844
rect 12068 11788 12078 11844
rect 17154 11788 17164 11844
rect 17220 11788 23548 11844
rect 23604 11788 23614 11844
rect 23772 11788 24220 11844
rect 24276 11788 24286 11844
rect 25890 11788 25900 11844
rect 25956 11788 28196 11844
rect 34962 11788 34972 11844
rect 35028 11788 35756 11844
rect 35812 11788 35822 11844
rect 35980 11788 40124 11844
rect 40180 11788 40190 11844
rect 40348 11788 42532 11844
rect 45910 11788 45948 11844
rect 46004 11788 46014 11844
rect 23772 11732 23828 11788
rect 24454 11732 24464 11788
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24728 11732 24738 11788
rect 28140 11732 28196 11788
rect 40348 11732 40404 11788
rect 44454 11732 44464 11788
rect 44520 11732 44568 11788
rect 44624 11732 44672 11788
rect 44728 11732 44738 11788
rect 57344 11732 57456 11760
rect 0 11676 1932 11732
rect 1988 11676 1998 11732
rect 9324 11676 18284 11732
rect 18340 11676 18350 11732
rect 20066 11676 20076 11732
rect 20132 11676 23828 11732
rect 24892 11676 27860 11732
rect 28140 11676 30380 11732
rect 30436 11676 30446 11732
rect 31938 11676 31948 11732
rect 32004 11676 40404 11732
rect 42018 11676 42028 11732
rect 42084 11676 42700 11732
rect 42756 11676 42766 11732
rect 43026 11676 43036 11732
rect 43092 11676 44156 11732
rect 44212 11676 44222 11732
rect 46834 11676 46844 11732
rect 46900 11676 46938 11732
rect 49186 11676 49196 11732
rect 49252 11676 57456 11732
rect 0 11648 112 11676
rect 24892 11620 24948 11676
rect 27804 11620 27860 11676
rect 57344 11648 57456 11676
rect 4610 11564 4620 11620
rect 4676 11564 5180 11620
rect 5236 11564 5246 11620
rect 6178 11564 6188 11620
rect 6244 11564 6748 11620
rect 6804 11564 6814 11620
rect 7746 11564 7756 11620
rect 7812 11564 8764 11620
rect 8820 11564 8830 11620
rect 14578 11564 14588 11620
rect 14644 11564 16716 11620
rect 16772 11564 16782 11620
rect 16930 11564 16940 11620
rect 16996 11564 24948 11620
rect 26002 11564 26012 11620
rect 26068 11564 26684 11620
rect 26740 11564 27580 11620
rect 27636 11564 27646 11620
rect 27804 11564 28812 11620
rect 28868 11564 28878 11620
rect 29026 11564 29036 11620
rect 29092 11564 33516 11620
rect 33572 11564 33582 11620
rect 36530 11564 36540 11620
rect 36596 11564 37324 11620
rect 37380 11564 37390 11620
rect 37986 11564 37996 11620
rect 38052 11564 44156 11620
rect 44212 11564 44222 11620
rect 46610 11564 46620 11620
rect 46676 11564 46714 11620
rect 46946 11564 46956 11620
rect 47012 11564 49084 11620
rect 49140 11564 49150 11620
rect 49522 11564 49532 11620
rect 49588 11564 50316 11620
rect 50372 11564 50382 11620
rect 51314 11564 51324 11620
rect 51380 11564 52556 11620
rect 52612 11564 52622 11620
rect 14130 11452 14140 11508
rect 14196 11452 28588 11508
rect 28644 11452 28654 11508
rect 28812 11452 31724 11508
rect 31780 11452 31790 11508
rect 32386 11452 32396 11508
rect 32452 11452 34524 11508
rect 34580 11452 34590 11508
rect 35970 11452 35980 11508
rect 36036 11452 38668 11508
rect 41234 11452 41244 11508
rect 41300 11452 41580 11508
rect 41636 11452 41916 11508
rect 41972 11452 44940 11508
rect 44996 11452 45006 11508
rect 46470 11452 46508 11508
rect 46564 11452 46574 11508
rect 48514 11452 48524 11508
rect 48580 11452 55020 11508
rect 55076 11452 55086 11508
rect 28812 11396 28868 11452
rect 38612 11396 38668 11452
rect 5282 11340 5292 11396
rect 5348 11340 19516 11396
rect 19572 11340 19582 11396
rect 21186 11340 21196 11396
rect 21252 11340 23100 11396
rect 23156 11340 23166 11396
rect 23324 11340 26908 11396
rect 26964 11340 26974 11396
rect 27570 11340 27580 11396
rect 27636 11340 28868 11396
rect 29026 11340 29036 11396
rect 29092 11340 31276 11396
rect 31332 11340 31342 11396
rect 31490 11340 31500 11396
rect 31556 11340 36316 11396
rect 36372 11340 36382 11396
rect 38612 11340 41804 11396
rect 41860 11340 42364 11396
rect 42420 11340 42430 11396
rect 42588 11340 44044 11396
rect 44100 11340 44110 11396
rect 45490 11340 45500 11396
rect 45556 11340 50428 11396
rect 50866 11340 50876 11396
rect 50932 11340 54348 11396
rect 54404 11340 54414 11396
rect 0 11284 112 11312
rect 23324 11284 23380 11340
rect 42588 11284 42644 11340
rect 0 11228 1820 11284
rect 1876 11228 1886 11284
rect 20178 11228 20188 11284
rect 20244 11228 23380 11284
rect 23986 11228 23996 11284
rect 24052 11228 28588 11284
rect 28644 11228 28654 11284
rect 31826 11228 31836 11284
rect 31892 11228 35308 11284
rect 35364 11228 35374 11284
rect 35522 11228 35532 11284
rect 35588 11228 36876 11284
rect 36932 11228 36942 11284
rect 39106 11228 39116 11284
rect 39172 11228 42644 11284
rect 43250 11228 43260 11284
rect 43316 11228 46060 11284
rect 46116 11228 46126 11284
rect 0 11200 112 11228
rect 50372 11172 50428 11340
rect 57344 11284 57456 11312
rect 55570 11228 55580 11284
rect 55636 11228 57456 11284
rect 57344 11200 57456 11228
rect 8418 11116 8428 11172
rect 8484 11116 24276 11172
rect 24434 11116 24444 11172
rect 24500 11116 31052 11172
rect 31108 11116 31118 11172
rect 33506 11116 33516 11172
rect 33572 11116 42700 11172
rect 42756 11116 42766 11172
rect 43596 11116 48860 11172
rect 48916 11116 48926 11172
rect 50372 11116 50764 11172
rect 50820 11116 50830 11172
rect 24220 11060 24276 11116
rect 43596 11060 43652 11116
rect 5506 11004 5516 11060
rect 5572 11004 12460 11060
rect 12516 11004 12526 11060
rect 13234 11004 13244 11060
rect 13300 11004 22204 11060
rect 22260 11004 22270 11060
rect 24220 11004 28028 11060
rect 28084 11004 28094 11060
rect 28354 11004 28364 11060
rect 28420 11004 32564 11060
rect 32722 11004 32732 11060
rect 32788 11004 43652 11060
rect 44146 11004 44156 11060
rect 44212 11004 46172 11060
rect 46228 11004 46238 11060
rect 49634 11004 49644 11060
rect 49700 11004 57036 11060
rect 57092 11004 57102 11060
rect 3794 10948 3804 11004
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 4068 10948 4078 11004
rect 23794 10948 23804 11004
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 24068 10948 24078 11004
rect 32508 10948 32564 11004
rect 43794 10948 43804 11004
rect 43860 10948 43908 11004
rect 43964 10948 44012 11004
rect 44068 10948 44078 11004
rect 5170 10892 5180 10948
rect 5236 10892 5628 10948
rect 5684 10892 5694 10948
rect 17938 10892 17948 10948
rect 18004 10892 21756 10948
rect 21812 10892 21822 10948
rect 26898 10892 26908 10948
rect 26964 10892 31948 10948
rect 32508 10892 38556 10948
rect 38612 10892 38622 10948
rect 44146 10892 44156 10948
rect 44212 10892 46956 10948
rect 47012 10892 47022 10948
rect 0 10836 112 10864
rect 31892 10836 31948 10892
rect 57344 10836 57456 10864
rect 0 10780 1148 10836
rect 1204 10780 1214 10836
rect 1474 10780 1484 10836
rect 1540 10780 5852 10836
rect 5908 10780 5918 10836
rect 8978 10780 8988 10836
rect 9044 10780 31500 10836
rect 31556 10780 31566 10836
rect 31892 10780 38780 10836
rect 38836 10780 38846 10836
rect 42578 10780 42588 10836
rect 42644 10780 55132 10836
rect 55188 10780 55198 10836
rect 55412 10780 57456 10836
rect 0 10752 112 10780
rect 55412 10724 55468 10780
rect 57344 10752 57456 10780
rect 2706 10668 2716 10724
rect 2772 10668 4172 10724
rect 4228 10668 4238 10724
rect 4386 10668 4396 10724
rect 4452 10668 11900 10724
rect 11956 10668 11966 10724
rect 18274 10668 18284 10724
rect 18340 10668 27692 10724
rect 27748 10668 27758 10724
rect 28578 10668 28588 10724
rect 28644 10668 29484 10724
rect 29540 10668 29550 10724
rect 29810 10668 29820 10724
rect 29876 10668 30828 10724
rect 30884 10668 30894 10724
rect 31042 10668 31052 10724
rect 31108 10668 31948 10724
rect 32004 10668 32014 10724
rect 32610 10668 32620 10724
rect 32676 10668 34804 10724
rect 34962 10668 34972 10724
rect 35028 10668 48188 10724
rect 48244 10668 48254 10724
rect 51986 10668 51996 10724
rect 52052 10668 55468 10724
rect 34748 10612 34804 10668
rect 2818 10556 2828 10612
rect 2884 10556 4956 10612
rect 5012 10556 5022 10612
rect 7410 10556 7420 10612
rect 7476 10556 10780 10612
rect 10836 10556 10846 10612
rect 10994 10556 11004 10612
rect 11060 10556 19404 10612
rect 19460 10556 19470 10612
rect 21970 10556 21980 10612
rect 22036 10556 27468 10612
rect 27524 10556 27534 10612
rect 29138 10556 29148 10612
rect 29204 10556 34524 10612
rect 34580 10556 34590 10612
rect 34748 10556 40236 10612
rect 40292 10556 40302 10612
rect 40674 10556 40684 10612
rect 40740 10556 41860 10612
rect 42242 10556 42252 10612
rect 42308 10556 43372 10612
rect 43428 10556 43438 10612
rect 44258 10556 44268 10612
rect 44324 10556 47068 10612
rect 47124 10556 47134 10612
rect 47506 10556 47516 10612
rect 47572 10556 52108 10612
rect 52164 10556 52174 10612
rect 41804 10500 41860 10556
rect 1922 10444 1932 10500
rect 1988 10444 2716 10500
rect 2772 10444 2782 10500
rect 3602 10444 3612 10500
rect 3668 10444 5180 10500
rect 5236 10444 5246 10500
rect 12114 10444 12124 10500
rect 12180 10444 14252 10500
rect 14308 10444 14318 10500
rect 14466 10444 14476 10500
rect 14532 10444 17164 10500
rect 17220 10444 17230 10500
rect 17378 10444 17388 10500
rect 17444 10444 21084 10500
rect 21140 10444 21150 10500
rect 22316 10444 22540 10500
rect 22596 10444 22606 10500
rect 22754 10444 22764 10500
rect 22820 10444 24892 10500
rect 24948 10444 24958 10500
rect 25330 10444 25340 10500
rect 25396 10444 27580 10500
rect 27636 10444 27646 10500
rect 27794 10444 27804 10500
rect 27860 10444 32396 10500
rect 32452 10444 32462 10500
rect 33842 10444 33852 10500
rect 33908 10444 38220 10500
rect 38276 10444 38286 10500
rect 39442 10444 39452 10500
rect 39508 10444 39900 10500
rect 39956 10444 40684 10500
rect 40740 10444 41580 10500
rect 41636 10444 41646 10500
rect 41804 10444 42252 10500
rect 42308 10444 42318 10500
rect 42476 10444 48300 10500
rect 48356 10444 48366 10500
rect 51426 10444 51436 10500
rect 51492 10444 51884 10500
rect 51940 10444 51950 10500
rect 53890 10444 53900 10500
rect 53956 10444 55804 10500
rect 55860 10444 55870 10500
rect 0 10388 112 10416
rect 22316 10388 22372 10444
rect 0 10332 2828 10388
rect 2884 10332 2894 10388
rect 11732 10332 20300 10388
rect 20356 10332 20366 10388
rect 20860 10332 22372 10388
rect 22978 10332 22988 10388
rect 23044 10332 27132 10388
rect 27188 10332 27198 10388
rect 27356 10332 28476 10388
rect 28532 10332 28542 10388
rect 28690 10332 28700 10388
rect 28756 10332 30492 10388
rect 30548 10332 30558 10388
rect 30818 10332 30828 10388
rect 30884 10332 35532 10388
rect 35588 10332 35598 10388
rect 36876 10332 39676 10388
rect 39732 10332 39742 10388
rect 40450 10332 40460 10388
rect 40516 10332 42252 10388
rect 42308 10332 42318 10388
rect 0 10304 112 10332
rect 11732 10276 11788 10332
rect 20860 10276 20916 10332
rect 10546 10220 10556 10276
rect 10612 10220 11788 10276
rect 13122 10220 13132 10276
rect 13188 10220 14476 10276
rect 14532 10220 14542 10276
rect 15698 10220 15708 10276
rect 15764 10220 17780 10276
rect 17938 10220 17948 10276
rect 18004 10220 18172 10276
rect 18228 10220 18238 10276
rect 19852 10220 20916 10276
rect 21074 10220 21084 10276
rect 21140 10220 23212 10276
rect 23268 10220 23278 10276
rect 23426 10220 23436 10276
rect 23492 10220 24220 10276
rect 24276 10220 24286 10276
rect 25106 10220 25116 10276
rect 25172 10220 26796 10276
rect 26852 10220 26862 10276
rect 4454 10164 4464 10220
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4728 10164 4738 10220
rect 17724 10164 17780 10220
rect 19852 10164 19908 10220
rect 24454 10164 24464 10220
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24728 10164 24738 10220
rect 27356 10164 27412 10332
rect 36876 10276 36932 10332
rect 42476 10276 42532 10444
rect 57344 10388 57456 10416
rect 42690 10332 42700 10388
rect 42756 10332 44828 10388
rect 44884 10332 44894 10388
rect 45378 10332 45388 10388
rect 45444 10332 51604 10388
rect 55458 10332 55468 10388
rect 55524 10332 57456 10388
rect 51548 10276 51604 10332
rect 57344 10304 57456 10332
rect 28130 10220 28140 10276
rect 28196 10220 34188 10276
rect 34244 10220 34254 10276
rect 34402 10220 34412 10276
rect 34468 10220 34748 10276
rect 34804 10220 34814 10276
rect 35186 10220 35196 10276
rect 35252 10220 36932 10276
rect 37314 10220 37324 10276
rect 37380 10220 40684 10276
rect 40740 10220 40750 10276
rect 40898 10220 40908 10276
rect 40964 10220 42532 10276
rect 46050 10220 46060 10276
rect 46116 10220 51324 10276
rect 51380 10220 51390 10276
rect 51538 10220 51548 10276
rect 51604 10220 51614 10276
rect 51762 10220 51772 10276
rect 51828 10220 54684 10276
rect 54740 10220 54750 10276
rect 44454 10164 44464 10220
rect 44520 10164 44568 10220
rect 44624 10164 44672 10220
rect 44728 10164 44738 10220
rect 1474 10108 1484 10164
rect 1540 10108 4340 10164
rect 4284 10052 4340 10108
rect 4844 10108 9212 10164
rect 9268 10108 9884 10164
rect 9940 10108 9950 10164
rect 11106 10108 11116 10164
rect 11172 10108 12124 10164
rect 12180 10108 12190 10164
rect 13346 10108 13356 10164
rect 13412 10108 15820 10164
rect 15876 10108 15886 10164
rect 17724 10108 19908 10164
rect 20066 10108 20076 10164
rect 20132 10108 23324 10164
rect 23380 10108 23390 10164
rect 24210 10108 24220 10164
rect 24276 10108 24332 10164
rect 24388 10108 24398 10164
rect 25218 10108 25228 10164
rect 25284 10108 27412 10164
rect 28242 10108 28252 10164
rect 28308 10108 30156 10164
rect 30212 10108 30222 10164
rect 30482 10108 30492 10164
rect 30548 10108 33180 10164
rect 33236 10108 33246 10164
rect 35308 10108 36988 10164
rect 37044 10108 37054 10164
rect 38210 10108 38220 10164
rect 38276 10108 41244 10164
rect 41300 10108 41310 10164
rect 41682 10108 41692 10164
rect 41748 10108 44268 10164
rect 44324 10108 44334 10164
rect 46946 10108 46956 10164
rect 47012 10108 49756 10164
rect 49812 10108 49822 10164
rect 54562 10108 54572 10164
rect 54628 10108 55468 10164
rect 4844 10052 4900 10108
rect 35308 10052 35364 10108
rect 4284 9996 4900 10052
rect 18834 9996 18844 10052
rect 18900 9996 22092 10052
rect 22148 9996 22158 10052
rect 22428 9996 22988 10052
rect 23044 9996 23054 10052
rect 23202 9996 23212 10052
rect 23268 9996 23996 10052
rect 24052 9996 26124 10052
rect 26180 9996 26190 10052
rect 26674 9996 26684 10052
rect 26740 9996 26908 10052
rect 26964 9996 26974 10052
rect 27234 9996 27244 10052
rect 27300 9996 28084 10052
rect 28242 9996 28252 10052
rect 28308 9996 35364 10052
rect 35522 9996 35532 10052
rect 35588 9996 38444 10052
rect 38500 9996 38510 10052
rect 40226 9996 40236 10052
rect 40292 9996 46396 10052
rect 46452 9996 46462 10052
rect 49074 9996 49084 10052
rect 49140 9996 55244 10052
rect 55300 9996 55310 10052
rect 0 9940 112 9968
rect 22428 9940 22484 9996
rect 28028 9940 28084 9996
rect 55412 9940 55468 10108
rect 57344 9940 57456 9968
rect 0 9884 5068 9940
rect 5124 9884 5134 9940
rect 17826 9884 17836 9940
rect 17892 9884 22484 9940
rect 22642 9884 22652 9940
rect 22708 9884 24388 9940
rect 24546 9884 24556 9940
rect 24612 9884 25340 9940
rect 25396 9884 25406 9940
rect 25554 9884 25564 9940
rect 25620 9884 27580 9940
rect 27636 9884 27646 9940
rect 28028 9884 33292 9940
rect 33348 9884 34076 9940
rect 34132 9884 35420 9940
rect 35476 9884 35756 9940
rect 35812 9884 35822 9940
rect 36530 9884 36540 9940
rect 36596 9884 43036 9940
rect 43092 9884 43102 9940
rect 50194 9884 50204 9940
rect 50260 9884 53788 9940
rect 53844 9884 53854 9940
rect 55412 9884 57456 9940
rect 0 9856 112 9884
rect 24332 9828 24388 9884
rect 57344 9856 57456 9884
rect 1586 9772 1596 9828
rect 1652 9772 7980 9828
rect 8036 9772 8046 9828
rect 10434 9772 10444 9828
rect 10500 9772 11788 9828
rect 11844 9772 11854 9828
rect 17714 9772 17724 9828
rect 17780 9772 18284 9828
rect 18340 9772 20188 9828
rect 20244 9772 20254 9828
rect 20738 9772 20748 9828
rect 20804 9772 23548 9828
rect 23604 9772 23614 9828
rect 24332 9772 26124 9828
rect 26180 9772 26190 9828
rect 28476 9772 50988 9828
rect 51044 9772 51054 9828
rect 6178 9660 6188 9716
rect 6244 9660 10108 9716
rect 10164 9660 10174 9716
rect 12002 9660 12012 9716
rect 12068 9660 20300 9716
rect 20356 9660 20366 9716
rect 20514 9660 20524 9716
rect 20580 9660 22652 9716
rect 22708 9660 22718 9716
rect 23090 9660 23100 9716
rect 23156 9660 28252 9716
rect 28308 9660 28318 9716
rect 28476 9604 28532 9772
rect 30594 9660 30604 9716
rect 30660 9660 53732 9716
rect 2258 9548 2268 9604
rect 2324 9548 11004 9604
rect 11060 9548 11070 9604
rect 12226 9548 12236 9604
rect 12292 9548 25228 9604
rect 25284 9548 25294 9604
rect 25564 9548 28532 9604
rect 28802 9548 28812 9604
rect 28868 9548 33516 9604
rect 33572 9548 33582 9604
rect 35970 9548 35980 9604
rect 36036 9548 36876 9604
rect 36932 9548 36942 9604
rect 37090 9548 37100 9604
rect 37156 9548 38780 9604
rect 38836 9548 38846 9604
rect 38994 9548 39004 9604
rect 39060 9548 49420 9604
rect 49476 9548 49486 9604
rect 0 9492 112 9520
rect 0 9436 3668 9492
rect 12002 9436 12012 9492
rect 12068 9436 12908 9492
rect 12964 9436 12974 9492
rect 13122 9436 13132 9492
rect 13188 9436 16604 9492
rect 16660 9436 16670 9492
rect 17938 9436 17948 9492
rect 18004 9436 22652 9492
rect 22708 9436 22718 9492
rect 24210 9436 24220 9492
rect 24276 9436 25340 9492
rect 25396 9436 25406 9492
rect 0 9408 112 9436
rect 1922 9324 1932 9380
rect 1988 9324 2380 9380
rect 2436 9324 2446 9380
rect 3612 9268 3668 9436
rect 3794 9380 3804 9436
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 4068 9380 4078 9436
rect 23794 9380 23804 9436
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 24068 9380 24078 9436
rect 25564 9380 25620 9548
rect 53676 9492 53732 9660
rect 57344 9492 57456 9520
rect 25778 9436 25788 9492
rect 25844 9436 27244 9492
rect 27300 9436 27310 9492
rect 27906 9436 27916 9492
rect 27972 9436 29820 9492
rect 29876 9436 29886 9492
rect 30258 9436 30268 9492
rect 30324 9436 40348 9492
rect 40404 9436 40414 9492
rect 48850 9436 48860 9492
rect 48916 9436 52332 9492
rect 52388 9436 52398 9492
rect 53666 9436 53676 9492
rect 53732 9436 53742 9492
rect 55122 9436 55132 9492
rect 55188 9436 57456 9492
rect 43794 9380 43804 9436
rect 43860 9380 43908 9436
rect 43964 9380 44012 9436
rect 44068 9380 44078 9436
rect 57344 9408 57456 9436
rect 10882 9324 10892 9380
rect 10948 9324 18284 9380
rect 18340 9324 18350 9380
rect 19282 9324 19292 9380
rect 19348 9324 23548 9380
rect 23604 9324 23614 9380
rect 24220 9324 25620 9380
rect 25778 9324 25788 9380
rect 25844 9324 33964 9380
rect 34020 9324 34030 9380
rect 34178 9324 34188 9380
rect 34244 9324 40124 9380
rect 40180 9324 40190 9380
rect 24220 9268 24276 9324
rect 802 9212 812 9268
rect 868 9212 3388 9268
rect 3612 9212 3836 9268
rect 3892 9212 3902 9268
rect 4060 9212 12572 9268
rect 12628 9212 12638 9268
rect 19394 9212 19404 9268
rect 19460 9212 21756 9268
rect 21812 9212 21822 9268
rect 22194 9212 22204 9268
rect 22260 9212 24276 9268
rect 24434 9212 24444 9268
rect 24500 9212 25116 9268
rect 25172 9212 25182 9268
rect 25442 9212 25452 9268
rect 25508 9212 28252 9268
rect 28308 9212 28318 9268
rect 31938 9212 31948 9268
rect 32004 9212 36876 9268
rect 36932 9212 36942 9268
rect 39554 9212 39564 9268
rect 39620 9212 42252 9268
rect 42308 9212 42318 9268
rect 43586 9212 43596 9268
rect 43652 9212 49980 9268
rect 50036 9212 50046 9268
rect 52994 9212 53004 9268
rect 53060 9212 54012 9268
rect 54068 9212 54078 9268
rect 3332 9156 3388 9212
rect 4060 9156 4116 9212
rect 3332 9100 4116 9156
rect 5618 9100 5628 9156
rect 5684 9100 5694 9156
rect 11890 9100 11900 9156
rect 11956 9100 18060 9156
rect 18116 9100 18126 9156
rect 18610 9100 18620 9156
rect 18676 9100 20860 9156
rect 20916 9100 20926 9156
rect 21746 9100 21756 9156
rect 21812 9100 26684 9156
rect 26740 9100 26750 9156
rect 26842 9100 26852 9156
rect 26908 9100 33740 9156
rect 33796 9100 33806 9156
rect 33954 9100 33964 9156
rect 34020 9100 37324 9156
rect 37380 9100 37390 9156
rect 38322 9100 38332 9156
rect 38388 9100 41356 9156
rect 41412 9100 41422 9156
rect 41906 9100 41916 9156
rect 41972 9100 45948 9156
rect 46004 9100 46014 9156
rect 47170 9100 47180 9156
rect 47236 9100 50428 9156
rect 51090 9100 51100 9156
rect 51156 9100 56364 9156
rect 56420 9100 56430 9156
rect 0 9044 112 9072
rect 5628 9044 5684 9100
rect 50372 9044 50428 9100
rect 57344 9044 57456 9072
rect 0 8988 1036 9044
rect 1092 8988 1102 9044
rect 5628 8988 17948 9044
rect 18004 8988 18014 9044
rect 18274 8988 18284 9044
rect 18340 8988 21308 9044
rect 21364 8988 21374 9044
rect 21634 8988 21644 9044
rect 21700 8988 22260 9044
rect 24098 8988 24108 9044
rect 24164 8988 25564 9044
rect 25620 8988 25630 9044
rect 25890 8988 25900 9044
rect 25956 8988 28924 9044
rect 28980 8988 28990 9044
rect 29148 8988 30828 9044
rect 30884 8988 30894 9044
rect 32610 8988 32620 9044
rect 32676 8988 33404 9044
rect 33460 8988 33470 9044
rect 34962 8988 34972 9044
rect 35028 8988 40012 9044
rect 40068 8988 40684 9044
rect 40740 8988 40750 9044
rect 41122 8988 41132 9044
rect 41188 8988 43148 9044
rect 43204 8988 43214 9044
rect 43372 8988 48972 9044
rect 49028 8988 49038 9044
rect 50372 8988 51996 9044
rect 52052 8988 52062 9044
rect 56130 8988 56140 9044
rect 56196 8988 57456 9044
rect 0 8960 112 8988
rect 22204 8932 22260 8988
rect 29148 8932 29204 8988
rect 43372 8932 43428 8988
rect 57344 8960 57456 8988
rect 3490 8876 3500 8932
rect 3556 8876 9660 8932
rect 9716 8876 9726 8932
rect 13794 8876 13804 8932
rect 13860 8876 21980 8932
rect 22036 8876 22046 8932
rect 22204 8876 25228 8932
rect 25284 8876 25294 8932
rect 26338 8876 26348 8932
rect 26404 8876 29204 8932
rect 30706 8876 30716 8932
rect 30772 8876 32508 8932
rect 32564 8876 33516 8932
rect 33572 8876 33582 8932
rect 33730 8876 33740 8932
rect 33796 8876 35364 8932
rect 36642 8876 36652 8932
rect 36708 8876 39564 8932
rect 39620 8876 39630 8932
rect 41794 8876 41804 8932
rect 41860 8876 43428 8932
rect 44268 8876 50204 8932
rect 50260 8876 50270 8932
rect 52098 8876 52108 8932
rect 52164 8876 55132 8932
rect 55188 8876 55198 8932
rect 35308 8820 35364 8876
rect 4386 8764 4396 8820
rect 4452 8764 6300 8820
rect 6356 8764 6366 8820
rect 7522 8764 7532 8820
rect 7588 8764 13692 8820
rect 13748 8764 13758 8820
rect 16482 8764 16492 8820
rect 16548 8764 17780 8820
rect 19954 8764 19964 8820
rect 20020 8764 21980 8820
rect 22036 8764 22046 8820
rect 23090 8764 23100 8820
rect 23156 8764 26908 8820
rect 26964 8764 26974 8820
rect 27122 8764 27132 8820
rect 27188 8764 32060 8820
rect 32116 8764 32126 8820
rect 33170 8764 33180 8820
rect 33236 8764 33628 8820
rect 33684 8764 33852 8820
rect 33908 8764 33918 8820
rect 34066 8764 34076 8820
rect 34132 8764 35252 8820
rect 35308 8764 39564 8820
rect 39620 8764 39630 8820
rect 39778 8764 39788 8820
rect 39844 8764 41468 8820
rect 41524 8764 41534 8820
rect 17724 8708 17780 8764
rect 35196 8708 35252 8764
rect 44268 8708 44324 8876
rect 48066 8764 48076 8820
rect 48132 8764 49084 8820
rect 49140 8764 49150 8820
rect 49634 8764 49644 8820
rect 49700 8764 50428 8820
rect 6402 8652 6412 8708
rect 6468 8652 17500 8708
rect 17556 8652 17566 8708
rect 17724 8652 22764 8708
rect 22820 8652 22830 8708
rect 25554 8652 25564 8708
rect 25620 8652 27468 8708
rect 27524 8652 27534 8708
rect 27682 8652 27692 8708
rect 27748 8652 29708 8708
rect 29764 8652 29774 8708
rect 31892 8652 34972 8708
rect 35028 8652 35038 8708
rect 35196 8652 44324 8708
rect 48402 8652 48412 8708
rect 48468 8652 50260 8708
rect 0 8596 112 8624
rect 4454 8596 4464 8652
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4728 8596 4738 8652
rect 24454 8596 24464 8652
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24728 8596 24738 8652
rect 31892 8596 31948 8652
rect 44454 8596 44464 8652
rect 44520 8596 44568 8652
rect 44624 8596 44672 8652
rect 44728 8596 44738 8652
rect 0 8540 2940 8596
rect 2996 8540 3006 8596
rect 9762 8540 9772 8596
rect 9828 8540 12684 8596
rect 12740 8540 12750 8596
rect 13010 8540 13020 8596
rect 13076 8540 14252 8596
rect 14308 8540 14318 8596
rect 15092 8540 22092 8596
rect 22148 8540 22158 8596
rect 22306 8540 22316 8596
rect 22372 8540 24332 8596
rect 24388 8540 24398 8596
rect 24882 8540 24892 8596
rect 24948 8540 28924 8596
rect 28980 8540 28990 8596
rect 30930 8540 30940 8596
rect 30996 8540 31948 8596
rect 32162 8540 32172 8596
rect 32228 8540 41916 8596
rect 41972 8540 41982 8596
rect 0 8512 112 8540
rect 15092 8484 15148 8540
rect 50204 8484 50260 8652
rect 50372 8596 50428 8764
rect 57344 8596 57456 8624
rect 50372 8540 53564 8596
rect 53620 8540 53630 8596
rect 54338 8540 54348 8596
rect 54404 8540 57456 8596
rect 57344 8512 57456 8540
rect 5394 8428 5404 8484
rect 5460 8428 13132 8484
rect 13188 8428 13198 8484
rect 13346 8428 13356 8484
rect 13412 8428 13422 8484
rect 13570 8428 13580 8484
rect 13636 8428 15148 8484
rect 15362 8428 15372 8484
rect 15428 8428 21532 8484
rect 21588 8428 21598 8484
rect 21868 8428 28364 8484
rect 28420 8428 28430 8484
rect 28588 8428 31276 8484
rect 31332 8428 31342 8484
rect 33506 8428 33516 8484
rect 33572 8428 33582 8484
rect 34962 8428 34972 8484
rect 35028 8428 37548 8484
rect 37604 8428 37614 8484
rect 37884 8428 38612 8484
rect 40226 8428 40236 8484
rect 40292 8428 49868 8484
rect 49924 8428 49934 8484
rect 50204 8428 52556 8484
rect 52612 8428 52622 8484
rect 13356 8372 13412 8428
rect 21868 8372 21924 8428
rect 28588 8372 28644 8428
rect 33516 8372 33572 8428
rect 37874 8372 37884 8428
rect 37940 8372 37950 8428
rect 38546 8372 38556 8428
rect 38612 8372 38622 8428
rect 4050 8316 4060 8372
rect 4116 8316 8428 8372
rect 8484 8316 8494 8372
rect 9762 8316 9772 8372
rect 9828 8316 13132 8372
rect 13188 8316 13198 8372
rect 13356 8316 21924 8372
rect 22166 8316 22204 8372
rect 22260 8316 22270 8372
rect 22754 8316 22764 8372
rect 22820 8316 24892 8372
rect 24948 8316 24958 8372
rect 25218 8316 25228 8372
rect 25284 8316 28028 8372
rect 28084 8316 28094 8372
rect 28588 8316 28700 8372
rect 28756 8316 28766 8372
rect 33516 8316 35588 8372
rect 35746 8316 35756 8372
rect 35812 8316 36428 8372
rect 36484 8316 36764 8372
rect 36820 8316 36830 8372
rect 38994 8316 39004 8372
rect 39060 8316 42252 8372
rect 42308 8316 42318 8372
rect 42466 8316 42476 8372
rect 42532 8316 45500 8372
rect 45556 8316 45566 8372
rect 50306 8316 50316 8372
rect 50372 8316 52220 8372
rect 52276 8316 52286 8372
rect 53330 8316 53340 8372
rect 53396 8316 55580 8372
rect 55636 8316 55646 8372
rect 35532 8260 35588 8316
rect 3154 8204 3164 8260
rect 3220 8204 7756 8260
rect 7812 8204 8652 8260
rect 8708 8204 8718 8260
rect 12114 8204 12124 8260
rect 12180 8204 13020 8260
rect 13076 8204 13580 8260
rect 13636 8204 13646 8260
rect 13794 8204 13804 8260
rect 13860 8204 14532 8260
rect 20290 8204 20300 8260
rect 20356 8204 22316 8260
rect 22372 8204 22382 8260
rect 22530 8204 22540 8260
rect 22596 8204 24220 8260
rect 24276 8204 24286 8260
rect 29474 8204 29484 8260
rect 29540 8204 35308 8260
rect 35364 8204 35374 8260
rect 35532 8204 37996 8260
rect 38052 8204 39340 8260
rect 39396 8204 39406 8260
rect 39554 8204 39564 8260
rect 39620 8204 40516 8260
rect 41010 8204 41020 8260
rect 41076 8204 41468 8260
rect 41524 8204 42140 8260
rect 42196 8204 42206 8260
rect 42914 8204 42924 8260
rect 42980 8204 52556 8260
rect 52612 8204 52622 8260
rect 0 8148 112 8176
rect 14476 8148 14532 8204
rect 40460 8148 40516 8204
rect 57344 8148 57456 8176
rect 0 8092 2604 8148
rect 2660 8092 2670 8148
rect 3490 8092 3500 8148
rect 3556 8092 10108 8148
rect 10164 8092 10174 8148
rect 10332 8092 14084 8148
rect 14466 8092 14476 8148
rect 14532 8092 15148 8148
rect 16146 8092 16156 8148
rect 16212 8092 21308 8148
rect 21364 8092 21374 8148
rect 21746 8092 21756 8148
rect 21812 8092 25004 8148
rect 25060 8092 25070 8148
rect 25228 8092 26236 8148
rect 26292 8092 30044 8148
rect 30100 8092 30110 8148
rect 32386 8092 32396 8148
rect 32452 8092 40236 8148
rect 40292 8092 40302 8148
rect 40460 8092 42588 8148
rect 42644 8092 42654 8148
rect 42914 8092 42924 8148
rect 42980 8092 46844 8148
rect 46900 8092 46910 8148
rect 55906 8092 55916 8148
rect 55972 8092 57456 8148
rect 0 8064 112 8092
rect 10332 8036 10388 8092
rect 242 7980 252 8036
rect 308 7980 4396 8036
rect 4452 7980 4462 8036
rect 6514 7980 6524 8036
rect 6580 7980 10388 8036
rect 12226 7980 12236 8036
rect 12292 7980 12796 8036
rect 12852 7980 12862 8036
rect 14028 7924 14084 8092
rect 15092 8036 15148 8092
rect 25228 8036 25284 8092
rect 57344 8064 57456 8092
rect 15092 7980 20412 8036
rect 20468 7980 20478 8036
rect 20626 7980 20636 8036
rect 20692 7980 24220 8036
rect 24276 7980 24286 8036
rect 24770 7980 24780 8036
rect 24836 7980 25284 8036
rect 25442 7980 25452 8036
rect 25508 7980 28700 8036
rect 28756 7980 28766 8036
rect 35074 7980 35084 8036
rect 35140 7980 36316 8036
rect 36372 7980 37100 8036
rect 37156 7980 37166 8036
rect 37538 7980 37548 8036
rect 37604 7980 54124 8036
rect 54180 7980 54190 8036
rect 6626 7868 6636 7924
rect 6692 7868 13748 7924
rect 14028 7868 21196 7924
rect 21252 7868 21262 7924
rect 21634 7868 21644 7924
rect 21700 7868 22540 7924
rect 22596 7868 22606 7924
rect 24780 7868 29596 7924
rect 29652 7868 29662 7924
rect 32050 7868 32060 7924
rect 32116 7868 33236 7924
rect 34962 7868 34972 7924
rect 35028 7868 40908 7924
rect 40964 7868 40974 7924
rect 41122 7868 41132 7924
rect 41188 7868 43596 7924
rect 43652 7868 43662 7924
rect 52994 7868 53004 7924
rect 53060 7868 57260 7924
rect 57316 7868 57326 7924
rect 3794 7812 3804 7868
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 4068 7812 4078 7868
rect 8316 7756 13468 7812
rect 13524 7756 13534 7812
rect 0 7700 112 7728
rect 8316 7700 8372 7756
rect 13692 7700 13748 7868
rect 23794 7812 23804 7868
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 24068 7812 24078 7868
rect 24780 7812 24836 7868
rect 33180 7812 33236 7868
rect 43794 7812 43804 7868
rect 43860 7812 43908 7868
rect 43964 7812 44012 7868
rect 44068 7812 44078 7868
rect 17042 7756 17052 7812
rect 17108 7756 23660 7812
rect 23716 7756 23726 7812
rect 24220 7756 24836 7812
rect 27122 7756 27132 7812
rect 27188 7756 31724 7812
rect 31780 7756 32956 7812
rect 33012 7756 33022 7812
rect 33180 7756 43260 7812
rect 43316 7756 43326 7812
rect 44156 7756 48076 7812
rect 48132 7756 48142 7812
rect 24220 7700 24276 7756
rect 44156 7700 44212 7756
rect 57344 7700 57456 7728
rect 0 7644 1036 7700
rect 1092 7644 1102 7700
rect 3154 7644 3164 7700
rect 3220 7644 8372 7700
rect 10322 7644 10332 7700
rect 10388 7644 12796 7700
rect 12852 7644 12862 7700
rect 13692 7644 24276 7700
rect 24434 7644 24444 7700
rect 24500 7644 25004 7700
rect 25060 7644 25070 7700
rect 25218 7644 25228 7700
rect 25284 7644 28924 7700
rect 28980 7644 28990 7700
rect 36082 7644 36092 7700
rect 36148 7644 37436 7700
rect 37492 7644 37884 7700
rect 37940 7644 37950 7700
rect 38108 7644 38892 7700
rect 38948 7644 38958 7700
rect 39106 7644 39116 7700
rect 39172 7644 44212 7700
rect 47058 7644 47068 7700
rect 47124 7644 52108 7700
rect 52164 7644 52174 7700
rect 56130 7644 56140 7700
rect 56196 7644 57456 7700
rect 0 7616 112 7644
rect 38108 7588 38164 7644
rect 57344 7616 57456 7644
rect 2370 7532 2380 7588
rect 2436 7532 10556 7588
rect 10612 7532 10622 7588
rect 12450 7532 12460 7588
rect 12516 7532 20188 7588
rect 20244 7532 20254 7588
rect 20972 7532 36540 7588
rect 36596 7532 36606 7588
rect 36978 7532 36988 7588
rect 37044 7532 38164 7588
rect 38770 7532 38780 7588
rect 38836 7532 42588 7588
rect 42644 7532 42654 7588
rect 43250 7532 43260 7588
rect 43316 7532 50092 7588
rect 50148 7532 50158 7588
rect 50530 7532 50540 7588
rect 50596 7532 52444 7588
rect 52500 7532 52510 7588
rect 4162 7420 4172 7476
rect 4228 7420 10332 7476
rect 10388 7420 10398 7476
rect 12002 7420 12012 7476
rect 12068 7420 12572 7476
rect 12628 7420 12638 7476
rect 12786 7420 12796 7476
rect 12852 7420 18732 7476
rect 18788 7420 18798 7476
rect 7858 7308 7868 7364
rect 7924 7308 8316 7364
rect 8372 7308 9324 7364
rect 9380 7308 9548 7364
rect 9604 7308 11452 7364
rect 11508 7308 11518 7364
rect 11666 7308 11676 7364
rect 11732 7308 17612 7364
rect 17668 7308 17678 7364
rect 18274 7308 18284 7364
rect 18340 7308 19740 7364
rect 19796 7308 19806 7364
rect 0 7252 112 7280
rect 20972 7252 21028 7532
rect 21858 7420 21868 7476
rect 21924 7420 29036 7476
rect 29092 7420 29102 7476
rect 29586 7420 29596 7476
rect 29652 7420 31500 7476
rect 31556 7420 31566 7476
rect 34290 7420 34300 7476
rect 34356 7420 36652 7476
rect 36708 7420 36718 7476
rect 36866 7420 36876 7476
rect 36932 7420 39116 7476
rect 39172 7420 39182 7476
rect 39442 7420 39452 7476
rect 39508 7420 43372 7476
rect 43428 7420 43438 7476
rect 43586 7420 43596 7476
rect 43652 7420 48300 7476
rect 48356 7420 48366 7476
rect 49186 7420 49196 7476
rect 49252 7420 50876 7476
rect 50932 7420 50942 7476
rect 21298 7308 21308 7364
rect 21364 7308 21644 7364
rect 21700 7308 21710 7364
rect 21970 7308 21980 7364
rect 22036 7308 26348 7364
rect 26404 7308 26414 7364
rect 28466 7308 28476 7364
rect 28532 7308 28924 7364
rect 28980 7308 38220 7364
rect 38276 7308 38286 7364
rect 38434 7308 38444 7364
rect 38500 7308 39508 7364
rect 39778 7308 39788 7364
rect 39844 7308 40572 7364
rect 40628 7308 40638 7364
rect 40786 7308 40796 7364
rect 40852 7308 41692 7364
rect 41748 7308 41758 7364
rect 42252 7308 51436 7364
rect 51492 7308 51502 7364
rect 39452 7252 39508 7308
rect 42252 7252 42308 7308
rect 57344 7252 57456 7280
rect 0 7196 1036 7252
rect 1092 7196 1102 7252
rect 1586 7196 1596 7252
rect 1652 7196 6188 7252
rect 6244 7196 6254 7252
rect 11442 7196 11452 7252
rect 11508 7196 12796 7252
rect 12852 7196 12862 7252
rect 13122 7196 13132 7252
rect 13188 7196 13468 7252
rect 13524 7196 21028 7252
rect 21186 7196 21196 7252
rect 21252 7196 25340 7252
rect 25396 7196 25406 7252
rect 25666 7196 25676 7252
rect 25732 7196 26460 7252
rect 26516 7196 26526 7252
rect 26852 7196 29260 7252
rect 29316 7196 29326 7252
rect 29484 7196 30940 7252
rect 30996 7196 31006 7252
rect 31154 7196 31164 7252
rect 31220 7196 33964 7252
rect 34020 7196 34030 7252
rect 35084 7196 39116 7252
rect 39172 7196 39182 7252
rect 39452 7196 39900 7252
rect 39956 7196 39966 7252
rect 40114 7196 40124 7252
rect 40180 7196 42308 7252
rect 43474 7196 43484 7252
rect 43540 7196 52108 7252
rect 52164 7196 52174 7252
rect 54562 7196 54572 7252
rect 54628 7196 57456 7252
rect 0 7168 112 7196
rect 26852 7140 26908 7196
rect 6626 7084 6636 7140
rect 6692 7084 21644 7140
rect 21700 7084 21710 7140
rect 22194 7084 22204 7140
rect 22260 7084 24220 7140
rect 24276 7084 24286 7140
rect 24882 7084 24892 7140
rect 24948 7084 26908 7140
rect 4454 7028 4464 7084
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4728 7028 4738 7084
rect 24454 7028 24464 7084
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 24728 7028 24738 7084
rect 29484 7028 29540 7196
rect 35084 7140 35140 7196
rect 57344 7168 57456 7196
rect 29698 7084 29708 7140
rect 29764 7084 35140 7140
rect 35298 7084 35308 7140
rect 35364 7084 37660 7140
rect 37716 7084 37726 7140
rect 37874 7084 37884 7140
rect 37940 7084 39452 7140
rect 39508 7084 39518 7140
rect 39666 7084 39676 7140
rect 39732 7084 41804 7140
rect 41860 7084 41870 7140
rect 42018 7084 42028 7140
rect 42084 7084 43036 7140
rect 43092 7084 43708 7140
rect 43764 7084 43774 7140
rect 45714 7084 45724 7140
rect 45780 7084 55356 7140
rect 55412 7084 55422 7140
rect 44454 7028 44464 7084
rect 44520 7028 44568 7084
rect 44624 7028 44672 7084
rect 44728 7028 44738 7084
rect 10434 6972 10444 7028
rect 10500 6972 17052 7028
rect 17108 6972 17118 7028
rect 17266 6972 17276 7028
rect 17332 6972 24388 7028
rect 24332 6916 24388 6972
rect 24892 6972 29540 7028
rect 30146 6972 30156 7028
rect 30212 6972 33852 7028
rect 33908 6972 33918 7028
rect 34738 6972 34748 7028
rect 34804 6972 40236 7028
rect 40292 6972 40302 7028
rect 40450 6972 40460 7028
rect 40516 6972 44268 7028
rect 44324 6972 44334 7028
rect 24892 6916 24948 6972
rect 11190 6860 11228 6916
rect 11284 6860 11294 6916
rect 11442 6860 11452 6916
rect 11508 6860 16156 6916
rect 16212 6860 16222 6916
rect 16818 6860 16828 6916
rect 16884 6860 23436 6916
rect 23492 6860 23502 6916
rect 23650 6860 23660 6916
rect 23716 6860 24108 6916
rect 24164 6860 24174 6916
rect 24332 6860 24948 6916
rect 25330 6860 25340 6916
rect 25396 6860 40236 6916
rect 40292 6860 40302 6916
rect 41234 6860 41244 6916
rect 41300 6860 45836 6916
rect 45892 6860 45902 6916
rect 46610 6860 46620 6916
rect 46676 6860 49868 6916
rect 49924 6860 49934 6916
rect 50082 6860 50092 6916
rect 50148 6860 50988 6916
rect 51044 6860 51054 6916
rect 0 6804 112 6832
rect 57344 6804 57456 6832
rect 0 6748 1820 6804
rect 1876 6748 1886 6804
rect 9874 6748 9884 6804
rect 9940 6748 10556 6804
rect 10612 6748 12236 6804
rect 12292 6748 12302 6804
rect 18386 6748 18396 6804
rect 18452 6748 18844 6804
rect 18900 6748 18910 6804
rect 20972 6748 30828 6804
rect 30884 6748 30894 6804
rect 31602 6748 31612 6804
rect 31668 6748 32620 6804
rect 32676 6748 32686 6804
rect 33394 6748 33404 6804
rect 33460 6748 34972 6804
rect 35028 6748 35038 6804
rect 35186 6748 35196 6804
rect 35252 6748 38444 6804
rect 38500 6748 38510 6804
rect 38882 6748 38892 6804
rect 38948 6748 39620 6804
rect 39890 6748 39900 6804
rect 39956 6748 41132 6804
rect 41188 6748 41198 6804
rect 42354 6748 42364 6804
rect 42420 6748 50428 6804
rect 56130 6748 56140 6804
rect 56196 6748 57456 6804
rect 0 6720 112 6748
rect 20972 6692 21028 6748
rect 39564 6692 39620 6748
rect 50372 6692 50428 6748
rect 57344 6720 57456 6748
rect 2482 6636 2492 6692
rect 2548 6636 9268 6692
rect 9426 6636 9436 6692
rect 9492 6636 10892 6692
rect 10948 6636 10958 6692
rect 11106 6636 11116 6692
rect 11172 6636 11788 6692
rect 11844 6636 11854 6692
rect 15092 6636 21028 6692
rect 22390 6636 22428 6692
rect 22484 6636 22494 6692
rect 23538 6636 23548 6692
rect 23604 6636 24332 6692
rect 24388 6636 24398 6692
rect 24770 6636 24780 6692
rect 24836 6636 25788 6692
rect 25844 6636 25854 6692
rect 26338 6636 26348 6692
rect 26404 6636 27692 6692
rect 27748 6636 29148 6692
rect 29204 6636 29214 6692
rect 29810 6636 29820 6692
rect 29876 6636 31276 6692
rect 31332 6636 31342 6692
rect 31490 6636 31500 6692
rect 31556 6636 35196 6692
rect 35252 6636 35262 6692
rect 36978 6636 36988 6692
rect 37044 6636 38332 6692
rect 38388 6636 38398 6692
rect 39564 6636 40460 6692
rect 40516 6636 40526 6692
rect 41346 6636 41356 6692
rect 41412 6636 42812 6692
rect 42868 6636 42878 6692
rect 43036 6636 43540 6692
rect 50372 6636 50540 6692
rect 50596 6636 50606 6692
rect 51090 6636 51100 6692
rect 51156 6636 52892 6692
rect 52948 6636 52958 6692
rect 9212 6580 9268 6636
rect 15092 6580 15148 6636
rect 43036 6580 43092 6636
rect 1362 6524 1372 6580
rect 1428 6524 3388 6580
rect 9212 6524 15148 6580
rect 18386 6524 18396 6580
rect 18452 6524 18620 6580
rect 18676 6524 18686 6580
rect 19842 6524 19852 6580
rect 19908 6524 20748 6580
rect 20804 6524 20814 6580
rect 22082 6524 22092 6580
rect 22148 6524 25340 6580
rect 25396 6524 25406 6580
rect 26226 6524 26236 6580
rect 26292 6524 27020 6580
rect 27076 6524 37212 6580
rect 37268 6524 37278 6580
rect 37762 6524 37772 6580
rect 37828 6524 40068 6580
rect 40226 6524 40236 6580
rect 40292 6524 43092 6580
rect 3332 6468 3388 6524
rect 40012 6468 40068 6524
rect 43484 6468 43540 6636
rect 43820 6524 47068 6580
rect 47124 6524 47134 6580
rect 47282 6524 47292 6580
rect 47348 6524 53228 6580
rect 53284 6524 53294 6580
rect 53554 6524 53564 6580
rect 53620 6524 53900 6580
rect 53956 6524 53966 6580
rect 43820 6468 43876 6524
rect 3332 6412 11228 6468
rect 11284 6412 11294 6468
rect 12674 6412 12684 6468
rect 12740 6412 17388 6468
rect 17444 6412 17454 6468
rect 17602 6412 17612 6468
rect 17668 6412 21196 6468
rect 21252 6412 21262 6468
rect 21970 6412 21980 6468
rect 22036 6412 28812 6468
rect 28868 6412 28878 6468
rect 29026 6412 29036 6468
rect 29092 6412 34860 6468
rect 34916 6412 34926 6468
rect 35074 6412 35084 6468
rect 35140 6412 38668 6468
rect 40012 6412 41468 6468
rect 41524 6412 42252 6468
rect 42308 6412 43148 6468
rect 43204 6412 43214 6468
rect 43484 6412 43876 6468
rect 44156 6412 55244 6468
rect 55300 6412 55310 6468
rect 0 6356 112 6384
rect 38612 6356 38668 6412
rect 0 6300 1036 6356
rect 1092 6300 1102 6356
rect 10098 6300 10108 6356
rect 10164 6300 16716 6356
rect 16772 6300 16782 6356
rect 19170 6300 19180 6356
rect 19236 6300 22652 6356
rect 22708 6300 22718 6356
rect 22978 6300 22988 6356
rect 23044 6300 23660 6356
rect 23716 6300 23726 6356
rect 24210 6300 24220 6356
rect 24276 6300 25452 6356
rect 25508 6300 25518 6356
rect 26450 6300 26460 6356
rect 26516 6300 28252 6356
rect 28308 6300 28318 6356
rect 28466 6300 28476 6356
rect 28532 6300 30380 6356
rect 30436 6300 30446 6356
rect 30594 6300 30604 6356
rect 30660 6300 35644 6356
rect 35700 6300 35710 6356
rect 38612 6300 42924 6356
rect 42980 6300 42990 6356
rect 0 6272 112 6300
rect 3794 6244 3804 6300
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 4068 6244 4078 6300
rect 23794 6244 23804 6300
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 24068 6244 24078 6300
rect 43794 6244 43804 6300
rect 43860 6244 43908 6300
rect 43964 6244 44012 6300
rect 44068 6244 44078 6300
rect 5058 6188 5068 6244
rect 5124 6188 13356 6244
rect 13412 6188 13422 6244
rect 18386 6188 18396 6244
rect 18452 6188 23548 6244
rect 23604 6188 23614 6244
rect 24882 6188 24892 6244
rect 24948 6188 26012 6244
rect 26068 6188 26078 6244
rect 26338 6188 26348 6244
rect 26404 6188 28476 6244
rect 28532 6188 28542 6244
rect 28690 6188 28700 6244
rect 28756 6188 31948 6244
rect 32004 6188 33628 6244
rect 33684 6188 33694 6244
rect 37202 6188 37212 6244
rect 37268 6188 37884 6244
rect 37940 6188 37950 6244
rect 38770 6188 38780 6244
rect 38836 6188 43596 6244
rect 43652 6188 43662 6244
rect 44156 6132 44212 6412
rect 57344 6356 57456 6384
rect 44370 6300 44380 6356
rect 44436 6300 48636 6356
rect 48692 6300 48702 6356
rect 55122 6300 55132 6356
rect 55188 6300 57456 6356
rect 57344 6272 57456 6300
rect 45938 6188 45948 6244
rect 46004 6188 47292 6244
rect 47348 6188 47358 6244
rect 52994 6188 53004 6244
rect 53060 6188 56700 6244
rect 56756 6188 56766 6244
rect 1922 6076 1932 6132
rect 1988 6076 1998 6132
rect 8194 6076 8204 6132
rect 8260 6076 12740 6132
rect 13346 6076 13356 6132
rect 13412 6076 14028 6132
rect 14084 6076 30156 6132
rect 30212 6076 30222 6132
rect 31826 6076 31836 6132
rect 31892 6076 32620 6132
rect 32676 6076 32686 6132
rect 34514 6076 34524 6132
rect 34580 6076 44212 6132
rect 44370 6076 44380 6132
rect 44436 6076 44828 6132
rect 44884 6076 44894 6132
rect 45276 6076 53452 6132
rect 53508 6076 53518 6132
rect 0 5908 112 5936
rect 1932 5908 1988 6076
rect 7298 5964 7308 6020
rect 7364 5964 12460 6020
rect 12516 5964 12526 6020
rect 12684 5908 12740 6076
rect 17490 5964 17500 6020
rect 17556 5964 22428 6020
rect 22484 5964 22494 6020
rect 23426 5964 23436 6020
rect 23492 5964 35308 6020
rect 35364 5964 35374 6020
rect 35522 5964 35532 6020
rect 35588 5964 41804 6020
rect 41860 5964 41870 6020
rect 42466 5964 42476 6020
rect 42532 5964 45052 6020
rect 45108 5964 45118 6020
rect 45276 5908 45332 6076
rect 48290 5964 48300 6020
rect 48356 5964 49420 6020
rect 49476 5964 49486 6020
rect 57344 5908 57456 5936
rect 0 5852 1988 5908
rect 3266 5852 3276 5908
rect 3332 5852 6748 5908
rect 6804 5852 8204 5908
rect 8260 5852 8270 5908
rect 10882 5852 10892 5908
rect 10948 5852 11676 5908
rect 11732 5852 11742 5908
rect 12684 5852 20524 5908
rect 20580 5852 20590 5908
rect 20850 5852 20860 5908
rect 20916 5852 22204 5908
rect 22260 5852 22270 5908
rect 22428 5852 24892 5908
rect 24948 5852 24958 5908
rect 25106 5852 25116 5908
rect 25172 5852 42588 5908
rect 42644 5852 42654 5908
rect 43362 5852 43372 5908
rect 43428 5852 45332 5908
rect 46834 5852 46844 5908
rect 46900 5852 48972 5908
rect 49028 5852 49038 5908
rect 54562 5852 54572 5908
rect 54628 5852 57456 5908
rect 0 5824 112 5852
rect 22428 5796 22484 5852
rect 57344 5824 57456 5852
rect 3042 5740 3052 5796
rect 3108 5740 11564 5796
rect 11620 5740 11630 5796
rect 20290 5740 20300 5796
rect 20356 5740 22484 5796
rect 22642 5740 22652 5796
rect 22708 5740 26796 5796
rect 26852 5740 26862 5796
rect 27794 5740 27804 5796
rect 27860 5740 29036 5796
rect 29092 5740 29102 5796
rect 29250 5740 29260 5796
rect 29316 5740 31948 5796
rect 32050 5740 32060 5796
rect 32116 5740 33180 5796
rect 33236 5740 33246 5796
rect 36642 5740 36652 5796
rect 36708 5740 44268 5796
rect 44324 5740 44334 5796
rect 44492 5740 54124 5796
rect 54180 5740 54190 5796
rect 31892 5684 31948 5740
rect 44492 5684 44548 5740
rect 3378 5628 3388 5684
rect 3444 5628 21532 5684
rect 21588 5628 21598 5684
rect 22082 5628 22092 5684
rect 22148 5628 24668 5684
rect 24724 5628 25004 5684
rect 25060 5628 25070 5684
rect 25218 5628 25228 5684
rect 25284 5628 30492 5684
rect 30548 5628 30558 5684
rect 31892 5628 38668 5684
rect 38724 5628 38734 5684
rect 40002 5628 40012 5684
rect 40068 5628 44548 5684
rect 44706 5628 44716 5684
rect 44772 5628 52556 5684
rect 52612 5628 52622 5684
rect 5170 5516 5180 5572
rect 5236 5516 5740 5572
rect 5796 5516 5806 5572
rect 12450 5516 12460 5572
rect 12516 5516 13244 5572
rect 13300 5516 13310 5572
rect 15586 5516 15596 5572
rect 15652 5516 23212 5572
rect 23268 5516 23278 5572
rect 25330 5516 25340 5572
rect 25396 5516 26796 5572
rect 26852 5516 26862 5572
rect 28354 5516 28364 5572
rect 28420 5516 30156 5572
rect 30212 5516 30222 5572
rect 30594 5516 30604 5572
rect 30660 5516 40124 5572
rect 40180 5516 40190 5572
rect 44818 5516 44828 5572
rect 44884 5516 47404 5572
rect 47460 5516 47470 5572
rect 0 5460 112 5488
rect 4454 5460 4464 5516
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4728 5460 4738 5516
rect 24454 5460 24464 5516
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24728 5460 24738 5516
rect 44454 5460 44464 5516
rect 44520 5460 44568 5516
rect 44624 5460 44672 5516
rect 44728 5460 44738 5516
rect 57344 5460 57456 5488
rect 0 5404 3164 5460
rect 3220 5404 3230 5460
rect 12898 5404 12908 5460
rect 12964 5404 21028 5460
rect 21522 5404 21532 5460
rect 21588 5404 24332 5460
rect 24388 5404 24398 5460
rect 25218 5404 25228 5460
rect 25284 5404 27244 5460
rect 27300 5404 27310 5460
rect 28690 5404 28700 5460
rect 28756 5404 31164 5460
rect 31220 5404 31230 5460
rect 31490 5404 31500 5460
rect 31556 5404 44324 5460
rect 56130 5404 56140 5460
rect 56196 5404 57456 5460
rect 0 5376 112 5404
rect 20972 5348 21028 5404
rect 44268 5348 44324 5404
rect 57344 5376 57456 5404
rect 2482 5292 2492 5348
rect 2548 5292 16604 5348
rect 16660 5292 16670 5348
rect 20972 5292 30156 5348
rect 30212 5292 30222 5348
rect 30482 5292 30492 5348
rect 30548 5292 31892 5348
rect 31948 5292 31958 5348
rect 32050 5292 32060 5348
rect 32116 5292 36988 5348
rect 37044 5292 37054 5348
rect 37202 5292 37212 5348
rect 37268 5292 42364 5348
rect 42420 5292 42430 5348
rect 44268 5292 55132 5348
rect 55188 5292 55198 5348
rect 10882 5180 10892 5236
rect 10948 5180 11900 5236
rect 11956 5180 11966 5236
rect 12114 5180 12124 5236
rect 12180 5180 13468 5236
rect 13524 5180 13534 5236
rect 20402 5180 20412 5236
rect 20468 5180 26572 5236
rect 26628 5180 26638 5236
rect 26786 5180 26796 5236
rect 26852 5180 29708 5236
rect 29764 5180 29774 5236
rect 30370 5180 30380 5236
rect 30436 5180 40460 5236
rect 40516 5180 40526 5236
rect 41906 5180 41916 5236
rect 41972 5180 44492 5236
rect 44548 5180 44558 5236
rect 45154 5180 45164 5236
rect 45220 5180 52108 5236
rect 52164 5180 52174 5236
rect 6178 5068 6188 5124
rect 6244 5068 6748 5124
rect 6804 5068 6814 5124
rect 12226 5068 12236 5124
rect 12292 5068 14140 5124
rect 14196 5068 14206 5124
rect 14364 5068 21644 5124
rect 21700 5068 21710 5124
rect 21858 5068 21868 5124
rect 21924 5068 22316 5124
rect 22372 5068 22382 5124
rect 22530 5068 22540 5124
rect 22596 5068 25228 5124
rect 25284 5068 25294 5124
rect 26908 5068 32172 5124
rect 32228 5068 32238 5124
rect 35252 5068 43484 5124
rect 43540 5068 43550 5124
rect 43698 5068 43708 5124
rect 43764 5068 45556 5124
rect 50082 5068 50092 5124
rect 50148 5068 51884 5124
rect 51940 5068 51950 5124
rect 54898 5068 54908 5124
rect 54964 5068 55468 5124
rect 0 5012 112 5040
rect 0 4956 5180 5012
rect 5236 4956 5246 5012
rect 5964 4956 6636 5012
rect 6692 4956 6702 5012
rect 11890 4956 11900 5012
rect 11956 4956 12348 5012
rect 12404 4956 12414 5012
rect 0 4928 112 4956
rect 5964 4900 6020 4956
rect 14364 4900 14420 5068
rect 26908 5012 26964 5068
rect 35252 5012 35308 5068
rect 45500 5012 45556 5068
rect 55412 5012 55468 5068
rect 57344 5012 57456 5040
rect 14690 4956 14700 5012
rect 14756 4956 15708 5012
rect 15764 4956 15774 5012
rect 16146 4956 16156 5012
rect 16212 4956 26964 5012
rect 29474 4956 29484 5012
rect 29540 4956 31892 5012
rect 31948 4956 31958 5012
rect 32050 4956 32060 5012
rect 32116 4956 32284 5012
rect 32340 4956 32350 5012
rect 34962 4956 34972 5012
rect 35028 4956 35308 5012
rect 37090 4956 37100 5012
rect 37156 4956 38220 5012
rect 38276 4956 38668 5012
rect 38724 4956 38734 5012
rect 42130 4956 42140 5012
rect 42196 4956 45276 5012
rect 45332 4956 45342 5012
rect 45500 4956 47180 5012
rect 47236 4956 47246 5012
rect 47394 4956 47404 5012
rect 47460 4956 53676 5012
rect 53732 4956 53742 5012
rect 55412 4956 57456 5012
rect 57344 4928 57456 4956
rect 1698 4844 1708 4900
rect 1764 4844 6020 4900
rect 6178 4844 6188 4900
rect 6244 4844 14420 4900
rect 17378 4844 17388 4900
rect 17444 4844 21868 4900
rect 21924 4844 21934 4900
rect 22764 4844 26684 4900
rect 26740 4844 26750 4900
rect 26898 4844 26908 4900
rect 26964 4844 35196 4900
rect 35252 4844 35262 4900
rect 35746 4844 35756 4900
rect 35812 4844 38108 4900
rect 38164 4844 39564 4900
rect 39620 4844 39630 4900
rect 40226 4844 40236 4900
rect 40292 4844 46284 4900
rect 46340 4844 46350 4900
rect 52322 4844 52332 4900
rect 52388 4844 54124 4900
rect 54180 4844 54190 4900
rect 12562 4732 12572 4788
rect 12628 4732 18956 4788
rect 19012 4732 19022 4788
rect 20066 4732 20076 4788
rect 20132 4732 22540 4788
rect 22596 4732 22606 4788
rect 3794 4676 3804 4732
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 4068 4676 4078 4732
rect 22764 4676 22820 4844
rect 24210 4732 24220 4788
rect 24276 4732 25788 4788
rect 25844 4732 25854 4788
rect 26002 4732 26012 4788
rect 26068 4732 32060 4788
rect 32116 4732 32126 4788
rect 32274 4732 32284 4788
rect 32340 4732 37996 4788
rect 38052 4732 38062 4788
rect 38210 4732 38220 4788
rect 38276 4732 41132 4788
rect 41188 4732 41198 4788
rect 41458 4732 41468 4788
rect 41524 4732 43484 4788
rect 43540 4732 43550 4788
rect 44146 4732 44156 4788
rect 44212 4732 48524 4788
rect 48580 4732 48590 4788
rect 23794 4676 23804 4732
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 24068 4676 24078 4732
rect 43794 4676 43804 4732
rect 43860 4676 43908 4732
rect 43964 4676 44012 4732
rect 44068 4676 44078 4732
rect 6402 4620 6412 4676
rect 6468 4620 13468 4676
rect 13524 4620 13534 4676
rect 13682 4620 13692 4676
rect 13748 4620 16828 4676
rect 16884 4620 16894 4676
rect 18284 4620 21532 4676
rect 21588 4620 21598 4676
rect 21746 4620 21756 4676
rect 21812 4620 22820 4676
rect 24322 4620 24332 4676
rect 24388 4620 26348 4676
rect 26404 4620 26414 4676
rect 26562 4620 26572 4676
rect 26628 4620 30044 4676
rect 30100 4620 30110 4676
rect 30482 4620 30492 4676
rect 30548 4620 42252 4676
rect 42308 4620 42318 4676
rect 46498 4620 46508 4676
rect 46564 4620 52556 4676
rect 52612 4620 52622 4676
rect 0 4564 112 4592
rect 0 4508 2268 4564
rect 2324 4508 2334 4564
rect 2482 4508 2492 4564
rect 2548 4508 6524 4564
rect 6580 4508 6590 4564
rect 6738 4508 6748 4564
rect 6804 4508 15148 4564
rect 15204 4508 15214 4564
rect 0 4480 112 4508
rect 18284 4452 18340 4620
rect 57344 4564 57456 4592
rect 20178 4508 20188 4564
rect 20244 4508 25340 4564
rect 25396 4508 25406 4564
rect 25564 4508 29932 4564
rect 29988 4508 29998 4564
rect 30146 4508 30156 4564
rect 30212 4508 36876 4564
rect 36932 4508 36942 4564
rect 37100 4508 44828 4564
rect 44884 4508 44894 4564
rect 45276 4508 53564 4564
rect 53620 4508 53630 4564
rect 54562 4508 54572 4564
rect 54628 4508 57456 4564
rect 6290 4396 6300 4452
rect 6356 4396 18340 4452
rect 18722 4396 18732 4452
rect 18788 4396 20076 4452
rect 20132 4396 20142 4452
rect 20962 4396 20972 4452
rect 21028 4396 24220 4452
rect 24276 4396 24286 4452
rect 25564 4340 25620 4508
rect 37100 4452 37156 4508
rect 45276 4452 45332 4508
rect 57344 4480 57456 4508
rect 25778 4396 25788 4452
rect 25844 4396 32060 4452
rect 32116 4396 32126 4452
rect 35298 4396 35308 4452
rect 35364 4396 37156 4452
rect 37874 4396 37884 4452
rect 37940 4396 41468 4452
rect 41524 4396 41534 4452
rect 41682 4396 41692 4452
rect 41748 4396 45332 4452
rect 45490 4396 45500 4452
rect 45556 4396 53116 4452
rect 53172 4396 53182 4452
rect 2594 4284 2604 4340
rect 2660 4284 6076 4340
rect 6132 4284 6142 4340
rect 15810 4284 15820 4340
rect 15876 4284 22092 4340
rect 22148 4284 22158 4340
rect 22390 4284 22428 4340
rect 22484 4284 22494 4340
rect 23650 4284 23660 4340
rect 23716 4284 25620 4340
rect 26674 4284 26684 4340
rect 26740 4284 27580 4340
rect 27636 4284 27646 4340
rect 27804 4284 45052 4340
rect 45108 4284 45118 4340
rect 46162 4284 46172 4340
rect 46228 4284 50428 4340
rect 52322 4284 52332 4340
rect 52388 4284 54236 4340
rect 54292 4284 54302 4340
rect 27804 4228 27860 4284
rect 50372 4228 50428 4284
rect 5282 4172 5292 4228
rect 5348 4172 9772 4228
rect 9828 4172 9838 4228
rect 10322 4172 10332 4228
rect 10388 4172 20972 4228
rect 21028 4172 21038 4228
rect 21186 4172 21196 4228
rect 21252 4172 25116 4228
rect 25172 4172 25182 4228
rect 25778 4172 25788 4228
rect 25844 4172 27860 4228
rect 29026 4172 29036 4228
rect 29092 4172 37828 4228
rect 37986 4172 37996 4228
rect 38052 4172 38780 4228
rect 38836 4172 38846 4228
rect 38994 4172 39004 4228
rect 39060 4172 48076 4228
rect 48132 4172 48142 4228
rect 50372 4172 52668 4228
rect 52724 4172 52734 4228
rect 0 4116 112 4144
rect 37772 4116 37828 4172
rect 57344 4116 57456 4144
rect 0 4060 812 4116
rect 868 4060 878 4116
rect 1474 4060 1484 4116
rect 1540 4060 15148 4116
rect 15250 4060 15260 4116
rect 15316 4060 18732 4116
rect 18788 4060 18798 4116
rect 18946 4060 18956 4116
rect 19012 4060 27188 4116
rect 27346 4060 27356 4116
rect 27412 4060 28588 4116
rect 28644 4060 30380 4116
rect 30436 4060 30446 4116
rect 30604 4060 32396 4116
rect 32452 4060 32462 4116
rect 34514 4060 34524 4116
rect 34580 4060 37436 4116
rect 37492 4060 37502 4116
rect 37772 4060 43372 4116
rect 43428 4060 43438 4116
rect 44258 4060 44268 4116
rect 44324 4060 55132 4116
rect 55188 4060 55198 4116
rect 56130 4060 56140 4116
rect 56196 4060 57456 4116
rect 0 4032 112 4060
rect 15092 4004 15148 4060
rect 27132 4004 27188 4060
rect 30604 4004 30660 4060
rect 57344 4032 57456 4060
rect 15092 3948 21756 4004
rect 21812 3948 21822 4004
rect 24882 3948 24892 4004
rect 24948 3948 25452 4004
rect 25508 3948 25518 4004
rect 27132 3948 30660 4004
rect 30818 3948 30828 4004
rect 30884 3948 34412 4004
rect 34468 3948 34478 4004
rect 35298 3948 35308 4004
rect 35364 3948 39116 4004
rect 39172 3948 39182 4004
rect 39666 3948 39676 4004
rect 39732 3948 44044 4004
rect 44100 3948 44110 4004
rect 4454 3892 4464 3948
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4728 3892 4738 3948
rect 24454 3892 24464 3948
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24728 3892 24738 3948
rect 44454 3892 44464 3948
rect 44520 3892 44568 3948
rect 44624 3892 44672 3948
rect 44728 3892 44738 3948
rect 7970 3836 7980 3892
rect 8036 3836 15820 3892
rect 15876 3836 15886 3892
rect 16034 3836 16044 3892
rect 16100 3836 19180 3892
rect 19236 3836 19246 3892
rect 20178 3836 20188 3892
rect 20244 3836 21644 3892
rect 21700 3836 21710 3892
rect 24892 3836 30604 3892
rect 30660 3836 30670 3892
rect 30930 3836 30940 3892
rect 30996 3836 34860 3892
rect 34916 3836 34926 3892
rect 35074 3836 35084 3892
rect 35140 3836 37044 3892
rect 37202 3836 37212 3892
rect 37268 3836 43260 3892
rect 43316 3836 43326 3892
rect 24892 3780 24948 3836
rect 1586 3724 1596 3780
rect 1652 3724 18788 3780
rect 19058 3724 19068 3780
rect 19124 3724 19628 3780
rect 19684 3724 24948 3780
rect 25330 3724 25340 3780
rect 25396 3724 29596 3780
rect 29652 3724 29662 3780
rect 30258 3724 30268 3780
rect 30324 3724 36932 3780
rect 0 3668 112 3696
rect 18732 3668 18788 3724
rect 0 3612 1652 3668
rect 13346 3612 13356 3668
rect 13412 3612 15036 3668
rect 15092 3612 15102 3668
rect 15250 3612 15260 3668
rect 15316 3612 17948 3668
rect 18004 3612 18014 3668
rect 18732 3612 28028 3668
rect 28084 3612 28094 3668
rect 28802 3612 28812 3668
rect 28868 3612 35196 3668
rect 35252 3612 35262 3668
rect 0 3584 112 3612
rect 1596 3332 1652 3612
rect 5058 3500 5068 3556
rect 5124 3500 5180 3556
rect 5236 3500 5246 3556
rect 14242 3500 14252 3556
rect 14308 3500 18172 3556
rect 18228 3500 18238 3556
rect 20066 3500 20076 3556
rect 20132 3500 21196 3556
rect 21252 3500 21262 3556
rect 21420 3500 21980 3556
rect 22036 3500 22046 3556
rect 23314 3500 23324 3556
rect 23380 3500 29820 3556
rect 29876 3500 29886 3556
rect 30258 3500 30268 3556
rect 30324 3500 36652 3556
rect 36708 3500 36718 3556
rect 21420 3444 21476 3500
rect 36876 3444 36932 3724
rect 36988 3668 37044 3836
rect 40338 3724 40348 3780
rect 40404 3724 44548 3780
rect 44818 3724 44828 3780
rect 44884 3724 54124 3780
rect 54180 3724 54190 3780
rect 44492 3668 44548 3724
rect 57344 3668 57456 3696
rect 36988 3612 44268 3668
rect 44324 3612 44334 3668
rect 44492 3612 50428 3668
rect 50484 3612 50494 3668
rect 54898 3612 54908 3668
rect 54964 3612 57456 3668
rect 57344 3584 57456 3612
rect 37650 3500 37660 3556
rect 37716 3500 41860 3556
rect 42018 3500 42028 3556
rect 42084 3500 47852 3556
rect 47908 3500 47918 3556
rect 48066 3500 48076 3556
rect 48132 3500 52220 3556
rect 52276 3500 52286 3556
rect 41804 3444 41860 3500
rect 5618 3388 5628 3444
rect 5684 3388 8428 3444
rect 9538 3388 9548 3444
rect 9604 3388 13524 3444
rect 15698 3388 15708 3444
rect 15764 3388 16884 3444
rect 18274 3388 18284 3444
rect 18340 3388 21476 3444
rect 21858 3388 21868 3444
rect 21924 3388 22652 3444
rect 22708 3388 22718 3444
rect 22866 3388 22876 3444
rect 22932 3388 28812 3444
rect 28868 3388 28878 3444
rect 29138 3388 29148 3444
rect 29204 3388 30828 3444
rect 30884 3388 30894 3444
rect 31892 3388 35532 3444
rect 35588 3388 35598 3444
rect 36876 3388 38724 3444
rect 41804 3388 45444 3444
rect 53554 3388 53564 3444
rect 53620 3388 57036 3444
rect 57092 3388 57102 3444
rect 8372 3332 8428 3388
rect 1596 3276 5068 3332
rect 5124 3276 5134 3332
rect 8372 3276 13244 3332
rect 13300 3276 13310 3332
rect 0 3220 112 3248
rect 13468 3220 13524 3388
rect 16828 3332 16884 3388
rect 31892 3332 31948 3388
rect 38668 3332 38724 3388
rect 45388 3332 45444 3388
rect 16828 3276 20188 3332
rect 21858 3276 21868 3332
rect 21924 3276 26012 3332
rect 26068 3276 26078 3332
rect 27458 3276 27468 3332
rect 27524 3276 28588 3332
rect 28644 3276 28654 3332
rect 29138 3276 29148 3332
rect 29204 3276 31948 3332
rect 35298 3276 35308 3332
rect 35364 3276 36204 3332
rect 36260 3276 36270 3332
rect 38668 3276 45164 3332
rect 45220 3276 45230 3332
rect 45388 3276 50652 3332
rect 50708 3276 50718 3332
rect 51314 3276 51324 3332
rect 51380 3276 52780 3332
rect 52836 3276 52846 3332
rect 20132 3220 20188 3276
rect 57344 3220 57456 3248
rect 0 3164 1372 3220
rect 1428 3164 1438 3220
rect 9090 3164 9100 3220
rect 9156 3164 10164 3220
rect 13468 3164 18396 3220
rect 18452 3164 18462 3220
rect 20132 3164 23100 3220
rect 23156 3164 23166 3220
rect 24322 3164 24332 3220
rect 24388 3164 27356 3220
rect 27412 3164 27422 3220
rect 27570 3164 27580 3220
rect 27636 3164 30156 3220
rect 30212 3164 30222 3220
rect 30594 3164 30604 3220
rect 30660 3164 33068 3220
rect 33124 3164 33134 3220
rect 33282 3164 33292 3220
rect 33348 3164 42476 3220
rect 42532 3164 42542 3220
rect 48066 3164 48076 3220
rect 48132 3164 52556 3220
rect 52612 3164 52622 3220
rect 54562 3164 54572 3220
rect 54628 3164 57456 3220
rect 0 3136 112 3164
rect 3794 3108 3804 3164
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 4068 3108 4078 3164
rect 10108 3108 10164 3164
rect 23794 3108 23804 3164
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 24068 3108 24078 3164
rect 43794 3108 43804 3164
rect 43860 3108 43908 3164
rect 43964 3108 44012 3164
rect 44068 3108 44078 3164
rect 57344 3136 57456 3164
rect 5730 3052 5740 3108
rect 5796 3052 9884 3108
rect 9940 3052 9950 3108
rect 10108 3052 23716 3108
rect 24210 3052 24220 3108
rect 24276 3052 25228 3108
rect 25284 3052 25294 3108
rect 25442 3052 25452 3108
rect 25508 3052 28140 3108
rect 28196 3052 28206 3108
rect 30034 3052 30044 3108
rect 30100 3052 31332 3108
rect 32050 3052 32060 3108
rect 32116 3052 38332 3108
rect 38388 3052 38398 3108
rect 38612 3052 40348 3108
rect 40404 3052 40414 3108
rect 41570 3052 41580 3108
rect 41636 3052 42700 3108
rect 42756 3052 42766 3108
rect 44818 3052 44828 3108
rect 44884 3052 53564 3108
rect 53620 3052 53630 3108
rect 23660 2996 23716 3052
rect 31276 2996 31332 3052
rect 38612 2996 38668 3052
rect 5170 2940 5180 2996
rect 5236 2940 9660 2996
rect 9716 2940 9726 2996
rect 12898 2940 12908 2996
rect 12964 2940 20636 2996
rect 20692 2940 20702 2996
rect 21970 2940 21980 2996
rect 22036 2940 23212 2996
rect 23268 2940 23278 2996
rect 23660 2940 26012 2996
rect 26068 2940 26078 2996
rect 28914 2940 28924 2996
rect 28980 2940 31052 2996
rect 31108 2940 31118 2996
rect 31276 2940 38668 2996
rect 42018 2940 42028 2996
rect 42084 2940 48748 2996
rect 48804 2940 48814 2996
rect 1250 2828 1260 2884
rect 1316 2828 5180 2884
rect 5236 2828 5246 2884
rect 5842 2828 5852 2884
rect 5908 2828 8428 2884
rect 9090 2828 9100 2884
rect 9156 2828 14140 2884
rect 14196 2828 14206 2884
rect 18162 2828 18172 2884
rect 18228 2828 23436 2884
rect 23492 2828 23502 2884
rect 23986 2828 23996 2884
rect 24052 2828 53340 2884
rect 53396 2828 53406 2884
rect 0 2772 112 2800
rect 8372 2772 8428 2828
rect 57344 2772 57456 2800
rect 0 2716 5404 2772
rect 5460 2716 5470 2772
rect 8372 2716 20132 2772
rect 20738 2716 20748 2772
rect 20804 2716 25956 2772
rect 27682 2716 27692 2772
rect 27748 2716 29260 2772
rect 29316 2716 29326 2772
rect 29810 2716 29820 2772
rect 29876 2716 30156 2772
rect 30212 2716 32844 2772
rect 32900 2716 32910 2772
rect 33058 2716 33068 2772
rect 33124 2716 38668 2772
rect 38724 2716 38734 2772
rect 40562 2716 40572 2772
rect 40628 2716 49028 2772
rect 51202 2716 51212 2772
rect 51268 2716 51996 2772
rect 52052 2716 52062 2772
rect 56130 2716 56140 2772
rect 56196 2716 57456 2772
rect 0 2688 112 2716
rect 20076 2660 20132 2716
rect 25900 2660 25956 2716
rect 48972 2660 49028 2716
rect 57344 2688 57456 2716
rect 6514 2604 6524 2660
rect 6580 2604 12124 2660
rect 12180 2604 12190 2660
rect 12338 2604 12348 2660
rect 12404 2604 14980 2660
rect 17154 2604 17164 2660
rect 17220 2604 19852 2660
rect 19908 2604 19918 2660
rect 20076 2604 20860 2660
rect 20916 2604 20926 2660
rect 21522 2604 21532 2660
rect 21588 2604 25676 2660
rect 25732 2604 25742 2660
rect 25900 2604 29148 2660
rect 29204 2604 29214 2660
rect 30258 2604 30268 2660
rect 30324 2604 33068 2660
rect 33124 2604 33134 2660
rect 33292 2604 40292 2660
rect 40450 2604 40460 2660
rect 40516 2604 48636 2660
rect 48692 2604 48702 2660
rect 48972 2604 52332 2660
rect 52388 2604 52398 2660
rect 52770 2604 52780 2660
rect 52836 2604 56924 2660
rect 56980 2604 56990 2660
rect 8372 2492 14756 2548
rect 8372 2436 8428 2492
rect 6066 2380 6076 2436
rect 6132 2380 8428 2436
rect 10770 2380 10780 2436
rect 10836 2380 12852 2436
rect 0 2324 112 2352
rect 4454 2324 4464 2380
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4728 2324 4738 2380
rect 0 2268 3444 2324
rect 0 2240 112 2268
rect 3388 2212 3444 2268
rect 3388 2156 5292 2212
rect 5348 2156 5358 2212
rect 12796 2100 12852 2380
rect 14700 2212 14756 2492
rect 14924 2324 14980 2604
rect 16930 2492 16940 2548
rect 16996 2492 20076 2548
rect 20132 2492 20142 2548
rect 20738 2492 20748 2548
rect 20804 2492 22764 2548
rect 22820 2492 22830 2548
rect 23426 2492 23436 2548
rect 23492 2492 24948 2548
rect 25554 2492 25564 2548
rect 25620 2492 28476 2548
rect 28532 2492 28542 2548
rect 28802 2492 28812 2548
rect 28868 2492 30604 2548
rect 30660 2492 30670 2548
rect 30930 2492 30940 2548
rect 30996 2492 32508 2548
rect 32564 2492 32574 2548
rect 24892 2436 24948 2492
rect 33292 2436 33348 2604
rect 40236 2548 40292 2604
rect 35634 2492 35644 2548
rect 35700 2492 40012 2548
rect 40068 2492 40078 2548
rect 40236 2492 41916 2548
rect 41972 2492 41982 2548
rect 42242 2492 42252 2548
rect 42308 2492 49868 2548
rect 49924 2492 49934 2548
rect 16818 2380 16828 2436
rect 16884 2380 21756 2436
rect 21812 2380 21822 2436
rect 22530 2380 22540 2436
rect 22596 2380 24332 2436
rect 24388 2380 24398 2436
rect 24892 2380 27804 2436
rect 27860 2380 27870 2436
rect 28018 2380 28028 2436
rect 28084 2380 30772 2436
rect 32274 2380 32284 2436
rect 32340 2380 33348 2436
rect 42242 2380 42252 2436
rect 42308 2380 44268 2436
rect 44324 2380 44334 2436
rect 24454 2324 24464 2380
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24728 2324 24738 2380
rect 30716 2324 30772 2380
rect 44454 2324 44464 2380
rect 44520 2324 44568 2380
rect 44624 2324 44672 2380
rect 44728 2324 44738 2380
rect 57344 2324 57456 2352
rect 14924 2268 24388 2324
rect 26786 2268 26796 2324
rect 26852 2268 30492 2324
rect 30548 2268 30558 2324
rect 30716 2268 34524 2324
rect 34580 2268 34590 2324
rect 54898 2268 54908 2324
rect 54964 2268 57456 2324
rect 24332 2212 24388 2268
rect 57344 2240 57456 2268
rect 14700 2156 24108 2212
rect 24164 2156 24174 2212
rect 24332 2156 36652 2212
rect 36708 2156 36988 2212
rect 37044 2156 37054 2212
rect 4274 2044 4284 2100
rect 4340 2044 12236 2100
rect 12292 2044 12302 2100
rect 12796 2044 26068 2100
rect 26012 1988 26068 2044
rect 26852 2044 27692 2100
rect 27748 2044 27758 2100
rect 29558 2044 29596 2100
rect 29652 2044 29662 2100
rect 29810 2044 29820 2100
rect 29876 2044 33068 2100
rect 33124 2044 33134 2100
rect 39106 2044 39116 2100
rect 39172 2044 51660 2100
rect 51716 2044 51726 2100
rect 51874 2044 51884 2100
rect 51940 2044 52220 2100
rect 52276 2044 52286 2100
rect 26852 1988 26908 2044
rect 8082 1932 8092 1988
rect 8148 1932 21980 1988
rect 22036 1932 22046 1988
rect 22418 1932 22428 1988
rect 22484 1932 23548 1988
rect 23604 1932 25116 1988
rect 25172 1932 25182 1988
rect 26012 1932 26908 1988
rect 27346 1932 27356 1988
rect 27412 1932 31164 1988
rect 31220 1932 31230 1988
rect 31378 1932 31388 1988
rect 31444 1932 34748 1988
rect 34804 1932 34814 1988
rect 38770 1932 38780 1988
rect 38836 1932 42924 1988
rect 42980 1932 42990 1988
rect 0 1876 112 1904
rect 57344 1876 57456 1904
rect 0 1820 9772 1876
rect 9828 1820 9838 1876
rect 13794 1820 13804 1876
rect 13860 1820 20748 1876
rect 20804 1820 20814 1876
rect 21634 1820 21644 1876
rect 21700 1820 25788 1876
rect 25844 1820 25854 1876
rect 26002 1820 26012 1876
rect 26068 1820 51436 1876
rect 51492 1820 51502 1876
rect 53554 1820 53564 1876
rect 53620 1820 57456 1876
rect 0 1792 112 1820
rect 57344 1792 57456 1820
rect 2044 1708 6188 1764
rect 6244 1708 6254 1764
rect 8372 1708 16828 1764
rect 16884 1708 16894 1764
rect 17042 1708 17052 1764
rect 17108 1708 23324 1764
rect 23380 1708 23390 1764
rect 23660 1708 31948 1764
rect 32274 1708 32284 1764
rect 32340 1708 34636 1764
rect 34692 1708 34702 1764
rect 35186 1708 35196 1764
rect 35252 1708 54124 1764
rect 54180 1708 54190 1764
rect 0 1428 112 1456
rect 2044 1428 2100 1708
rect 8372 1652 8428 1708
rect 4946 1596 4956 1652
rect 5012 1596 8428 1652
rect 9986 1596 9996 1652
rect 10052 1596 16492 1652
rect 16548 1596 16558 1652
rect 16706 1596 16716 1652
rect 16772 1596 21644 1652
rect 21700 1596 21710 1652
rect 3794 1540 3804 1596
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 4068 1540 4078 1596
rect 23660 1540 23716 1708
rect 24322 1596 24332 1652
rect 24388 1596 26180 1652
rect 28242 1596 28252 1652
rect 28308 1596 30940 1652
rect 30996 1596 31006 1652
rect 23794 1540 23804 1596
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 24068 1540 24078 1596
rect 15138 1484 15148 1540
rect 15204 1484 23716 1540
rect 26124 1428 26180 1596
rect 26338 1484 26348 1540
rect 26404 1484 30268 1540
rect 30324 1484 30334 1540
rect 0 1372 2100 1428
rect 2258 1372 2268 1428
rect 2324 1372 9548 1428
rect 9604 1372 9614 1428
rect 11554 1372 11564 1428
rect 11620 1372 17052 1428
rect 17108 1372 17118 1428
rect 17266 1372 17276 1428
rect 17332 1372 20412 1428
rect 20468 1372 20478 1428
rect 23538 1372 23548 1428
rect 23604 1372 25900 1428
rect 25956 1372 25966 1428
rect 26124 1372 31724 1428
rect 31780 1372 31790 1428
rect 0 1344 112 1372
rect 31892 1316 31948 1708
rect 33618 1596 33628 1652
rect 33684 1596 36764 1652
rect 36820 1596 36830 1652
rect 45266 1596 45276 1652
rect 45332 1596 49308 1652
rect 49364 1596 49374 1652
rect 43794 1540 43804 1596
rect 43860 1540 43908 1596
rect 43964 1540 44012 1596
rect 44068 1540 44078 1596
rect 32050 1484 32060 1540
rect 32116 1484 33404 1540
rect 33460 1484 33470 1540
rect 35746 1484 35756 1540
rect 35812 1484 42028 1540
rect 42084 1484 42094 1540
rect 45714 1484 45724 1540
rect 45780 1484 51548 1540
rect 51604 1484 51614 1540
rect 57344 1428 57456 1456
rect 33730 1372 33740 1428
rect 33796 1372 35084 1428
rect 35140 1372 35150 1428
rect 38658 1372 38668 1428
rect 38724 1372 44044 1428
rect 44100 1372 44110 1428
rect 44258 1372 44268 1428
rect 44324 1372 52108 1428
rect 52164 1372 52174 1428
rect 53554 1372 53564 1428
rect 53620 1372 57456 1428
rect 57344 1344 57456 1372
rect 4162 1260 4172 1316
rect 4228 1260 9100 1316
rect 9156 1260 9166 1316
rect 14914 1260 14924 1316
rect 14980 1260 21868 1316
rect 21924 1260 21934 1316
rect 22082 1260 22092 1316
rect 22148 1260 29036 1316
rect 29092 1260 29102 1316
rect 31892 1260 50988 1316
rect 51044 1260 51054 1316
rect 5058 1148 5068 1204
rect 5124 1148 16940 1204
rect 16996 1148 17006 1204
rect 21522 1148 21532 1204
rect 21588 1148 26796 1204
rect 26852 1148 26862 1204
rect 31154 1148 31164 1204
rect 31220 1148 35420 1204
rect 35476 1148 35486 1204
rect 35634 1148 35644 1204
rect 35700 1148 55132 1204
rect 55188 1148 55198 1204
rect 13906 1036 13916 1092
rect 13972 1036 25956 1092
rect 26114 1036 26124 1092
rect 26180 1036 48412 1092
rect 48468 1036 48478 1092
rect 48626 1036 48636 1092
rect 48692 1036 55804 1092
rect 55860 1036 55870 1092
rect 0 980 112 1008
rect 25900 980 25956 1036
rect 57344 980 57456 1008
rect 0 924 1260 980
rect 1316 924 1326 980
rect 8372 924 22876 980
rect 22932 924 22942 980
rect 23202 924 23212 980
rect 23268 924 25060 980
rect 25900 924 30548 980
rect 30706 924 30716 980
rect 30772 924 35644 980
rect 35700 924 35710 980
rect 36978 924 36988 980
rect 37044 924 49756 980
rect 49812 924 49822 980
rect 51986 924 51996 980
rect 52052 924 57456 980
rect 0 896 112 924
rect 8372 868 8428 924
rect 25004 868 25060 924
rect 30492 868 30548 924
rect 57344 896 57456 924
rect 8082 812 8092 868
rect 8148 812 8428 868
rect 9650 812 9660 868
rect 9716 812 17164 868
rect 17220 812 17230 868
rect 22642 812 22652 868
rect 22708 812 24332 868
rect 24388 812 24398 868
rect 25004 812 29820 868
rect 29876 812 29886 868
rect 30492 812 33740 868
rect 33796 812 33806 868
rect 34850 812 34860 868
rect 34916 812 38780 868
rect 38836 812 38846 868
rect 48514 812 48524 868
rect 48580 812 53788 868
rect 53844 812 53854 868
rect 4454 756 4464 812
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4728 756 4738 812
rect 24454 756 24464 812
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24728 756 24738 812
rect 44454 756 44464 812
rect 44520 756 44568 812
rect 44624 756 44672 812
rect 44728 756 44738 812
rect 5954 700 5964 756
rect 6020 700 15148 756
rect 15204 700 15214 756
rect 24882 700 24892 756
rect 24948 700 29988 756
rect 31938 700 31948 756
rect 32004 700 44324 756
rect 49746 700 49756 756
rect 49812 700 54460 756
rect 54516 700 54526 756
rect 29932 644 29988 700
rect 44268 644 44324 700
rect 9874 588 9884 644
rect 9940 588 28476 644
rect 28532 588 28542 644
rect 29932 588 34972 644
rect 35028 588 35038 644
rect 38434 588 38444 644
rect 38500 588 43708 644
rect 43764 588 43774 644
rect 44268 588 45612 644
rect 45668 588 45678 644
rect 48402 588 48412 644
rect 48468 588 53676 644
rect 53732 588 53742 644
rect 0 532 112 560
rect 57344 532 57456 560
rect 0 476 5628 532
rect 5684 476 5694 532
rect 12786 476 12796 532
rect 12852 476 16716 532
rect 16772 476 16782 532
rect 20514 476 20524 532
rect 20580 476 31388 532
rect 31444 476 31454 532
rect 38658 476 38668 532
rect 38724 476 47404 532
rect 47460 476 47470 532
rect 57026 476 57036 532
rect 57092 476 57456 532
rect 0 448 112 476
rect 57344 448 57456 476
rect 10210 364 10220 420
rect 10276 364 14084 420
rect 16818 364 16828 420
rect 16884 364 29148 420
rect 29204 364 29214 420
rect 44034 364 44044 420
rect 44100 364 49644 420
rect 49700 364 49710 420
rect 14028 308 14084 364
rect 2146 252 2156 308
rect 2212 252 13804 308
rect 13860 252 13870 308
rect 14028 252 17276 308
rect 17332 252 17342 308
rect 22978 252 22988 308
rect 23044 252 24892 308
rect 24948 252 24958 308
rect 26012 252 38556 308
rect 38612 252 38622 308
rect 26012 196 26068 252
rect 9426 140 9436 196
rect 9492 140 10108 196
rect 10164 140 10174 196
rect 11442 140 11452 196
rect 11508 140 11900 196
rect 11956 140 11966 196
rect 13458 140 13468 196
rect 13524 140 14140 196
rect 14196 140 14206 196
rect 15474 140 15484 196
rect 15540 140 15820 196
rect 15876 140 15886 196
rect 17490 140 17500 196
rect 17556 140 17566 196
rect 18610 140 18620 196
rect 18676 140 26068 196
rect 29586 140 29596 196
rect 29652 140 31948 196
rect 32004 140 32014 196
rect 42130 140 42140 196
rect 42196 140 47740 196
rect 47796 140 47806 196
rect 0 84 112 112
rect 17500 84 17556 140
rect 57344 84 57456 112
rect 0 28 5068 84
rect 5124 28 5134 84
rect 17500 28 20300 84
rect 20356 28 20366 84
rect 21746 28 21756 84
rect 21812 28 32284 84
rect 32340 28 32350 84
rect 56914 28 56924 84
rect 56980 28 57456 84
rect 0 0 112 28
rect 57344 0 57456 28
<< via3 >>
rect 25340 14140 25396 14196
rect 28476 14140 28532 14196
rect 28700 14140 28756 14196
rect 34748 14140 34804 14196
rect 24220 14028 24276 14084
rect 25228 13916 25284 13972
rect 25452 13916 25508 13972
rect 40236 13916 40292 13972
rect 21980 13804 22036 13860
rect 26236 13804 26292 13860
rect 27244 13804 27300 13860
rect 34748 13804 34804 13860
rect 27692 13692 27748 13748
rect 28588 13692 28644 13748
rect 18508 13580 18564 13636
rect 28924 13580 28980 13636
rect 33404 13468 33460 13524
rect 37660 13468 37716 13524
rect 24220 13356 24276 13412
rect 4464 13300 4520 13356
rect 4568 13300 4624 13356
rect 4672 13300 4728 13356
rect 24464 13300 24520 13356
rect 24568 13300 24624 13356
rect 24672 13300 24728 13356
rect 44464 13300 44520 13356
rect 44568 13300 44624 13356
rect 44672 13300 44728 13356
rect 29484 13244 29540 13300
rect 23548 13132 23604 13188
rect 25788 13132 25844 13188
rect 32732 13132 32788 13188
rect 18508 13020 18564 13076
rect 33516 13020 33572 13076
rect 33852 12908 33908 12964
rect 23548 12796 23604 12852
rect 26236 12796 26292 12852
rect 33292 12796 33348 12852
rect 24220 12684 24276 12740
rect 32732 12684 32788 12740
rect 3804 12516 3860 12572
rect 3908 12516 3964 12572
rect 4012 12516 4068 12572
rect 17948 12572 18004 12628
rect 24892 12572 24948 12628
rect 25228 12572 25284 12628
rect 33180 12572 33236 12628
rect 23804 12516 23860 12572
rect 23908 12516 23964 12572
rect 24012 12516 24068 12572
rect 43804 12516 43860 12572
rect 43908 12516 43964 12572
rect 44012 12516 44068 12572
rect 21532 12348 21588 12404
rect 33292 12460 33348 12516
rect 25788 12348 25844 12404
rect 18396 12124 18452 12180
rect 17948 12012 18004 12068
rect 21980 12012 22036 12068
rect 4464 11732 4520 11788
rect 4568 11732 4624 11788
rect 4672 11732 4728 11788
rect 24220 11788 24276 11844
rect 45948 11788 46004 11844
rect 24464 11732 24520 11788
rect 24568 11732 24624 11788
rect 24672 11732 24728 11788
rect 44464 11732 44520 11788
rect 44568 11732 44624 11788
rect 44672 11732 44728 11788
rect 30380 11676 30436 11732
rect 44156 11676 44212 11732
rect 46844 11676 46900 11732
rect 46620 11564 46676 11620
rect 46956 11564 47012 11620
rect 32396 11452 32452 11508
rect 46508 11452 46564 11508
rect 27580 11340 27636 11396
rect 28588 11228 28644 11284
rect 35308 11228 35364 11284
rect 31052 11116 31108 11172
rect 42700 11116 42756 11172
rect 44156 11004 44212 11060
rect 3804 10948 3860 11004
rect 3908 10948 3964 11004
rect 4012 10948 4068 11004
rect 23804 10948 23860 11004
rect 23908 10948 23964 11004
rect 24012 10948 24068 11004
rect 43804 10948 43860 11004
rect 43908 10948 43964 11004
rect 44012 10948 44068 11004
rect 21756 10892 21812 10948
rect 46956 10892 47012 10948
rect 38780 10780 38836 10836
rect 42588 10780 42644 10836
rect 31052 10668 31108 10724
rect 31948 10668 32004 10724
rect 11004 10556 11060 10612
rect 34524 10556 34580 10612
rect 40684 10556 40740 10612
rect 25340 10444 25396 10500
rect 27580 10444 27636 10500
rect 27804 10444 27860 10500
rect 33852 10444 33908 10500
rect 38220 10444 38276 10500
rect 42252 10444 42308 10500
rect 30492 10332 30548 10388
rect 10556 10220 10612 10276
rect 25116 10220 25172 10276
rect 4464 10164 4520 10220
rect 4568 10164 4624 10220
rect 4672 10164 4728 10220
rect 24464 10164 24520 10220
rect 24568 10164 24624 10220
rect 24672 10164 24728 10220
rect 42700 10332 42756 10388
rect 40684 10220 40740 10276
rect 44464 10164 44520 10220
rect 44568 10164 44624 10220
rect 44672 10164 44728 10220
rect 24220 10108 24276 10164
rect 30492 10108 30548 10164
rect 41692 10108 41748 10164
rect 26684 9996 26740 10052
rect 28252 9996 28308 10052
rect 22652 9884 22708 9940
rect 25340 9884 25396 9940
rect 28252 9660 28308 9716
rect 11004 9548 11060 9604
rect 13132 9436 13188 9492
rect 22652 9436 22708 9492
rect 25340 9436 25396 9492
rect 3804 9380 3860 9436
rect 3908 9380 3964 9436
rect 4012 9380 4068 9436
rect 23804 9380 23860 9436
rect 23908 9380 23964 9436
rect 24012 9380 24068 9436
rect 43804 9380 43860 9436
rect 43908 9380 43964 9436
rect 44012 9380 44068 9436
rect 25788 9324 25844 9380
rect 33964 9324 34020 9380
rect 22204 9212 22260 9268
rect 25116 9212 25172 9268
rect 31948 9212 32004 9268
rect 36876 9212 36932 9268
rect 39564 9212 39620 9268
rect 42252 9212 42308 9268
rect 21756 9100 21812 9156
rect 26684 9100 26740 9156
rect 26852 9100 26908 9156
rect 33740 9100 33796 9156
rect 33964 9100 34020 9156
rect 41916 9100 41972 9156
rect 45948 9100 46004 9156
rect 21980 8876 22036 8932
rect 33740 8876 33796 8932
rect 41804 8876 41860 8932
rect 39564 8764 39620 8820
rect 25564 8652 25620 8708
rect 4464 8596 4520 8652
rect 4568 8596 4624 8652
rect 4672 8596 4728 8652
rect 24464 8596 24520 8652
rect 24568 8596 24624 8652
rect 24672 8596 24728 8652
rect 44464 8596 44520 8652
rect 44568 8596 44624 8652
rect 44672 8596 44728 8652
rect 22092 8540 22148 8596
rect 22316 8540 22372 8596
rect 24892 8540 24948 8596
rect 13132 8428 13188 8484
rect 13580 8428 13636 8484
rect 28364 8428 28420 8484
rect 34972 8428 35028 8484
rect 22204 8316 22260 8372
rect 24892 8316 24948 8372
rect 42476 8316 42532 8372
rect 22540 8204 22596 8260
rect 39564 8204 39620 8260
rect 25004 8092 25060 8148
rect 42924 8092 42980 8148
rect 24220 7980 24276 8036
rect 25452 7980 25508 8036
rect 22540 7868 22596 7924
rect 29596 7868 29652 7924
rect 41132 7868 41188 7924
rect 43596 7868 43652 7924
rect 3804 7812 3860 7868
rect 3908 7812 3964 7868
rect 4012 7812 4068 7868
rect 23804 7812 23860 7868
rect 23908 7812 23964 7868
rect 24012 7812 24068 7868
rect 43804 7812 43860 7868
rect 43908 7812 43964 7868
rect 44012 7812 44068 7868
rect 25004 7644 25060 7700
rect 38892 7644 38948 7700
rect 39116 7644 39172 7700
rect 10556 7532 10612 7588
rect 20188 7532 20244 7588
rect 36988 7532 37044 7588
rect 50092 7532 50148 7588
rect 12796 7420 12852 7476
rect 11452 7308 11508 7364
rect 21868 7420 21924 7476
rect 31500 7420 31556 7476
rect 36876 7420 36932 7476
rect 39116 7420 39172 7476
rect 43596 7420 43652 7476
rect 38444 7308 38500 7364
rect 40796 7308 40852 7364
rect 41692 7308 41748 7364
rect 12796 7196 12852 7252
rect 30940 7196 30996 7252
rect 39900 7196 39956 7252
rect 22204 7084 22260 7140
rect 24892 7084 24948 7140
rect 4464 7028 4520 7084
rect 4568 7028 4624 7084
rect 4672 7028 4728 7084
rect 24464 7028 24520 7084
rect 24568 7028 24624 7084
rect 24672 7028 24728 7084
rect 37660 7084 37716 7140
rect 44464 7028 44520 7084
rect 44568 7028 44624 7084
rect 44672 7028 44728 7084
rect 40236 6972 40292 7028
rect 11228 6860 11284 6916
rect 11452 6860 11508 6916
rect 23436 6860 23492 6916
rect 23660 6860 23716 6916
rect 46620 6860 46676 6916
rect 50092 6860 50148 6916
rect 34972 6748 35028 6804
rect 35196 6748 35252 6804
rect 38444 6748 38500 6804
rect 38892 6748 38948 6804
rect 22428 6636 22484 6692
rect 31500 6636 31556 6692
rect 18396 6524 18452 6580
rect 22092 6524 22148 6580
rect 25340 6524 25396 6580
rect 40236 6524 40292 6580
rect 47292 6524 47348 6580
rect 11228 6412 11284 6468
rect 21980 6412 22036 6468
rect 23660 6300 23716 6356
rect 28252 6300 28308 6356
rect 28476 6300 28532 6356
rect 42924 6300 42980 6356
rect 3804 6244 3860 6300
rect 3908 6244 3964 6300
rect 4012 6244 4068 6300
rect 23804 6244 23860 6300
rect 23908 6244 23964 6300
rect 24012 6244 24068 6300
rect 43804 6244 43860 6300
rect 43908 6244 43964 6300
rect 44012 6244 44068 6300
rect 5068 6188 5124 6244
rect 13356 6188 13412 6244
rect 18396 6188 18452 6244
rect 24892 6188 24948 6244
rect 28700 6188 28756 6244
rect 38780 6188 38836 6244
rect 47292 6188 47348 6244
rect 34524 6076 34580 6132
rect 44828 6076 44884 6132
rect 23436 5964 23492 6020
rect 41804 5964 41860 6020
rect 42476 5964 42532 6020
rect 20860 5852 20916 5908
rect 22204 5852 22260 5908
rect 24892 5852 24948 5908
rect 42588 5852 42644 5908
rect 46844 5852 46900 5908
rect 21532 5628 21588 5684
rect 25228 5628 25284 5684
rect 38668 5628 38724 5684
rect 25340 5516 25396 5572
rect 26796 5516 26852 5572
rect 30604 5516 30660 5572
rect 44828 5516 44884 5572
rect 4464 5460 4520 5516
rect 4568 5460 4624 5516
rect 4672 5460 4728 5516
rect 24464 5460 24520 5516
rect 24568 5460 24624 5516
rect 24672 5460 24728 5516
rect 44464 5460 44520 5516
rect 44568 5460 44624 5516
rect 44672 5460 44728 5516
rect 30156 5292 30212 5348
rect 31892 5292 31948 5348
rect 6748 5068 6804 5124
rect 21644 5068 21700 5124
rect 25228 5068 25284 5124
rect 29484 4956 29540 5012
rect 31892 4956 31948 5012
rect 32060 4956 32116 5012
rect 21868 4844 21924 4900
rect 26684 4844 26740 4900
rect 26908 4844 26964 4900
rect 35196 4844 35252 4900
rect 18956 4732 19012 4788
rect 20076 4732 20132 4788
rect 3804 4676 3860 4732
rect 3908 4676 3964 4732
rect 4012 4676 4068 4732
rect 24220 4732 24276 4788
rect 25788 4732 25844 4788
rect 32284 4732 32340 4788
rect 38220 4732 38276 4788
rect 41468 4732 41524 4788
rect 23804 4676 23860 4732
rect 23908 4676 23964 4732
rect 24012 4676 24068 4732
rect 43804 4676 43860 4732
rect 43908 4676 43964 4732
rect 44012 4676 44068 4732
rect 21756 4620 21812 4676
rect 30044 4620 30100 4676
rect 46508 4620 46564 4676
rect 6748 4508 6804 4564
rect 44828 4508 44884 4564
rect 18732 4396 18788 4452
rect 20076 4396 20132 4452
rect 24220 4396 24276 4452
rect 25788 4396 25844 4452
rect 35308 4396 35364 4452
rect 41468 4396 41524 4452
rect 22428 4284 22484 4340
rect 25788 4172 25844 4228
rect 38780 4172 38836 4228
rect 48076 4172 48132 4228
rect 15260 4060 15316 4116
rect 18732 4060 18788 4116
rect 18956 4060 19012 4116
rect 32396 4060 32452 4116
rect 44268 4060 44324 4116
rect 30828 3948 30884 4004
rect 4464 3892 4520 3948
rect 4568 3892 4624 3948
rect 4672 3892 4728 3948
rect 24464 3892 24520 3948
rect 24568 3892 24624 3948
rect 24672 3892 24728 3948
rect 44464 3892 44520 3948
rect 44568 3892 44624 3948
rect 44672 3892 44728 3948
rect 20188 3836 20244 3892
rect 21644 3836 21700 3892
rect 30940 3836 30996 3892
rect 30268 3724 30324 3780
rect 15036 3612 15092 3668
rect 28812 3612 28868 3668
rect 5180 3500 5236 3556
rect 36652 3500 36708 3556
rect 44828 3724 44884 3780
rect 44268 3612 44324 3668
rect 48076 3500 48132 3556
rect 21868 3388 21924 3444
rect 30828 3388 30884 3444
rect 29148 3276 29204 3332
rect 18396 3164 18452 3220
rect 27356 3164 27412 3220
rect 33292 3164 33348 3220
rect 42476 3164 42532 3220
rect 3804 3108 3860 3164
rect 3908 3108 3964 3164
rect 4012 3108 4068 3164
rect 23804 3108 23860 3164
rect 23908 3108 23964 3164
rect 24012 3108 24068 3164
rect 43804 3108 43860 3164
rect 43908 3108 43964 3164
rect 44012 3108 44068 3164
rect 26012 2940 26068 2996
rect 5180 2828 5236 2884
rect 33068 2716 33124 2772
rect 20860 2604 20916 2660
rect 29148 2604 29204 2660
rect 4464 2324 4520 2380
rect 4568 2324 4624 2380
rect 4672 2324 4728 2380
rect 20748 2492 20804 2548
rect 41916 2492 41972 2548
rect 27804 2380 27860 2436
rect 28028 2380 28084 2436
rect 42252 2380 42308 2436
rect 24464 2324 24520 2380
rect 24568 2324 24624 2380
rect 24672 2324 24728 2380
rect 44464 2324 44520 2380
rect 44568 2324 44624 2380
rect 44672 2324 44728 2380
rect 27692 2044 27748 2100
rect 29596 2044 29652 2100
rect 29820 2044 29876 2100
rect 33068 2044 33124 2100
rect 21980 1932 22036 1988
rect 27356 1932 27412 1988
rect 20748 1820 20804 1876
rect 25788 1820 25844 1876
rect 26012 1820 26068 1876
rect 3804 1540 3860 1596
rect 3908 1540 3964 1596
rect 4012 1540 4068 1596
rect 23804 1540 23860 1596
rect 23908 1540 23964 1596
rect 24012 1540 24068 1596
rect 15148 1484 15204 1540
rect 17276 1372 17332 1428
rect 43804 1540 43860 1596
rect 43908 1540 43964 1596
rect 44012 1540 44068 1596
rect 38668 1372 38724 1428
rect 35644 1148 35700 1204
rect 48412 1036 48468 1092
rect 30716 924 30772 980
rect 35644 924 35700 980
rect 29820 812 29876 868
rect 4464 756 4520 812
rect 4568 756 4624 812
rect 4672 756 4728 812
rect 24464 756 24520 812
rect 24568 756 24624 812
rect 24672 756 24728 812
rect 44464 756 44520 812
rect 44568 756 44624 812
rect 44672 756 44728 812
rect 15148 700 15204 756
rect 24892 700 24948 756
rect 48412 588 48468 644
rect 17276 252 17332 308
rect 24892 252 24948 308
rect 5068 28 5124 84
<< metal4 >>
rect 3776 12572 4096 14224
rect 3776 12516 3804 12572
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 4068 12516 4096 12572
rect 3776 11004 4096 12516
rect 3776 10948 3804 11004
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 4068 10948 4096 11004
rect 3776 9436 4096 10948
rect 3776 9380 3804 9436
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 4068 9380 4096 9436
rect 3776 7868 4096 9380
rect 3776 7812 3804 7868
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 4068 7812 4096 7868
rect 3776 6300 4096 7812
rect 3776 6244 3804 6300
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 4068 6244 4096 6300
rect 3776 4732 4096 6244
rect 3776 4676 3804 4732
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 4068 4676 4096 4732
rect 3776 3164 4096 4676
rect 3776 3108 3804 3164
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 4068 3108 4096 3164
rect 3776 1596 4096 3108
rect 3776 1540 3804 1596
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 4068 1540 4096 1596
rect 3776 0 4096 1540
rect 4436 13356 4756 14224
rect 21980 13860 22036 13870
rect 4436 13300 4464 13356
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4728 13300 4756 13356
rect 4436 11788 4756 13300
rect 18508 13636 18564 13646
rect 18508 13076 18564 13580
rect 18508 13010 18564 13020
rect 17948 12628 18004 12638
rect 17948 12068 18004 12572
rect 21532 12404 21588 12414
rect 17948 12002 18004 12012
rect 18396 12180 18452 12190
rect 4436 11732 4464 11788
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4728 11732 4756 11788
rect 4436 10220 4756 11732
rect 11004 10612 11060 10622
rect 4436 10164 4464 10220
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4728 10164 4756 10220
rect 4436 8652 4756 10164
rect 4436 8596 4464 8652
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4728 8596 4756 8652
rect 4436 7084 4756 8596
rect 10556 10276 10612 10286
rect 10556 7588 10612 10220
rect 11004 9604 11060 10556
rect 11004 9538 11060 9548
rect 13132 9492 13188 9502
rect 13132 8484 13188 9436
rect 13132 8418 13188 8428
rect 13580 8484 13636 8494
rect 13580 8398 13636 8428
rect 10556 7522 10612 7532
rect 13356 8342 13636 8398
rect 12796 7476 12852 7486
rect 4436 7028 4464 7084
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4728 7028 4756 7084
rect 4436 5516 4756 7028
rect 11452 7364 11508 7374
rect 11228 6916 11284 6926
rect 11228 6468 11284 6860
rect 11452 6916 11508 7308
rect 12796 7252 12852 7420
rect 12796 7186 12852 7196
rect 11452 6850 11508 6860
rect 11228 6402 11284 6412
rect 4436 5460 4464 5516
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4728 5460 4756 5516
rect 4436 3948 4756 5460
rect 4436 3892 4464 3948
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4728 3892 4756 3948
rect 4436 2380 4756 3892
rect 4436 2324 4464 2380
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4728 2324 4756 2380
rect 4436 812 4756 2324
rect 4436 756 4464 812
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4728 756 4756 812
rect 4436 0 4756 756
rect 5068 6244 5124 6254
rect 5068 84 5124 6188
rect 13356 6244 13412 8342
rect 18396 6580 18452 12124
rect 18396 6514 18452 6524
rect 20188 7588 20244 7598
rect 13356 6178 13412 6188
rect 18396 6244 18452 6254
rect 6748 5124 6804 5134
rect 6748 4564 6804 5068
rect 6748 4498 6804 4508
rect 15260 4116 15316 4126
rect 15260 3718 15316 4060
rect 15036 3668 15316 3718
rect 15092 3662 15316 3668
rect 15036 3602 15092 3612
rect 5180 3556 5236 3566
rect 5180 2884 5236 3500
rect 18396 3220 18452 6188
rect 18956 4788 19012 4798
rect 18732 4452 18788 4462
rect 18732 4116 18788 4396
rect 18732 4050 18788 4060
rect 18956 4116 19012 4732
rect 20076 4788 20132 4798
rect 20076 4452 20132 4732
rect 20076 4386 20132 4396
rect 18956 4050 19012 4060
rect 20188 3892 20244 7532
rect 20188 3826 20244 3836
rect 20860 5908 20916 5918
rect 18396 3154 18452 3164
rect 5180 2818 5236 2828
rect 20860 2660 20916 5852
rect 21532 5684 21588 12348
rect 21980 12068 22036 13804
rect 23548 13188 23604 13198
rect 23548 12852 23604 13132
rect 23548 12786 23604 12796
rect 21980 12002 22036 12012
rect 23776 12572 24096 14224
rect 24220 14084 24276 14094
rect 24220 13412 24276 14028
rect 24220 13346 24276 13356
rect 24436 13356 24756 14224
rect 25340 14196 25396 14206
rect 28476 14196 28532 14206
rect 25396 14140 25508 14158
rect 25340 14102 25508 14140
rect 24436 13300 24464 13356
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24728 13300 24756 13356
rect 23776 12516 23804 12572
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 24068 12516 24096 12572
rect 23776 11004 24096 12516
rect 24220 12740 24276 12750
rect 24220 11844 24276 12684
rect 24220 11778 24276 11788
rect 24436 11788 24756 13300
rect 25228 13972 25284 13982
rect 21756 10948 21812 10958
rect 21756 9156 21812 10892
rect 23776 10948 23804 11004
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 24068 10948 24096 11004
rect 22652 9940 22708 9950
rect 22652 9492 22708 9884
rect 22652 9426 22708 9436
rect 23776 9436 24096 10948
rect 24436 11732 24464 11788
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24728 11732 24756 11788
rect 24436 10220 24756 11732
rect 23776 9380 23804 9436
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 24068 9380 24096 9436
rect 21756 9090 21812 9100
rect 22204 9268 22260 9278
rect 21980 8932 22036 8942
rect 21532 5618 21588 5628
rect 21868 7476 21924 7486
rect 21644 5124 21700 5134
rect 21644 4978 21700 5068
rect 21644 4922 21812 4978
rect 21756 4676 21812 4922
rect 21868 4900 21924 7420
rect 21980 6468 22036 8876
rect 22092 8596 22148 8606
rect 22092 6580 22148 8540
rect 22204 8372 22260 9212
rect 22204 8306 22260 8316
rect 22316 8596 22372 8606
rect 22092 6514 22148 6524
rect 22204 7140 22260 7150
rect 21980 6402 22036 6412
rect 22204 6238 22260 7084
rect 21868 4834 21924 4844
rect 21980 6182 22260 6238
rect 21756 4610 21812 4620
rect 21644 3892 21700 3902
rect 21644 3358 21700 3836
rect 21868 3444 21924 3454
rect 21868 3358 21924 3388
rect 21644 3302 21924 3358
rect 20860 2594 20916 2604
rect 20748 2548 20804 2558
rect 20748 1876 20804 2492
rect 21980 1988 22036 6182
rect 22316 6058 22372 8540
rect 22540 8260 22596 8270
rect 22540 7924 22596 8204
rect 22540 7858 22596 7868
rect 23776 7868 24096 9380
rect 24220 10164 24276 10174
rect 24220 8036 24276 10108
rect 24220 7970 24276 7980
rect 24436 10164 24464 10220
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24728 10164 24756 10220
rect 24436 8652 24756 10164
rect 24436 8596 24464 8652
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24728 8596 24756 8652
rect 23776 7812 23804 7868
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 24068 7812 24096 7868
rect 23436 6916 23492 6926
rect 22204 6002 22372 6058
rect 22428 6692 22484 6702
rect 22204 5908 22260 6002
rect 22204 5842 22260 5852
rect 22428 4340 22484 6636
rect 23436 6020 23492 6860
rect 23660 6916 23716 6926
rect 23660 6356 23716 6860
rect 23660 6290 23716 6300
rect 23776 6300 24096 7812
rect 23436 5954 23492 5964
rect 23776 6244 23804 6300
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 24068 6244 24096 6300
rect 22428 4274 22484 4284
rect 23776 4732 24096 6244
rect 24436 7084 24756 8596
rect 24892 12628 24948 12638
rect 24892 8596 24948 12572
rect 25228 12628 25284 13916
rect 25452 13972 25508 14102
rect 25452 13906 25508 13916
rect 26236 13860 26292 13870
rect 25228 12562 25284 12572
rect 25788 13188 25844 13198
rect 25788 12404 25844 13132
rect 26236 12852 26292 13804
rect 27244 13860 27300 13870
rect 27244 13798 27300 13804
rect 27244 13748 27748 13798
rect 27244 13742 27692 13748
rect 27692 13682 27748 13692
rect 28476 13618 28532 14140
rect 28700 14196 28756 14206
rect 28700 13798 28756 14140
rect 28588 13748 28756 13798
rect 34748 14196 34804 14206
rect 34748 13860 34804 14140
rect 34748 13794 34804 13804
rect 40236 13972 40292 13982
rect 28644 13742 28756 13748
rect 28588 13682 28644 13692
rect 28924 13636 28980 13646
rect 28476 13580 28924 13618
rect 28476 13562 28980 13580
rect 33404 13524 33460 13534
rect 26236 12786 26292 12796
rect 29484 13300 29540 13310
rect 25788 12338 25844 12348
rect 27580 11396 27636 11406
rect 25340 10500 25396 10510
rect 25116 10276 25172 10286
rect 25116 9268 25172 10220
rect 25340 9940 25396 10444
rect 27580 10500 27636 11340
rect 28588 11284 28644 11294
rect 27580 10434 27636 10444
rect 27804 10500 27860 10510
rect 25340 9874 25396 9884
rect 26684 10052 26740 10062
rect 25340 9492 25396 9502
rect 25396 9436 25844 9478
rect 25340 9422 25844 9436
rect 25788 9380 25844 9422
rect 25788 9314 25844 9324
rect 25116 9202 25172 9212
rect 26684 9156 26740 9996
rect 26852 9156 26908 9166
rect 26684 9090 26740 9100
rect 26796 9100 26852 9118
rect 26796 9062 26908 9100
rect 24892 8530 24948 8540
rect 25564 8708 25620 8718
rect 24436 7028 24464 7084
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 24728 7028 24756 7084
rect 24892 8372 24948 8382
rect 24892 7140 24948 8316
rect 25004 8148 25060 8158
rect 25004 8038 25060 8092
rect 25452 8038 25508 8046
rect 25004 8036 25508 8038
rect 25004 7982 25452 8036
rect 25452 7970 25508 7980
rect 25004 7700 25060 7710
rect 25564 7678 25620 8652
rect 25060 7644 25620 7678
rect 25004 7622 25620 7644
rect 24892 7074 24948 7084
rect 24436 5516 24756 7028
rect 25340 6580 25396 6590
rect 24892 6244 24948 6254
rect 24892 5908 24948 6188
rect 24892 5842 24948 5852
rect 24436 5460 24464 5516
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24728 5460 24756 5516
rect 23776 4676 23804 4732
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 24068 4676 24096 4732
rect 21980 1922 22036 1932
rect 23776 3164 24096 4676
rect 24220 4788 24276 4798
rect 24220 4452 24276 4732
rect 24220 4386 24276 4396
rect 23776 3108 23804 3164
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 24068 3108 24096 3164
rect 20748 1810 20804 1820
rect 23776 1596 24096 3108
rect 15148 1540 15204 1550
rect 15148 756 15204 1484
rect 23776 1540 23804 1596
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 24068 1540 24096 1596
rect 15148 690 15204 700
rect 17276 1428 17332 1438
rect 17276 308 17332 1372
rect 17276 242 17332 252
rect 5068 18 5124 28
rect 23776 0 24096 1540
rect 24436 3948 24756 5460
rect 25228 5684 25284 5694
rect 25228 5124 25284 5628
rect 25340 5572 25396 6524
rect 26796 5698 26852 9062
rect 25340 5506 25396 5516
rect 26684 5642 26852 5698
rect 25228 5058 25284 5068
rect 26684 4900 26740 5642
rect 26796 5572 26852 5582
rect 26796 5158 26852 5516
rect 26796 5102 26964 5158
rect 26684 4834 26740 4844
rect 26908 4900 26964 5102
rect 26908 4834 26964 4844
rect 25788 4788 25844 4798
rect 25788 4452 25844 4732
rect 25788 4386 25844 4396
rect 24436 3892 24464 3948
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24728 3892 24756 3948
rect 24436 2380 24756 3892
rect 24436 2324 24464 2380
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24728 2324 24756 2380
rect 24436 812 24756 2324
rect 25788 4228 25844 4238
rect 25788 1876 25844 4172
rect 27356 3220 27412 3230
rect 25788 1810 25844 1820
rect 26012 2996 26068 3006
rect 26012 1876 26068 2940
rect 27356 1988 27412 3164
rect 27804 2436 27860 10444
rect 28252 10052 28308 10062
rect 28252 9716 28308 9996
rect 28252 9650 28308 9660
rect 28364 8522 28532 8578
rect 28364 8484 28420 8522
rect 28364 8418 28420 8428
rect 28252 6356 28308 6366
rect 28252 6058 28308 6300
rect 28476 6356 28532 8522
rect 28588 6418 28644 11228
rect 28588 6362 28868 6418
rect 28476 6290 28532 6300
rect 28700 6244 28756 6254
rect 28700 6058 28756 6188
rect 28252 6002 28756 6058
rect 28812 3668 28868 6362
rect 29484 5012 29540 13244
rect 32732 13188 32788 13198
rect 32732 12740 32788 13132
rect 33404 13078 33460 13468
rect 37660 13524 37716 13534
rect 33516 13078 33572 13086
rect 33404 13076 33572 13078
rect 33404 13022 33516 13076
rect 33516 13010 33572 13020
rect 33852 12964 33908 12974
rect 32732 12674 32788 12684
rect 33292 12852 33348 12862
rect 33180 12628 33236 12638
rect 30380 11732 30436 11742
rect 29484 4946 29540 4956
rect 29596 7924 29652 7934
rect 28812 3602 28868 3612
rect 29148 3332 29204 3342
rect 29148 2660 29204 3276
rect 29148 2594 29204 2604
rect 27804 2370 27860 2380
rect 28028 2436 28084 2446
rect 28028 2278 28084 2380
rect 27692 2222 28084 2278
rect 27692 2100 27748 2222
rect 27692 2034 27748 2044
rect 29596 2100 29652 7868
rect 30380 5698 30436 11676
rect 32396 11508 32452 11518
rect 31052 11172 31108 11182
rect 31052 10724 31108 11116
rect 31052 10658 31108 10668
rect 31948 10724 32004 10734
rect 30492 10388 30548 10398
rect 30492 10164 30548 10332
rect 30492 10098 30548 10108
rect 31948 9268 32004 10668
rect 31948 9202 32004 9212
rect 31500 7476 31556 7486
rect 30940 7252 30996 7262
rect 30380 5642 30772 5698
rect 30604 5572 30660 5582
rect 30044 5516 30604 5518
rect 30044 5462 30660 5516
rect 30044 4676 30100 5462
rect 30156 5348 30212 5358
rect 30212 5292 30324 5338
rect 30156 5282 30324 5292
rect 30044 4610 30100 4620
rect 30268 3780 30324 5282
rect 30268 3714 30324 3724
rect 29596 2034 29652 2044
rect 29820 2100 29876 2110
rect 27356 1922 27412 1932
rect 26012 1810 26068 1820
rect 24436 756 24464 812
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24728 756 24756 812
rect 29820 868 29876 2044
rect 30716 980 30772 5642
rect 30828 4004 30884 4014
rect 30828 3444 30884 3948
rect 30940 3892 30996 7196
rect 31500 6692 31556 7420
rect 31500 6626 31556 6636
rect 31892 5348 31948 5358
rect 31948 5292 32116 5338
rect 31892 5282 32116 5292
rect 31892 5012 31948 5022
rect 32060 5012 32116 5282
rect 31948 4956 32004 4978
rect 31892 4922 32004 4956
rect 32060 4946 32116 4956
rect 31948 4798 32004 4922
rect 31948 4788 32340 4798
rect 31948 4742 32284 4788
rect 32284 4722 32340 4732
rect 32396 4116 32452 11452
rect 33180 7498 33236 12572
rect 33292 12516 33348 12796
rect 33292 12450 33348 12460
rect 33852 10500 33908 12908
rect 35308 11284 35364 11294
rect 33852 10434 33908 10444
rect 34524 10612 34580 10622
rect 33964 9380 34020 9390
rect 33740 9156 33796 9166
rect 33740 8932 33796 9100
rect 33964 9156 34020 9324
rect 33964 9090 34020 9100
rect 33740 8866 33796 8876
rect 33180 7442 33348 7498
rect 32396 4050 32452 4060
rect 30940 3826 30996 3836
rect 30828 3378 30884 3388
rect 33292 3220 33348 7442
rect 34524 6132 34580 10556
rect 34972 8484 35028 8494
rect 34972 6804 35028 8428
rect 34972 6738 35028 6748
rect 35196 6804 35252 6814
rect 34524 6066 34580 6076
rect 35196 4900 35252 6748
rect 35196 4834 35252 4844
rect 35308 4452 35364 11228
rect 36876 9268 36932 9278
rect 36876 7476 36932 9212
rect 36876 7410 36932 7420
rect 36988 7588 37044 7598
rect 35308 4386 35364 4396
rect 36652 3556 36708 3566
rect 36988 3538 37044 7532
rect 37660 7140 37716 13468
rect 38780 10836 38836 10846
rect 37660 7074 37716 7084
rect 38220 10500 38276 10510
rect 38220 4788 38276 10444
rect 38444 7364 38500 7374
rect 38444 6804 38500 7308
rect 38444 6738 38500 6748
rect 38780 6244 38836 10780
rect 39564 9268 39620 9278
rect 39564 8820 39620 9212
rect 39564 8754 39620 8764
rect 39564 8260 39620 8270
rect 38892 7700 38948 7710
rect 38892 6804 38948 7644
rect 39116 7700 39172 7710
rect 39116 7476 39172 7644
rect 39116 7410 39172 7420
rect 38892 6738 38948 6748
rect 38780 6178 38836 6188
rect 38220 4722 38276 4732
rect 38668 5684 38724 5694
rect 36708 3500 37044 3538
rect 36652 3482 37044 3500
rect 33292 3154 33348 3164
rect 33068 2772 33124 2782
rect 33068 2100 33124 2716
rect 33068 2034 33124 2044
rect 38668 1428 38724 5628
rect 39564 4258 39620 8204
rect 40236 8038 40292 13916
rect 43776 12572 44096 14224
rect 43776 12516 43804 12572
rect 43860 12516 43908 12572
rect 43964 12516 44012 12572
rect 44068 12516 44096 12572
rect 42700 11172 42756 11182
rect 42588 10836 42644 10846
rect 40684 10612 40740 10622
rect 40684 10276 40740 10556
rect 42252 10500 42308 10510
rect 42252 10378 42308 10444
rect 42252 10322 42532 10378
rect 40684 10210 40740 10220
rect 41692 10164 41748 10174
rect 40236 7982 41188 8038
rect 41132 7924 41188 7982
rect 41132 7858 41188 7868
rect 40796 7364 40852 7374
rect 39900 7308 40796 7318
rect 39900 7262 40852 7308
rect 41692 7364 41748 10108
rect 42252 9268 42308 9278
rect 41916 9156 41972 9166
rect 41692 7298 41748 7308
rect 41804 8932 41860 8942
rect 39900 7252 39956 7262
rect 39900 7186 39956 7196
rect 40236 7028 40292 7038
rect 40236 6580 40292 6972
rect 40236 6514 40292 6524
rect 41804 6020 41860 8876
rect 41804 5954 41860 5964
rect 41468 4788 41524 4798
rect 41468 4452 41524 4732
rect 41468 4386 41524 4396
rect 38780 4228 39620 4258
rect 38836 4202 39620 4228
rect 38780 4162 38836 4172
rect 41916 2548 41972 9100
rect 41916 2482 41972 2492
rect 42252 2436 42308 9212
rect 42476 8372 42532 10322
rect 42476 8306 42532 8316
rect 42476 6020 42532 6030
rect 42476 3220 42532 5964
rect 42588 5908 42644 10780
rect 42700 10388 42756 11116
rect 42700 10322 42756 10332
rect 43776 11004 44096 12516
rect 44436 13356 44756 14224
rect 44436 13300 44464 13356
rect 44520 13300 44568 13356
rect 44624 13300 44672 13356
rect 44728 13300 44756 13356
rect 44436 11788 44756 13300
rect 43776 10948 43804 11004
rect 43860 10948 43908 11004
rect 43964 10948 44012 11004
rect 44068 10948 44096 11004
rect 44156 11732 44212 11742
rect 44156 11060 44212 11676
rect 44156 10994 44212 11004
rect 44436 11732 44464 11788
rect 44520 11732 44568 11788
rect 44624 11732 44672 11788
rect 44728 11732 44756 11788
rect 43776 9436 44096 10948
rect 43776 9380 43804 9436
rect 43860 9380 43908 9436
rect 43964 9380 44012 9436
rect 44068 9380 44096 9436
rect 42924 8148 42980 8158
rect 42924 6356 42980 8092
rect 43596 7924 43652 7934
rect 43596 7476 43652 7868
rect 43596 7410 43652 7420
rect 43776 7868 44096 9380
rect 43776 7812 43804 7868
rect 43860 7812 43908 7868
rect 43964 7812 44012 7868
rect 44068 7812 44096 7868
rect 42924 6290 42980 6300
rect 43776 6300 44096 7812
rect 42588 5842 42644 5852
rect 43776 6244 43804 6300
rect 43860 6244 43908 6300
rect 43964 6244 44012 6300
rect 44068 6244 44096 6300
rect 42476 3154 42532 3164
rect 43776 4732 44096 6244
rect 43776 4676 43804 4732
rect 43860 4676 43908 4732
rect 43964 4676 44012 4732
rect 44068 4676 44096 4732
rect 43776 3164 44096 4676
rect 44436 10220 44756 11732
rect 44436 10164 44464 10220
rect 44520 10164 44568 10220
rect 44624 10164 44672 10220
rect 44728 10164 44756 10220
rect 44436 8652 44756 10164
rect 45948 11844 46004 11854
rect 45948 9156 46004 11788
rect 46844 11732 46900 11742
rect 46620 11620 46676 11630
rect 45948 9090 46004 9100
rect 46508 11508 46564 11518
rect 44436 8596 44464 8652
rect 44520 8596 44568 8652
rect 44624 8596 44672 8652
rect 44728 8596 44756 8652
rect 44436 7084 44756 8596
rect 44436 7028 44464 7084
rect 44520 7028 44568 7084
rect 44624 7028 44672 7084
rect 44728 7028 44756 7084
rect 44436 5516 44756 7028
rect 44436 5460 44464 5516
rect 44520 5460 44568 5516
rect 44624 5460 44672 5516
rect 44728 5460 44756 5516
rect 44828 6132 44884 6142
rect 44828 5572 44884 6076
rect 44828 5506 44884 5516
rect 44268 4116 44324 4126
rect 44268 3668 44324 4060
rect 44268 3602 44324 3612
rect 44436 3948 44756 5460
rect 46508 4676 46564 11452
rect 46620 6916 46676 11564
rect 46620 6850 46676 6860
rect 46844 5908 46900 11676
rect 46956 11620 47012 11630
rect 46956 10948 47012 11564
rect 46956 10882 47012 10892
rect 50092 7588 50148 7598
rect 50092 6916 50148 7532
rect 50092 6850 50148 6860
rect 47292 6580 47348 6590
rect 47292 6244 47348 6524
rect 47292 6178 47348 6188
rect 46844 5842 46900 5852
rect 46508 4610 46564 4620
rect 44436 3892 44464 3948
rect 44520 3892 44568 3948
rect 44624 3892 44672 3948
rect 44728 3892 44756 3948
rect 42252 2370 42308 2380
rect 43776 3108 43804 3164
rect 43860 3108 43908 3164
rect 43964 3108 44012 3164
rect 44068 3108 44096 3164
rect 38668 1362 38724 1372
rect 43776 1596 44096 3108
rect 43776 1540 43804 1596
rect 43860 1540 43908 1596
rect 43964 1540 44012 1596
rect 44068 1540 44096 1596
rect 30716 914 30772 924
rect 35644 1204 35700 1214
rect 35644 980 35700 1148
rect 35644 914 35700 924
rect 29820 802 29876 812
rect 24436 0 24756 756
rect 24892 756 24948 766
rect 24892 308 24948 700
rect 24892 242 24948 252
rect 43776 0 44096 1540
rect 44436 2380 44756 3892
rect 44828 4564 44884 4574
rect 44828 3780 44884 4508
rect 44828 3714 44884 3724
rect 48076 4228 48132 4238
rect 48076 3556 48132 4172
rect 48076 3490 48132 3500
rect 44436 2324 44464 2380
rect 44520 2324 44568 2380
rect 44624 2324 44672 2380
rect 44728 2324 44756 2380
rect 44436 812 44756 2324
rect 44436 756 44464 812
rect 44520 756 44568 812
rect 44624 756 44672 812
rect 44728 756 44756 812
rect 44436 0 44756 756
rect 48412 1092 48468 1102
rect 48412 644 48468 1036
rect 48412 578 48468 588
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _043_
timestamp 1486834041
transform 1 0 41440 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _044_
timestamp 1486834041
transform 1 0 40544 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _045_
timestamp 1486834041
transform -1 0 42784 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _046_
timestamp 1486834041
transform -1 0 39760 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _047_
timestamp 1486834041
transform 1 0 38528 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _048_
timestamp 1486834041
transform -1 0 19264 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _049_
timestamp 1486834041
transform 1 0 18144 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _050_
timestamp 1486834041
transform -1 0 27552 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _051_
timestamp 1486834041
transform 1 0 26656 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _052_
timestamp 1486834041
transform 1 0 10416 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _053_
timestamp 1486834041
transform -1 0 11872 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _054_
timestamp 1486834041
transform -1 0 39312 0 -1 8624
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _055_
timestamp 1486834041
transform -1 0 42448 0 -1 8624
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _056_
timestamp 1486834041
transform -1 0 36960 0 -1 8624
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _057_
timestamp 1486834041
transform 1 0 39424 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _058_
timestamp 1486834041
transform 1 0 42560 0 -1 7056
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _059_
timestamp 1486834041
transform 1 0 40992 0 1 10192
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _060_
timestamp 1486834041
transform -1 0 40992 0 1 10192
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _061_
timestamp 1486834041
transform -1 0 41440 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _062_
timestamp 1486834041
transform -1 0 43792 0 1 8624
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _063_
timestamp 1486834041
transform 1 0 40880 0 -1 7056
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _064_
timestamp 1486834041
transform 1 0 40656 0 -1 11760
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _065_
timestamp 1486834041
transform -1 0 39760 0 1 5488
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _066_
timestamp 1486834041
transform -1 0 39872 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _067_
timestamp 1486834041
transform 1 0 36176 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _068_
timestamp 1486834041
transform -1 0 37520 0 1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _069_
timestamp 1486834041
transform -1 0 38864 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _070_
timestamp 1486834041
transform 1 0 17696 0 1 3920
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _071_
timestamp 1486834041
transform -1 0 18928 0 1 10192
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _072_
timestamp 1486834041
transform 1 0 18256 0 -1 8624
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _073_
timestamp 1486834041
transform 1 0 18256 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _074_
timestamp 1486834041
transform 1 0 20832 0 1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _075_
timestamp 1486834041
transform -1 0 20160 0 1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _076_
timestamp 1486834041
transform 1 0 18592 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _077_
timestamp 1486834041
transform 1 0 26432 0 1 5488
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _078_
timestamp 1486834041
transform 1 0 28336 0 1 7056
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _079_
timestamp 1486834041
transform 1 0 28336 0 1 3920
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _080_
timestamp 1486834041
transform -1 0 27776 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _081_
timestamp 1486834041
transform 1 0 28784 0 1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _082_
timestamp 1486834041
transform -1 0 30128 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _083_
timestamp 1486834041
transform 1 0 28560 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _084_
timestamp 1486834041
transform 1 0 10752 0 1 8624
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _085_
timestamp 1486834041
transform 1 0 12544 0 -1 8624
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _086_
timestamp 1486834041
transform -1 0 12432 0 1 7056
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _087_
timestamp 1486834041
transform 1 0 10864 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _088_
timestamp 1486834041
transform 1 0 12320 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _089_
timestamp 1486834041
transform -1 0 12320 0 -1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _090_
timestamp 1486834041
transform 1 0 11760 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _091_
timestamp 1486834041
transform 1 0 22064 0 -1 5488
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _092_
timestamp 1486834041
transform 1 0 32368 0 1 5488
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _093_
timestamp 1486834041
transform 1 0 26432 0 -1 10192
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _094_
timestamp 1486834041
transform 1 0 31136 0 1 8624
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _095_
timestamp 1486834041
transform 1 0 29680 0 1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _096_
timestamp 1486834041
transform 1 0 25872 0 1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _097_
timestamp 1486834041
transform 1 0 30128 0 1 5488
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _098_
timestamp 1486834041
transform 1 0 21056 0 1 3920
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _099_
timestamp 1486834041
transform 1 0 9184 0 1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _100_
timestamp 1486834041
transform 1 0 7952 0 1 7056
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _101_
timestamp 1486834041
transform 1 0 8960 0 1 3920
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _102_
timestamp 1486834041
transform 1 0 24416 0 -1 7056
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _103_
timestamp 1486834041
transform 1 0 24976 0 1 2352
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _104_
timestamp 1486834041
transform 1 0 24416 0 -1 2352
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _105_
timestamp 1486834041
transform 1 0 7504 0 1 5488
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _106_
timestamp 1486834041
transform 1 0 20944 0 -1 7056
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _107_
timestamp 1486834041
transform 1 0 15792 0 1 7056
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _108_
timestamp 1486834041
transform 1 0 34048 0 -1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _109_
timestamp 1486834041
transform 1 0 33824 0 -1 5488
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _110_
timestamp 1486834041
transform 1 0 36288 0 1 2352
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _111_
timestamp 1486834041
transform 1 0 35392 0 -1 3920
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _112_
timestamp 1486834041
transform 1 0 37520 0 1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _113_
timestamp 1486834041
transform 1 0 33040 0 1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _115_
timestamp 1486834041
transform 1 0 50288 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _116_
timestamp 1486834041
transform 1 0 45808 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _117_
timestamp 1486834041
transform 1 0 4816 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _118_
timestamp 1486834041
transform 1 0 51856 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _119_
timestamp 1486834041
transform 1 0 9744 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _120_
timestamp 1486834041
transform 1 0 23296 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _121_
timestamp 1486834041
transform 1 0 25200 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _122_
timestamp 1486834041
transform 1 0 13104 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _123_
timestamp 1486834041
transform 1 0 31136 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _124_
timestamp 1486834041
transform 1 0 44912 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _125_
timestamp 1486834041
transform 1 0 40992 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _126_
timestamp 1486834041
transform 1 0 23184 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _127_
timestamp 1486834041
transform 1 0 13216 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _128_
timestamp 1486834041
transform 1 0 29904 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _129_
timestamp 1486834041
transform 1 0 27440 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _130_
timestamp 1486834041
transform 1 0 30800 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _131_
timestamp 1486834041
transform 1 0 21392 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _132_
timestamp 1486834041
transform 1 0 9072 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _133_
timestamp 1486834041
transform 1 0 7616 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _134_
timestamp 1486834041
transform 1 0 9184 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _135_
timestamp 1486834041
transform 1 0 24528 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _136_
timestamp 1486834041
transform 1 0 25424 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _137_
timestamp 1486834041
transform 1 0 23296 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _138_
timestamp 1486834041
transform 1 0 6608 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _139_
timestamp 1486834041
transform 1 0 21504 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _140_
timestamp 1486834041
transform 1 0 16576 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _141_
timestamp 1486834041
transform 1 0 34272 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _142_
timestamp 1486834041
transform 1 0 34272 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _143_
timestamp 1486834041
transform 1 0 36512 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _144_
timestamp 1486834041
transform 1 0 35056 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _145_
timestamp 1486834041
transform 1 0 38304 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _146_
timestamp 1486834041
transform 1 0 33376 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _147_
timestamp 1486834041
transform 1 0 36176 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _148_
timestamp 1486834041
transform 1 0 51520 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _149_
timestamp 1486834041
transform 1 0 49728 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _150_
timestamp 1486834041
transform 1 0 46256 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _151_
timestamp 1486834041
transform 1 0 49840 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _152_
timestamp 1486834041
transform 1 0 49616 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _153_
timestamp 1486834041
transform 1 0 45360 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _154_
timestamp 1486834041
transform 1 0 46816 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _155_
timestamp 1486834041
transform 1 0 50400 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _156_
timestamp 1486834041
transform 1 0 39872 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _157_
timestamp 1486834041
transform 1 0 50624 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _158_
timestamp 1486834041
transform 1 0 48384 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _159_
timestamp 1486834041
transform 1 0 47712 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _160_
timestamp 1486834041
transform -1 0 38640 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _161_
timestamp 1486834041
transform 1 0 51296 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _162_
timestamp 1486834041
transform -1 0 42336 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _163_
timestamp 1486834041
transform 1 0 54320 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _164_
timestamp 1486834041
transform -1 0 32144 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _165_
timestamp 1486834041
transform -1 0 4256 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _166_
timestamp 1486834041
transform -1 0 13664 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _167_
timestamp 1486834041
transform -1 0 31920 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _168_
timestamp 1486834041
transform 1 0 26544 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _169_
timestamp 1486834041
transform -1 0 32032 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _170_
timestamp 1486834041
transform -1 0 22064 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _171_
timestamp 1486834041
transform 1 0 32144 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _172_
timestamp 1486834041
transform -1 0 18816 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _173_
timestamp 1486834041
transform -1 0 21616 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _174_
timestamp 1486834041
transform -1 0 20272 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _175_
timestamp 1486834041
transform -1 0 38864 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _176_
timestamp 1486834041
transform -1 0 24192 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _177_
timestamp 1486834041
transform 1 0 32368 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _178_
timestamp 1486834041
transform -1 0 15904 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _179_
timestamp 1486834041
transform -1 0 35280 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _180_
timestamp 1486834041
transform -1 0 22288 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _181_
timestamp 1486834041
transform -1 0 30352 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _182_
timestamp 1486834041
transform -1 0 14224 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _183_
timestamp 1486834041
transform -1 0 37072 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _184_
timestamp 1486834041
transform -1 0 21280 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _185_
timestamp 1486834041
transform -1 0 28896 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _186_
timestamp 1486834041
transform -1 0 12432 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _187_
timestamp 1486834041
transform 1 0 52528 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _188_
timestamp 1486834041
transform 1 0 50736 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _189_
timestamp 1486834041
transform 1 0 46816 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _190_
timestamp 1486834041
transform 1 0 44352 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _191_
timestamp 1486834041
transform 1 0 45696 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _192_
timestamp 1486834041
transform 1 0 50736 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _193_
timestamp 1486834041
transform 1 0 49168 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _194_
timestamp 1486834041
transform -1 0 5712 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _195_
timestamp 1486834041
transform -1 0 42560 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _196_
timestamp 1486834041
transform -1 0 18704 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _197_
timestamp 1486834041
transform -1 0 26432 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _198_
timestamp 1486834041
transform 1 0 11424 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _199_
timestamp 1486834041
transform -1 0 43344 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _200_
timestamp 1486834041
transform -1 0 19824 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _201_
timestamp 1486834041
transform -1 0 29232 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _202_
timestamp 1486834041
transform 1 0 12768 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _203_
timestamp 1486834041
transform -1 0 47600 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _204_
timestamp 1486834041
transform 1 0 48832 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _205_
timestamp 1486834041
transform -1 0 46816 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _206_
timestamp 1486834041
transform 1 0 51520 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _207_
timestamp 1486834041
transform 1 0 53088 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _208_
timestamp 1486834041
transform 1 0 48272 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _209_
timestamp 1486834041
transform 1 0 47600 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _210_
timestamp 1486834041
transform 1 0 49728 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _211_
timestamp 1486834041
transform -1 0 42112 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _212_
timestamp 1486834041
transform -1 0 18144 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _213_
timestamp 1486834041
transform -1 0 28784 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _214_
timestamp 1486834041
transform 1 0 13328 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _215_
timestamp 1486834041
transform -1 0 43008 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _216_
timestamp 1486834041
transform 1 0 18144 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _217_
timestamp 1486834041
transform -1 0 29680 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _218_
timestamp 1486834041
transform 1 0 14224 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _219_
timestamp 1486834041
transform -1 0 49616 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout5
timestamp 1486834041
transform 1 0 25872 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout6
timestamp 1486834041
transform 1 0 26096 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2
timestamp 1486834041
transform 1 0 896 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6
timestamp 1486834041
transform 1 0 1344 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15
timestamp 1486834041
transform 1 0 2352 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23
timestamp 1486834041
transform 1 0 3248 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33
timestamp 1486834041
transform 1 0 4368 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36
timestamp 1486834041
transform 1 0 4704 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70
timestamp 1486834041
transform 1 0 8512 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78
timestamp 1486834041
transform 1 0 9408 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_93
timestamp 1486834041
transform 1 0 11088 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_101
timestamp 1486834041
transform 1 0 11984 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_104
timestamp 1486834041
transform 1 0 12320 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_112
timestamp 1486834041
transform 1 0 13216 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_114
timestamp 1486834041
transform 1 0 13440 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_129
timestamp 1486834041
transform 1 0 15120 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_133
timestamp 1486834041
transform 1 0 15568 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_135
timestamp 1486834041
transform 1 0 15792 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_138
timestamp 1486834041
transform 1 0 16128 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_172
timestamp 1486834041
transform 1 0 19936 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_206
timestamp 1486834041
transform 1 0 23744 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_214
timestamp 1486834041
transform 1 0 24640 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_218
timestamp 1486834041
transform 1 0 25088 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_220
timestamp 1486834041
transform 1 0 25312 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_229
timestamp 1486834041
transform 1 0 26320 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_237
timestamp 1486834041
transform 1 0 27216 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_240
timestamp 1486834041
transform 1 0 27552 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_274
timestamp 1486834041
transform 1 0 31360 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_308
timestamp 1486834041
transform 1 0 35168 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_342
timestamp 1486834041
transform 1 0 38976 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_376
timestamp 1486834041
transform 1 0 42784 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_410
timestamp 1486834041
transform 1 0 46592 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_444
timestamp 1486834041
transform 1 0 50400 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_478
timestamp 1486834041
transform 1 0 54208 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_482
timestamp 1486834041
transform 1 0 54656 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_484
timestamp 1486834041
transform 1 0 54880 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_2
timestamp 1486834041
transform 1 0 896 0 -1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_66
timestamp 1486834041
transform 1 0 8064 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_72
timestamp 1486834041
transform 1 0 8736 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_88
timestamp 1486834041
transform 1 0 10528 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_96
timestamp 1486834041
transform 1 0 11424 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_111
timestamp 1486834041
transform 1 0 13104 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_127
timestamp 1486834041
transform 1 0 14896 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_135
timestamp 1486834041
transform 1 0 15792 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_139
timestamp 1486834041
transform 1 0 16240 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_142
timestamp 1486834041
transform 1 0 16576 0 -1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_174
timestamp 1486834041
transform 1 0 20160 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_190
timestamp 1486834041
transform 1 0 21952 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_198
timestamp 1486834041
transform 1 0 22848 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_232
timestamp 1486834041
transform 1 0 26656 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_240
timestamp 1486834041
transform 1 0 27552 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_252
timestamp 1486834041
transform 1 0 28896 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_256
timestamp 1486834041
transform 1 0 29344 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_265
timestamp 1486834041
transform 1 0 30352 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_273
timestamp 1486834041
transform 1 0 31248 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_277
timestamp 1486834041
transform 1 0 31696 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_279
timestamp 1486834041
transform 1 0 31920 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_282
timestamp 1486834041
transform 1 0 32256 0 -1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_314
timestamp 1486834041
transform 1 0 35840 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_318
timestamp 1486834041
transform 1 0 36288 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_328
timestamp 1486834041
transform 1 0 37408 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_330
timestamp 1486834041
transform 1 0 37632 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_339
timestamp 1486834041
transform 1 0 38640 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_347
timestamp 1486834041
transform 1 0 39536 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_349
timestamp 1486834041
transform 1 0 39760 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_352
timestamp 1486834041
transform 1 0 40096 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_368
timestamp 1486834041
transform 1 0 41888 0 -1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_400
timestamp 1486834041
transform 1 0 45472 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_408
timestamp 1486834041
transform 1 0 46368 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_422
timestamp 1486834041
transform 1 0 47936 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_430
timestamp 1486834041
transform 1 0 48832 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_437
timestamp 1486834041
transform 1 0 49616 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_492
timestamp 1486834041
transform 1 0 55776 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_496
timestamp 1486834041
transform 1 0 56224 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_498
timestamp 1486834041
transform 1 0 56448 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_2
timestamp 1486834041
transform 1 0 896 0 1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1486834041
transform 1 0 4480 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_37
timestamp 1486834041
transform 1 0 4816 0 1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_101
timestamp 1486834041
transform 1 0 11984 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_107
timestamp 1486834041
transform 1 0 12656 0 1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_171
timestamp 1486834041
transform 1 0 19824 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_177
timestamp 1486834041
transform 1 0 20496 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_193
timestamp 1486834041
transform 1 0 22288 0 1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_209
timestamp 1486834041
transform 1 0 24080 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_237
timestamp 1486834041
transform 1 0 27216 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_247
timestamp 1486834041
transform 1 0 28336 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_291
timestamp 1486834041
transform 1 0 33264 0 1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_317
timestamp 1486834041
transform 1 0 36176 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_338
timestamp 1486834041
transform 1 0 38528 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_346
timestamp 1486834041
transform 1 0 39424 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_358
timestamp 1486834041
transform 1 0 40768 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_362
timestamp 1486834041
transform 1 0 41216 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_372
timestamp 1486834041
transform 1 0 42336 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_380
timestamp 1486834041
transform 1 0 43232 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_384
timestamp 1486834041
transform 1 0 43680 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_387
timestamp 1486834041
transform 1 0 44016 0 1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_419
timestamp 1486834041
transform 1 0 47600 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_428
timestamp 1486834041
transform 1 0 48608 0 1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_444
timestamp 1486834041
transform 1 0 50400 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_446
timestamp 1486834041
transform 1 0 50624 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_2
timestamp 1486834041
transform 1 0 896 0 -1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_66
timestamp 1486834041
transform 1 0 8064 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_72
timestamp 1486834041
transform 1 0 8736 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_84
timestamp 1486834041
transform 1 0 10080 0 -1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_116
timestamp 1486834041
transform 1 0 13664 0 -1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_132
timestamp 1486834041
transform 1 0 15456 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_142
timestamp 1486834041
transform 1 0 16576 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_150
timestamp 1486834041
transform 1 0 17472 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_152
timestamp 1486834041
transform 1 0 17696 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_161
timestamp 1486834041
transform 1 0 18704 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_171
timestamp 1486834041
transform 1 0 19824 0 -1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_203
timestamp 1486834041
transform 1 0 23408 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_207
timestamp 1486834041
transform 1 0 23856 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_209
timestamp 1486834041
transform 1 0 24080 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_212
timestamp 1486834041
transform 1 0 24416 0 -1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_228
timestamp 1486834041
transform 1 0 26208 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_240
timestamp 1486834041
transform 1 0 27552 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_248
timestamp 1486834041
transform 1 0 28448 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_263
timestamp 1486834041
transform 1 0 30128 0 -1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_279
timestamp 1486834041
transform 1 0 31920 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_282
timestamp 1486834041
transform 1 0 32256 0 -1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_298
timestamp 1486834041
transform 1 0 34048 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_306
timestamp 1486834041
transform 1 0 34944 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_330
timestamp 1486834041
transform 1 0 37632 0 -1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_346
timestamp 1486834041
transform 1 0 39424 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_352
timestamp 1486834041
transform 1 0 40096 0 -1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_416
timestamp 1486834041
transform 1 0 47264 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_422
timestamp 1486834041
transform 1 0 47936 0 -1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_492
timestamp 1486834041
transform 1 0 55776 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_496
timestamp 1486834041
transform 1 0 56224 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_498
timestamp 1486834041
transform 1 0 56448 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_10
timestamp 1486834041
transform 1 0 1792 0 1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_26
timestamp 1486834041
transform 1 0 3584 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1486834041
transform 1 0 4480 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_37
timestamp 1486834041
transform 1 0 4816 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_69
timestamp 1486834041
transform 1 0 8400 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_73
timestamp 1486834041
transform 1 0 8848 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_94
timestamp 1486834041
transform 1 0 11200 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_96
timestamp 1486834041
transform 1 0 11424 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_107
timestamp 1486834041
transform 1 0 12656 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_111
timestamp 1486834041
transform 1 0 13104 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_121
timestamp 1486834041
transform 1 0 14224 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_125
timestamp 1486834041
transform 1 0 14672 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_127
timestamp 1486834041
transform 1 0 14896 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_136
timestamp 1486834041
transform 1 0 15904 0 1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_167
timestamp 1486834041
transform 1 0 19376 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_177
timestamp 1486834041
transform 1 0 20496 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_181
timestamp 1486834041
transform 1 0 20944 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_202
timestamp 1486834041
transform 1 0 23296 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_242
timestamp 1486834041
transform 1 0 27776 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_244
timestamp 1486834041
transform 1 0 28000 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_252
timestamp 1486834041
transform 1 0 28896 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_284
timestamp 1486834041
transform 1 0 32480 0 1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_308
timestamp 1486834041
transform 1 0 35168 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_312
timestamp 1486834041
transform 1 0 35616 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_314
timestamp 1486834041
transform 1 0 35840 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_317
timestamp 1486834041
transform 1 0 36176 0 1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_333
timestamp 1486834041
transform 1 0 37968 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_341
timestamp 1486834041
transform 1 0 38864 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_349
timestamp 1486834041
transform 1 0 39760 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_381
timestamp 1486834041
transform 1 0 43344 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_387
timestamp 1486834041
transform 1 0 44016 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_389
timestamp 1486834041
transform 1 0 44240 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_398
timestamp 1486834041
transform 1 0 45248 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_430
timestamp 1486834041
transform 1 0 48832 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_446
timestamp 1486834041
transform 1 0 50624 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_454
timestamp 1486834041
transform 1 0 51520 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_457
timestamp 1486834041
transform 1 0 51856 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_461
timestamp 1486834041
transform 1 0 52304 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_18
timestamp 1486834041
transform 1 0 2688 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_50
timestamp 1486834041
transform 1 0 6272 0 -1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_66
timestamp 1486834041
transform 1 0 8064 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_72
timestamp 1486834041
transform 1 0 8736 0 -1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_88
timestamp 1486834041
transform 1 0 10528 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_96
timestamp 1486834041
transform 1 0 11424 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_136
timestamp 1486834041
transform 1 0 15904 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_142
timestamp 1486834041
transform 1 0 16576 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_174
timestamp 1486834041
transform 1 0 20160 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_182
timestamp 1486834041
transform 1 0 21056 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_206
timestamp 1486834041
transform 1 0 23744 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_212
timestamp 1486834041
transform 1 0 24416 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_244
timestamp 1486834041
transform 1 0 28000 0 -1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_260
timestamp 1486834041
transform 1 0 29792 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_268
timestamp 1486834041
transform 1 0 30688 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_277
timestamp 1486834041
transform 1 0 31696 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_279
timestamp 1486834041
transform 1 0 31920 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_282
timestamp 1486834041
transform 1 0 32256 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_290
timestamp 1486834041
transform 1 0 33152 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_294
timestamp 1486834041
transform 1 0 33600 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_316
timestamp 1486834041
transform 1 0 36064 0 -1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_332
timestamp 1486834041
transform 1 0 37856 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_336
timestamp 1486834041
transform 1 0 38304 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_352
timestamp 1486834041
transform 1 0 40096 0 -1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_416
timestamp 1486834041
transform 1 0 47264 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_422
timestamp 1486834041
transform 1 0 47936 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_454
timestamp 1486834041
transform 1 0 51520 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_456
timestamp 1486834041
transform 1 0 51744 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_465
timestamp 1486834041
transform 1 0 52752 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_467
timestamp 1486834041
transform 1 0 52976 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_492
timestamp 1486834041
transform 1 0 55776 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_496
timestamp 1486834041
transform 1 0 56224 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_498
timestamp 1486834041
transform 1 0 56448 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_18
timestamp 1486834041
transform 1 0 2688 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1486834041
transform 1 0 4480 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_37
timestamp 1486834041
transform 1 0 4816 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_81
timestamp 1486834041
transform 1 0 9744 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_89
timestamp 1486834041
transform 1 0 10640 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_93
timestamp 1486834041
transform 1 0 11088 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_95
timestamp 1486834041
transform 1 0 11312 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_100
timestamp 1486834041
transform 1 0 11872 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_104
timestamp 1486834041
transform 1 0 12320 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_107
timestamp 1486834041
transform 1 0 12656 0 1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_171
timestamp 1486834041
transform 1 0 19824 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_177
timestamp 1486834041
transform 1 0 20496 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_185
timestamp 1486834041
transform 1 0 21392 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_194
timestamp 1486834041
transform 1 0 22400 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_210
timestamp 1486834041
transform 1 0 24192 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_212
timestamp 1486834041
transform 1 0 24416 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_221
timestamp 1486834041
transform 1 0 25424 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_255
timestamp 1486834041
transform 1 0 29232 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_298
timestamp 1486834041
transform 1 0 34048 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_314
timestamp 1486834041
transform 1 0 35840 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_317
timestamp 1486834041
transform 1 0 36176 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_321
timestamp 1486834041
transform 1 0 36624 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_329
timestamp 1486834041
transform 1 0 37520 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_341
timestamp 1486834041
transform 1 0 38864 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_343
timestamp 1486834041
transform 1 0 39088 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_349
timestamp 1486834041
transform 1 0 39760 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_365
timestamp 1486834041
transform 1 0 41552 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_374
timestamp 1486834041
transform 1 0 42560 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_382
timestamp 1486834041
transform 1 0 43456 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_384
timestamp 1486834041
transform 1 0 43680 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_387
timestamp 1486834041
transform 1 0 44016 0 1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_419
timestamp 1486834041
transform 1 0 47600 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_427
timestamp 1486834041
transform 1 0 48496 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_429
timestamp 1486834041
transform 1 0 48720 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_438
timestamp 1486834041
transform 1 0 49728 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_454
timestamp 1486834041
transform 1 0 51520 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_26
timestamp 1486834041
transform 1 0 3584 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_58
timestamp 1486834041
transform 1 0 7168 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_66
timestamp 1486834041
transform 1 0 8064 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_72
timestamp 1486834041
transform 1 0 8736 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_80
timestamp 1486834041
transform 1 0 9632 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_84
timestamp 1486834041
transform 1 0 10080 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_86
timestamp 1486834041
transform 1 0 10304 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_107
timestamp 1486834041
transform 1 0 12656 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_139
timestamp 1486834041
transform 1 0 16240 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_150
timestamp 1486834041
transform 1 0 17472 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_154
timestamp 1486834041
transform 1 0 17920 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_156
timestamp 1486834041
transform 1 0 18144 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_165
timestamp 1486834041
transform 1 0 19152 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_201
timestamp 1486834041
transform 1 0 23184 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_209
timestamp 1486834041
transform 1 0 24080 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_232
timestamp 1486834041
transform 1 0 26656 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_264
timestamp 1486834041
transform 1 0 30240 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_282
timestamp 1486834041
transform 1 0 32256 0 -1 7056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_346
timestamp 1486834041
transform 1 0 39424 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_352
timestamp 1486834041
transform 1 0 40096 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_356
timestamp 1486834041
transform 1 0 40544 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_358
timestamp 1486834041
transform 1 0 40768 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_389
timestamp 1486834041
transform 1 0 44240 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_397
timestamp 1486834041
transform 1 0 45136 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_401
timestamp 1486834041
transform 1 0 45584 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_410
timestamp 1486834041
transform 1 0 46592 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_418
timestamp 1486834041
transform 1 0 47488 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_422
timestamp 1486834041
transform 1 0 47936 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_438
timestamp 1486834041
transform 1 0 49728 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_442
timestamp 1486834041
transform 1 0 50176 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_460
timestamp 1486834041
transform 1 0 52192 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_492
timestamp 1486834041
transform 1 0 55776 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_496
timestamp 1486834041
transform 1 0 56224 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_498
timestamp 1486834041
transform 1 0 56448 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1486834041
transform 1 0 4480 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_37
timestamp 1486834041
transform 1 0 4816 0 1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_53
timestamp 1486834041
transform 1 0 6608 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_61
timestamp 1486834041
transform 1 0 7504 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_85
timestamp 1486834041
transform 1 0 10192 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_93
timestamp 1486834041
transform 1 0 11088 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_97
timestamp 1486834041
transform 1 0 11536 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_99
timestamp 1486834041
transform 1 0 11760 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_107
timestamp 1486834041
transform 1 0 12656 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_111
timestamp 1486834041
transform 1 0 13104 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_121
timestamp 1486834041
transform 1 0 14224 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_129
timestamp 1486834041
transform 1 0 15120 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_133
timestamp 1486834041
transform 1 0 15568 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_155
timestamp 1486834041
transform 1 0 18032 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_174
timestamp 1486834041
transform 1 0 20160 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_177
timestamp 1486834041
transform 1 0 20496 0 1 7056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_241
timestamp 1486834041
transform 1 0 27664 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_262
timestamp 1486834041
transform 1 0 30016 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_294
timestamp 1486834041
transform 1 0 33600 0 1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_310
timestamp 1486834041
transform 1 0 35392 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_314
timestamp 1486834041
transform 1 0 35840 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_349
timestamp 1486834041
transform 1 0 39760 0 1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_365
timestamp 1486834041
transform 1 0 41552 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_381
timestamp 1486834041
transform 1 0 43344 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_387
timestamp 1486834041
transform 1 0 44016 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_419
timestamp 1486834041
transform 1 0 47600 0 1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_435
timestamp 1486834041
transform 1 0 49392 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_40
timestamp 1486834041
transform 1 0 5152 0 -1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_56
timestamp 1486834041
transform 1 0 6944 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_60
timestamp 1486834041
transform 1 0 7392 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_72
timestamp 1486834041
transform 1 0 8736 0 -1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_104
timestamp 1486834041
transform 1 0 12320 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_129
timestamp 1486834041
transform 1 0 15120 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_137
timestamp 1486834041
transform 1 0 16016 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_139
timestamp 1486834041
transform 1 0 16240 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_142
timestamp 1486834041
transform 1 0 16576 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_150
timestamp 1486834041
transform 1 0 17472 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_154
timestamp 1486834041
transform 1 0 17920 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_156
timestamp 1486834041
transform 1 0 18144 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_166
timestamp 1486834041
transform 1 0 19264 0 -1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_198
timestamp 1486834041
transform 1 0 22848 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_206
timestamp 1486834041
transform 1 0 23744 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_212
timestamp 1486834041
transform 1 0 24416 0 -1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_228
timestamp 1486834041
transform 1 0 26208 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_236
timestamp 1486834041
transform 1 0 27104 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_240
timestamp 1486834041
transform 1 0 27552 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_242
timestamp 1486834041
transform 1 0 27776 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_259
timestamp 1486834041
transform 1 0 29680 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_267
timestamp 1486834041
transform 1 0 30576 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_279
timestamp 1486834041
transform 1 0 31920 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_282
timestamp 1486834041
transform 1 0 32256 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_290
timestamp 1486834041
transform 1 0 33152 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_300
timestamp 1486834041
transform 1 0 34272 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_324
timestamp 1486834041
transform 1 0 36960 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_328
timestamp 1486834041
transform 1 0 37408 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_345
timestamp 1486834041
transform 1 0 39312 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_349
timestamp 1486834041
transform 1 0 39760 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_352
timestamp 1486834041
transform 1 0 40096 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_373
timestamp 1486834041
transform 1 0 42448 0 -1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_405
timestamp 1486834041
transform 1 0 46032 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_413
timestamp 1486834041
transform 1 0 46928 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_417
timestamp 1486834041
transform 1 0 47376 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_419
timestamp 1486834041
transform 1 0 47600 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_422
timestamp 1486834041
transform 1 0 47936 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_430
timestamp 1486834041
transform 1 0 48832 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_434
timestamp 1486834041
transform 1 0 49280 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_436
timestamp 1486834041
transform 1 0 49504 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_445
timestamp 1486834041
transform 1 0 50512 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_447
timestamp 1486834041
transform 1 0 50736 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_492
timestamp 1486834041
transform 1 0 55776 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_496
timestamp 1486834041
transform 1 0 56224 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_498
timestamp 1486834041
transform 1 0 56448 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_2
timestamp 1486834041
transform 1 0 896 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_4
timestamp 1486834041
transform 1 0 1120 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_53
timestamp 1486834041
transform 1 0 6608 0 1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_69
timestamp 1486834041
transform 1 0 8400 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_77
timestamp 1486834041
transform 1 0 9296 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_89
timestamp 1486834041
transform 1 0 10640 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_107
timestamp 1486834041
transform 1 0 12656 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_116
timestamp 1486834041
transform 1 0 13664 0 1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_148
timestamp 1486834041
transform 1 0 17248 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_152
timestamp 1486834041
transform 1 0 17696 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_162
timestamp 1486834041
transform 1 0 18816 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_170
timestamp 1486834041
transform 1 0 19712 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_174
timestamp 1486834041
transform 1 0 20160 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_177
timestamp 1486834041
transform 1 0 20496 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_179
timestamp 1486834041
transform 1 0 20720 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_212
timestamp 1486834041
transform 1 0 24416 0 1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_228
timestamp 1486834041
transform 1 0 26208 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_230
timestamp 1486834041
transform 1 0 26432 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_239
timestamp 1486834041
transform 1 0 27440 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_243
timestamp 1486834041
transform 1 0 27888 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_247
timestamp 1486834041
transform 1 0 28336 0 1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_263
timestamp 1486834041
transform 1 0 30128 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_271
timestamp 1486834041
transform 1 0 31024 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_287
timestamp 1486834041
transform 1 0 32816 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_309
timestamp 1486834041
transform 1 0 35280 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_313
timestamp 1486834041
transform 1 0 35728 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_325
timestamp 1486834041
transform 1 0 37072 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_341
timestamp 1486834041
transform 1 0 38864 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_345
timestamp 1486834041
transform 1 0 39312 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_354
timestamp 1486834041
transform 1 0 40320 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_360
timestamp 1486834041
transform 1 0 40992 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_387
timestamp 1486834041
transform 1 0 44016 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_395
timestamp 1486834041
transform 1 0 44912 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_407
timestamp 1486834041
transform 1 0 46256 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_415
timestamp 1486834041
transform 1 0 47152 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_2
timestamp 1486834041
transform 1 0 896 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_6
timestamp 1486834041
transform 1 0 1344 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_8
timestamp 1486834041
transform 1 0 1568 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_23
timestamp 1486834041
transform 1 0 3248 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_27
timestamp 1486834041
transform 1 0 3696 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_43
timestamp 1486834041
transform 1 0 5488 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_47
timestamp 1486834041
transform 1 0 5936 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_63
timestamp 1486834041
transform 1 0 7728 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_67
timestamp 1486834041
transform 1 0 8176 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_69
timestamp 1486834041
transform 1 0 8400 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_72
timestamp 1486834041
transform 1 0 8736 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_74
timestamp 1486834041
transform 1 0 8960 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_103
timestamp 1486834041
transform 1 0 12208 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_107
timestamp 1486834041
transform 1 0 12656 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_116
timestamp 1486834041
transform 1 0 13664 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_131
timestamp 1486834041
transform 1 0 15344 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_139
timestamp 1486834041
transform 1 0 16240 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_142
timestamp 1486834041
transform 1 0 16576 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_146
timestamp 1486834041
transform 1 0 17024 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_164
timestamp 1486834041
transform 1 0 19040 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_172
timestamp 1486834041
transform 1 0 19936 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_184
timestamp 1486834041
transform 1 0 21280 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_193
timestamp 1486834041
transform 1 0 22288 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_201
timestamp 1486834041
transform 1 0 23184 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_212
timestamp 1486834041
transform 1 0 24416 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_216
timestamp 1486834041
transform 1 0 24864 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_225
timestamp 1486834041
transform 1 0 25872 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_229
timestamp 1486834041
transform 1 0 26320 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_245
timestamp 1486834041
transform 1 0 28112 0 -1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_269
timestamp 1486834041
transform 1 0 30800 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_277
timestamp 1486834041
transform 1 0 31696 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_279
timestamp 1486834041
transform 1 0 31920 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_282
timestamp 1486834041
transform 1 0 32256 0 -1 10192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_346
timestamp 1486834041
transform 1 0 39424 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_352
timestamp 1486834041
transform 1 0 40096 0 -1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_368
timestamp 1486834041
transform 1 0 41888 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_376
timestamp 1486834041
transform 1 0 42784 0 -1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_392
timestamp 1486834041
transform 1 0 44576 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_400
timestamp 1486834041
transform 1 0 45472 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_404
timestamp 1486834041
transform 1 0 45920 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_406
timestamp 1486834041
transform 1 0 46144 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_415
timestamp 1486834041
transform 1 0 47152 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_419
timestamp 1486834041
transform 1 0 47600 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_422
timestamp 1486834041
transform 1 0 47936 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_492
timestamp 1486834041
transform 1 0 55776 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_496
timestamp 1486834041
transform 1 0 56224 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_498
timestamp 1486834041
transform 1 0 56448 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_2
timestamp 1486834041
transform 1 0 896 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_6
timestamp 1486834041
transform 1 0 1344 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_45
timestamp 1486834041
transform 1 0 5712 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_47
timestamp 1486834041
transform 1 0 5936 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_104
timestamp 1486834041
transform 1 0 12320 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_107
timestamp 1486834041
transform 1 0 12656 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_111
timestamp 1486834041
transform 1 0 13104 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_163
timestamp 1486834041
transform 1 0 18928 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_177
timestamp 1486834041
transform 1 0 20496 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_195
timestamp 1486834041
transform 1 0 22512 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_199
timestamp 1486834041
transform 1 0 22960 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_247
timestamp 1486834041
transform 1 0 28336 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_255
timestamp 1486834041
transform 1 0 29232 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_279
timestamp 1486834041
transform 1 0 31920 0 1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_295
timestamp 1486834041
transform 1 0 33712 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_299
timestamp 1486834041
transform 1 0 34160 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_308
timestamp 1486834041
transform 1 0 35168 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_312
timestamp 1486834041
transform 1 0 35616 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_314
timestamp 1486834041
transform 1 0 35840 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_317
timestamp 1486834041
transform 1 0 36176 0 1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_349
timestamp 1486834041
transform 1 0 39760 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_353
timestamp 1486834041
transform 1 0 40208 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_375
timestamp 1486834041
transform 1 0 42672 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_383
timestamp 1486834041
transform 1 0 43568 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_387
timestamp 1486834041
transform 1 0 44016 0 1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_403
timestamp 1486834041
transform 1 0 45808 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_10
timestamp 1486834041
transform 1 0 1792 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_72
timestamp 1486834041
transform 1 0 8736 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_74
timestamp 1486834041
transform 1 0 8960 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_83
timestamp 1486834041
transform 1 0 9968 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_142
timestamp 1486834041
transform 1 0 16576 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_199
timestamp 1486834041
transform 1 0 22960 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_201
timestamp 1486834041
transform 1 0 23184 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_212
timestamp 1486834041
transform 1 0 24416 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_216
timestamp 1486834041
transform 1 0 24864 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_247
timestamp 1486834041
transform 1 0 28336 0 -1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_263
timestamp 1486834041
transform 1 0 30128 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_271
timestamp 1486834041
transform 1 0 31024 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_290
timestamp 1486834041
transform 1 0 33152 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_334
timestamp 1486834041
transform 1 0 38080 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_344
timestamp 1486834041
transform 1 0 39200 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_348
timestamp 1486834041
transform 1 0 39648 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_352
timestamp 1486834041
transform 1 0 40096 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_356
timestamp 1486834041
transform 1 0 40544 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_372
timestamp 1486834041
transform 1 0 42336 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_397
timestamp 1486834041
transform 1 0 45136 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_401
timestamp 1486834041
transform 1 0 45584 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_403
timestamp 1486834041
transform 1 0 45808 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_422
timestamp 1486834041
transform 1 0 47936 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_487
timestamp 1486834041
transform 1 0 55216 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_489
timestamp 1486834041
transform 1 0 55440 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_492
timestamp 1486834041
transform 1 0 55776 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_496
timestamp 1486834041
transform 1 0 56224 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_498
timestamp 1486834041
transform 1 0 56448 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_2
timestamp 1486834041
transform 1 0 896 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_6
timestamp 1486834041
transform 1 0 1344 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_45
timestamp 1486834041
transform 1 0 5712 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_107
timestamp 1486834041
transform 1 0 12656 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_177
timestamp 1486834041
transform 1 0 20496 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_241
timestamp 1486834041
transform 1 0 27664 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_247
timestamp 1486834041
transform 1 0 28336 0 1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_263
timestamp 1486834041
transform 1 0 30128 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_313
timestamp 1486834041
transform 1 0 35728 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_325
timestamp 1486834041
transform 1 0 37072 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_349
timestamp 1486834041
transform 1 0 39760 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_357
timestamp 1486834041
transform 1 0 40656 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_361
timestamp 1486834041
transform 1 0 41104 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_378
timestamp 1486834041
transform 1 0 43008 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_382
timestamp 1486834041
transform 1 0 43456 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_384
timestamp 1486834041
transform 1 0 43680 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_411
timestamp 1486834041
transform 1 0 46704 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_451
timestamp 1486834041
transform 1 0 51184 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_2
timestamp 1486834041
transform 1 0 896 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_36
timestamp 1486834041
transform 1 0 4704 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_70
timestamp 1486834041
transform 1 0 8512 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_104
timestamp 1486834041
transform 1 0 12320 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_138
timestamp 1486834041
transform 1 0 16128 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_172
timestamp 1486834041
transform 1 0 19936 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_220
timestamp 1486834041
transform 1 0 25312 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_240
timestamp 1486834041
transform 1 0 27552 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_257
timestamp 1486834041
transform 1 0 29456 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_269
timestamp 1486834041
transform 1 0 30800 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_271
timestamp 1486834041
transform 1 0 31024 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_342
timestamp 1486834041
transform 1 0 38976 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_350
timestamp 1486834041
transform 1 0 39872 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_354
timestamp 1486834041
transform 1 0 40320 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_356
timestamp 1486834041
transform 1 0 40544 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_373
timestamp 1486834041
transform 1 0 42448 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_392
timestamp 1486834041
transform 1 0 44576 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_410
timestamp 1486834041
transform 1 0 46592 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_439
timestamp 1486834041
transform 1 0 49840 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_441
timestamp 1486834041
transform 1 0 50064 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_472
timestamp 1486834041
transform 1 0 53536 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_492
timestamp 1486834041
transform 1 0 55776 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_496
timestamp 1486834041
transform 1 0 56224 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_498
timestamp 1486834041
transform 1 0 56448 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input1
timestamp 1486834041
transform 1 0 3472 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input2
timestamp 1486834041
transform 1 0 1792 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input3
timestamp 1486834041
transform 1 0 896 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input4
timestamp 1486834041
transform 1 0 1792 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input5
timestamp 1486834041
transform 1 0 896 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input6
timestamp 1486834041
transform 1 0 896 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input7
timestamp 1486834041
transform 1 0 2464 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input8
timestamp 1486834041
transform 1 0 2800 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input9
timestamp 1486834041
transform 1 0 896 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input10
timestamp 1486834041
transform 1 0 3696 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input11
timestamp 1486834041
transform 1 0 4816 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input12
timestamp 1486834041
transform 1 0 2688 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input13
timestamp 1486834041
transform 1 0 896 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input14
timestamp 1486834041
transform 1 0 1792 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input15
timestamp 1486834041
transform 1 0 2688 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input16
timestamp 1486834041
transform 1 0 4256 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input17
timestamp 1486834041
transform 1 0 3584 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input18
timestamp 1486834041
transform 1 0 896 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input19
timestamp 1486834041
transform 1 0 5712 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input20
timestamp 1486834041
transform 1 0 1792 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input21
timestamp 1486834041
transform 1 0 1456 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input22
timestamp 1486834041
transform -1 0 24976 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input23
timestamp 1486834041
transform 1 0 24976 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input24
timestamp 1486834041
transform 1 0 24976 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input25
timestamp 1486834041
transform -1 0 25872 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input26
timestamp 1486834041
transform 1 0 29904 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input27
timestamp 1486834041
transform 1 0 30352 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input28
timestamp 1486834041
transform 1 0 31360 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input29
timestamp 1486834041
transform 1 0 32256 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input30
timestamp 1486834041
transform 1 0 33152 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input31
timestamp 1486834041
transform 1 0 32256 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input32
timestamp 1486834041
transform 1 0 33040 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input33
timestamp 1486834041
transform 1 0 34048 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input34
timestamp 1486834041
transform 1 0 28560 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input35
timestamp 1486834041
transform -1 0 26432 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input36
timestamp 1486834041
transform -1 0 27328 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input37
timestamp 1486834041
transform 1 0 27664 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input38
timestamp 1486834041
transform 1 0 33936 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input39
timestamp 1486834041
transform 1 0 35168 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input40
timestamp 1486834041
transform 1 0 34832 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input41
timestamp 1486834041
transform 1 0 36064 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input42
timestamp 1486834041
transform 1 0 36960 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input43
timestamp 1486834041
transform 1 0 37856 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input44
timestamp 1486834041
transform 1 0 36288 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input45
timestamp 1486834041
transform 1 0 37184 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input46
timestamp 1486834041
transform 1 0 40656 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input47
timestamp 1486834041
transform 1 0 41552 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input48
timestamp 1486834041
transform 1 0 42784 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input49
timestamp 1486834041
transform 1 0 43680 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input50
timestamp 1486834041
transform 1 0 42448 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input51
timestamp 1486834041
transform 1 0 44016 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input52
timestamp 1486834041
transform 1 0 43344 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input53
timestamp 1486834041
transform 1 0 44240 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output54
timestamp 1486834041
transform -1 0 15120 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output55
timestamp 1486834041
transform 1 0 51856 0 1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output56
timestamp 1486834041
transform 1 0 53424 0 1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output57
timestamp 1486834041
transform 1 0 53984 0 -1 5488
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output58
timestamp 1486834041
transform 1 0 54992 0 1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output59
timestamp 1486834041
transform 1 0 53424 0 1 5488
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output60
timestamp 1486834041
transform 1 0 53984 0 -1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output61
timestamp 1486834041
transform 1 0 54992 0 1 5488
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output62
timestamp 1486834041
transform 1 0 53424 0 1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output63
timestamp 1486834041
transform 1 0 54992 0 1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output64
timestamp 1486834041
transform 1 0 54992 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output65
timestamp 1486834041
transform 1 0 53424 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output66
timestamp 1486834041
transform 1 0 52416 0 -1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output67
timestamp 1486834041
transform 1 0 54992 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output68
timestamp 1486834041
transform 1 0 53984 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output69
timestamp 1486834041
transform 1 0 53424 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output70
timestamp 1486834041
transform 1 0 53984 0 -1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output71
timestamp 1486834041
transform 1 0 50848 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output72
timestamp 1486834041
transform 1 0 52416 0 -1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output73
timestamp 1486834041
transform 1 0 48048 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output74
timestamp 1486834041
transform 1 0 51856 0 1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output75
timestamp 1486834041
transform 1 0 50848 0 -1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output76
timestamp 1486834041
transform 1 0 48496 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output77
timestamp 1486834041
transform 1 0 50848 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output78
timestamp 1486834041
transform 1 0 49280 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output79
timestamp 1486834041
transform 1 0 50064 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output80
timestamp 1486834041
transform 1 0 52416 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output81
timestamp 1486834041
transform 1 0 52416 0 -1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output82
timestamp 1486834041
transform 1 0 53984 0 -1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output83
timestamp 1486834041
transform 1 0 54992 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output84
timestamp 1486834041
transform 1 0 53424 0 1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output85
timestamp 1486834041
transform 1 0 53984 0 -1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output86
timestamp 1486834041
transform 1 0 54992 0 1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output87
timestamp 1486834041
transform 1 0 48272 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output88
timestamp 1486834041
transform 1 0 52752 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output89
timestamp 1486834041
transform 1 0 54992 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output90
timestamp 1486834041
transform 1 0 52416 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output91
timestamp 1486834041
transform 1 0 51856 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output92
timestamp 1486834041
transform -1 0 51632 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output93
timestamp 1486834041
transform 1 0 46704 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output94
timestamp 1486834041
transform -1 0 48720 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output95
timestamp 1486834041
transform 1 0 52416 0 -1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output96
timestamp 1486834041
transform 1 0 44800 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output97
timestamp 1486834041
transform 1 0 51856 0 1 5488
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output98
timestamp 1486834041
transform -1 0 50288 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output99
timestamp 1486834041
transform 1 0 50400 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output100
timestamp 1486834041
transform 1 0 49616 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output101
timestamp 1486834041
transform 1 0 51968 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output102
timestamp 1486834041
transform 1 0 51856 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output103
timestamp 1486834041
transform 1 0 51184 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output104
timestamp 1486834041
transform 1 0 51856 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output105
timestamp 1486834041
transform 1 0 53424 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output106
timestamp 1486834041
transform 1 0 54208 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output107
timestamp 1486834041
transform -1 0 2464 0 -1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output108
timestamp 1486834041
transform -1 0 2800 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output109
timestamp 1486834041
transform -1 0 3248 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output110
timestamp 1486834041
transform -1 0 3024 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output111
timestamp 1486834041
transform -1 0 3808 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output112
timestamp 1486834041
transform -1 0 4592 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output113
timestamp 1486834041
transform -1 0 3024 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output114
timestamp 1486834041
transform -1 0 5488 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output115
timestamp 1486834041
transform -1 0 2912 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output116
timestamp 1486834041
transform -1 0 4592 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output117
timestamp 1486834041
transform -1 0 5376 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output118
timestamp 1486834041
transform -1 0 4480 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output119
timestamp 1486834041
transform -1 0 7728 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output120
timestamp 1486834041
transform -1 0 7616 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output121
timestamp 1486834041
transform -1 0 6944 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output122
timestamp 1486834041
transform -1 0 6720 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output123
timestamp 1486834041
transform -1 0 9184 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output124
timestamp 1486834041
transform -1 0 7728 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output125
timestamp 1486834041
transform -1 0 8512 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output126
timestamp 1486834041
transform -1 0 10640 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output127
timestamp 1486834041
transform -1 0 8288 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output128
timestamp 1486834041
transform -1 0 14784 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output129
timestamp 1486834041
transform 1 0 14112 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output130
timestamp 1486834041
transform -1 0 14336 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output131
timestamp 1486834041
transform -1 0 16352 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output132
timestamp 1486834041
transform -1 0 15568 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output133
timestamp 1486834041
transform 1 0 15680 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output134
timestamp 1486834041
transform -1 0 9296 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output135
timestamp 1486834041
transform -1 0 12208 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output136
timestamp 1486834041
transform -1 0 10864 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output137
timestamp 1486834041
transform -1 0 11648 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output138
timestamp 1486834041
transform -1 0 10528 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output139
timestamp 1486834041
transform -1 0 13216 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output140
timestamp 1486834041
transform 1 0 10864 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output141
timestamp 1486834041
transform -1 0 12096 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output142
timestamp 1486834041
transform -1 0 15344 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output143
timestamp 1486834041
transform -1 0 15904 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output144
timestamp 1486834041
transform -1 0 22960 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output145
timestamp 1486834041
transform 1 0 20384 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output146
timestamp 1486834041
transform -1 0 23184 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output147
timestamp 1486834041
transform 1 0 21952 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output148
timestamp 1486834041
transform -1 0 24752 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output149
timestamp 1486834041
transform 1 0 23744 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output150
timestamp 1486834041
transform -1 0 17136 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output151
timestamp 1486834041
transform -1 0 18256 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output152
timestamp 1486834041
transform -1 0 18704 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output153
timestamp 1486834041
transform -1 0 18144 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output154
timestamp 1486834041
transform -1 0 19824 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output155
timestamp 1486834041
transform -1 0 20272 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output156
timestamp 1486834041
transform -1 0 19712 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output157
timestamp 1486834041
transform -1 0 21392 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output158
timestamp 1486834041
transform 1 0 20944 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output159
timestamp 1486834041
transform -1 0 6720 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output160
timestamp 1486834041
transform -1 0 8288 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output161
timestamp 1486834041
transform -1 0 11088 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output162
timestamp 1486834041
transform -1 0 13104 0 -1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output163
timestamp 1486834041
transform -1 0 48272 0 1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_16
timestamp 1486834041
transform 1 0 672 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1486834041
transform -1 0 56784 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_17
timestamp 1486834041
transform 1 0 672 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1486834041
transform -1 0 56784 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_18
timestamp 1486834041
transform 1 0 672 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1486834041
transform -1 0 56784 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_19
timestamp 1486834041
transform 1 0 672 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1486834041
transform -1 0 56784 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_20
timestamp 1486834041
transform 1 0 672 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1486834041
transform -1 0 56784 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_21
timestamp 1486834041
transform 1 0 672 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1486834041
transform -1 0 56784 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_22
timestamp 1486834041
transform 1 0 672 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1486834041
transform -1 0 56784 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_23
timestamp 1486834041
transform 1 0 672 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1486834041
transform -1 0 56784 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_24
timestamp 1486834041
transform 1 0 672 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1486834041
transform -1 0 56784 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_25
timestamp 1486834041
transform 1 0 672 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1486834041
transform -1 0 56784 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_26
timestamp 1486834041
transform 1 0 672 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1486834041
transform -1 0 56784 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_27
timestamp 1486834041
transform 1 0 672 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1486834041
transform -1 0 56784 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_28
timestamp 1486834041
transform 1 0 672 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1486834041
transform -1 0 56784 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_29
timestamp 1486834041
transform 1 0 672 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1486834041
transform -1 0 56784 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_30
timestamp 1486834041
transform 1 0 672 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1486834041
transform -1 0 56784 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_31
timestamp 1486834041
transform 1 0 672 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1486834041
transform -1 0 56784 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  S_WARMBOOT_164
timestamp 1486834041
transform -1 0 25200 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_32
timestamp 1486834041
transform 1 0 4480 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_33
timestamp 1486834041
transform 1 0 8288 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_34
timestamp 1486834041
transform 1 0 12096 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_35
timestamp 1486834041
transform 1 0 15904 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_36
timestamp 1486834041
transform 1 0 19712 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_37
timestamp 1486834041
transform 1 0 23520 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_38
timestamp 1486834041
transform 1 0 27328 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_39
timestamp 1486834041
transform 1 0 31136 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_40
timestamp 1486834041
transform 1 0 34944 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_41
timestamp 1486834041
transform 1 0 38752 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_42
timestamp 1486834041
transform 1 0 42560 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_43
timestamp 1486834041
transform 1 0 46368 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_44
timestamp 1486834041
transform 1 0 50176 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_45
timestamp 1486834041
transform 1 0 53984 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_46
timestamp 1486834041
transform 1 0 8512 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_47
timestamp 1486834041
transform 1 0 16352 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_48
timestamp 1486834041
transform 1 0 24192 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_49
timestamp 1486834041
transform 1 0 32032 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_50
timestamp 1486834041
transform 1 0 39872 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_51
timestamp 1486834041
transform 1 0 47712 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_52
timestamp 1486834041
transform 1 0 55552 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_53
timestamp 1486834041
transform 1 0 4592 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_54
timestamp 1486834041
transform 1 0 12432 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_55
timestamp 1486834041
transform 1 0 20272 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_56
timestamp 1486834041
transform 1 0 28112 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_57
timestamp 1486834041
transform 1 0 35952 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_58
timestamp 1486834041
transform 1 0 43792 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_59
timestamp 1486834041
transform 1 0 51632 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_60
timestamp 1486834041
transform 1 0 8512 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_61
timestamp 1486834041
transform 1 0 16352 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_62
timestamp 1486834041
transform 1 0 24192 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_63
timestamp 1486834041
transform 1 0 32032 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_64
timestamp 1486834041
transform 1 0 39872 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_65
timestamp 1486834041
transform 1 0 47712 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_66
timestamp 1486834041
transform 1 0 55552 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_67
timestamp 1486834041
transform 1 0 4592 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_68
timestamp 1486834041
transform 1 0 12432 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_69
timestamp 1486834041
transform 1 0 20272 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_70
timestamp 1486834041
transform 1 0 28112 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_71
timestamp 1486834041
transform 1 0 35952 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_72
timestamp 1486834041
transform 1 0 43792 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_73
timestamp 1486834041
transform 1 0 51632 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_74
timestamp 1486834041
transform 1 0 8512 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_75
timestamp 1486834041
transform 1 0 16352 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_76
timestamp 1486834041
transform 1 0 24192 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_77
timestamp 1486834041
transform 1 0 32032 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_78
timestamp 1486834041
transform 1 0 39872 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_79
timestamp 1486834041
transform 1 0 47712 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_80
timestamp 1486834041
transform 1 0 55552 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_81
timestamp 1486834041
transform 1 0 4592 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_82
timestamp 1486834041
transform 1 0 12432 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_83
timestamp 1486834041
transform 1 0 20272 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_84
timestamp 1486834041
transform 1 0 28112 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_85
timestamp 1486834041
transform 1 0 35952 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_86
timestamp 1486834041
transform 1 0 43792 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_87
timestamp 1486834041
transform 1 0 51632 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_88
timestamp 1486834041
transform 1 0 8512 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_89
timestamp 1486834041
transform 1 0 16352 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_90
timestamp 1486834041
transform 1 0 24192 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_91
timestamp 1486834041
transform 1 0 32032 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_92
timestamp 1486834041
transform 1 0 39872 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_93
timestamp 1486834041
transform 1 0 47712 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_94
timestamp 1486834041
transform 1 0 55552 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_95
timestamp 1486834041
transform 1 0 4592 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_96
timestamp 1486834041
transform 1 0 12432 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_97
timestamp 1486834041
transform 1 0 20272 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_98
timestamp 1486834041
transform 1 0 28112 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_99
timestamp 1486834041
transform 1 0 35952 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_100
timestamp 1486834041
transform 1 0 43792 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_101
timestamp 1486834041
transform 1 0 51632 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_102
timestamp 1486834041
transform 1 0 8512 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_103
timestamp 1486834041
transform 1 0 16352 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_104
timestamp 1486834041
transform 1 0 24192 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_105
timestamp 1486834041
transform 1 0 32032 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_106
timestamp 1486834041
transform 1 0 39872 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_107
timestamp 1486834041
transform 1 0 47712 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_108
timestamp 1486834041
transform 1 0 55552 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_109
timestamp 1486834041
transform 1 0 4592 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_110
timestamp 1486834041
transform 1 0 12432 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_111
timestamp 1486834041
transform 1 0 20272 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_112
timestamp 1486834041
transform 1 0 28112 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_113
timestamp 1486834041
transform 1 0 35952 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_114
timestamp 1486834041
transform 1 0 43792 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_115
timestamp 1486834041
transform 1 0 51632 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_116
timestamp 1486834041
transform 1 0 8512 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_117
timestamp 1486834041
transform 1 0 16352 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_118
timestamp 1486834041
transform 1 0 24192 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_119
timestamp 1486834041
transform 1 0 32032 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_120
timestamp 1486834041
transform 1 0 39872 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_121
timestamp 1486834041
transform 1 0 47712 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_122
timestamp 1486834041
transform 1 0 55552 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_123
timestamp 1486834041
transform 1 0 4592 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_124
timestamp 1486834041
transform 1 0 12432 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_125
timestamp 1486834041
transform 1 0 20272 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_126
timestamp 1486834041
transform 1 0 28112 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_127
timestamp 1486834041
transform 1 0 35952 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_128
timestamp 1486834041
transform 1 0 43792 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_129
timestamp 1486834041
transform 1 0 51632 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_130
timestamp 1486834041
transform 1 0 8512 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_131
timestamp 1486834041
transform 1 0 16352 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_132
timestamp 1486834041
transform 1 0 24192 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_133
timestamp 1486834041
transform 1 0 32032 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_134
timestamp 1486834041
transform 1 0 39872 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_135
timestamp 1486834041
transform 1 0 47712 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_136
timestamp 1486834041
transform 1 0 55552 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_137
timestamp 1486834041
transform 1 0 4592 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_138
timestamp 1486834041
transform 1 0 12432 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_139
timestamp 1486834041
transform 1 0 20272 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_140
timestamp 1486834041
transform 1 0 28112 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_141
timestamp 1486834041
transform 1 0 35952 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_142
timestamp 1486834041
transform 1 0 43792 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_143
timestamp 1486834041
transform 1 0 51632 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_144
timestamp 1486834041
transform 1 0 4480 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_145
timestamp 1486834041
transform 1 0 8288 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_146
timestamp 1486834041
transform 1 0 12096 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_147
timestamp 1486834041
transform 1 0 15904 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_148
timestamp 1486834041
transform 1 0 19712 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_149
timestamp 1486834041
transform 1 0 23520 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_150
timestamp 1486834041
transform 1 0 27328 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_151
timestamp 1486834041
transform 1 0 31136 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_152
timestamp 1486834041
transform 1 0 34944 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_153
timestamp 1486834041
transform 1 0 38752 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_154
timestamp 1486834041
transform 1 0 42560 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_155
timestamp 1486834041
transform 1 0 46368 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_156
timestamp 1486834041
transform 1 0 50176 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_157
timestamp 1486834041
transform 1 0 53984 0 -1 13328
box -86 -86 310 870
<< labels >>
flabel metal2 s 13440 0 13552 112 0 FreeSans 448 0 0 0 BOOT_top
port 0 nsew signal output
flabel metal2 s 3360 0 3472 112 0 FreeSans 448 0 0 0 CONFIGURED_top
port 1 nsew signal input
flabel metal2 s 23968 14112 24080 14224 0 FreeSans 448 0 0 0 Co
port 2 nsew signal output
flabel metal3 s 0 0 112 112 0 FreeSans 448 0 0 0 FrameData[0]
port 3 nsew signal input
flabel metal3 s 0 4480 112 4592 0 FreeSans 448 0 0 0 FrameData[10]
port 4 nsew signal input
flabel metal3 s 0 4928 112 5040 0 FreeSans 448 0 0 0 FrameData[11]
port 5 nsew signal input
flabel metal3 s 0 5376 112 5488 0 FreeSans 448 0 0 0 FrameData[12]
port 6 nsew signal input
flabel metal3 s 0 5824 112 5936 0 FreeSans 448 0 0 0 FrameData[13]
port 7 nsew signal input
flabel metal3 s 0 6272 112 6384 0 FreeSans 448 0 0 0 FrameData[14]
port 8 nsew signal input
flabel metal3 s 0 6720 112 6832 0 FreeSans 448 0 0 0 FrameData[15]
port 9 nsew signal input
flabel metal3 s 0 7168 112 7280 0 FreeSans 448 0 0 0 FrameData[16]
port 10 nsew signal input
flabel metal3 s 0 7616 112 7728 0 FreeSans 448 0 0 0 FrameData[17]
port 11 nsew signal input
flabel metal3 s 0 8064 112 8176 0 FreeSans 448 0 0 0 FrameData[18]
port 12 nsew signal input
flabel metal3 s 0 8512 112 8624 0 FreeSans 448 0 0 0 FrameData[19]
port 13 nsew signal input
flabel metal3 s 0 448 112 560 0 FreeSans 448 0 0 0 FrameData[1]
port 14 nsew signal input
flabel metal3 s 0 8960 112 9072 0 FreeSans 448 0 0 0 FrameData[20]
port 15 nsew signal input
flabel metal3 s 0 9408 112 9520 0 FreeSans 448 0 0 0 FrameData[21]
port 16 nsew signal input
flabel metal3 s 0 9856 112 9968 0 FreeSans 448 0 0 0 FrameData[22]
port 17 nsew signal input
flabel metal3 s 0 10304 112 10416 0 FreeSans 448 0 0 0 FrameData[23]
port 18 nsew signal input
flabel metal3 s 0 10752 112 10864 0 FreeSans 448 0 0 0 FrameData[24]
port 19 nsew signal input
flabel metal3 s 0 11200 112 11312 0 FreeSans 448 0 0 0 FrameData[25]
port 20 nsew signal input
flabel metal3 s 0 11648 112 11760 0 FreeSans 448 0 0 0 FrameData[26]
port 21 nsew signal input
flabel metal3 s 0 12096 112 12208 0 FreeSans 448 0 0 0 FrameData[27]
port 22 nsew signal input
flabel metal3 s 0 12544 112 12656 0 FreeSans 448 0 0 0 FrameData[28]
port 23 nsew signal input
flabel metal3 s 0 12992 112 13104 0 FreeSans 448 0 0 0 FrameData[29]
port 24 nsew signal input
flabel metal3 s 0 896 112 1008 0 FreeSans 448 0 0 0 FrameData[2]
port 25 nsew signal input
flabel metal3 s 0 13440 112 13552 0 FreeSans 448 0 0 0 FrameData[30]
port 26 nsew signal input
flabel metal3 s 0 13888 112 14000 0 FreeSans 448 0 0 0 FrameData[31]
port 27 nsew signal input
flabel metal3 s 0 1344 112 1456 0 FreeSans 448 0 0 0 FrameData[3]
port 28 nsew signal input
flabel metal3 s 0 1792 112 1904 0 FreeSans 448 0 0 0 FrameData[4]
port 29 nsew signal input
flabel metal3 s 0 2240 112 2352 0 FreeSans 448 0 0 0 FrameData[5]
port 30 nsew signal input
flabel metal3 s 0 2688 112 2800 0 FreeSans 448 0 0 0 FrameData[6]
port 31 nsew signal input
flabel metal3 s 0 3136 112 3248 0 FreeSans 448 0 0 0 FrameData[7]
port 32 nsew signal input
flabel metal3 s 0 3584 112 3696 0 FreeSans 448 0 0 0 FrameData[8]
port 33 nsew signal input
flabel metal3 s 0 4032 112 4144 0 FreeSans 448 0 0 0 FrameData[9]
port 34 nsew signal input
flabel metal3 s 57344 0 57456 112 0 FreeSans 448 0 0 0 FrameData_O[0]
port 35 nsew signal output
flabel metal3 s 57344 4480 57456 4592 0 FreeSans 448 0 0 0 FrameData_O[10]
port 36 nsew signal output
flabel metal3 s 57344 4928 57456 5040 0 FreeSans 448 0 0 0 FrameData_O[11]
port 37 nsew signal output
flabel metal3 s 57344 5376 57456 5488 0 FreeSans 448 0 0 0 FrameData_O[12]
port 38 nsew signal output
flabel metal3 s 57344 5824 57456 5936 0 FreeSans 448 0 0 0 FrameData_O[13]
port 39 nsew signal output
flabel metal3 s 57344 6272 57456 6384 0 FreeSans 448 0 0 0 FrameData_O[14]
port 40 nsew signal output
flabel metal3 s 57344 6720 57456 6832 0 FreeSans 448 0 0 0 FrameData_O[15]
port 41 nsew signal output
flabel metal3 s 57344 7168 57456 7280 0 FreeSans 448 0 0 0 FrameData_O[16]
port 42 nsew signal output
flabel metal3 s 57344 7616 57456 7728 0 FreeSans 448 0 0 0 FrameData_O[17]
port 43 nsew signal output
flabel metal3 s 57344 8064 57456 8176 0 FreeSans 448 0 0 0 FrameData_O[18]
port 44 nsew signal output
flabel metal3 s 57344 8512 57456 8624 0 FreeSans 448 0 0 0 FrameData_O[19]
port 45 nsew signal output
flabel metal3 s 57344 448 57456 560 0 FreeSans 448 0 0 0 FrameData_O[1]
port 46 nsew signal output
flabel metal3 s 57344 8960 57456 9072 0 FreeSans 448 0 0 0 FrameData_O[20]
port 47 nsew signal output
flabel metal3 s 57344 9408 57456 9520 0 FreeSans 448 0 0 0 FrameData_O[21]
port 48 nsew signal output
flabel metal3 s 57344 9856 57456 9968 0 FreeSans 448 0 0 0 FrameData_O[22]
port 49 nsew signal output
flabel metal3 s 57344 10304 57456 10416 0 FreeSans 448 0 0 0 FrameData_O[23]
port 50 nsew signal output
flabel metal3 s 57344 10752 57456 10864 0 FreeSans 448 0 0 0 FrameData_O[24]
port 51 nsew signal output
flabel metal3 s 57344 11200 57456 11312 0 FreeSans 448 0 0 0 FrameData_O[25]
port 52 nsew signal output
flabel metal3 s 57344 11648 57456 11760 0 FreeSans 448 0 0 0 FrameData_O[26]
port 53 nsew signal output
flabel metal3 s 57344 12096 57456 12208 0 FreeSans 448 0 0 0 FrameData_O[27]
port 54 nsew signal output
flabel metal3 s 57344 12544 57456 12656 0 FreeSans 448 0 0 0 FrameData_O[28]
port 55 nsew signal output
flabel metal3 s 57344 12992 57456 13104 0 FreeSans 448 0 0 0 FrameData_O[29]
port 56 nsew signal output
flabel metal3 s 57344 896 57456 1008 0 FreeSans 448 0 0 0 FrameData_O[2]
port 57 nsew signal output
flabel metal3 s 57344 13440 57456 13552 0 FreeSans 448 0 0 0 FrameData_O[30]
port 58 nsew signal output
flabel metal3 s 57344 13888 57456 14000 0 FreeSans 448 0 0 0 FrameData_O[31]
port 59 nsew signal output
flabel metal3 s 57344 1344 57456 1456 0 FreeSans 448 0 0 0 FrameData_O[3]
port 60 nsew signal output
flabel metal3 s 57344 1792 57456 1904 0 FreeSans 448 0 0 0 FrameData_O[4]
port 61 nsew signal output
flabel metal3 s 57344 2240 57456 2352 0 FreeSans 448 0 0 0 FrameData_O[5]
port 62 nsew signal output
flabel metal3 s 57344 2688 57456 2800 0 FreeSans 448 0 0 0 FrameData_O[6]
port 63 nsew signal output
flabel metal3 s 57344 3136 57456 3248 0 FreeSans 448 0 0 0 FrameData_O[7]
port 64 nsew signal output
flabel metal3 s 57344 3584 57456 3696 0 FreeSans 448 0 0 0 FrameData_O[8]
port 65 nsew signal output
flabel metal3 s 57344 4032 57456 4144 0 FreeSans 448 0 0 0 FrameData_O[9]
port 66 nsew signal output
flabel metal2 s 17472 0 17584 112 0 FreeSans 448 0 0 0 FrameStrobe[0]
port 67 nsew signal input
flabel metal2 s 37632 0 37744 112 0 FreeSans 448 0 0 0 FrameStrobe[10]
port 68 nsew signal input
flabel metal2 s 39648 0 39760 112 0 FreeSans 448 0 0 0 FrameStrobe[11]
port 69 nsew signal input
flabel metal2 s 41664 0 41776 112 0 FreeSans 448 0 0 0 FrameStrobe[12]
port 70 nsew signal input
flabel metal2 s 43680 0 43792 112 0 FreeSans 448 0 0 0 FrameStrobe[13]
port 71 nsew signal input
flabel metal2 s 45696 0 45808 112 0 FreeSans 448 0 0 0 FrameStrobe[14]
port 72 nsew signal input
flabel metal2 s 47712 0 47824 112 0 FreeSans 448 0 0 0 FrameStrobe[15]
port 73 nsew signal input
flabel metal2 s 49728 0 49840 112 0 FreeSans 448 0 0 0 FrameStrobe[16]
port 74 nsew signal input
flabel metal2 s 51744 0 51856 112 0 FreeSans 448 0 0 0 FrameStrobe[17]
port 75 nsew signal input
flabel metal2 s 53760 0 53872 112 0 FreeSans 448 0 0 0 FrameStrobe[18]
port 76 nsew signal input
flabel metal2 s 55776 0 55888 112 0 FreeSans 448 0 0 0 FrameStrobe[19]
port 77 nsew signal input
flabel metal2 s 19488 0 19600 112 0 FreeSans 448 0 0 0 FrameStrobe[1]
port 78 nsew signal input
flabel metal2 s 21504 0 21616 112 0 FreeSans 448 0 0 0 FrameStrobe[2]
port 79 nsew signal input
flabel metal2 s 23520 0 23632 112 0 FreeSans 448 0 0 0 FrameStrobe[3]
port 80 nsew signal input
flabel metal2 s 25536 0 25648 112 0 FreeSans 448 0 0 0 FrameStrobe[4]
port 81 nsew signal input
flabel metal2 s 27552 0 27664 112 0 FreeSans 448 0 0 0 FrameStrobe[5]
port 82 nsew signal input
flabel metal2 s 29568 0 29680 112 0 FreeSans 448 0 0 0 FrameStrobe[6]
port 83 nsew signal input
flabel metal2 s 31584 0 31696 112 0 FreeSans 448 0 0 0 FrameStrobe[7]
port 84 nsew signal input
flabel metal2 s 33600 0 33712 112 0 FreeSans 448 0 0 0 FrameStrobe[8]
port 85 nsew signal input
flabel metal2 s 35616 0 35728 112 0 FreeSans 448 0 0 0 FrameStrobe[9]
port 86 nsew signal input
flabel metal2 s 48160 14112 48272 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[0]
port 87 nsew signal output
flabel metal2 s 52640 14112 52752 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[10]
port 88 nsew signal output
flabel metal2 s 53088 14112 53200 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[11]
port 89 nsew signal output
flabel metal2 s 53536 14112 53648 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[12]
port 90 nsew signal output
flabel metal2 s 53984 14112 54096 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[13]
port 91 nsew signal output
flabel metal2 s 54432 14112 54544 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[14]
port 92 nsew signal output
flabel metal2 s 54880 14112 54992 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[15]
port 93 nsew signal output
flabel metal2 s 55328 14112 55440 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[16]
port 94 nsew signal output
flabel metal2 s 55776 14112 55888 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[17]
port 95 nsew signal output
flabel metal2 s 56224 14112 56336 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[18]
port 96 nsew signal output
flabel metal2 s 56672 14112 56784 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[19]
port 97 nsew signal output
flabel metal2 s 48608 14112 48720 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[1]
port 98 nsew signal output
flabel metal2 s 49056 14112 49168 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[2]
port 99 nsew signal output
flabel metal2 s 49504 14112 49616 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[3]
port 100 nsew signal output
flabel metal2 s 49952 14112 50064 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[4]
port 101 nsew signal output
flabel metal2 s 50400 14112 50512 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[5]
port 102 nsew signal output
flabel metal2 s 50848 14112 50960 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[6]
port 103 nsew signal output
flabel metal2 s 51296 14112 51408 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[7]
port 104 nsew signal output
flabel metal2 s 51744 14112 51856 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[8]
port 105 nsew signal output
flabel metal2 s 52192 14112 52304 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[9]
port 106 nsew signal output
flabel metal2 s 672 14112 784 14224 0 FreeSans 448 0 0 0 N1BEG[0]
port 107 nsew signal output
flabel metal2 s 1120 14112 1232 14224 0 FreeSans 448 0 0 0 N1BEG[1]
port 108 nsew signal output
flabel metal2 s 1568 14112 1680 14224 0 FreeSans 448 0 0 0 N1BEG[2]
port 109 nsew signal output
flabel metal2 s 2016 14112 2128 14224 0 FreeSans 448 0 0 0 N1BEG[3]
port 110 nsew signal output
flabel metal2 s 2464 14112 2576 14224 0 FreeSans 448 0 0 0 N2BEG[0]
port 111 nsew signal output
flabel metal2 s 2912 14112 3024 14224 0 FreeSans 448 0 0 0 N2BEG[1]
port 112 nsew signal output
flabel metal2 s 3360 14112 3472 14224 0 FreeSans 448 0 0 0 N2BEG[2]
port 113 nsew signal output
flabel metal2 s 3808 14112 3920 14224 0 FreeSans 448 0 0 0 N2BEG[3]
port 114 nsew signal output
flabel metal2 s 4256 14112 4368 14224 0 FreeSans 448 0 0 0 N2BEG[4]
port 115 nsew signal output
flabel metal2 s 4704 14112 4816 14224 0 FreeSans 448 0 0 0 N2BEG[5]
port 116 nsew signal output
flabel metal2 s 5152 14112 5264 14224 0 FreeSans 448 0 0 0 N2BEG[6]
port 117 nsew signal output
flabel metal2 s 5600 14112 5712 14224 0 FreeSans 448 0 0 0 N2BEG[7]
port 118 nsew signal output
flabel metal2 s 6048 14112 6160 14224 0 FreeSans 448 0 0 0 N2BEGb[0]
port 119 nsew signal output
flabel metal2 s 6496 14112 6608 14224 0 FreeSans 448 0 0 0 N2BEGb[1]
port 120 nsew signal output
flabel metal2 s 6944 14112 7056 14224 0 FreeSans 448 0 0 0 N2BEGb[2]
port 121 nsew signal output
flabel metal2 s 7392 14112 7504 14224 0 FreeSans 448 0 0 0 N2BEGb[3]
port 122 nsew signal output
flabel metal2 s 7840 14112 7952 14224 0 FreeSans 448 0 0 0 N2BEGb[4]
port 123 nsew signal output
flabel metal2 s 8288 14112 8400 14224 0 FreeSans 448 0 0 0 N2BEGb[5]
port 124 nsew signal output
flabel metal2 s 8736 14112 8848 14224 0 FreeSans 448 0 0 0 N2BEGb[6]
port 125 nsew signal output
flabel metal2 s 9184 14112 9296 14224 0 FreeSans 448 0 0 0 N2BEGb[7]
port 126 nsew signal output
flabel metal2 s 9632 14112 9744 14224 0 FreeSans 448 0 0 0 N4BEG[0]
port 127 nsew signal output
flabel metal2 s 14112 14112 14224 14224 0 FreeSans 448 0 0 0 N4BEG[10]
port 128 nsew signal output
flabel metal2 s 14560 14112 14672 14224 0 FreeSans 448 0 0 0 N4BEG[11]
port 129 nsew signal output
flabel metal2 s 15008 14112 15120 14224 0 FreeSans 448 0 0 0 N4BEG[12]
port 130 nsew signal output
flabel metal2 s 15456 14112 15568 14224 0 FreeSans 448 0 0 0 N4BEG[13]
port 131 nsew signal output
flabel metal2 s 15904 14112 16016 14224 0 FreeSans 448 0 0 0 N4BEG[14]
port 132 nsew signal output
flabel metal2 s 16352 14112 16464 14224 0 FreeSans 448 0 0 0 N4BEG[15]
port 133 nsew signal output
flabel metal2 s 10080 14112 10192 14224 0 FreeSans 448 0 0 0 N4BEG[1]
port 134 nsew signal output
flabel metal2 s 10528 14112 10640 14224 0 FreeSans 448 0 0 0 N4BEG[2]
port 135 nsew signal output
flabel metal2 s 10976 14112 11088 14224 0 FreeSans 448 0 0 0 N4BEG[3]
port 136 nsew signal output
flabel metal2 s 11424 14112 11536 14224 0 FreeSans 448 0 0 0 N4BEG[4]
port 137 nsew signal output
flabel metal2 s 11872 14112 11984 14224 0 FreeSans 448 0 0 0 N4BEG[5]
port 138 nsew signal output
flabel metal2 s 12320 14112 12432 14224 0 FreeSans 448 0 0 0 N4BEG[6]
port 139 nsew signal output
flabel metal2 s 12768 14112 12880 14224 0 FreeSans 448 0 0 0 N4BEG[7]
port 140 nsew signal output
flabel metal2 s 13216 14112 13328 14224 0 FreeSans 448 0 0 0 N4BEG[8]
port 141 nsew signal output
flabel metal2 s 13664 14112 13776 14224 0 FreeSans 448 0 0 0 N4BEG[9]
port 142 nsew signal output
flabel metal2 s 16800 14112 16912 14224 0 FreeSans 448 0 0 0 NN4BEG[0]
port 143 nsew signal output
flabel metal2 s 21280 14112 21392 14224 0 FreeSans 448 0 0 0 NN4BEG[10]
port 144 nsew signal output
flabel metal2 s 21728 14112 21840 14224 0 FreeSans 448 0 0 0 NN4BEG[11]
port 145 nsew signal output
flabel metal2 s 22176 14112 22288 14224 0 FreeSans 448 0 0 0 NN4BEG[12]
port 146 nsew signal output
flabel metal2 s 22624 14112 22736 14224 0 FreeSans 448 0 0 0 NN4BEG[13]
port 147 nsew signal output
flabel metal2 s 23072 14112 23184 14224 0 FreeSans 448 0 0 0 NN4BEG[14]
port 148 nsew signal output
flabel metal2 s 23520 14112 23632 14224 0 FreeSans 448 0 0 0 NN4BEG[15]
port 149 nsew signal output
flabel metal2 s 17248 14112 17360 14224 0 FreeSans 448 0 0 0 NN4BEG[1]
port 150 nsew signal output
flabel metal2 s 17696 14112 17808 14224 0 FreeSans 448 0 0 0 NN4BEG[2]
port 151 nsew signal output
flabel metal2 s 18144 14112 18256 14224 0 FreeSans 448 0 0 0 NN4BEG[3]
port 152 nsew signal output
flabel metal2 s 18592 14112 18704 14224 0 FreeSans 448 0 0 0 NN4BEG[4]
port 153 nsew signal output
flabel metal2 s 19040 14112 19152 14224 0 FreeSans 448 0 0 0 NN4BEG[5]
port 154 nsew signal output
flabel metal2 s 19488 14112 19600 14224 0 FreeSans 448 0 0 0 NN4BEG[6]
port 155 nsew signal output
flabel metal2 s 19936 14112 20048 14224 0 FreeSans 448 0 0 0 NN4BEG[7]
port 156 nsew signal output
flabel metal2 s 20384 14112 20496 14224 0 FreeSans 448 0 0 0 NN4BEG[8]
port 157 nsew signal output
flabel metal2 s 20832 14112 20944 14224 0 FreeSans 448 0 0 0 NN4BEG[9]
port 158 nsew signal output
flabel metal2 s 1344 0 1456 112 0 FreeSans 448 0 0 0 RESET_top
port 159 nsew signal input
flabel metal2 s 24416 14112 24528 14224 0 FreeSans 448 0 0 0 S1END[0]
port 160 nsew signal input
flabel metal2 s 24864 14112 24976 14224 0 FreeSans 448 0 0 0 S1END[1]
port 161 nsew signal input
flabel metal2 s 25312 14112 25424 14224 0 FreeSans 448 0 0 0 S1END[2]
port 162 nsew signal input
flabel metal2 s 25760 14112 25872 14224 0 FreeSans 448 0 0 0 S1END[3]
port 163 nsew signal input
flabel metal2 s 29792 14112 29904 14224 0 FreeSans 448 0 0 0 S2END[0]
port 164 nsew signal input
flabel metal2 s 30240 14112 30352 14224 0 FreeSans 448 0 0 0 S2END[1]
port 165 nsew signal input
flabel metal2 s 30688 14112 30800 14224 0 FreeSans 448 0 0 0 S2END[2]
port 166 nsew signal input
flabel metal2 s 31136 14112 31248 14224 0 FreeSans 448 0 0 0 S2END[3]
port 167 nsew signal input
flabel metal2 s 31584 14112 31696 14224 0 FreeSans 448 0 0 0 S2END[4]
port 168 nsew signal input
flabel metal2 s 32032 14112 32144 14224 0 FreeSans 448 0 0 0 S2END[5]
port 169 nsew signal input
flabel metal2 s 32480 14112 32592 14224 0 FreeSans 448 0 0 0 S2END[6]
port 170 nsew signal input
flabel metal2 s 32928 14112 33040 14224 0 FreeSans 448 0 0 0 S2END[7]
port 171 nsew signal input
flabel metal2 s 26208 14112 26320 14224 0 FreeSans 448 0 0 0 S2MID[0]
port 172 nsew signal input
flabel metal2 s 26656 14112 26768 14224 0 FreeSans 448 0 0 0 S2MID[1]
port 173 nsew signal input
flabel metal2 s 27104 14112 27216 14224 0 FreeSans 448 0 0 0 S2MID[2]
port 174 nsew signal input
flabel metal2 s 27552 14112 27664 14224 0 FreeSans 448 0 0 0 S2MID[3]
port 175 nsew signal input
flabel metal2 s 28000 14112 28112 14224 0 FreeSans 448 0 0 0 S2MID[4]
port 176 nsew signal input
flabel metal2 s 28448 14112 28560 14224 0 FreeSans 448 0 0 0 S2MID[5]
port 177 nsew signal input
flabel metal2 s 28896 14112 29008 14224 0 FreeSans 448 0 0 0 S2MID[6]
port 178 nsew signal input
flabel metal2 s 29344 14112 29456 14224 0 FreeSans 448 0 0 0 S2MID[7]
port 179 nsew signal input
flabel metal2 s 33376 14112 33488 14224 0 FreeSans 448 0 0 0 S4END[0]
port 180 nsew signal input
flabel metal2 s 37856 14112 37968 14224 0 FreeSans 448 0 0 0 S4END[10]
port 181 nsew signal input
flabel metal2 s 38304 14112 38416 14224 0 FreeSans 448 0 0 0 S4END[11]
port 182 nsew signal input
flabel metal2 s 38752 14112 38864 14224 0 FreeSans 448 0 0 0 S4END[12]
port 183 nsew signal input
flabel metal2 s 39200 14112 39312 14224 0 FreeSans 448 0 0 0 S4END[13]
port 184 nsew signal input
flabel metal2 s 39648 14112 39760 14224 0 FreeSans 448 0 0 0 S4END[14]
port 185 nsew signal input
flabel metal2 s 40096 14112 40208 14224 0 FreeSans 448 0 0 0 S4END[15]
port 186 nsew signal input
flabel metal2 s 33824 14112 33936 14224 0 FreeSans 448 0 0 0 S4END[1]
port 187 nsew signal input
flabel metal2 s 34272 14112 34384 14224 0 FreeSans 448 0 0 0 S4END[2]
port 188 nsew signal input
flabel metal2 s 34720 14112 34832 14224 0 FreeSans 448 0 0 0 S4END[3]
port 189 nsew signal input
flabel metal2 s 35168 14112 35280 14224 0 FreeSans 448 0 0 0 S4END[4]
port 190 nsew signal input
flabel metal2 s 35616 14112 35728 14224 0 FreeSans 448 0 0 0 S4END[5]
port 191 nsew signal input
flabel metal2 s 36064 14112 36176 14224 0 FreeSans 448 0 0 0 S4END[6]
port 192 nsew signal input
flabel metal2 s 36512 14112 36624 14224 0 FreeSans 448 0 0 0 S4END[7]
port 193 nsew signal input
flabel metal2 s 36960 14112 37072 14224 0 FreeSans 448 0 0 0 S4END[8]
port 194 nsew signal input
flabel metal2 s 37408 14112 37520 14224 0 FreeSans 448 0 0 0 S4END[9]
port 195 nsew signal input
flabel metal2 s 5376 0 5488 112 0 FreeSans 448 0 0 0 SLOT_top0
port 196 nsew signal output
flabel metal2 s 7392 0 7504 112 0 FreeSans 448 0 0 0 SLOT_top1
port 197 nsew signal output
flabel metal2 s 9408 0 9520 112 0 FreeSans 448 0 0 0 SLOT_top2
port 198 nsew signal output
flabel metal2 s 11424 0 11536 112 0 FreeSans 448 0 0 0 SLOT_top3
port 199 nsew signal output
flabel metal2 s 40544 14112 40656 14224 0 FreeSans 448 0 0 0 SS4END[0]
port 200 nsew signal input
flabel metal2 s 45024 14112 45136 14224 0 FreeSans 448 0 0 0 SS4END[10]
port 201 nsew signal input
flabel metal2 s 45472 14112 45584 14224 0 FreeSans 448 0 0 0 SS4END[11]
port 202 nsew signal input
flabel metal2 s 45920 14112 46032 14224 0 FreeSans 448 0 0 0 SS4END[12]
port 203 nsew signal input
flabel metal2 s 46368 14112 46480 14224 0 FreeSans 448 0 0 0 SS4END[13]
port 204 nsew signal input
flabel metal2 s 46816 14112 46928 14224 0 FreeSans 448 0 0 0 SS4END[14]
port 205 nsew signal input
flabel metal2 s 47264 14112 47376 14224 0 FreeSans 448 0 0 0 SS4END[15]
port 206 nsew signal input
flabel metal2 s 40992 14112 41104 14224 0 FreeSans 448 0 0 0 SS4END[1]
port 207 nsew signal input
flabel metal2 s 41440 14112 41552 14224 0 FreeSans 448 0 0 0 SS4END[2]
port 208 nsew signal input
flabel metal2 s 41888 14112 42000 14224 0 FreeSans 448 0 0 0 SS4END[3]
port 209 nsew signal input
flabel metal2 s 42336 14112 42448 14224 0 FreeSans 448 0 0 0 SS4END[4]
port 210 nsew signal input
flabel metal2 s 42784 14112 42896 14224 0 FreeSans 448 0 0 0 SS4END[5]
port 211 nsew signal input
flabel metal2 s 43232 14112 43344 14224 0 FreeSans 448 0 0 0 SS4END[6]
port 212 nsew signal input
flabel metal2 s 43680 14112 43792 14224 0 FreeSans 448 0 0 0 SS4END[7]
port 213 nsew signal input
flabel metal2 s 44128 14112 44240 14224 0 FreeSans 448 0 0 0 SS4END[8]
port 214 nsew signal input
flabel metal2 s 44576 14112 44688 14224 0 FreeSans 448 0 0 0 SS4END[9]
port 215 nsew signal input
flabel metal2 s 15456 0 15568 112 0 FreeSans 448 0 0 0 UserCLK
port 216 nsew signal input
flabel metal2 s 47712 14112 47824 14224 0 FreeSans 448 0 0 0 UserCLKo
port 217 nsew signal output
flabel metal4 s 3776 0 4096 14224 0 FreeSans 1472 90 0 0 VDD
port 218 nsew power bidirectional
flabel metal4 s 3776 0 4096 56 0 FreeSans 368 0 0 0 VDD
port 218 nsew power bidirectional
flabel metal4 s 3776 14168 4096 14224 0 FreeSans 368 0 0 0 VDD
port 218 nsew power bidirectional
flabel metal4 s 23776 0 24096 14224 0 FreeSans 1472 90 0 0 VDD
port 218 nsew power bidirectional
flabel metal4 s 23776 0 24096 56 0 FreeSans 368 0 0 0 VDD
port 218 nsew power bidirectional
flabel metal4 s 23776 14168 24096 14224 0 FreeSans 368 0 0 0 VDD
port 218 nsew power bidirectional
flabel metal4 s 43776 0 44096 14224 0 FreeSans 1472 90 0 0 VDD
port 218 nsew power bidirectional
flabel metal4 s 43776 0 44096 56 0 FreeSans 368 0 0 0 VDD
port 218 nsew power bidirectional
flabel metal4 s 43776 14168 44096 14224 0 FreeSans 368 0 0 0 VDD
port 218 nsew power bidirectional
flabel metal4 s 4436 0 4756 14224 0 FreeSans 1472 90 0 0 VSS
port 219 nsew ground bidirectional
flabel metal4 s 4436 0 4756 56 0 FreeSans 368 0 0 0 VSS
port 219 nsew ground bidirectional
flabel metal4 s 4436 14168 4756 14224 0 FreeSans 368 0 0 0 VSS
port 219 nsew ground bidirectional
flabel metal4 s 24436 0 24756 14224 0 FreeSans 1472 90 0 0 VSS
port 219 nsew ground bidirectional
flabel metal4 s 24436 0 24756 56 0 FreeSans 368 0 0 0 VSS
port 219 nsew ground bidirectional
flabel metal4 s 24436 14168 24756 14224 0 FreeSans 368 0 0 0 VSS
port 219 nsew ground bidirectional
flabel metal4 s 44436 0 44756 14224 0 FreeSans 1472 90 0 0 VSS
port 219 nsew ground bidirectional
flabel metal4 s 44436 0 44756 56 0 FreeSans 368 0 0 0 VSS
port 219 nsew ground bidirectional
flabel metal4 s 44436 14168 44756 14224 0 FreeSans 368 0 0 0 VSS
port 219 nsew ground bidirectional
rlabel metal1 28728 12544 28728 12544 0 VDD
rlabel metal1 28728 13328 28728 13328 0 VSS
rlabel metal2 13496 126 13496 126 0 BOOT_top
rlabel metal2 3416 518 3416 518 0 CONFIGURED_top
rlabel metal3 2590 56 2590 56 0 FrameData[0]
rlabel metal3 1190 4536 1190 4536 0 FrameData[10]
rlabel metal2 9688 1904 9688 1904 0 FrameData[11]
rlabel metal3 1638 5432 1638 5432 0 FrameData[12]
rlabel metal3 1022 5880 1022 5880 0 FrameData[13]
rlabel metal2 1064 6104 1064 6104 0 FrameData[14]
rlabel metal3 966 6776 966 6776 0 FrameData[15]
rlabel metal3 574 7224 574 7224 0 FrameData[16]
rlabel metal2 1064 7560 1064 7560 0 FrameData[17]
rlabel metal3 1358 8120 1358 8120 0 FrameData[18]
rlabel metal3 1526 8568 1526 8568 0 FrameData[19]
rlabel metal3 2870 504 2870 504 0 FrameData[1]
rlabel metal3 574 9016 574 9016 0 FrameData[20]
rlabel metal2 3864 9128 3864 9128 0 FrameData[21]
rlabel metal2 5096 10248 5096 10248 0 FrameData[22]
rlabel metal3 1470 10360 1470 10360 0 FrameData[23]
rlabel metal3 630 10808 630 10808 0 FrameData[24]
rlabel metal2 1848 5880 1848 5880 0 FrameData[25]
rlabel metal2 2800 6888 2800 6888 0 FrameData[26]
rlabel metal3 182 12152 182 12152 0 FrameData[27]
rlabel metal2 3696 7448 3696 7448 0 FrameData[28]
rlabel metal2 1008 4312 1008 4312 0 FrameData[29]
rlabel metal3 686 952 686 952 0 FrameData[2]
rlabel metal2 1512 12152 1512 12152 0 FrameData[30]
rlabel metal3 1246 13944 1246 13944 0 FrameData[31]
rlabel metal3 1078 1400 1078 1400 0 FrameData[3]
rlabel metal3 4942 1848 4942 1848 0 FrameData[4]
rlabel metal3 1750 2296 1750 2296 0 FrameData[5]
rlabel metal3 2758 2744 2758 2744 0 FrameData[6]
rlabel metal3 742 3192 742 3192 0 FrameData[7]
rlabel metal3 854 3640 854 3640 0 FrameData[8]
rlabel metal3 462 4088 462 4088 0 FrameData[9]
rlabel metal3 57162 56 57162 56 0 FrameData_O[0]
rlabel metal3 55986 4536 55986 4536 0 FrameData_O[10]
rlabel metal3 55188 5096 55188 5096 0 FrameData_O[11]
rlabel metal2 56168 4984 56168 4984 0 FrameData_O[12]
rlabel metal2 54600 5936 54600 5936 0 FrameData_O[13]
rlabel metal2 55160 6384 55160 6384 0 FrameData_O[14]
rlabel metal2 56168 6440 56168 6440 0 FrameData_O[15]
rlabel metal2 54600 7392 54600 7392 0 FrameData_O[16]
rlabel metal3 56770 7672 56770 7672 0 FrameData_O[17]
rlabel metal3 56658 8120 56658 8120 0 FrameData_O[18]
rlabel metal2 54376 8736 54376 8736 0 FrameData_O[19]
rlabel metal3 57218 504 57218 504 0 FrameData_O[1]
rlabel metal3 56770 9016 56770 9016 0 FrameData_O[20]
rlabel metal2 55160 9520 55160 9520 0 FrameData_O[21]
rlabel metal2 54600 10416 54600 10416 0 FrameData_O[22]
rlabel metal2 55160 8232 55160 8232 0 FrameData_O[23]
rlabel metal2 52024 10192 52024 10192 0 FrameData_O[24]
rlabel metal3 54488 8344 54488 8344 0 FrameData_O[25]
rlabel metal2 49224 11480 49224 11480 0 FrameData_O[26]
rlabel metal2 53032 7784 53032 7784 0 FrameData_O[27]
rlabel metal3 53256 10248 53256 10248 0 FrameData_O[28]
rlabel metal3 57218 13048 57218 13048 0 FrameData_O[29]
rlabel metal2 52024 1120 52024 1120 0 FrameData_O[2]
rlabel metal2 53816 11704 53816 11704 0 FrameData_O[30]
rlabel metal3 56882 13944 56882 13944 0 FrameData_O[31]
rlabel metal3 55482 1400 55482 1400 0 FrameData_O[3]
rlabel metal3 55482 1848 55482 1848 0 FrameData_O[4]
rlabel metal2 54936 2184 54936 2184 0 FrameData_O[5]
rlabel metal2 56168 2072 56168 2072 0 FrameData_O[6]
rlabel metal2 54600 3080 54600 3080 0 FrameData_O[7]
rlabel metal3 56154 3640 56154 3640 0 FrameData_O[8]
rlabel metal2 56168 3528 56168 3528 0 FrameData_O[9]
rlabel metal2 17528 126 17528 126 0 FrameStrobe[0]
rlabel metal3 48048 3304 48048 3304 0 FrameStrobe[10]
rlabel metal3 41888 3976 41888 3976 0 FrameStrobe[11]
rlabel metal2 41720 966 41720 966 0 FrameStrobe[12]
rlabel metal2 43736 350 43736 350 0 FrameStrobe[13]
rlabel metal2 45752 798 45752 798 0 FrameStrobe[14]
rlabel metal2 47768 126 47768 126 0 FrameStrobe[15]
rlabel metal2 49784 406 49784 406 0 FrameStrobe[16]
rlabel metal2 51800 1806 51800 1806 0 FrameStrobe[17]
rlabel metal3 29288 5544 29288 5544 0 FrameStrobe[18]
rlabel metal3 29456 6328 29456 6328 0 FrameStrobe[19]
rlabel metal2 29624 5600 29624 5600 0 FrameStrobe[1]
rlabel metal2 21560 630 21560 630 0 FrameStrobe[2]
rlabel metal2 23576 742 23576 742 0 FrameStrobe[3]
rlabel metal2 25592 1302 25592 1302 0 FrameStrobe[4]
rlabel metal3 33544 4536 33544 4536 0 FrameStrobe[5]
rlabel metal3 44296 672 44296 672 0 FrameStrobe[6]
rlabel metal3 32144 6776 32144 6776 0 FrameStrobe[7]
rlabel metal2 37016 4760 37016 4760 0 FrameStrobe[8]
rlabel metal2 35672 1302 35672 1302 0 FrameStrobe[9]
rlabel metal2 48216 13650 48216 13650 0 FrameStrobe_O[0]
rlabel metal2 52696 13538 52696 13538 0 FrameStrobe_O[10]
rlabel metal2 53144 13762 53144 13762 0 FrameStrobe_O[11]
rlabel metal2 53648 9688 53648 9688 0 FrameStrobe_O[12]
rlabel metal3 53536 9240 53536 9240 0 FrameStrobe_O[13]
rlabel metal2 54488 13202 54488 13202 0 FrameStrobe_O[14]
rlabel metal2 54936 13930 54936 13930 0 FrameStrobe_O[15]
rlabel metal2 55384 13538 55384 13538 0 FrameStrobe_O[16]
rlabel metal3 53760 6552 53760 6552 0 FrameStrobe_O[17]
rlabel metal2 56280 13482 56280 13482 0 FrameStrobe_O[18]
rlabel metal2 53032 6160 53032 6160 0 FrameStrobe_O[19]
rlabel metal2 49112 12656 49112 12656 0 FrameStrobe_O[1]
rlabel metal2 51128 13328 51128 13328 0 FrameStrobe_O[2]
rlabel metal3 49952 11592 49952 11592 0 FrameStrobe_O[3]
rlabel metal2 50008 13594 50008 13594 0 FrameStrobe_O[4]
rlabel metal2 50456 13258 50456 13258 0 FrameStrobe_O[5]
rlabel metal2 50904 13426 50904 13426 0 FrameStrobe_O[6]
rlabel metal2 51352 12866 51352 12866 0 FrameStrobe_O[7]
rlabel metal2 51800 13706 51800 13706 0 FrameStrobe_O[8]
rlabel metal2 52248 13650 52248 13650 0 FrameStrobe_O[9]
rlabel metal2 31976 9632 31976 9632 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit13.Q
rlabel metal2 27832 10080 27832 10080 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit14.Q
rlabel metal3 32648 5768 32648 5768 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit15.Q
rlabel metal2 23016 4872 23016 4872 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit16.Q
rlabel metal2 12152 9576 12152 9576 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit17.Q
rlabel metal2 12208 7224 12208 7224 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit18.Q
rlabel metal3 11424 5208 11424 5208 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit19.Q
rlabel metal2 29176 7000 29176 7000 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit20.Q
rlabel metal3 29512 4088 29512 4088 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit21.Q
rlabel metal2 29736 4480 29736 4480 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit22.Q
rlabel metal2 17976 10360 17976 10360 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit23.Q
rlabel metal2 22680 7952 22680 7952 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit24.Q
rlabel metal2 18032 7336 18032 7336 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit25.Q
rlabel metal2 36848 7448 36848 7448 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit26.Q
rlabel metal2 38024 6720 38024 6720 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit27.Q
rlabel metal2 37128 5320 37128 5320 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit28.Q
rlabel metal2 37912 7952 37912 7952 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit29.Q
rlabel metal3 40096 10472 40096 10472 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit30.Q
rlabel metal3 40376 9016 40376 9016 0 Inst_S_WARMBOOT_ConfigMem.Inst_frame0_bit31.Q
rlabel metal2 31640 8316 31640 8316 0 Inst_S_WARMBOOT_switch_matrix.N1BEG0
rlabel metal2 26712 9296 26712 9296 0 Inst_S_WARMBOOT_switch_matrix.N1BEG1
rlabel metal2 31864 6384 31864 6384 0 Inst_S_WARMBOOT_switch_matrix.N1BEG2
rlabel metal3 22120 5096 22120 5096 0 Inst_S_WARMBOOT_switch_matrix.N1BEG3
rlabel metal2 728 12866 728 12866 0 N1BEG[0]
rlabel metal2 2128 9240 2128 9240 0 N1BEG[1]
rlabel metal2 1624 13034 1624 13034 0 N1BEG[2]
rlabel metal2 2072 12418 2072 12418 0 N1BEG[3]
rlabel metal2 2520 12698 2520 12698 0 N2BEG[0]
rlabel metal2 2968 13146 2968 13146 0 N2BEG[1]
rlabel metal2 3416 13258 3416 13258 0 N2BEG[2]
rlabel metal2 3864 13426 3864 13426 0 N2BEG[3]
rlabel metal2 2184 13272 2184 13272 0 N2BEG[4]
rlabel metal2 4760 13818 4760 13818 0 N2BEG[5]
rlabel metal3 4928 11592 4928 11592 0 N2BEG[6]
rlabel metal2 5656 13650 5656 13650 0 N2BEG[7]
rlabel metal2 6104 13034 6104 13034 0 N2BEGb[0]
rlabel metal2 6440 11984 6440 11984 0 N2BEGb[1]
rlabel metal3 6496 11592 6496 11592 0 N2BEGb[2]
rlabel metal3 6720 13160 6720 13160 0 N2BEGb[3]
rlabel metal2 7952 10808 7952 10808 0 N2BEGb[4]
rlabel metal2 8344 12978 8344 12978 0 N2BEGb[5]
rlabel metal3 8288 11592 8288 11592 0 N2BEGb[6]
rlabel metal2 9240 13538 9240 13538 0 N2BEGb[7]
rlabel metal2 7560 13272 7560 13272 0 N4BEG[0]
rlabel metal2 14056 12376 14056 12376 0 N4BEG[10]
rlabel metal2 14616 13202 14616 13202 0 N4BEG[11]
rlabel metal2 13384 13104 13384 13104 0 N4BEG[12]
rlabel metal2 15512 12698 15512 12698 0 N4BEG[13]
rlabel metal2 15960 13258 15960 13258 0 N4BEG[14]
rlabel metal2 16408 13930 16408 13930 0 N4BEG[15]
rlabel metal2 10136 13706 10136 13706 0 N4BEG[1]
rlabel metal2 10584 11914 10584 11914 0 N4BEG[2]
rlabel metal2 11032 13594 11032 13594 0 N4BEG[3]
rlabel metal2 10920 12040 10920 12040 0 N4BEG[4]
rlabel metal3 10864 13160 10864 13160 0 N4BEG[5]
rlabel metal2 12376 12698 12376 12698 0 N4BEG[6]
rlabel metal3 12432 12376 12432 12376 0 N4BEG[7]
rlabel metal2 11368 13216 11368 13216 0 N4BEG[8]
rlabel metal2 13720 13202 13720 13202 0 N4BEG[9]
rlabel metal2 16856 13594 16856 13594 0 NN4BEG[0]
rlabel metal2 21336 13426 21336 13426 0 NN4BEG[10]
rlabel metal2 21672 12824 21672 12824 0 NN4BEG[11]
rlabel metal2 22232 13202 22232 13202 0 NN4BEG[12]
rlabel metal2 22680 13650 22680 13650 0 NN4BEG[13]
rlabel metal2 23576 12656 23576 12656 0 NN4BEG[14]
rlabel metal2 23576 13650 23576 13650 0 NN4BEG[15]
rlabel metal2 17304 13258 17304 13258 0 NN4BEG[1]
rlabel metal2 17528 12096 17528 12096 0 NN4BEG[2]
rlabel metal2 18200 13258 18200 13258 0 NN4BEG[3]
rlabel metal3 18032 13160 18032 13160 0 NN4BEG[4]
rlabel metal2 19096 12866 19096 12866 0 NN4BEG[5]
rlabel metal2 19544 13650 19544 13650 0 NN4BEG[6]
rlabel metal3 19488 13160 19488 13160 0 NN4BEG[7]
rlabel metal2 20440 12810 20440 12810 0 NN4BEG[8]
rlabel metal2 20888 13314 20888 13314 0 NN4BEG[9]
rlabel metal2 1400 518 1400 518 0 RESET_top
rlabel metal2 24696 11032 24696 11032 0 S1END[0]
rlabel metal2 25088 10024 25088 10024 0 S1END[1]
rlabel metal2 25256 11424 25256 11424 0 S1END[2]
rlabel metal2 25816 12866 25816 12866 0 S1END[3]
rlabel metal2 29848 13650 29848 13650 0 S2END[0]
rlabel metal2 30520 12432 30520 12432 0 S2END[1]
rlabel metal2 30744 13650 30744 13650 0 S2END[2]
rlabel metal2 31192 13090 31192 13090 0 S2END[3]
rlabel metal2 31640 13594 31640 13594 0 S2END[4]
rlabel metal2 32088 12866 32088 12866 0 S2END[5]
rlabel metal3 32872 12152 32872 12152 0 S2END[6]
rlabel metal2 32984 13650 32984 13650 0 S2END[7]
rlabel metal2 28728 13384 28728 13384 0 S2MID[0]
rlabel metal2 26712 13650 26712 13650 0 S2MID[1]
rlabel metal2 27160 13650 27160 13650 0 S2MID[2]
rlabel metal2 27608 13650 27608 13650 0 S2MID[3]
rlabel metal2 28056 13818 28056 13818 0 S2MID[4]
rlabel metal2 28504 13146 28504 13146 0 S2MID[5]
rlabel metal2 28952 14042 28952 14042 0 S2MID[6]
rlabel metal2 29400 13146 29400 13146 0 S2MID[7]
rlabel metal3 33768 12152 33768 12152 0 S4END[0]
rlabel metal2 37912 13538 37912 13538 0 S4END[10]
rlabel metal2 38360 13146 38360 13146 0 S4END[11]
rlabel metal2 44520 4760 44520 4760 0 S4END[12]
rlabel metal2 47152 1960 47152 1960 0 S4END[13]
rlabel metal2 50848 2744 50848 2744 0 S4END[14]
rlabel metal3 51548 4200 51548 4200 0 S4END[15]
rlabel metal2 33880 13874 33880 13874 0 S4END[1]
rlabel metal3 34664 12152 34664 12152 0 S4END[2]
rlabel metal2 34776 13650 34776 13650 0 S4END[3]
rlabel metal2 35224 13818 35224 13818 0 S4END[4]
rlabel metal2 35672 13874 35672 13874 0 S4END[5]
rlabel metal2 36120 12866 36120 12866 0 S4END[6]
rlabel metal2 36568 12866 36568 12866 0 S4END[7]
rlabel metal3 7140 2856 7140 2856 0 S4END[8]
rlabel metal2 37464 13986 37464 13986 0 S4END[9]
rlabel metal2 5432 686 5432 686 0 SLOT_top0
rlabel metal2 7448 686 7448 686 0 SLOT_top1
rlabel metal2 9464 126 9464 126 0 SLOT_top2
rlabel metal2 11480 126 11480 126 0 SLOT_top3
rlabel metal2 40600 13650 40600 13650 0 SS4END[0]
rlabel metal2 48440 10528 48440 10528 0 SS4END[10]
rlabel metal2 53256 5936 53256 5936 0 SS4END[11]
rlabel metal2 51688 8568 51688 8568 0 SS4END[12]
rlabel metal2 46312 12152 46312 12152 0 SS4END[13]
rlabel metal2 46816 13160 46816 13160 0 SS4END[14]
rlabel metal2 47320 12362 47320 12362 0 SS4END[15]
rlabel metal2 41048 13650 41048 13650 0 SS4END[1]
rlabel metal2 41496 13874 41496 13874 0 SS4END[2]
rlabel metal2 41944 13650 41944 13650 0 SS4END[3]
rlabel metal2 42392 12866 42392 12866 0 SS4END[4]
rlabel metal3 43512 12152 43512 12152 0 SS4END[5]
rlabel metal2 43288 12866 43288 12866 0 SS4END[6]
rlabel metal2 43736 13426 43736 13426 0 SS4END[7]
rlabel metal2 49896 5600 49896 5600 0 SS4END[8]
rlabel metal2 47712 10472 47712 10472 0 SS4END[9]
rlabel metal3 26936 5040 26936 5040 0 UserCLK
rlabel metal2 47824 8904 47824 8904 0 UserCLKo
rlabel metal3 28056 3304 28056 3304 0 _000_
rlabel metal2 29960 2968 29960 2968 0 _001_
rlabel metal2 29288 3472 29288 3472 0 _002_
rlabel metal2 11032 7728 11032 7728 0 _003_
rlabel metal2 12264 7728 12264 7728 0 _004_
rlabel metal2 12152 6720 12152 6720 0 _005_
rlabel metal3 11480 6664 11480 6664 0 _006_
rlabel metal2 12152 5096 12152 5096 0 _007_
rlabel metal3 12152 4984 12152 4984 0 _008_
rlabel metal2 41608 8008 41608 8008 0 _009_
rlabel metal2 40824 8512 40824 8512 0 _010_
rlabel metal2 42504 9240 42504 9240 0 _011_
rlabel metal2 39480 4816 39480 4816 0 _012_
rlabel metal2 38976 5096 38976 5096 0 _013_
rlabel metal2 18760 6888 18760 6888 0 _014_
rlabel metal2 18872 6720 18872 6720 0 _015_
rlabel metal2 27272 3976 27272 3976 0 _016_
rlabel metal2 26992 3752 26992 3752 0 _017_
rlabel metal2 11256 6552 11256 6552 0 _018_
rlabel metal2 11592 6384 11592 6384 0 _019_
rlabel metal3 40656 8344 40656 8344 0 _020_
rlabel metal2 41944 8372 41944 8372 0 _021_
rlabel metal2 36680 8624 36680 8624 0 _022_
rlabel metal3 40656 8792 40656 8792 0 _023_
rlabel metal3 42112 6664 42112 6664 0 _024_
rlabel metal2 41048 10472 41048 10472 0 _025_
rlabel metal3 41384 10360 41384 10360 0 _026_
rlabel metal2 41160 8680 41160 8680 0 _027_
rlabel metal2 39816 5936 39816 5936 0 _028_
rlabel metal2 39592 6384 39592 6384 0 _029_
rlabel metal2 38472 5712 38472 5712 0 _030_
rlabel metal2 39424 5320 39424 5320 0 _031_
rlabel metal2 37352 6664 37352 6664 0 _032_
rlabel metal2 38136 5824 38136 5824 0 _033_
rlabel metal2 17976 5600 17976 5600 0 _034_
rlabel metal2 18424 9352 18424 9352 0 _035_
rlabel metal2 18928 7448 18928 7448 0 _036_
rlabel metal2 18648 7168 18648 7168 0 _037_
rlabel metal2 19992 8232 19992 8232 0 _038_
rlabel metal2 19656 7504 19656 7504 0 _039_
rlabel metal2 26712 4984 26712 4984 0 _040_
rlabel metal2 28560 4312 28560 4312 0 _041_
rlabel metal2 28952 3808 28952 3808 0 _042_
rlabel metal4 29512 9128 29512 9128 0 net1
rlabel metal2 9688 6552 9688 6552 0 net10
rlabel metal3 52080 2072 52080 2072 0 net100
rlabel metal2 50680 8960 50680 8960 0 net101
rlabel metal2 46984 10024 46984 10024 0 net102
rlabel metal3 51520 7560 51520 7560 0 net103
rlabel metal2 52248 10248 52248 10248 0 net104
rlabel metal2 51352 10808 51352 10808 0 net105
rlabel metal2 47544 10920 47544 10920 0 net106
rlabel metal3 52024 6664 52024 6664 0 net107
rlabel metal3 49000 2688 49000 2688 0 net108
rlabel metal2 28728 8176 28728 8176 0 net109
rlabel metal2 1624 10528 1624 10528 0 net11
rlabel metal2 2576 7560 2576 7560 0 net110
rlabel metal2 29848 5096 29848 5096 0 net111
rlabel metal2 18312 12040 18312 12040 0 net112
rlabel metal2 9912 1848 9912 1848 0 net113
rlabel metal2 11928 9912 11928 9912 0 net114
rlabel metal2 2856 12432 2856 12432 0 net115
rlabel metal2 19544 11032 19544 11032 0 net116
rlabel metal2 2744 11816 2744 11816 0 net117
rlabel metal2 20776 11536 20776 11536 0 net118
rlabel metal2 26264 1512 26264 1512 0 net119
rlabel metal3 23632 2632 23632 2632 0 net12
rlabel metal2 15176 4480 15176 4480 0 net120
rlabel metal2 21784 1232 21784 1232 0 net121
rlabel metal2 21448 13216 21448 13216 0 net122
rlabel metal3 13720 7784 13720 7784 0 net123
rlabel metal2 13496 4536 13496 4536 0 net124
rlabel metal2 31528 11088 31528 11088 0 net125
rlabel metal2 20664 11704 20664 11704 0 net126
rlabel metal2 25480 3220 25480 3220 0 net127
rlabel metal2 11816 5432 11816 5432 0 net128
rlabel metal3 15064 1960 15064 1960 0 net129
rlabel metal3 23016 1960 23016 1960 0 net13
rlabel metal2 23016 6720 23016 6720 0 net130
rlabel metal3 13216 10472 13216 10472 0 net131
rlabel metal2 28616 12488 28616 12488 0 net132
rlabel metal2 19208 3640 19208 3640 0 net133
rlabel metal2 28504 6104 28504 6104 0 net134
rlabel metal2 15848 10304 15848 10304 0 net135
rlabel metal3 23688 3024 23688 3024 0 net136
rlabel metal3 22624 2968 22624 2968 0 net137
rlabel metal2 21672 1736 21672 1736 0 net138
rlabel metal2 17640 6888 17640 6888 0 net139
rlabel metal2 3304 6720 3304 6720 0 net14
rlabel metal4 30072 5069 30072 5069 0 net140
rlabel metal2 23464 2688 23464 2688 0 net141
rlabel metal3 8064 12264 8064 12264 0 net142
rlabel metal3 27384 10248 27384 10248 0 net143
rlabel metal3 16632 3640 16632 3640 0 net144
rlabel metal3 23968 280 23968 280 0 net145
rlabel metal2 25256 8400 25256 8400 0 net146
rlabel metal2 14056 8456 14056 8456 0 net147
rlabel metal2 30240 9464 30240 9464 0 net148
rlabel metal2 18872 9968 18872 9968 0 net149
rlabel metal2 1736 4984 1736 4984 0 net15
rlabel metal2 28952 8456 28952 8456 0 net150
rlabel metal2 23800 13552 23800 13552 0 net151
rlabel metal3 27832 11648 27832 11648 0 net152
rlabel metal2 27160 9576 27160 9576 0 net153
rlabel metal3 26040 224 26040 224 0 net154
rlabel metal2 26936 10472 26936 10472 0 net155
rlabel metal3 23352 2744 23352 2744 0 net156
rlabel metal3 31444 8568 31444 8568 0 net157
rlabel metal2 30016 4536 30016 4536 0 net158
rlabel metal4 28280 9856 28280 9856 0 net159
rlabel metal2 2520 5544 2520 5544 0 net16
rlabel metal2 17416 10192 17416 10192 0 net160
rlabel metal2 6552 1904 6552 1904 0 net161
rlabel metal2 8120 952 8120 952 0 net162
rlabel metal2 18760 7336 18760 7336 0 net163
rlabel metal2 12936 2520 12936 2520 0 net164
rlabel metal3 48608 8792 48608 8792 0 net165
rlabel metal2 24864 11928 24864 11928 0 net166
rlabel metal4 27272 13801 27272 13801 0 net17
rlabel metal3 30016 3416 30016 3416 0 net18
rlabel metal3 24360 2240 24360 2240 0 net19
rlabel metal2 30240 10472 30240 10472 0 net2
rlabel metal2 1624 3976 1624 3976 0 net20
rlabel metal3 23464 2408 23464 2408 0 net21
rlabel metal2 2520 4760 2520 4760 0 net22
rlabel metal2 2184 672 2184 672 0 net23
rlabel metal2 23240 5376 23240 5376 0 net24
rlabel metal4 28280 6179 28280 6179 0 net25
rlabel metal2 25592 9856 25592 9856 0 net26
rlabel metal2 30744 10584 30744 10584 0 net27
rlabel metal2 30632 12432 30632 12432 0 net28
rlabel metal2 28952 2912 28952 2912 0 net29
rlabel metal2 1624 6608 1624 6608 0 net3
rlabel metal2 21112 10136 21112 10136 0 net30
rlabel metal3 36288 8344 36288 8344 0 net31
rlabel metal2 30184 6552 30184 6552 0 net32
rlabel metal3 31360 2744 31360 2744 0 net33
rlabel metal2 27496 11984 27496 11984 0 net34
rlabel metal3 36736 8008 36736 8008 0 net35
rlabel metal2 26936 9296 26936 9296 0 net36
rlabel metal2 25480 11032 25480 11032 0 net37
rlabel metal3 25088 10024 25088 10024 0 net38
rlabel metal2 28392 11928 28392 11928 0 net39
rlabel metal2 2520 7000 2520 7000 0 net4
rlabel metal4 18984 4424 18984 4424 0 net40
rlabel metal2 29064 6160 29064 6160 0 net41
rlabel metal2 30632 5096 30632 5096 0 net42
rlabel metal2 36792 12712 36792 12712 0 net43
rlabel metal3 26040 2016 26040 2016 0 net44
rlabel metal2 27048 6328 27048 6328 0 net45
rlabel metal3 29176 8960 29176 8960 0 net46
rlabel metal2 37800 8904 37800 8904 0 net47
rlabel metal4 28504 13879 28504 13879 0 net48
rlabel metal2 29512 7784 29512 7784 0 net49
rlabel metal2 30072 8260 30072 8260 0 net5
rlabel metal2 26936 12712 26936 12712 0 net50
rlabel metal2 42728 12488 42728 12488 0 net51
rlabel metal2 36568 8736 36568 8736 0 net52
rlabel metal2 28952 7392 28952 7392 0 net53
rlabel metal2 27720 9688 27720 9688 0 net54
rlabel metal2 41944 11704 41944 11704 0 net55
rlabel metal2 21896 2296 21896 2296 0 net56
rlabel metal3 51632 2744 51632 2744 0 net57
rlabel metal2 53592 4424 53592 4424 0 net58
rlabel metal3 53256 4872 53256 4872 0 net59
rlabel metal2 24864 1960 24864 1960 0 net6
rlabel metal3 25928 1008 25928 1008 0 net60
rlabel metal3 53704 9576 53704 9576 0 net61
rlabel metal2 54152 6216 54152 6216 0 net62
rlabel metal2 31528 5320 31528 5320 0 net63
rlabel metal2 22120 1960 22120 1960 0 net64
rlabel metal2 29064 7560 29064 7560 0 net65
rlabel metal3 53648 8904 53648 8904 0 net66
rlabel metal2 29288 6496 29288 6496 0 net67
rlabel metal2 52584 4144 52584 4144 0 net68
rlabel metal2 55160 10696 55160 10696 0 net69
rlabel metal2 1512 5320 1512 5320 0 net7
rlabel metal4 48440 840 48440 840 0 net70
rlabel metal2 24024 2464 24024 2464 0 net71
rlabel metal4 21784 3330 21784 3330 0 net72
rlabel metal3 28504 9688 28504 9688 0 net73
rlabel metal3 29512 7112 29512 7112 0 net74
rlabel metal2 48216 11032 48216 11032 0 net75
rlabel metal2 52136 7336 52136 7336 0 net76
rlabel metal2 51016 7560 51016 7560 0 net77
rlabel metal2 42056 2240 42056 2240 0 net78
rlabel metal3 23688 1624 23688 1624 0 net79
rlabel metal2 1624 7980 1624 7980 0 net8
rlabel metal2 39032 10416 39032 10416 0 net80
rlabel metal3 34664 8792 34664 8792 0 net81
rlabel metal2 52528 1176 52528 1176 0 net82
rlabel metal3 50344 3192 50344 3192 0 net83
rlabel metal4 28728 6390 28728 6390 0 net84
rlabel metal4 30576 5670 30576 5670 0 net85
rlabel metal3 49224 3080 49224 3080 0 net86
rlabel metal2 54152 3696 54152 3696 0 net87
rlabel metal2 55384 4928 55384 4928 0 net88
rlabel metal3 42616 12208 42616 12208 0 net89
rlabel metal2 8680 7784 8680 7784 0 net9
rlabel metal3 52080 3304 52080 3304 0 net90
rlabel metal2 55272 11088 55272 11088 0 net91
rlabel metal2 52584 9128 52584 9128 0 net92
rlabel metal3 51212 9016 51212 9016 0 net93
rlabel metal3 51688 10472 51688 10472 0 net94
rlabel metal2 41608 2968 41608 2968 0 net95
rlabel metal2 48552 11760 48552 11760 0 net96
rlabel metal2 52584 6160 52584 6160 0 net97
rlabel metal2 35336 6552 35336 6552 0 net98
rlabel via3 30184 5315 30184 5315 0 net99
<< properties >>
string FIXED_BBOX 0 0 57456 14224
<< end >>
