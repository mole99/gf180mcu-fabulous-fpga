magic
tech gf180mcuD
magscale 1 10
timestamp 1764324464
<< metal1 >>
rect 672 113706 31024 113740
rect 672 113654 4466 113706
rect 4518 113654 4570 113706
rect 4622 113654 4674 113706
rect 4726 113654 24466 113706
rect 24518 113654 24570 113706
rect 24622 113654 24674 113706
rect 24726 113654 31024 113706
rect 672 113620 31024 113654
rect 4846 113538 4898 113550
rect 1474 113486 1486 113538
rect 1538 113486 1550 113538
rect 5170 113486 5182 113538
rect 5234 113486 5246 113538
rect 14690 113486 14702 113538
rect 14754 113486 14766 113538
rect 15362 113486 15374 113538
rect 15426 113486 15438 113538
rect 18498 113486 18510 113538
rect 18562 113486 18574 113538
rect 19170 113486 19182 113538
rect 19234 113486 19246 113538
rect 22306 113486 22318 113538
rect 22370 113486 22382 113538
rect 22978 113486 22990 113538
rect 23042 113486 23054 113538
rect 24546 113486 24558 113538
rect 24610 113486 24622 113538
rect 25442 113486 25454 113538
rect 25506 113486 25518 113538
rect 26114 113486 26126 113538
rect 26178 113486 26190 113538
rect 26786 113486 26798 113538
rect 26850 113486 26862 113538
rect 27682 113486 27694 113538
rect 27746 113486 27758 113538
rect 28354 113486 28366 113538
rect 28418 113486 28430 113538
rect 29026 113486 29038 113538
rect 29090 113486 29102 113538
rect 29810 113486 29822 113538
rect 29874 113486 29886 113538
rect 4846 113474 4898 113486
rect 5854 113426 5906 113438
rect 12574 113426 12626 113438
rect 2930 113374 2942 113426
rect 2994 113374 3006 113426
rect 5506 113374 5518 113426
rect 5570 113374 5582 113426
rect 6850 113374 6862 113426
rect 6914 113374 6926 113426
rect 9650 113374 9662 113426
rect 9714 113374 9726 113426
rect 11554 113374 11566 113426
rect 11618 113374 11630 113426
rect 13682 113374 13694 113426
rect 13746 113374 13758 113426
rect 17602 113374 17614 113426
rect 17666 113374 17678 113426
rect 21298 113374 21310 113426
rect 21362 113374 21374 113426
rect 23874 113374 23886 113426
rect 23938 113374 23950 113426
rect 5854 113362 5906 113374
rect 12574 113362 12626 113374
rect 15038 113314 15090 113326
rect 18846 113314 18898 113326
rect 1250 113262 1262 113314
rect 1314 113262 1326 113314
rect 6290 113262 6302 113314
rect 6354 113262 6366 113314
rect 11778 113262 11790 113314
rect 11842 113262 11854 113314
rect 15586 113262 15598 113314
rect 15650 113262 15662 113314
rect 15038 113250 15090 113262
rect 18846 113250 18898 113262
rect 19518 113314 19570 113326
rect 24222 113314 24274 113326
rect 25790 113314 25842 113326
rect 22530 113262 22542 113314
rect 22594 113262 22606 113314
rect 23202 113262 23214 113314
rect 23266 113262 23278 113314
rect 24770 113262 24782 113314
rect 24834 113262 24846 113314
rect 26338 113262 26350 113314
rect 26402 113262 26414 113314
rect 27010 113262 27022 113314
rect 27074 113262 27086 113314
rect 27906 113262 27918 113314
rect 27970 113262 27982 113314
rect 28578 113262 28590 113314
rect 28642 113262 28654 113314
rect 29250 113262 29262 113314
rect 29314 113262 29326 113314
rect 30034 113262 30046 113314
rect 30098 113262 30110 113314
rect 19518 113250 19570 113262
rect 24222 113250 24274 113262
rect 25790 113250 25842 113262
rect 11230 113202 11282 113214
rect 25230 113202 25282 113214
rect 2594 113150 2606 113202
rect 2658 113150 2670 113202
rect 9202 113150 9214 113202
rect 9266 113150 9278 113202
rect 14130 113150 14142 113202
rect 14194 113150 14206 113202
rect 17938 113150 17950 113202
rect 18002 113150 18014 113202
rect 21746 113150 21758 113202
rect 21810 113150 21822 113202
rect 11230 113138 11282 113150
rect 25230 113138 25282 113150
rect 4174 113090 4226 113102
rect 4174 113026 4226 113038
rect 7982 113090 8034 113102
rect 7982 113026 8034 113038
rect 10782 113090 10834 113102
rect 10782 113026 10834 113038
rect 16382 113090 16434 113102
rect 16382 113026 16434 113038
rect 20190 113090 20242 113102
rect 20190 113026 20242 113038
rect 672 112922 31024 112956
rect 672 112870 3806 112922
rect 3858 112870 3910 112922
rect 3962 112870 4014 112922
rect 4066 112870 23806 112922
rect 23858 112870 23910 112922
rect 23962 112870 24014 112922
rect 24066 112870 31024 112922
rect 672 112836 31024 112870
rect 16706 112590 16718 112642
rect 16770 112590 16782 112642
rect 18946 112590 18958 112642
rect 19010 112590 19022 112642
rect 15150 112530 15202 112542
rect 2706 112478 2718 112530
rect 2770 112478 2782 112530
rect 8418 112478 8430 112530
rect 8482 112478 8494 112530
rect 10770 112478 10782 112530
rect 10834 112478 10846 112530
rect 14466 112478 14478 112530
rect 14530 112478 14542 112530
rect 23538 112478 23550 112530
rect 23602 112478 23614 112530
rect 24210 112478 24222 112530
rect 24274 112478 24286 112530
rect 25778 112478 25790 112530
rect 25842 112478 25854 112530
rect 15150 112466 15202 112478
rect 11566 112418 11618 112430
rect 27470 112418 27522 112430
rect 1474 112366 1486 112418
rect 1538 112366 1550 112418
rect 6066 112366 6078 112418
rect 6130 112366 6142 112418
rect 10210 112366 10222 112418
rect 10274 112366 10286 112418
rect 12226 112366 12238 112418
rect 12290 112366 12302 112418
rect 16370 112366 16382 112418
rect 16434 112366 16446 112418
rect 18610 112366 18622 112418
rect 18674 112366 18686 112418
rect 19506 112366 19518 112418
rect 19570 112366 19582 112418
rect 20626 112366 20638 112418
rect 20690 112366 20702 112418
rect 21298 112366 21310 112418
rect 21362 112366 21374 112418
rect 21970 112366 21982 112418
rect 22034 112366 22046 112418
rect 23314 112366 23326 112418
rect 23378 112366 23390 112418
rect 23986 112366 23998 112418
rect 24050 112366 24062 112418
rect 24658 112366 24670 112418
rect 24722 112366 24734 112418
rect 25554 112366 25566 112418
rect 25618 112366 25630 112418
rect 26450 112366 26462 112418
rect 26514 112366 26526 112418
rect 27122 112366 27134 112418
rect 27186 112366 27198 112418
rect 28466 112366 28478 112418
rect 28530 112366 28542 112418
rect 29138 112366 29150 112418
rect 29202 112366 29214 112418
rect 29810 112366 29822 112418
rect 29874 112366 29886 112418
rect 11566 112354 11618 112366
rect 27470 112354 27522 112366
rect 1150 112306 1202 112318
rect 1150 112242 1202 112254
rect 1822 112306 1874 112318
rect 4286 112306 4338 112318
rect 2146 112254 2158 112306
rect 2210 112254 2222 112306
rect 3154 112254 3166 112306
rect 3218 112254 3230 112306
rect 1822 112242 1874 112254
rect 4286 112242 4338 112254
rect 5070 112306 5122 112318
rect 5742 112306 5794 112318
rect 5394 112254 5406 112306
rect 5458 112254 5470 112306
rect 5070 112242 5122 112254
rect 5742 112242 5794 112254
rect 6862 112306 6914 112318
rect 9102 112306 9154 112318
rect 11902 112306 11954 112318
rect 7970 112254 7982 112306
rect 8034 112254 8046 112306
rect 11218 112254 11230 112306
rect 11282 112254 11294 112306
rect 6862 112242 6914 112254
rect 9102 112242 9154 112254
rect 11902 112242 11954 112254
rect 12910 112306 12962 112318
rect 17390 112306 17442 112318
rect 14018 112254 14030 112306
rect 14082 112254 14094 112306
rect 12910 112242 12962 112254
rect 17390 112242 17442 112254
rect 19854 112306 19906 112318
rect 19854 112242 19906 112254
rect 20974 112306 21026 112318
rect 20974 112242 21026 112254
rect 21646 112306 21698 112318
rect 21646 112242 21698 112254
rect 22318 112306 22370 112318
rect 22990 112306 23042 112318
rect 22642 112254 22654 112306
rect 22706 112254 22718 112306
rect 22318 112242 22370 112254
rect 22990 112242 23042 112254
rect 25006 112306 25058 112318
rect 25006 112242 25058 112254
rect 25342 112306 25394 112318
rect 25342 112242 25394 112254
rect 26238 112306 26290 112318
rect 26238 112242 26290 112254
rect 26798 112306 26850 112318
rect 26798 112242 26850 112254
rect 28814 112306 28866 112318
rect 28814 112242 28866 112254
rect 29486 112306 29538 112318
rect 29486 112242 29538 112254
rect 30158 112306 30210 112318
rect 30158 112242 30210 112254
rect 672 112138 31024 112172
rect 672 112086 4466 112138
rect 4518 112086 4570 112138
rect 4622 112086 4674 112138
rect 4726 112086 24466 112138
rect 24518 112086 24570 112138
rect 24622 112086 24674 112138
rect 24726 112086 31024 112138
rect 672 112052 31024 112086
rect 21198 111970 21250 111982
rect 8082 111918 8094 111970
rect 8146 111918 8158 111970
rect 9202 111918 9214 111970
rect 9266 111918 9278 111970
rect 10882 111918 10894 111970
rect 10946 111918 10958 111970
rect 21198 111906 21250 111918
rect 21870 111970 21922 111982
rect 22866 111918 22878 111970
rect 22930 111918 22942 111970
rect 24882 111918 24894 111970
rect 24946 111918 24958 111970
rect 26562 111918 26574 111970
rect 26626 111918 26638 111970
rect 27234 111918 27246 111970
rect 27298 111918 27310 111970
rect 27570 111918 27582 111970
rect 27634 111918 27646 111970
rect 28242 111918 28254 111970
rect 28306 111918 28318 111970
rect 28914 111918 28926 111970
rect 28978 111918 28990 111970
rect 29922 111918 29934 111970
rect 29986 111918 29998 111970
rect 21870 111906 21922 111918
rect 5070 111858 5122 111870
rect 29262 111858 29314 111870
rect 1586 111806 1598 111858
rect 1650 111806 1662 111858
rect 3826 111806 3838 111858
rect 3890 111806 3902 111858
rect 6178 111806 6190 111858
rect 6242 111806 6254 111858
rect 12450 111806 12462 111858
rect 12514 111806 12526 111858
rect 14914 111806 14926 111858
rect 14978 111806 14990 111858
rect 17938 111806 17950 111858
rect 18002 111806 18014 111858
rect 20178 111806 20190 111858
rect 20242 111806 20254 111858
rect 21522 111806 21534 111858
rect 21586 111806 21598 111858
rect 22194 111806 22206 111858
rect 22258 111806 22270 111858
rect 23650 111806 23662 111858
rect 23714 111806 23726 111858
rect 25554 111806 25566 111858
rect 25618 111806 25630 111858
rect 30594 111806 30606 111858
rect 30658 111806 30670 111858
rect 5070 111794 5122 111806
rect 29262 111794 29314 111806
rect 7758 111746 7810 111758
rect 10558 111746 10610 111758
rect 22542 111746 22594 111758
rect 5618 111694 5630 111746
rect 5682 111694 5694 111746
rect 8978 111694 8990 111746
rect 9042 111694 9054 111746
rect 12002 111694 12014 111746
rect 12066 111694 12078 111746
rect 14354 111694 14366 111746
rect 14418 111694 14430 111746
rect 20738 111694 20750 111746
rect 20802 111694 20814 111746
rect 7758 111682 7810 111694
rect 10558 111682 10610 111694
rect 22542 111682 22594 111694
rect 23326 111746 23378 111758
rect 23326 111682 23378 111694
rect 24558 111746 24610 111758
rect 24558 111682 24610 111694
rect 25230 111746 25282 111758
rect 25230 111682 25282 111694
rect 26014 111746 26066 111758
rect 26014 111682 26066 111694
rect 26238 111746 26290 111758
rect 29598 111746 29650 111758
rect 27010 111694 27022 111746
rect 27074 111694 27086 111746
rect 27794 111694 27806 111746
rect 27858 111694 27870 111746
rect 28466 111694 28478 111746
rect 28530 111694 28542 111746
rect 26238 111682 26290 111694
rect 29598 111682 29650 111694
rect 30270 111746 30322 111758
rect 30270 111682 30322 111694
rect 9662 111634 9714 111646
rect 1250 111582 1262 111634
rect 1314 111582 1326 111634
rect 3490 111582 3502 111634
rect 3554 111582 3566 111634
rect 9662 111570 9714 111582
rect 9998 111634 10050 111646
rect 9998 111570 10050 111582
rect 11230 111634 11282 111646
rect 11230 111570 11282 111582
rect 11566 111634 11618 111646
rect 18386 111582 18398 111634
rect 18450 111582 18462 111634
rect 11566 111570 11618 111582
rect 2830 111522 2882 111534
rect 2830 111458 2882 111470
rect 7310 111522 7362 111534
rect 7310 111458 7362 111470
rect 13582 111522 13634 111534
rect 13582 111458 13634 111470
rect 16046 111522 16098 111534
rect 16046 111458 16098 111470
rect 16830 111522 16882 111534
rect 16830 111458 16882 111470
rect 19070 111522 19122 111534
rect 19070 111458 19122 111470
rect 672 111354 31024 111388
rect 672 111302 3806 111354
rect 3858 111302 3910 111354
rect 3962 111302 4014 111354
rect 4066 111302 23806 111354
rect 23858 111302 23910 111354
rect 23962 111302 24014 111354
rect 24066 111302 31024 111354
rect 672 111268 31024 111302
rect 9662 111074 9714 111086
rect 9662 111010 9714 111022
rect 11566 111074 11618 111086
rect 19506 111022 19518 111074
rect 19570 111022 19582 111074
rect 11566 111010 11618 111022
rect 7534 110962 7586 110974
rect 9998 110962 10050 110974
rect 1250 110910 1262 110962
rect 1314 110910 1326 110962
rect 5506 110910 5518 110962
rect 5570 110910 5582 110962
rect 6402 110910 6414 110962
rect 6466 110910 6478 110962
rect 6850 110910 6862 110962
rect 6914 110910 6926 110962
rect 8082 110910 8094 110962
rect 8146 110910 8158 110962
rect 9090 110910 9102 110962
rect 9154 110910 9166 110962
rect 7534 110898 7586 110910
rect 9998 110898 10050 110910
rect 10558 110962 10610 110974
rect 10558 110898 10610 110910
rect 10894 110962 10946 110974
rect 15150 110962 15202 110974
rect 17950 110962 18002 110974
rect 21310 110962 21362 110974
rect 12002 110910 12014 110962
rect 12066 110910 12078 110962
rect 13570 110910 13582 110962
rect 13634 110910 13646 110962
rect 15810 110910 15822 110962
rect 15874 110910 15886 110962
rect 20850 110910 20862 110962
rect 20914 110910 20926 110962
rect 10894 110898 10946 110910
rect 15150 110898 15202 110910
rect 17950 110898 18002 110910
rect 21310 110898 21362 110910
rect 21982 110962 22034 110974
rect 23326 110962 23378 110974
rect 22754 110910 22766 110962
rect 22818 110910 22830 110962
rect 21982 110898 22034 110910
rect 23326 110898 23378 110910
rect 23998 110962 24050 110974
rect 23998 110898 24050 110910
rect 24670 110962 24722 110974
rect 24670 110898 24722 110910
rect 26126 110962 26178 110974
rect 26126 110898 26178 110910
rect 30270 110962 30322 110974
rect 30270 110898 30322 110910
rect 6078 110850 6130 110862
rect 1586 110798 1598 110850
rect 1650 110798 1662 110850
rect 3714 110798 3726 110850
rect 3778 110798 3790 110850
rect 4386 110798 4398 110850
rect 4450 110798 4462 110850
rect 10210 110798 10222 110850
rect 10274 110798 10286 110850
rect 19058 110798 19070 110850
rect 19122 110798 19134 110850
rect 20626 110798 20638 110850
rect 20690 110798 20702 110850
rect 22306 110798 22318 110850
rect 22370 110798 22382 110850
rect 22978 110798 22990 110850
rect 23042 110798 23054 110850
rect 23650 110798 23662 110850
rect 23714 110798 23726 110850
rect 24322 110798 24334 110850
rect 24386 110798 24398 110850
rect 24994 110798 25006 110850
rect 25058 110798 25070 110850
rect 25666 110798 25678 110850
rect 25730 110798 25742 110850
rect 26786 110798 26798 110850
rect 26850 110798 26862 110850
rect 27458 110798 27470 110850
rect 27522 110798 27534 110850
rect 29810 110798 29822 110850
rect 29874 110798 29886 110850
rect 6078 110786 6130 110798
rect 2830 110738 2882 110750
rect 2830 110674 2882 110686
rect 3390 110738 3442 110750
rect 3390 110674 3442 110686
rect 4062 110738 4114 110750
rect 17390 110738 17442 110750
rect 25342 110738 25394 110750
rect 5730 110686 5742 110738
rect 5794 110686 5806 110738
rect 7074 110686 7086 110738
rect 7138 110686 7150 110738
rect 11218 110686 11230 110738
rect 11282 110686 11294 110738
rect 12226 110686 12238 110738
rect 12290 110686 12302 110738
rect 14018 110686 14030 110738
rect 14082 110686 14094 110738
rect 16258 110686 16270 110738
rect 16322 110686 16334 110738
rect 21634 110686 21646 110738
rect 21698 110686 21710 110738
rect 4062 110674 4114 110686
rect 17390 110674 17442 110686
rect 25342 110674 25394 110686
rect 26462 110738 26514 110750
rect 26462 110674 26514 110686
rect 27134 110738 27186 110750
rect 27134 110674 27186 110686
rect 29486 110738 29538 110750
rect 30594 110686 30606 110738
rect 30658 110686 30670 110738
rect 29486 110674 29538 110686
rect 672 110570 31024 110604
rect 672 110518 4466 110570
rect 4518 110518 4570 110570
rect 4622 110518 4674 110570
rect 4726 110518 24466 110570
rect 24518 110518 24570 110570
rect 24622 110518 24674 110570
rect 24726 110518 31024 110570
rect 672 110484 31024 110518
rect 19966 110402 20018 110414
rect 1698 110350 1710 110402
rect 1762 110350 1774 110402
rect 9986 110350 9998 110402
rect 10050 110350 10062 110402
rect 13906 110350 13918 110402
rect 13970 110350 13982 110402
rect 18946 110350 18958 110402
rect 19010 110350 19022 110402
rect 19966 110338 20018 110350
rect 20302 110402 20354 110414
rect 20302 110338 20354 110350
rect 21646 110402 21698 110414
rect 27022 110402 27074 110414
rect 21970 110350 21982 110402
rect 22034 110350 22046 110402
rect 22642 110350 22654 110402
rect 22706 110350 22718 110402
rect 23874 110350 23886 110402
rect 23938 110350 23950 110402
rect 24882 110350 24894 110402
rect 24946 110350 24958 110402
rect 25554 110350 25566 110402
rect 25618 110350 25630 110402
rect 27346 110350 27358 110402
rect 27410 110350 27422 110402
rect 21646 110338 21698 110350
rect 27022 110338 27074 110350
rect 25230 110290 25282 110302
rect 27694 110290 27746 110302
rect 2706 110238 2718 110290
rect 2770 110238 2782 110290
rect 4610 110238 4622 110290
rect 4674 110238 4686 110290
rect 4946 110238 4958 110290
rect 5010 110238 5022 110290
rect 6626 110238 6638 110290
rect 6690 110238 6702 110290
rect 9202 110238 9214 110290
rect 9266 110238 9278 110290
rect 11330 110238 11342 110290
rect 11394 110238 11406 110290
rect 17938 110238 17950 110290
rect 18002 110238 18014 110290
rect 19618 110238 19630 110290
rect 19682 110238 19694 110290
rect 20626 110238 20638 110290
rect 20690 110238 20702 110290
rect 20962 110238 20974 110290
rect 21026 110238 21038 110290
rect 26562 110238 26574 110290
rect 26626 110238 26638 110290
rect 30594 110238 30606 110290
rect 30658 110238 30670 110290
rect 25230 110226 25282 110238
rect 27694 110226 27746 110238
rect 1374 110178 1426 110190
rect 1374 110114 1426 110126
rect 8878 110178 8930 110190
rect 8878 110114 8930 110126
rect 10334 110178 10386 110190
rect 14590 110178 14642 110190
rect 19294 110178 19346 110190
rect 22318 110178 22370 110190
rect 10882 110126 10894 110178
rect 10946 110126 10958 110178
rect 13346 110126 13358 110178
rect 13410 110126 13422 110178
rect 13682 110126 13694 110178
rect 13746 110126 13758 110178
rect 15026 110126 15038 110178
rect 15090 110126 15102 110178
rect 15922 110126 15934 110178
rect 15986 110126 15998 110178
rect 21186 110126 21198 110178
rect 21250 110126 21262 110178
rect 10334 110114 10386 110126
rect 14590 110114 14642 110126
rect 19294 110114 19346 110126
rect 22318 110114 22370 110126
rect 23550 110178 23602 110190
rect 30270 110178 30322 110190
rect 24658 110126 24670 110178
rect 24722 110126 24734 110178
rect 26338 110126 26350 110178
rect 26402 110126 26414 110178
rect 23550 110114 23602 110126
rect 30270 110114 30322 110126
rect 5630 110066 5682 110078
rect 9550 110066 9602 110078
rect 2258 110014 2270 110066
rect 2322 110014 2334 110066
rect 6290 110014 6302 110066
rect 6354 110014 6366 110066
rect 5630 110002 5682 110014
rect 9550 110002 9602 110014
rect 12910 110066 12962 110078
rect 25902 110066 25954 110078
rect 18386 110014 18398 110066
rect 18450 110014 18462 110066
rect 12910 110002 12962 110014
rect 25902 110002 25954 110014
rect 26798 110066 26850 110078
rect 26798 110002 26850 110014
rect 3838 109954 3890 109966
rect 3838 109890 3890 109902
rect 5294 109954 5346 109966
rect 5294 109890 5346 109902
rect 7870 109954 7922 109966
rect 7870 109890 7922 109902
rect 12462 109954 12514 109966
rect 12462 109890 12514 109902
rect 16830 109954 16882 109966
rect 16830 109890 16882 109902
rect 672 109786 31024 109820
rect 672 109734 3806 109786
rect 3858 109734 3910 109786
rect 3962 109734 4014 109786
rect 4066 109734 23806 109786
rect 23858 109734 23910 109786
rect 23962 109734 24014 109786
rect 24066 109734 31024 109786
rect 672 109700 31024 109734
rect 6078 109506 6130 109518
rect 1250 109454 1262 109506
rect 1314 109454 1326 109506
rect 13458 109454 13470 109506
rect 13522 109454 13534 109506
rect 6078 109442 6130 109454
rect 11118 109394 11170 109406
rect 17166 109394 17218 109406
rect 19070 109394 19122 109406
rect 29486 109394 29538 109406
rect 4162 109342 4174 109394
rect 4226 109342 4238 109394
rect 6514 109342 6526 109394
rect 6578 109342 6590 109394
rect 6850 109342 6862 109394
rect 6914 109342 6926 109394
rect 7634 109342 7646 109394
rect 7698 109342 7710 109394
rect 8082 109342 8094 109394
rect 8146 109342 8158 109394
rect 9090 109342 9102 109394
rect 9154 109342 9166 109394
rect 9874 109342 9886 109394
rect 9938 109342 9950 109394
rect 15922 109342 15934 109394
rect 15986 109342 15998 109394
rect 16370 109342 16382 109394
rect 16434 109342 16446 109394
rect 17490 109342 17502 109394
rect 17554 109342 17566 109394
rect 18610 109342 18622 109394
rect 18674 109342 18686 109394
rect 19842 109342 19854 109394
rect 19906 109342 19918 109394
rect 22978 109342 22990 109394
rect 23042 109342 23054 109394
rect 11118 109330 11170 109342
rect 17166 109330 17218 109342
rect 19070 109330 19122 109342
rect 29486 109330 29538 109342
rect 3726 109282 3778 109294
rect 5742 109282 5794 109294
rect 12126 109282 12178 109294
rect 15038 109282 15090 109294
rect 1586 109230 1598 109282
rect 1650 109230 1662 109282
rect 3378 109230 3390 109282
rect 3442 109230 3454 109282
rect 4386 109230 4398 109282
rect 4450 109230 4462 109282
rect 5394 109230 5406 109282
rect 5458 109230 5470 109282
rect 7074 109230 7086 109282
rect 7138 109230 7150 109282
rect 11442 109230 11454 109282
rect 11506 109230 11518 109282
rect 11778 109230 11790 109282
rect 11842 109230 11854 109282
rect 13906 109230 13918 109282
rect 13970 109230 13982 109282
rect 3726 109218 3778 109230
rect 5742 109218 5794 109230
rect 12126 109218 12178 109230
rect 15038 109218 15090 109230
rect 15486 109282 15538 109294
rect 26798 109282 26850 109294
rect 19394 109230 19406 109282
rect 19458 109230 19470 109282
rect 23202 109230 23214 109282
rect 23266 109230 23278 109282
rect 29810 109230 29822 109282
rect 29874 109230 29886 109282
rect 15486 109218 15538 109230
rect 26798 109218 26850 109230
rect 2830 109170 2882 109182
rect 10782 109170 10834 109182
rect 23550 109170 23602 109182
rect 9650 109118 9662 109170
rect 9714 109118 9726 109170
rect 16482 109118 16494 109170
rect 16546 109118 16558 109170
rect 20066 109118 20078 109170
rect 20130 109118 20142 109170
rect 2830 109106 2882 109118
rect 10782 109106 10834 109118
rect 23550 109106 23602 109118
rect 25230 109170 25282 109182
rect 25230 109106 25282 109118
rect 26126 109170 26178 109182
rect 26126 109106 26178 109118
rect 27022 109170 27074 109182
rect 27022 109106 27074 109118
rect 672 109002 31024 109036
rect 672 108950 4466 109002
rect 4518 108950 4570 109002
rect 4622 108950 4674 109002
rect 4726 108950 24466 109002
rect 24518 108950 24570 109002
rect 24622 108950 24674 109002
rect 24726 108950 31024 109002
rect 672 108916 31024 108950
rect 10222 108834 10274 108846
rect 3378 108782 3390 108834
rect 3442 108782 3454 108834
rect 9202 108782 9214 108834
rect 9266 108782 9278 108834
rect 9538 108782 9550 108834
rect 9602 108782 9614 108834
rect 10546 108782 10558 108834
rect 10610 108782 10622 108834
rect 14802 108782 14814 108834
rect 14866 108782 14878 108834
rect 10222 108770 10274 108782
rect 6190 108722 6242 108734
rect 23438 108722 23490 108734
rect 30270 108722 30322 108734
rect 5730 108670 5742 108722
rect 5794 108670 5806 108722
rect 11890 108670 11902 108722
rect 11954 108670 11966 108722
rect 16146 108670 16158 108722
rect 16210 108670 16222 108722
rect 17938 108670 17950 108722
rect 18002 108670 18014 108722
rect 29810 108670 29822 108722
rect 29874 108670 29886 108722
rect 30594 108670 30606 108722
rect 30658 108670 30670 108722
rect 6190 108658 6242 108670
rect 23438 108658 23490 108670
rect 30270 108658 30322 108670
rect 2942 108610 2994 108622
rect 8878 108610 8930 108622
rect 1250 108558 1262 108610
rect 1314 108558 1326 108610
rect 2258 108558 2270 108610
rect 2322 108558 2334 108610
rect 3490 108558 3502 108610
rect 3554 108558 3566 108610
rect 3938 108558 3950 108610
rect 4002 108558 4014 108610
rect 5058 108558 5070 108610
rect 5122 108558 5134 108610
rect 5618 108558 5630 108610
rect 5682 108558 5694 108610
rect 6738 108558 6750 108610
rect 6802 108558 6814 108610
rect 7858 108558 7870 108610
rect 7922 108558 7934 108610
rect 2942 108546 2994 108558
rect 8878 108546 8930 108558
rect 9886 108610 9938 108622
rect 15822 108610 15874 108622
rect 11218 108558 11230 108610
rect 11282 108558 11294 108610
rect 11666 108558 11678 108610
rect 11730 108558 11742 108610
rect 12450 108558 12462 108610
rect 12514 108558 12526 108610
rect 12898 108558 12910 108610
rect 12962 108558 12974 108610
rect 13906 108558 13918 108610
rect 13970 108558 13982 108610
rect 15026 108558 15038 108610
rect 15090 108558 15102 108610
rect 18498 108558 18510 108610
rect 18562 108558 18574 108610
rect 29586 108558 29598 108610
rect 29650 108558 29662 108610
rect 9886 108546 9938 108558
rect 15822 108546 15874 108558
rect 4398 108498 4450 108510
rect 4398 108434 4450 108446
rect 4734 108498 4786 108510
rect 4734 108434 4786 108446
rect 8318 108498 8370 108510
rect 8318 108434 8370 108446
rect 10894 108498 10946 108510
rect 10894 108434 10946 108446
rect 15374 108498 15426 108510
rect 15374 108434 15426 108446
rect 25118 108498 25170 108510
rect 25118 108434 25170 108446
rect 26126 108498 26178 108510
rect 26126 108434 26178 108446
rect 16830 108386 16882 108398
rect 16830 108322 16882 108334
rect 672 108218 31024 108252
rect 672 108166 3806 108218
rect 3858 108166 3910 108218
rect 3962 108166 4014 108218
rect 4066 108166 23806 108218
rect 23858 108166 23910 108218
rect 23962 108166 24014 108218
rect 24066 108166 31024 108218
rect 672 108132 31024 108166
rect 25118 107938 25170 107950
rect 6290 107886 6302 107938
rect 6354 107886 6366 107938
rect 25118 107874 25170 107886
rect 2942 107826 2994 107838
rect 1250 107774 1262 107826
rect 1314 107774 1326 107826
rect 2370 107774 2382 107826
rect 2434 107774 2446 107826
rect 3602 107774 3614 107826
rect 3666 107774 3678 107826
rect 4050 107774 4062 107826
rect 4114 107774 4126 107826
rect 5170 107774 5182 107826
rect 5234 107774 5246 107826
rect 9314 107774 9326 107826
rect 9378 107774 9390 107826
rect 9762 107774 9774 107826
rect 9826 107774 9838 107826
rect 10994 107774 11006 107826
rect 11058 107774 11070 107826
rect 12002 107774 12014 107826
rect 12066 107774 12078 107826
rect 13458 107774 13470 107826
rect 13522 107774 13534 107826
rect 14242 107774 14254 107826
rect 14306 107774 14318 107826
rect 15138 107774 15150 107826
rect 15202 107774 15214 107826
rect 15586 107774 15598 107826
rect 15650 107774 15662 107826
rect 16818 107774 16830 107826
rect 16882 107774 16894 107826
rect 17714 107774 17726 107826
rect 17778 107774 17790 107826
rect 30370 107774 30382 107826
rect 30434 107774 30446 107826
rect 2942 107762 2994 107774
rect 4398 107714 4450 107726
rect 7870 107714 7922 107726
rect 8990 107714 9042 107726
rect 3378 107662 3390 107714
rect 3442 107662 3454 107714
rect 5394 107662 5406 107714
rect 5458 107662 5470 107714
rect 8642 107662 8654 107714
rect 8706 107662 8718 107714
rect 4398 107650 4450 107662
rect 7870 107650 7922 107662
rect 8990 107650 9042 107662
rect 10446 107714 10498 107726
rect 14702 107714 14754 107726
rect 16158 107714 16210 107726
rect 13682 107662 13694 107714
rect 13746 107662 13758 107714
rect 14018 107662 14030 107714
rect 14082 107662 14094 107714
rect 15698 107662 15710 107714
rect 15762 107662 15774 107714
rect 10446 107650 10498 107662
rect 14702 107650 14754 107662
rect 16158 107650 16210 107662
rect 8318 107602 8370 107614
rect 6738 107550 6750 107602
rect 6802 107550 6814 107602
rect 9986 107550 9998 107602
rect 10050 107550 10062 107602
rect 30594 107550 30606 107602
rect 30658 107550 30670 107602
rect 8318 107538 8370 107550
rect 672 107434 31024 107468
rect 672 107382 4466 107434
rect 4518 107382 4570 107434
rect 4622 107382 4674 107434
rect 4726 107382 24466 107434
rect 24518 107382 24570 107434
rect 24622 107382 24674 107434
rect 24726 107382 31024 107434
rect 672 107348 31024 107382
rect 25118 107266 25170 107278
rect 1138 107214 1150 107266
rect 1202 107214 1214 107266
rect 7298 107214 7310 107266
rect 7362 107214 7374 107266
rect 10098 107214 10110 107266
rect 10162 107214 10174 107266
rect 12674 107214 12686 107266
rect 12738 107214 12750 107266
rect 14018 107214 14030 107266
rect 14082 107214 14094 107266
rect 25118 107202 25170 107214
rect 4050 107102 4062 107154
rect 4114 107102 4126 107154
rect 5394 107102 5406 107154
rect 5458 107102 5470 107154
rect 17938 107102 17950 107154
rect 18002 107102 18014 107154
rect 30594 107102 30606 107154
rect 30658 107102 30670 107154
rect 1486 107042 1538 107054
rect 3390 107042 3442 107054
rect 5742 107042 5794 107054
rect 16830 107042 16882 107054
rect 1922 106990 1934 107042
rect 1986 106990 1998 107042
rect 2818 106990 2830 107042
rect 2882 106990 2894 107042
rect 4162 106990 4174 107042
rect 4226 106990 4238 107042
rect 4722 106990 4734 107042
rect 4786 106990 4798 107042
rect 9874 106990 9886 107042
rect 9938 106990 9950 107042
rect 13794 106990 13806 107042
rect 13858 106990 13870 107042
rect 1486 106978 1538 106990
rect 3390 106978 3442 106990
rect 5742 106978 5794 106990
rect 16830 106978 16882 106990
rect 30270 107042 30322 107054
rect 30270 106978 30322 106990
rect 5070 106930 5122 106942
rect 8318 106930 8370 106942
rect 7746 106878 7758 106930
rect 7810 106878 7822 106930
rect 5070 106866 5122 106878
rect 8318 106866 8370 106878
rect 8878 106930 8930 106942
rect 8878 106866 8930 106878
rect 9550 106930 9602 106942
rect 9550 106866 9602 106878
rect 10782 106930 10834 106942
rect 14590 106930 14642 106942
rect 13122 106878 13134 106930
rect 13186 106878 13198 106930
rect 18386 106878 18398 106930
rect 18450 106878 18462 106930
rect 10782 106866 10834 106878
rect 14590 106866 14642 106878
rect 6190 106818 6242 106830
rect 6190 106754 6242 106766
rect 11566 106818 11618 106830
rect 11566 106754 11618 106766
rect 672 106650 31024 106684
rect 672 106598 3806 106650
rect 3858 106598 3910 106650
rect 3962 106598 4014 106650
rect 4066 106598 23806 106650
rect 23858 106598 23910 106650
rect 23962 106598 24014 106650
rect 24066 106598 31024 106650
rect 672 106564 31024 106598
rect 15150 106370 15202 106382
rect 5394 106318 5406 106370
rect 5458 106318 5470 106370
rect 15150 106306 15202 106318
rect 2942 106258 2994 106270
rect 1250 106206 1262 106258
rect 1314 106206 1326 106258
rect 2146 106206 2158 106258
rect 2210 106206 2222 106258
rect 3602 106206 3614 106258
rect 3666 106206 3678 106258
rect 4050 106206 4062 106258
rect 4114 106206 4126 106258
rect 7634 106206 7646 106258
rect 7698 106206 7710 106258
rect 13010 106206 13022 106258
rect 13074 106206 13086 106258
rect 16706 106206 16718 106258
rect 16770 106206 16782 106258
rect 2942 106194 2994 106206
rect 4398 106146 4450 106158
rect 9986 106094 9998 106146
rect 10050 106094 10062 106146
rect 13346 106094 13358 106146
rect 13410 106094 13422 106146
rect 29810 106094 29822 106146
rect 29874 106094 29886 106146
rect 4398 106082 4450 106094
rect 6974 106034 7026 106046
rect 9214 106034 9266 106046
rect 3378 105982 3390 106034
rect 3442 105982 3454 106034
rect 5842 105982 5854 106034
rect 5906 105982 5918 106034
rect 8082 105982 8094 106034
rect 8146 105982 8158 106034
rect 6974 105970 7026 105982
rect 9214 105970 9266 105982
rect 9662 106034 9714 106046
rect 10670 106034 10722 106046
rect 10322 105982 10334 106034
rect 10386 105982 10398 106034
rect 9662 105970 9714 105982
rect 10670 105970 10722 105982
rect 11118 106034 11170 106046
rect 11118 105970 11170 105982
rect 14590 106034 14642 106046
rect 29486 106034 29538 106046
rect 16258 105982 16270 106034
rect 16322 105982 16334 106034
rect 14590 105970 14642 105982
rect 29486 105970 29538 105982
rect 672 105866 31024 105900
rect 672 105814 4466 105866
rect 4518 105814 4570 105866
rect 4622 105814 4674 105866
rect 4726 105814 24466 105866
rect 24518 105814 24570 105866
rect 24622 105814 24674 105866
rect 24726 105814 31024 105866
rect 672 105780 31024 105814
rect 16046 105698 16098 105710
rect 9202 105646 9214 105698
rect 9266 105646 9278 105698
rect 11106 105646 11118 105698
rect 11170 105646 11182 105698
rect 22082 105646 22094 105698
rect 22146 105646 22158 105698
rect 16046 105634 16098 105646
rect 19070 105586 19122 105598
rect 30270 105586 30322 105598
rect 1586 105534 1598 105586
rect 1650 105534 1662 105586
rect 2594 105534 2606 105586
rect 2658 105534 2670 105586
rect 4722 105534 4734 105586
rect 4786 105534 4798 105586
rect 6962 105534 6974 105586
rect 7026 105534 7038 105586
rect 13346 105534 13358 105586
rect 13410 105534 13422 105586
rect 14914 105534 14926 105586
rect 14978 105534 14990 105586
rect 19394 105534 19406 105586
rect 19458 105534 19470 105586
rect 30594 105534 30606 105586
rect 30658 105534 30670 105586
rect 19070 105522 19122 105534
rect 30270 105522 30322 105534
rect 1262 105474 1314 105486
rect 8978 105422 8990 105474
rect 9042 105422 9054 105474
rect 11330 105422 11342 105474
rect 11394 105422 11406 105474
rect 14354 105422 14366 105474
rect 14418 105422 14430 105474
rect 21858 105422 21870 105474
rect 21922 105422 21934 105474
rect 1262 105410 1314 105422
rect 9662 105362 9714 105374
rect 2146 105310 2158 105362
rect 2210 105310 2222 105362
rect 4386 105310 4398 105362
rect 4450 105310 4462 105362
rect 6626 105310 6638 105362
rect 6690 105310 6702 105362
rect 13682 105310 13694 105362
rect 13746 105310 13758 105362
rect 9662 105298 9714 105310
rect 3726 105250 3778 105262
rect 3726 105186 3778 105198
rect 5966 105250 6018 105262
rect 5966 105186 6018 105198
rect 8206 105250 8258 105262
rect 8206 105186 8258 105198
rect 12126 105250 12178 105262
rect 12126 105186 12178 105198
rect 672 105082 31024 105116
rect 672 105030 3806 105082
rect 3858 105030 3910 105082
rect 3962 105030 4014 105082
rect 4066 105030 23806 105082
rect 23858 105030 23910 105082
rect 23962 105030 24014 105082
rect 24066 105030 31024 105082
rect 672 104996 31024 105030
rect 11666 104862 11678 104914
rect 11730 104862 11742 104914
rect 6078 104802 6130 104814
rect 1250 104750 1262 104802
rect 1314 104750 1326 104802
rect 6078 104738 6130 104750
rect 12798 104802 12850 104814
rect 16594 104750 16606 104802
rect 16658 104750 16670 104802
rect 12798 104738 12850 104750
rect 7534 104690 7586 104702
rect 14478 104690 14530 104702
rect 3490 104638 3502 104690
rect 3554 104638 3566 104690
rect 4274 104638 4286 104690
rect 4338 104638 4350 104690
rect 5058 104638 5070 104690
rect 5122 104638 5134 104690
rect 6402 104638 6414 104690
rect 6466 104638 6478 104690
rect 6962 104638 6974 104690
rect 7026 104638 7038 104690
rect 8082 104638 8094 104690
rect 8146 104638 8158 104690
rect 9202 104638 9214 104690
rect 9266 104638 9278 104690
rect 11554 104638 11566 104690
rect 11618 104638 11630 104690
rect 13122 104638 13134 104690
rect 13186 104638 13198 104690
rect 13570 104638 13582 104690
rect 13634 104638 13646 104690
rect 15026 104638 15038 104690
rect 15090 104638 15102 104690
rect 15810 104638 15822 104690
rect 15874 104638 15886 104690
rect 7534 104626 7586 104638
rect 14478 104626 14530 104638
rect 12238 104578 12290 104590
rect 1698 104526 1710 104578
rect 1762 104526 1774 104578
rect 3714 104526 3726 104578
rect 3778 104526 3790 104578
rect 4050 104526 4062 104578
rect 4114 104526 4126 104578
rect 5282 104526 5294 104578
rect 5346 104526 5358 104578
rect 7074 104526 7086 104578
rect 7138 104526 7150 104578
rect 12002 104526 12014 104578
rect 12066 104526 12078 104578
rect 16930 104526 16942 104578
rect 16994 104526 17006 104578
rect 12238 104514 12290 104526
rect 2830 104466 2882 104478
rect 2830 104402 2882 104414
rect 9662 104466 9714 104478
rect 9662 104402 9714 104414
rect 11118 104466 11170 104478
rect 11118 104402 11170 104414
rect 11454 104466 11506 104478
rect 18174 104466 18226 104478
rect 13794 104414 13806 104466
rect 13858 104414 13870 104466
rect 11454 104402 11506 104414
rect 18174 104402 18226 104414
rect 30270 104466 30322 104478
rect 30594 104414 30606 104466
rect 30658 104414 30670 104466
rect 30270 104402 30322 104414
rect 672 104298 31024 104332
rect 672 104246 4466 104298
rect 4518 104246 4570 104298
rect 4622 104246 4674 104298
rect 4726 104246 24466 104298
rect 24518 104246 24570 104298
rect 24622 104246 24674 104298
rect 24726 104246 31024 104298
rect 672 104212 31024 104246
rect 12350 104130 12402 104142
rect 20526 104130 20578 104142
rect 14242 104078 14254 104130
rect 14306 104078 14318 104130
rect 20850 104078 20862 104130
rect 20914 104078 20926 104130
rect 12350 104066 12402 104078
rect 20526 104066 20578 104078
rect 12574 104018 12626 104030
rect 1586 103966 1598 104018
rect 1650 103966 1662 104018
rect 2594 103966 2606 104018
rect 2658 103966 2670 104018
rect 4722 103966 4734 104018
rect 4786 103966 4798 104018
rect 7074 103966 7086 104018
rect 7138 103966 7150 104018
rect 11442 103966 11454 104018
rect 11506 103966 11518 104018
rect 12574 103954 12626 103966
rect 12686 104018 12738 104030
rect 12686 103954 12738 103966
rect 15262 104018 15314 104030
rect 18946 103966 18958 104018
rect 19010 103966 19022 104018
rect 15262 103954 15314 103966
rect 15598 103906 15650 103918
rect 18510 103906 18562 103918
rect 1362 103854 1374 103906
rect 1426 103854 1438 103906
rect 15810 103854 15822 103906
rect 15874 103854 15886 103906
rect 16818 103854 16830 103906
rect 16882 103854 16894 103906
rect 17714 103854 17726 103906
rect 17778 103854 17790 103906
rect 19058 103854 19070 103906
rect 19122 103854 19134 103906
rect 19506 103854 19518 103906
rect 19570 103854 19582 103906
rect 15598 103842 15650 103854
rect 18510 103842 18562 103854
rect 19966 103794 20018 103806
rect 2146 103742 2158 103794
rect 2210 103742 2222 103794
rect 4386 103742 4398 103794
rect 4450 103742 4462 103794
rect 6626 103742 6638 103794
rect 6690 103742 6702 103794
rect 11890 103742 11902 103794
rect 11954 103742 11966 103794
rect 14690 103742 14702 103794
rect 14754 103742 14766 103794
rect 19966 103730 20018 103742
rect 3726 103682 3778 103694
rect 3726 103618 3778 103630
rect 5966 103682 6018 103694
rect 5966 103618 6018 103630
rect 8206 103682 8258 103694
rect 8206 103618 8258 103630
rect 10334 103682 10386 103694
rect 10334 103618 10386 103630
rect 13134 103682 13186 103694
rect 13134 103618 13186 103630
rect 15374 103682 15426 103694
rect 15374 103618 15426 103630
rect 672 103514 31024 103548
rect 672 103462 3806 103514
rect 3858 103462 3910 103514
rect 3962 103462 4014 103514
rect 4066 103462 23806 103514
rect 23858 103462 23910 103514
rect 23962 103462 24014 103514
rect 24066 103462 31024 103514
rect 672 103428 31024 103462
rect 11678 103346 11730 103358
rect 11678 103282 11730 103294
rect 12238 103346 12290 103358
rect 12238 103282 12290 103294
rect 12798 103346 12850 103358
rect 12798 103282 12850 103294
rect 18734 103346 18786 103358
rect 18734 103282 18786 103294
rect 6302 103234 6354 103246
rect 12126 103234 12178 103246
rect 1250 103182 1262 103234
rect 1314 103182 1326 103234
rect 10098 103182 10110 103234
rect 10162 103182 10174 103234
rect 6302 103170 6354 103182
rect 12126 103170 12178 103182
rect 12910 103234 12962 103246
rect 12910 103170 12962 103182
rect 3390 103122 3442 103134
rect 7982 103122 8034 103134
rect 19182 103122 19234 103134
rect 5058 103070 5070 103122
rect 5122 103070 5134 103122
rect 6738 103070 6750 103122
rect 6802 103070 6814 103122
rect 7186 103070 7198 103122
rect 7250 103070 7262 103122
rect 8530 103070 8542 103122
rect 8594 103070 8606 103122
rect 9314 103070 9326 103122
rect 9378 103070 9390 103122
rect 13122 103070 13134 103122
rect 13186 103070 13198 103122
rect 13682 103070 13694 103122
rect 13746 103070 13758 103122
rect 17042 103070 17054 103122
rect 17106 103070 17118 103122
rect 3390 103058 3442 103070
rect 7982 103058 8034 103070
rect 19182 103058 19234 103070
rect 1586 102958 1598 103010
rect 1650 102958 1662 103010
rect 3714 102958 3726 103010
rect 3778 102958 3790 103010
rect 4386 102958 4398 103010
rect 4450 102958 4462 103010
rect 5954 102958 5966 103010
rect 6018 102958 6030 103010
rect 7298 102958 7310 103010
rect 7362 102958 7374 103010
rect 17602 102958 17614 103010
rect 17666 102958 17678 103010
rect 2830 102898 2882 102910
rect 2830 102834 2882 102846
rect 4062 102898 4114 102910
rect 5630 102898 5682 102910
rect 15262 102898 15314 102910
rect 5282 102846 5294 102898
rect 5346 102846 5358 102898
rect 10546 102846 10558 102898
rect 10610 102846 10622 102898
rect 14130 102846 14142 102898
rect 14194 102846 14206 102898
rect 4062 102834 4114 102846
rect 5630 102834 5682 102846
rect 15262 102834 15314 102846
rect 16606 102898 16658 102910
rect 30270 102898 30322 102910
rect 19506 102846 19518 102898
rect 19570 102846 19582 102898
rect 30594 102846 30606 102898
rect 30658 102846 30670 102898
rect 16606 102834 16658 102846
rect 30270 102834 30322 102846
rect 672 102730 31024 102764
rect 672 102678 4466 102730
rect 4518 102678 4570 102730
rect 4622 102678 4674 102730
rect 4726 102678 24466 102730
rect 24518 102678 24570 102730
rect 24622 102678 24674 102730
rect 24726 102678 31024 102730
rect 672 102644 31024 102678
rect 7086 102450 7138 102462
rect 8318 102450 8370 102462
rect 1698 102398 1710 102450
rect 1762 102398 1774 102450
rect 6066 102398 6078 102450
rect 6130 102398 6142 102450
rect 7970 102398 7982 102450
rect 8034 102398 8046 102450
rect 7086 102386 7138 102398
rect 8318 102386 8370 102398
rect 9102 102450 9154 102462
rect 12910 102450 12962 102462
rect 30270 102450 30322 102462
rect 10098 102398 10110 102450
rect 10162 102398 10174 102450
rect 11330 102398 11342 102450
rect 11394 102398 11406 102450
rect 13906 102398 13918 102450
rect 13970 102398 13982 102450
rect 17602 102398 17614 102450
rect 17666 102398 17678 102450
rect 30594 102398 30606 102450
rect 30658 102398 30670 102450
rect 9102 102386 9154 102398
rect 12910 102386 12962 102398
rect 30270 102386 30322 102398
rect 5406 102338 5458 102350
rect 14590 102338 14642 102350
rect 17278 102338 17330 102350
rect 1250 102286 1262 102338
rect 1314 102286 1326 102338
rect 3938 102286 3950 102338
rect 4002 102286 4014 102338
rect 4834 102286 4846 102338
rect 4898 102286 4910 102338
rect 6178 102286 6190 102338
rect 6242 102286 6254 102338
rect 6626 102286 6638 102338
rect 6690 102286 6702 102338
rect 10210 102286 10222 102338
rect 10274 102286 10286 102338
rect 13234 102286 13246 102338
rect 13298 102286 13310 102338
rect 13682 102286 13694 102338
rect 13746 102286 13758 102338
rect 15138 102286 15150 102338
rect 15202 102286 15214 102338
rect 16034 102286 16046 102338
rect 16098 102286 16110 102338
rect 5406 102274 5458 102286
rect 14590 102274 14642 102286
rect 17278 102274 17330 102286
rect 10882 102174 10894 102226
rect 10946 102174 10958 102226
rect 2942 102114 2994 102126
rect 2942 102050 2994 102062
rect 9438 102114 9490 102126
rect 9438 102050 9490 102062
rect 12462 102114 12514 102126
rect 12462 102050 12514 102062
rect 672 101946 31024 101980
rect 672 101894 3806 101946
rect 3858 101894 3910 101946
rect 3962 101894 4014 101946
rect 4066 101894 23806 101946
rect 23858 101894 23910 101946
rect 23962 101894 24014 101946
rect 24066 101894 31024 101946
rect 672 101860 31024 101894
rect 13246 101666 13298 101678
rect 13246 101602 13298 101614
rect 2942 101554 2994 101566
rect 14926 101554 14978 101566
rect 1362 101502 1374 101554
rect 1426 101502 1438 101554
rect 2146 101502 2158 101554
rect 2210 101502 2222 101554
rect 3490 101502 3502 101554
rect 3554 101502 3566 101554
rect 4050 101502 4062 101554
rect 4114 101502 4126 101554
rect 5170 101502 5182 101554
rect 5234 101502 5246 101554
rect 5842 101502 5854 101554
rect 5906 101502 5918 101554
rect 8978 101502 8990 101554
rect 9042 101502 9054 101554
rect 9538 101502 9550 101554
rect 9602 101502 9614 101554
rect 10658 101502 10670 101554
rect 10722 101502 10734 101554
rect 11666 101502 11678 101554
rect 11730 101502 11742 101554
rect 13570 101502 13582 101554
rect 13634 101502 13646 101554
rect 14018 101502 14030 101554
rect 14082 101502 14094 101554
rect 15250 101502 15262 101554
rect 15314 101502 15326 101554
rect 16258 101502 16270 101554
rect 16322 101502 16334 101554
rect 2942 101490 2994 101502
rect 14926 101490 14978 101502
rect 4398 101442 4450 101454
rect 8654 101442 8706 101454
rect 10110 101442 10162 101454
rect 3378 101390 3390 101442
rect 3442 101390 3454 101442
rect 5394 101390 5406 101442
rect 5458 101390 5470 101442
rect 9650 101390 9662 101442
rect 9714 101390 9726 101442
rect 4398 101378 4450 101390
rect 8654 101378 8706 101390
rect 10110 101378 10162 101390
rect 7534 101330 7586 101342
rect 6402 101278 6414 101330
rect 6466 101278 6478 101330
rect 14242 101278 14254 101330
rect 14306 101278 14318 101330
rect 7534 101266 7586 101278
rect 672 101162 31024 101196
rect 672 101110 4466 101162
rect 4518 101110 4570 101162
rect 4622 101110 4674 101162
rect 4726 101110 24466 101162
rect 24518 101110 24570 101162
rect 24622 101110 24674 101162
rect 24726 101110 31024 101162
rect 672 101076 31024 101110
rect 2370 100942 2382 100994
rect 2434 100942 2446 100994
rect 6974 100882 7026 100894
rect 5954 100830 5966 100882
rect 6018 100830 6030 100882
rect 7298 100830 7310 100882
rect 7362 100830 7374 100882
rect 10546 100830 10558 100882
rect 10610 100830 10622 100882
rect 14242 100830 14254 100882
rect 14306 100830 14318 100882
rect 17602 100830 17614 100882
rect 17666 100830 17678 100882
rect 29810 100830 29822 100882
rect 29874 100830 29886 100882
rect 30594 100830 30606 100882
rect 30658 100830 30670 100882
rect 6974 100818 7026 100830
rect 5294 100770 5346 100782
rect 7646 100770 7698 100782
rect 11230 100770 11282 100782
rect 15486 100770 15538 100782
rect 2818 100718 2830 100770
rect 2882 100718 2894 100770
rect 3826 100718 3838 100770
rect 3890 100718 3902 100770
rect 4722 100718 4734 100770
rect 4786 100718 4798 100770
rect 6178 100718 6190 100770
rect 6242 100718 6254 100770
rect 6626 100718 6638 100770
rect 6690 100718 6702 100770
rect 9874 100718 9886 100770
rect 9938 100718 9950 100770
rect 10322 100718 10334 100770
rect 10386 100718 10398 100770
rect 11554 100718 11566 100770
rect 11618 100718 11630 100770
rect 12562 100718 12574 100770
rect 12626 100718 12638 100770
rect 13906 100718 13918 100770
rect 13970 100718 13982 100770
rect 5294 100706 5346 100718
rect 7646 100706 7698 100718
rect 11230 100706 11282 100718
rect 15486 100706 15538 100718
rect 17278 100770 17330 100782
rect 17278 100706 17330 100718
rect 29486 100770 29538 100782
rect 29486 100706 29538 100718
rect 30270 100770 30322 100782
rect 30270 100706 30322 100718
rect 9550 100658 9602 100670
rect 9550 100594 9602 100606
rect 1262 100546 1314 100558
rect 1262 100482 1314 100494
rect 672 100378 31024 100412
rect 672 100326 3806 100378
rect 3858 100326 3910 100378
rect 3962 100326 4014 100378
rect 4066 100326 23806 100378
rect 23858 100326 23910 100378
rect 23962 100326 24014 100378
rect 24066 100326 31024 100378
rect 672 100292 31024 100326
rect 12910 100210 12962 100222
rect 12910 100146 12962 100158
rect 8990 100098 9042 100110
rect 5170 100046 5182 100098
rect 5234 100046 5246 100098
rect 14466 100046 14478 100098
rect 14530 100046 14542 100098
rect 8990 100034 9042 100046
rect 2942 99986 2994 99998
rect 10670 99986 10722 99998
rect 1250 99934 1262 99986
rect 1314 99934 1326 99986
rect 2146 99934 2158 99986
rect 2210 99934 2222 99986
rect 3602 99934 3614 99986
rect 3666 99934 3678 99986
rect 4050 99934 4062 99986
rect 4114 99934 4126 99986
rect 9314 99934 9326 99986
rect 9378 99934 9390 99986
rect 9874 99934 9886 99986
rect 9938 99934 9950 99986
rect 11218 99934 11230 99986
rect 11282 99934 11294 99986
rect 12114 99934 12126 99986
rect 12178 99934 12190 99986
rect 17154 99934 17166 99986
rect 17218 99934 17230 99986
rect 2942 99922 2994 99934
rect 10670 99922 10722 99934
rect 4398 99874 4450 99886
rect 5618 99822 5630 99874
rect 5682 99822 5694 99874
rect 9986 99822 9998 99874
rect 10050 99822 10062 99874
rect 17714 99822 17726 99874
rect 17778 99822 17790 99874
rect 22530 99822 22542 99874
rect 22594 99822 22606 99874
rect 4398 99810 4450 99822
rect 6750 99762 6802 99774
rect 18846 99762 18898 99774
rect 3378 99710 3390 99762
rect 3442 99710 3454 99762
rect 14018 99710 14030 99762
rect 14082 99710 14094 99762
rect 6750 99698 6802 99710
rect 18846 99698 18898 99710
rect 22206 99762 22258 99774
rect 22206 99698 22258 99710
rect 30270 99762 30322 99774
rect 30594 99710 30606 99762
rect 30658 99710 30670 99762
rect 30270 99698 30322 99710
rect 672 99594 31024 99628
rect 672 99542 4466 99594
rect 4518 99542 4570 99594
rect 4622 99542 4674 99594
rect 4726 99542 24466 99594
rect 24518 99542 24570 99594
rect 24622 99542 24674 99594
rect 24726 99542 31024 99594
rect 672 99508 31024 99542
rect 18958 99426 19010 99438
rect 14802 99374 14814 99426
rect 14866 99374 14878 99426
rect 18958 99362 19010 99374
rect 30270 99314 30322 99326
rect 1922 99262 1934 99314
rect 1986 99262 1998 99314
rect 4386 99262 4398 99314
rect 4450 99262 4462 99314
rect 6626 99262 6638 99314
rect 6690 99262 6702 99314
rect 10882 99262 10894 99314
rect 10946 99262 10958 99314
rect 17378 99262 17390 99314
rect 17442 99262 17454 99314
rect 19282 99262 19294 99314
rect 19346 99262 19358 99314
rect 30594 99262 30606 99314
rect 30658 99262 30670 99314
rect 30270 99250 30322 99262
rect 3166 99202 3218 99214
rect 8318 99202 8370 99214
rect 3826 99150 3838 99202
rect 3890 99150 3902 99202
rect 10210 99156 10222 99208
rect 10274 99156 10286 99208
rect 10770 99150 10782 99202
rect 10834 99150 10846 99202
rect 11442 99150 11454 99202
rect 11506 99150 11518 99202
rect 11890 99150 11902 99202
rect 11954 99150 11966 99202
rect 12898 99150 12910 99202
rect 12962 99150 12974 99202
rect 16930 99150 16942 99202
rect 16994 99150 17006 99202
rect 3166 99138 3218 99150
rect 8318 99138 8370 99150
rect 7758 99090 7810 99102
rect 1586 99038 1598 99090
rect 1650 99038 1662 99090
rect 6178 99038 6190 99090
rect 6242 99038 6254 99090
rect 7758 99026 7810 99038
rect 9886 99090 9938 99102
rect 14354 99038 14366 99090
rect 14418 99038 14430 99090
rect 9886 99026 9938 99038
rect 5518 98978 5570 98990
rect 5518 98914 5570 98926
rect 8206 98978 8258 98990
rect 8206 98914 8258 98926
rect 15934 98978 15986 98990
rect 15934 98914 15986 98926
rect 18510 98978 18562 98990
rect 18510 98914 18562 98926
rect 672 98810 31024 98844
rect 672 98758 3806 98810
rect 3858 98758 3910 98810
rect 3962 98758 4014 98810
rect 4066 98758 23806 98810
rect 23858 98758 23910 98810
rect 23962 98758 24014 98810
rect 24066 98758 31024 98810
rect 672 98724 31024 98758
rect 11342 98642 11394 98654
rect 11342 98578 11394 98590
rect 18846 98530 18898 98542
rect 1810 98478 1822 98530
rect 1874 98478 1886 98530
rect 5282 98478 5294 98530
rect 5346 98478 5358 98530
rect 9762 98478 9774 98530
rect 9826 98478 9838 98530
rect 18846 98466 18898 98478
rect 19966 98530 20018 98542
rect 19966 98466 20018 98478
rect 16830 98418 16882 98430
rect 19182 98418 19234 98430
rect 7410 98366 7422 98418
rect 7474 98366 7486 98418
rect 13010 98366 13022 98418
rect 13074 98366 13086 98418
rect 15586 98366 15598 98418
rect 15650 98366 15662 98418
rect 16034 98366 16046 98418
rect 16098 98366 16110 98418
rect 17154 98366 17166 98418
rect 17218 98366 17230 98418
rect 18162 98366 18174 98418
rect 18226 98366 18238 98418
rect 18946 98366 18958 98418
rect 19010 98366 19022 98418
rect 19282 98366 19294 98418
rect 19346 98366 19358 98418
rect 16830 98354 16882 98366
rect 19182 98354 19234 98366
rect 4174 98306 4226 98318
rect 4174 98242 4226 98254
rect 4286 98306 4338 98318
rect 15150 98306 15202 98318
rect 18734 98306 18786 98318
rect 5730 98254 5742 98306
rect 5794 98254 5806 98306
rect 7970 98254 7982 98306
rect 8034 98254 8046 98306
rect 10098 98254 10110 98306
rect 10162 98254 10174 98306
rect 13570 98254 13582 98306
rect 13634 98254 13646 98306
rect 16146 98254 16158 98306
rect 16210 98254 16222 98306
rect 4286 98242 4338 98254
rect 15150 98242 15202 98254
rect 18734 98242 18786 98254
rect 3390 98194 3442 98206
rect 2258 98142 2270 98194
rect 2322 98142 2334 98194
rect 3390 98130 3442 98142
rect 4510 98194 4562 98206
rect 4510 98130 4562 98142
rect 6862 98194 6914 98206
rect 6862 98130 6914 98142
rect 9102 98194 9154 98206
rect 9102 98130 9154 98142
rect 14702 98194 14754 98206
rect 14702 98130 14754 98142
rect 19854 98194 19906 98206
rect 19854 98130 19906 98142
rect 672 98026 31024 98060
rect 672 97974 4466 98026
rect 4518 97974 4570 98026
rect 4622 97974 4674 98026
rect 4726 97974 24466 98026
rect 24518 97974 24570 98026
rect 24622 97974 24674 98026
rect 24726 97974 31024 98026
rect 672 97940 31024 97974
rect 8094 97858 8146 97870
rect 16830 97858 16882 97870
rect 1698 97806 1710 97858
rect 1762 97806 1774 97858
rect 11778 97806 11790 97858
rect 11842 97806 11854 97858
rect 14914 97806 14926 97858
rect 14978 97806 14990 97858
rect 8094 97794 8146 97806
rect 16830 97794 16882 97806
rect 19070 97858 19122 97870
rect 21970 97806 21982 97858
rect 22034 97806 22046 97858
rect 19070 97794 19122 97806
rect 4062 97746 4114 97758
rect 30270 97746 30322 97758
rect 5058 97694 5070 97746
rect 5122 97694 5134 97746
rect 10210 97694 10222 97746
rect 10274 97694 10286 97746
rect 18050 97694 18062 97746
rect 18114 97694 18126 97746
rect 29810 97694 29822 97746
rect 29874 97694 29886 97746
rect 30594 97694 30606 97746
rect 30658 97694 30670 97746
rect 4062 97682 4114 97694
rect 30270 97682 30322 97694
rect 7758 97634 7810 97646
rect 1138 97582 1150 97634
rect 1202 97582 1214 97634
rect 4386 97582 4398 97634
rect 4450 97582 4462 97634
rect 4834 97582 4846 97634
rect 4898 97582 4910 97634
rect 5618 97582 5630 97634
rect 5682 97582 5694 97634
rect 6178 97582 6190 97634
rect 6242 97582 6254 97634
rect 7074 97582 7086 97634
rect 7138 97582 7150 97634
rect 7758 97570 7810 97582
rect 7982 97634 8034 97646
rect 19182 97634 19234 97646
rect 29486 97634 29538 97646
rect 8194 97582 8206 97634
rect 8258 97582 8270 97634
rect 10546 97582 10558 97634
rect 10610 97582 10622 97634
rect 11330 97582 11342 97634
rect 11394 97582 11406 97634
rect 18386 97582 18398 97634
rect 18450 97582 18462 97634
rect 21746 97582 21758 97634
rect 21810 97582 21822 97634
rect 7982 97570 8034 97582
rect 19182 97570 19234 97582
rect 29486 97570 29538 97582
rect 8990 97522 9042 97534
rect 14466 97470 14478 97522
rect 14530 97470 14542 97522
rect 8990 97458 9042 97470
rect 2830 97410 2882 97422
rect 2830 97346 2882 97358
rect 12910 97410 12962 97422
rect 12910 97346 12962 97358
rect 16046 97410 16098 97422
rect 16046 97346 16098 97358
rect 19070 97410 19122 97422
rect 19070 97346 19122 97358
rect 19406 97410 19458 97422
rect 19406 97346 19458 97358
rect 672 97242 31024 97276
rect 672 97190 3806 97242
rect 3858 97190 3910 97242
rect 3962 97190 4014 97242
rect 4066 97190 23806 97242
rect 23858 97190 23910 97242
rect 23962 97190 24014 97242
rect 24066 97190 31024 97242
rect 672 97156 31024 97190
rect 18286 97074 18338 97086
rect 18286 97010 18338 97022
rect 18622 97074 18674 97086
rect 18622 97010 18674 97022
rect 14702 96962 14754 96974
rect 5506 96910 5518 96962
rect 5570 96910 5582 96962
rect 7746 96910 7758 96962
rect 7810 96910 7822 96962
rect 9986 96910 9998 96962
rect 10050 96910 10062 96962
rect 14702 96898 14754 96910
rect 11566 96850 11618 96862
rect 13694 96850 13746 96862
rect 16158 96850 16210 96862
rect 19518 96850 19570 96862
rect 2706 96798 2718 96850
rect 2770 96798 2782 96850
rect 13010 96798 13022 96850
rect 13074 96798 13086 96850
rect 15026 96798 15038 96850
rect 15090 96798 15102 96850
rect 15474 96798 15486 96850
rect 15538 96798 15550 96850
rect 16930 96798 16942 96850
rect 16994 96798 17006 96850
rect 17714 96798 17726 96850
rect 17778 96798 17790 96850
rect 18610 96798 18622 96850
rect 18674 96798 18686 96850
rect 22306 96798 22318 96850
rect 22370 96798 22382 96850
rect 11566 96786 11618 96798
rect 13694 96786 13746 96798
rect 16158 96786 16210 96798
rect 19518 96786 19570 96798
rect 8194 96686 8206 96738
rect 8258 96686 8270 96738
rect 12898 96686 12910 96738
rect 12962 96686 12974 96738
rect 4286 96626 4338 96638
rect 7086 96626 7138 96638
rect 3154 96574 3166 96626
rect 3218 96574 3230 96626
rect 5954 96574 5966 96626
rect 6018 96574 6030 96626
rect 4286 96562 4338 96574
rect 7086 96562 7138 96574
rect 9326 96626 9378 96638
rect 14030 96626 14082 96638
rect 20750 96626 20802 96638
rect 30270 96626 30322 96638
rect 10434 96574 10446 96626
rect 10498 96574 10510 96626
rect 15698 96574 15710 96626
rect 15762 96574 15774 96626
rect 19842 96574 19854 96626
rect 19906 96574 19918 96626
rect 21858 96574 21870 96626
rect 21922 96574 21934 96626
rect 30594 96574 30606 96626
rect 30658 96574 30670 96626
rect 9326 96562 9378 96574
rect 14030 96562 14082 96574
rect 20750 96562 20802 96574
rect 30270 96562 30322 96574
rect 672 96458 31024 96492
rect 672 96406 4466 96458
rect 4518 96406 4570 96458
rect 4622 96406 4674 96458
rect 4726 96406 24466 96458
rect 24518 96406 24570 96458
rect 24622 96406 24674 96458
rect 24726 96406 31024 96458
rect 672 96372 31024 96406
rect 8094 96290 8146 96302
rect 16830 96290 16882 96302
rect 29486 96290 29538 96302
rect 11442 96238 11454 96290
rect 11506 96238 11518 96290
rect 19954 96238 19966 96290
rect 20018 96238 20030 96290
rect 22194 96238 22206 96290
rect 22258 96238 22270 96290
rect 29810 96238 29822 96290
rect 29874 96238 29886 96290
rect 8094 96226 8146 96238
rect 16830 96226 16882 96238
rect 29486 96226 29538 96238
rect 7310 96178 7362 96190
rect 1698 96126 1710 96178
rect 1762 96126 1774 96178
rect 4722 96126 4734 96178
rect 4786 96126 4798 96178
rect 7310 96114 7362 96126
rect 17054 96178 17106 96190
rect 17054 96114 17106 96126
rect 17166 96178 17218 96190
rect 18946 96126 18958 96178
rect 19010 96126 19022 96178
rect 17166 96114 17218 96126
rect 5406 96066 5458 96078
rect 7646 96066 7698 96078
rect 4162 96014 4174 96066
rect 4226 96014 4238 96066
rect 4610 96014 4622 96066
rect 4674 96014 4686 96066
rect 5730 96014 5742 96066
rect 5794 96014 5806 96066
rect 6738 96014 6750 96066
rect 6802 96014 6814 96066
rect 5406 96002 5458 96014
rect 7646 96002 7698 96014
rect 7758 96066 7810 96078
rect 12126 96066 12178 96078
rect 18622 96066 18674 96078
rect 7858 96014 7870 96066
rect 7922 96014 7934 96066
rect 10882 96014 10894 96066
rect 10946 96014 10958 96066
rect 11218 96014 11230 96066
rect 11282 96014 11294 96066
rect 12450 96014 12462 96066
rect 12514 96014 12526 96066
rect 13458 96014 13470 96066
rect 13522 96014 13534 96066
rect 7758 96002 7810 96014
rect 12126 96002 12178 96014
rect 18622 96002 18674 96014
rect 3726 95954 3778 95966
rect 1362 95902 1374 95954
rect 1426 95902 1438 95954
rect 3726 95890 3778 95902
rect 10446 95954 10498 95966
rect 19506 95902 19518 95954
rect 19570 95902 19582 95954
rect 21746 95902 21758 95954
rect 21810 95902 21822 95954
rect 10446 95890 10498 95902
rect 2942 95842 2994 95854
rect 2942 95778 2994 95790
rect 21086 95842 21138 95854
rect 21086 95778 21138 95790
rect 23326 95842 23378 95854
rect 23326 95778 23378 95790
rect 672 95674 31024 95708
rect 672 95622 3806 95674
rect 3858 95622 3910 95674
rect 3962 95622 4014 95674
rect 4066 95622 23806 95674
rect 23858 95622 23910 95674
rect 23962 95622 24014 95674
rect 24066 95622 31024 95674
rect 672 95588 31024 95622
rect 12910 95506 12962 95518
rect 12910 95442 12962 95454
rect 7074 95342 7086 95394
rect 7138 95342 7150 95394
rect 14466 95342 14478 95394
rect 14530 95342 14542 95394
rect 2494 95282 2546 95294
rect 9550 95282 9602 95294
rect 1474 95230 1486 95282
rect 1538 95230 1550 95282
rect 1922 95230 1934 95282
rect 1986 95230 1998 95282
rect 3042 95230 3054 95282
rect 3106 95230 3118 95282
rect 4162 95230 4174 95282
rect 4226 95230 4238 95282
rect 8530 95230 8542 95282
rect 8594 95230 8606 95282
rect 8866 95230 8878 95282
rect 8930 95230 8942 95282
rect 10322 95230 10334 95282
rect 10386 95230 10398 95282
rect 11106 95230 11118 95282
rect 11170 95230 11182 95282
rect 18386 95230 18398 95282
rect 18450 95230 18462 95282
rect 21074 95230 21086 95282
rect 21138 95230 21150 95282
rect 21410 95230 21422 95282
rect 21474 95230 21486 95282
rect 22194 95230 22206 95282
rect 22258 95230 22270 95282
rect 22866 95230 22878 95282
rect 22930 95230 22942 95282
rect 23762 95230 23774 95282
rect 23826 95230 23838 95282
rect 2494 95218 2546 95230
rect 9550 95218 9602 95230
rect 1038 95170 1090 95182
rect 8094 95170 8146 95182
rect 20638 95170 20690 95182
rect 6626 95118 6638 95170
rect 6690 95118 6702 95170
rect 14130 95118 14142 95170
rect 14194 95118 14206 95170
rect 1038 95106 1090 95118
rect 8094 95106 8146 95118
rect 20638 95106 20690 95118
rect 5518 95058 5570 95070
rect 19966 95058 20018 95070
rect 30270 95058 30322 95070
rect 2034 95006 2046 95058
rect 2098 95006 2110 95058
rect 9090 95006 9102 95058
rect 9154 95006 9166 95058
rect 18834 95006 18846 95058
rect 18898 95006 18910 95058
rect 21634 95006 21646 95058
rect 21698 95006 21710 95058
rect 30594 95006 30606 95058
rect 30658 95006 30670 95058
rect 5518 94994 5570 95006
rect 19966 94994 20018 95006
rect 30270 94994 30322 95006
rect 672 94890 31024 94924
rect 672 94838 4466 94890
rect 4518 94838 4570 94890
rect 4622 94838 4674 94890
rect 4726 94838 24466 94890
rect 24518 94838 24570 94890
rect 24622 94838 24674 94890
rect 24726 94838 31024 94890
rect 672 94804 31024 94838
rect 16830 94722 16882 94734
rect 6626 94670 6638 94722
rect 6690 94670 6702 94722
rect 12002 94670 12014 94722
rect 12066 94670 12078 94722
rect 18162 94670 18174 94722
rect 18226 94670 18238 94722
rect 23650 94670 23662 94722
rect 23714 94670 23726 94722
rect 16830 94658 16882 94670
rect 1822 94610 1874 94622
rect 23326 94610 23378 94622
rect 2818 94558 2830 94610
rect 2882 94558 2894 94610
rect 9202 94558 9214 94610
rect 9266 94558 9278 94610
rect 9650 94558 9662 94610
rect 9714 94558 9726 94610
rect 14802 94558 14814 94610
rect 14866 94558 14878 94610
rect 17154 94558 17166 94610
rect 17218 94558 17230 94610
rect 20738 94558 20750 94610
rect 20802 94558 20814 94610
rect 30594 94558 30606 94610
rect 30658 94558 30670 94610
rect 1822 94546 1874 94558
rect 23326 94546 23378 94558
rect 12686 94498 12738 94510
rect 2258 94446 2270 94498
rect 2322 94446 2334 94498
rect 2706 94446 2718 94498
rect 2770 94446 2782 94498
rect 3378 94446 3390 94498
rect 3442 94446 3454 94498
rect 4050 94446 4062 94498
rect 4114 94446 4126 94498
rect 4834 94446 4846 94498
rect 4898 94446 4910 94498
rect 7074 94446 7086 94498
rect 7138 94446 7150 94498
rect 11442 94446 11454 94498
rect 11506 94446 11518 94498
rect 11890 94446 11902 94498
rect 11954 94446 11966 94498
rect 13010 94446 13022 94498
rect 13074 94446 13086 94498
rect 13234 94446 13246 94498
rect 13298 94446 13310 94498
rect 14130 94446 14142 94498
rect 14194 94446 14206 94498
rect 14690 94446 14702 94498
rect 14754 94446 14766 94498
rect 20178 94446 20190 94498
rect 20242 94446 20254 94498
rect 20514 94446 20526 94498
rect 20578 94446 20590 94498
rect 21298 94446 21310 94498
rect 21362 94446 21374 94498
rect 21858 94446 21870 94498
rect 21922 94446 21934 94498
rect 22754 94446 22766 94498
rect 22818 94446 22830 94498
rect 30370 94446 30382 94498
rect 30434 94446 30446 94498
rect 12686 94434 12738 94446
rect 11006 94386 11058 94398
rect 11006 94322 11058 94334
rect 15822 94386 15874 94398
rect 19742 94386 19794 94398
rect 17714 94334 17726 94386
rect 17778 94334 17790 94386
rect 15822 94322 15874 94334
rect 19742 94322 19794 94334
rect 5518 94274 5570 94286
rect 5518 94210 5570 94222
rect 9886 94274 9938 94286
rect 9886 94210 9938 94222
rect 10222 94274 10274 94286
rect 10222 94210 10274 94222
rect 15486 94274 15538 94286
rect 15486 94210 15538 94222
rect 19294 94274 19346 94286
rect 19294 94210 19346 94222
rect 672 94106 31024 94140
rect 672 94054 3806 94106
rect 3858 94054 3910 94106
rect 3962 94054 4014 94106
rect 4066 94054 23806 94106
rect 23858 94054 23910 94106
rect 23962 94054 24014 94106
rect 24066 94054 31024 94106
rect 672 94020 31024 94054
rect 4398 93826 4450 93838
rect 4398 93762 4450 93774
rect 8542 93826 8594 93838
rect 22754 93774 22766 93826
rect 22818 93774 22830 93826
rect 8542 93762 8594 93774
rect 2942 93714 2994 93726
rect 10222 93714 10274 93726
rect 15150 93714 15202 93726
rect 17054 93714 17106 93726
rect 1250 93662 1262 93714
rect 1314 93662 1326 93714
rect 2146 93662 2158 93714
rect 2210 93662 2222 93714
rect 3490 93662 3502 93714
rect 3554 93662 3566 93714
rect 3938 93662 3950 93714
rect 4002 93662 4014 93714
rect 5730 93662 5742 93714
rect 5794 93662 5806 93714
rect 8978 93662 8990 93714
rect 9042 93662 9054 93714
rect 9314 93662 9326 93714
rect 9378 93662 9390 93714
rect 10770 93662 10782 93714
rect 10834 93662 10846 93714
rect 11554 93662 11566 93714
rect 11618 93662 11630 93714
rect 13570 93662 13582 93714
rect 13634 93662 13646 93714
rect 16034 93662 16046 93714
rect 16098 93662 16110 93714
rect 16370 93662 16382 93714
rect 16434 93662 16446 93714
rect 17826 93662 17838 93714
rect 17890 93662 17902 93714
rect 18610 93662 18622 93714
rect 18674 93662 18686 93714
rect 26898 93662 26910 93714
rect 26962 93662 26974 93714
rect 2942 93650 2994 93662
rect 10222 93650 10274 93662
rect 15150 93650 15202 93662
rect 17054 93650 17106 93662
rect 15598 93602 15650 93614
rect 6066 93550 6078 93602
rect 6130 93550 6142 93602
rect 9538 93550 9550 93602
rect 9602 93550 9614 93602
rect 15598 93538 15650 93550
rect 7310 93490 7362 93502
rect 19182 93490 19234 93502
rect 3378 93438 3390 93490
rect 3442 93438 3454 93490
rect 14018 93438 14030 93490
rect 14082 93438 14094 93490
rect 16594 93438 16606 93490
rect 16658 93438 16670 93490
rect 19506 93438 19518 93490
rect 19570 93438 19582 93490
rect 7310 93426 7362 93438
rect 19182 93426 19234 93438
rect 672 93322 31024 93356
rect 672 93270 4466 93322
rect 4518 93270 4570 93322
rect 4622 93270 4674 93322
rect 4726 93270 24466 93322
rect 24518 93270 24570 93322
rect 24622 93270 24674 93322
rect 24726 93270 31024 93322
rect 672 93236 31024 93270
rect 8206 93154 8258 93166
rect 13806 93154 13858 93166
rect 30270 93154 30322 93166
rect 7074 93102 7086 93154
rect 7138 93102 7150 93154
rect 9874 93102 9886 93154
rect 9938 93102 9950 93154
rect 17602 93102 17614 93154
rect 17666 93102 17678 93154
rect 8206 93090 8258 93102
rect 13806 93090 13858 93102
rect 30270 93090 30322 93102
rect 1038 93042 1090 93054
rect 2494 93042 2546 93054
rect 8878 93042 8930 93054
rect 19742 93042 19794 93054
rect 21198 93042 21250 93054
rect 2034 92990 2046 93042
rect 2098 92990 2110 93042
rect 4946 92990 4958 93042
rect 5010 92990 5022 93042
rect 5282 92990 5294 93042
rect 5346 92990 5358 93042
rect 12898 92990 12910 93042
rect 12962 92990 12974 93042
rect 14802 92990 14814 93042
rect 14866 92990 14878 93042
rect 17490 92990 17502 93042
rect 17554 92990 17566 93042
rect 20738 92990 20750 93042
rect 20802 92990 20814 93042
rect 24658 92990 24670 93042
rect 24722 92990 24734 93042
rect 30594 92990 30606 93042
rect 30658 92990 30670 93042
rect 1038 92978 1090 92990
rect 2494 92978 2546 92990
rect 8878 92978 8930 92990
rect 19742 92978 19794 92990
rect 21198 92978 21250 92990
rect 5630 92930 5682 92942
rect 1474 92878 1486 92930
rect 1538 92878 1550 92930
rect 1922 92878 1934 92930
rect 1986 92878 1998 92930
rect 3042 92878 3054 92930
rect 3106 92878 3118 92930
rect 4162 92878 4174 92930
rect 4226 92878 4238 92930
rect 6626 92878 6638 92930
rect 6690 92878 6702 92930
rect 9314 92878 9326 92930
rect 9378 92878 9390 92930
rect 9650 92878 9662 92930
rect 9714 92878 9726 92930
rect 10434 92878 10446 92930
rect 10498 92878 10510 92930
rect 10882 92878 10894 92930
rect 10946 92878 10958 92930
rect 11890 92878 11902 92930
rect 11954 92878 11966 92930
rect 12674 92878 12686 92930
rect 12738 92878 12750 92930
rect 14466 92878 14478 92930
rect 14530 92878 14542 92930
rect 17042 92878 17054 92930
rect 17106 92878 17118 92930
rect 20178 92878 20190 92930
rect 20242 92878 20254 92930
rect 20514 92878 20526 92930
rect 20578 92878 20590 92930
rect 21858 92878 21870 92930
rect 21922 92878 21934 92930
rect 22754 92878 22766 92930
rect 22818 92878 22830 92930
rect 24882 92878 24894 92930
rect 24946 92878 24958 92930
rect 5630 92866 5682 92878
rect 5966 92818 6018 92830
rect 5966 92754 6018 92766
rect 13470 92706 13522 92718
rect 13470 92642 13522 92654
rect 16046 92706 16098 92718
rect 16046 92642 16098 92654
rect 18734 92706 18786 92718
rect 18734 92642 18786 92654
rect 25454 92706 25506 92718
rect 25454 92642 25506 92654
rect 25790 92706 25842 92718
rect 25790 92642 25842 92654
rect 672 92538 31024 92572
rect 672 92486 3806 92538
rect 3858 92486 3910 92538
rect 3962 92486 4014 92538
rect 4066 92486 23806 92538
rect 23858 92486 23910 92538
rect 23962 92486 24014 92538
rect 24066 92486 31024 92538
rect 672 92452 31024 92486
rect 5070 92370 5122 92382
rect 5070 92306 5122 92318
rect 8206 92258 8258 92270
rect 5394 92206 5406 92258
rect 5458 92206 5470 92258
rect 8206 92194 8258 92206
rect 15598 92258 15650 92270
rect 15598 92194 15650 92206
rect 9662 92146 9714 92158
rect 17054 92146 17106 92158
rect 22094 92146 22146 92158
rect 2706 92094 2718 92146
rect 2770 92094 2782 92146
rect 6178 92094 6190 92146
rect 6242 92094 6254 92146
rect 8530 92094 8542 92146
rect 8594 92094 8606 92146
rect 8978 92094 8990 92146
rect 9042 92094 9054 92146
rect 10210 92094 10222 92146
rect 10274 92094 10286 92146
rect 10434 92094 10446 92146
rect 10498 92094 10510 92146
rect 11218 92094 11230 92146
rect 11282 92094 11294 92146
rect 13570 92094 13582 92146
rect 13634 92094 13646 92146
rect 15922 92094 15934 92146
rect 15986 92094 15998 92146
rect 16370 92094 16382 92146
rect 16434 92094 16446 92146
rect 17826 92094 17838 92146
rect 17890 92094 17902 92146
rect 18610 92094 18622 92146
rect 18674 92094 18686 92146
rect 21074 92094 21086 92146
rect 21138 92094 21150 92146
rect 21410 92094 21422 92146
rect 21474 92094 21486 92146
rect 22642 92094 22654 92146
rect 22706 92094 22718 92146
rect 22866 92094 22878 92146
rect 22930 92094 22942 92146
rect 23650 92094 23662 92146
rect 23714 92094 23726 92146
rect 9662 92082 9714 92094
rect 17054 92082 17106 92094
rect 22094 92082 22146 92094
rect 20638 92034 20690 92046
rect 2258 91982 2270 92034
rect 2322 91982 2334 92034
rect 6626 91982 6638 92034
rect 6690 91982 6702 92034
rect 9202 91982 9214 92034
rect 9266 91982 9278 92034
rect 14018 91982 14030 92034
rect 14082 91982 14094 92034
rect 21634 91982 21646 92034
rect 21698 91982 21710 92034
rect 20638 91970 20690 91982
rect 1150 91922 1202 91934
rect 1150 91858 1202 91870
rect 5294 91922 5346 91934
rect 5294 91858 5346 91870
rect 7758 91922 7810 91934
rect 7758 91858 7810 91870
rect 15150 91922 15202 91934
rect 19182 91922 19234 91934
rect 30270 91922 30322 91934
rect 16594 91870 16606 91922
rect 16658 91870 16670 91922
rect 19506 91870 19518 91922
rect 19570 91870 19582 91922
rect 30594 91870 30606 91922
rect 30658 91870 30670 91922
rect 15150 91858 15202 91870
rect 19182 91858 19234 91870
rect 30270 91858 30322 91870
rect 672 91754 31024 91788
rect 672 91702 4466 91754
rect 4518 91702 4570 91754
rect 4622 91702 4674 91754
rect 4726 91702 24466 91754
rect 24518 91702 24570 91754
rect 24622 91702 24674 91754
rect 24726 91702 31024 91754
rect 672 91668 31024 91702
rect 8206 91586 8258 91598
rect 7074 91534 7086 91586
rect 7138 91534 7150 91586
rect 13906 91534 13918 91586
rect 13970 91534 13982 91586
rect 8206 91522 8258 91534
rect 12910 91474 12962 91486
rect 1698 91422 1710 91474
rect 1762 91422 1774 91474
rect 4610 91422 4622 91474
rect 4674 91422 4686 91474
rect 10882 91422 10894 91474
rect 10946 91422 10958 91474
rect 17714 91422 17726 91474
rect 17778 91422 17790 91474
rect 21522 91422 21534 91474
rect 21586 91422 21598 91474
rect 30594 91422 30606 91474
rect 30658 91422 30670 91474
rect 12910 91410 12962 91422
rect 12126 91362 12178 91374
rect 14366 91362 14418 91374
rect 18174 91362 18226 91374
rect 30270 91362 30322 91374
rect 6514 91310 6526 91362
rect 6578 91310 6590 91362
rect 13346 91310 13358 91362
rect 13410 91310 13422 91362
rect 13794 91310 13806 91362
rect 13858 91310 13870 91362
rect 14914 91310 14926 91362
rect 14978 91310 14990 91362
rect 15922 91310 15934 91362
rect 15986 91310 15998 91362
rect 17042 91310 17054 91362
rect 17106 91310 17118 91362
rect 17490 91310 17502 91362
rect 17554 91310 17566 91362
rect 18722 91310 18734 91362
rect 18786 91310 18798 91362
rect 19730 91310 19742 91362
rect 19794 91310 19806 91362
rect 21074 91310 21086 91362
rect 21138 91310 21150 91362
rect 12126 91298 12178 91310
rect 14366 91298 14418 91310
rect 18174 91298 18226 91310
rect 30270 91298 30322 91310
rect 16718 91250 16770 91262
rect 1250 91198 1262 91250
rect 1314 91198 1326 91250
rect 4946 91198 4958 91250
rect 5010 91198 5022 91250
rect 10546 91198 10558 91250
rect 10610 91198 10622 91250
rect 16718 91186 16770 91198
rect 2830 91138 2882 91150
rect 2830 91074 2882 91086
rect 3390 91138 3442 91150
rect 3390 91074 3442 91086
rect 22766 91138 22818 91150
rect 22766 91074 22818 91086
rect 672 90970 31024 91004
rect 672 90918 3806 90970
rect 3858 90918 3910 90970
rect 3962 90918 4014 90970
rect 4066 90918 23806 90970
rect 23858 90918 23910 90970
rect 23962 90918 24014 90970
rect 24066 90918 31024 90970
rect 672 90884 31024 90918
rect 9998 90802 10050 90814
rect 9998 90738 10050 90750
rect 15262 90802 15314 90814
rect 15262 90738 15314 90750
rect 6078 90690 6130 90702
rect 2706 90638 2718 90690
rect 2770 90638 2782 90690
rect 6078 90626 6130 90638
rect 22318 90690 22370 90702
rect 22318 90626 22370 90638
rect 7534 90578 7586 90590
rect 17166 90578 17218 90590
rect 6514 90526 6526 90578
rect 6578 90526 6590 90578
rect 6850 90526 6862 90578
rect 6914 90526 6926 90578
rect 8082 90526 8094 90578
rect 8146 90526 8158 90578
rect 9202 90526 9214 90578
rect 9266 90526 9278 90578
rect 11666 90526 11678 90578
rect 11730 90526 11742 90578
rect 13570 90526 13582 90578
rect 13634 90526 13646 90578
rect 16034 90526 16046 90578
rect 16098 90526 16110 90578
rect 16482 90526 16494 90578
rect 16546 90526 16558 90578
rect 17714 90526 17726 90578
rect 17778 90526 17790 90578
rect 18834 90526 18846 90578
rect 18898 90526 18910 90578
rect 7534 90514 7586 90526
rect 17166 90514 17218 90526
rect 12798 90466 12850 90478
rect 15710 90466 15762 90478
rect 7074 90414 7086 90466
rect 7138 90414 7150 90466
rect 13122 90414 13134 90466
rect 13186 90414 13198 90466
rect 21522 90414 21534 90466
rect 21586 90414 21598 90466
rect 22082 90414 22094 90466
rect 22146 90414 22158 90466
rect 12798 90402 12850 90414
rect 15710 90402 15762 90414
rect 1150 90354 1202 90366
rect 22654 90354 22706 90366
rect 2258 90302 2270 90354
rect 2322 90302 2334 90354
rect 11106 90302 11118 90354
rect 11170 90302 11182 90354
rect 14130 90302 14142 90354
rect 14194 90302 14206 90354
rect 16706 90302 16718 90354
rect 16770 90302 16782 90354
rect 1150 90290 1202 90302
rect 22654 90290 22706 90302
rect 672 90186 31024 90220
rect 672 90134 4466 90186
rect 4518 90134 4570 90186
rect 4622 90134 4674 90186
rect 4726 90134 24466 90186
rect 24518 90134 24570 90186
rect 24622 90134 24674 90186
rect 24726 90134 31024 90186
rect 672 90100 31024 90134
rect 12238 90018 12290 90030
rect 4050 89966 4062 90018
rect 4114 89966 4126 90018
rect 13906 89966 13918 90018
rect 13970 89966 13982 90018
rect 12238 89954 12290 89966
rect 4510 89906 4562 89918
rect 14366 89906 14418 89918
rect 30270 89906 30322 89918
rect 1586 89854 1598 89906
rect 1650 89854 1662 89906
rect 6738 89854 6750 89906
rect 6802 89854 6814 89906
rect 7186 89854 7198 89906
rect 7250 89854 7262 89906
rect 10098 89854 10110 89906
rect 10162 89854 10174 89906
rect 12562 89854 12574 89906
rect 12626 89854 12638 89906
rect 18274 89854 18286 89906
rect 18338 89854 18350 89906
rect 19506 89854 19518 89906
rect 19570 89854 19582 89906
rect 30594 89854 30606 89906
rect 30658 89854 30670 89906
rect 4510 89842 4562 89854
rect 14366 89842 14418 89854
rect 30270 89842 30322 89854
rect 2270 89794 2322 89806
rect 14590 89794 14642 89806
rect 20190 89794 20242 89806
rect 1474 89742 1486 89794
rect 1538 89742 1550 89794
rect 3490 89742 3502 89794
rect 3554 89742 3566 89794
rect 3826 89742 3838 89794
rect 3890 89742 3902 89794
rect 5282 89742 5294 89794
rect 5346 89742 5358 89794
rect 6178 89742 6190 89794
rect 6242 89742 6254 89794
rect 13234 89742 13246 89794
rect 13298 89742 13310 89794
rect 13794 89742 13806 89794
rect 13858 89742 13870 89794
rect 15026 89742 15038 89794
rect 15090 89742 15102 89794
rect 16034 89742 16046 89794
rect 16098 89742 16110 89794
rect 18722 89742 18734 89794
rect 18786 89742 18798 89794
rect 19394 89742 19406 89794
rect 19458 89742 19470 89794
rect 2270 89730 2322 89742
rect 14590 89730 14642 89742
rect 20190 89730 20242 89742
rect 3054 89682 3106 89694
rect 3054 89618 3106 89630
rect 7534 89682 7586 89694
rect 12910 89682 12962 89694
rect 9650 89630 9662 89682
rect 9714 89630 9726 89682
rect 7534 89618 7586 89630
rect 12910 89618 12962 89630
rect 2606 89570 2658 89582
rect 2606 89506 2658 89518
rect 7870 89570 7922 89582
rect 7870 89506 7922 89518
rect 11230 89570 11282 89582
rect 11230 89506 11282 89518
rect 17166 89570 17218 89582
rect 17166 89506 17218 89518
rect 20526 89570 20578 89582
rect 20526 89506 20578 89518
rect 672 89402 31024 89436
rect 672 89350 3806 89402
rect 3858 89350 3910 89402
rect 3962 89350 4014 89402
rect 4066 89350 23806 89402
rect 23858 89350 23910 89402
rect 23962 89350 24014 89402
rect 24066 89350 31024 89402
rect 672 89316 31024 89350
rect 14590 89234 14642 89246
rect 14590 89170 14642 89182
rect 18174 89234 18226 89246
rect 18174 89170 18226 89182
rect 5854 89122 5906 89134
rect 9650 89070 9662 89122
rect 9714 89070 9726 89122
rect 13010 89070 13022 89122
rect 13074 89070 13086 89122
rect 5854 89058 5906 89070
rect 7310 89010 7362 89022
rect 2594 88958 2606 89010
rect 2658 88958 2670 89010
rect 6178 88958 6190 89010
rect 6242 88958 6254 89010
rect 6626 88958 6638 89010
rect 6690 88958 6702 89010
rect 8082 88958 8094 89010
rect 8146 88958 8158 89010
rect 8978 88958 8990 89010
rect 9042 88958 9054 89010
rect 17490 88958 17502 89010
rect 17554 88958 17566 89010
rect 21410 88958 21422 89010
rect 21474 88958 21486 89010
rect 7310 88946 7362 88958
rect 3154 88846 3166 88898
rect 3218 88846 3230 88898
rect 6850 88846 6862 88898
rect 6914 88846 6926 88898
rect 9986 88846 9998 88898
rect 10050 88846 10062 88898
rect 13346 88846 13358 88898
rect 13410 88846 13422 88898
rect 17378 88846 17390 88898
rect 17442 88846 17454 88898
rect 21970 88846 21982 88898
rect 22034 88846 22046 88898
rect 4286 88786 4338 88798
rect 4286 88722 4338 88734
rect 11230 88786 11282 88798
rect 11230 88722 11282 88734
rect 18510 88786 18562 88798
rect 18510 88722 18562 88734
rect 23102 88786 23154 88798
rect 23102 88722 23154 88734
rect 30270 88786 30322 88798
rect 30594 88734 30606 88786
rect 30658 88734 30670 88786
rect 30270 88722 30322 88734
rect 672 88618 31024 88652
rect 672 88566 4466 88618
rect 4518 88566 4570 88618
rect 4622 88566 4674 88618
rect 4726 88566 24466 88618
rect 24518 88566 24570 88618
rect 24622 88566 24674 88618
rect 24726 88566 31024 88618
rect 672 88532 31024 88566
rect 1698 88398 1710 88450
rect 1762 88398 1774 88450
rect 21746 88398 21758 88450
rect 21810 88398 21822 88450
rect 29810 88398 29822 88450
rect 29874 88398 29886 88450
rect 4274 88286 4286 88338
rect 4338 88286 4350 88338
rect 11442 88286 11454 88338
rect 11506 88286 11518 88338
rect 13682 88286 13694 88338
rect 13746 88286 13758 88338
rect 18386 88286 18398 88338
rect 18450 88286 18462 88338
rect 29486 88226 29538 88238
rect 3602 88174 3614 88226
rect 3666 88174 3678 88226
rect 4050 88174 4062 88226
rect 4114 88174 4126 88226
rect 4834 88174 4846 88226
rect 4898 88174 4910 88226
rect 5282 88174 5294 88226
rect 5346 88174 5358 88226
rect 6402 88174 6414 88226
rect 6466 88174 6478 88226
rect 13234 88174 13246 88226
rect 13298 88174 13310 88226
rect 21186 88174 21198 88226
rect 21250 88174 21262 88226
rect 29486 88162 29538 88174
rect 3278 88114 3330 88126
rect 1250 88062 1262 88114
rect 1314 88062 1326 88114
rect 3278 88050 3330 88062
rect 7310 88114 7362 88126
rect 10994 88062 11006 88114
rect 11058 88062 11070 88114
rect 18050 88062 18062 88114
rect 18114 88062 18126 88114
rect 7310 88050 7362 88062
rect 2830 88002 2882 88014
rect 2830 87938 2882 87950
rect 12574 88002 12626 88014
rect 12574 87938 12626 87950
rect 14814 88002 14866 88014
rect 14814 87938 14866 87950
rect 19630 88002 19682 88014
rect 19630 87938 19682 87950
rect 22878 88002 22930 88014
rect 22878 87938 22930 87950
rect 672 87834 31024 87868
rect 672 87782 3806 87834
rect 3858 87782 3910 87834
rect 3962 87782 4014 87834
rect 4066 87782 23806 87834
rect 23858 87782 23910 87834
rect 23962 87782 24014 87834
rect 24066 87782 31024 87834
rect 672 87748 31024 87782
rect 12238 87554 12290 87566
rect 1810 87502 1822 87554
rect 1874 87502 1886 87554
rect 6290 87502 6302 87554
rect 6354 87502 6366 87554
rect 13122 87502 13134 87554
rect 13186 87502 13198 87554
rect 22306 87502 22318 87554
rect 22370 87502 22382 87554
rect 12238 87490 12290 87502
rect 10782 87442 10834 87454
rect 14702 87442 14754 87454
rect 22878 87442 22930 87454
rect 9090 87390 9102 87442
rect 9154 87390 9166 87442
rect 10098 87390 10110 87442
rect 10162 87390 10174 87442
rect 11442 87390 11454 87442
rect 11506 87390 11518 87442
rect 11778 87390 11790 87442
rect 11842 87390 11854 87442
rect 18274 87390 18286 87442
rect 18338 87390 18350 87442
rect 10782 87378 10834 87390
rect 14702 87378 14754 87390
rect 22878 87378 22930 87390
rect 30270 87442 30322 87454
rect 30270 87378 30322 87390
rect 2146 87278 2158 87330
rect 2210 87278 2222 87330
rect 6626 87278 6638 87330
rect 6690 87278 6702 87330
rect 11218 87278 11230 87330
rect 11282 87278 11294 87330
rect 21858 87278 21870 87330
rect 21922 87278 21934 87330
rect 23202 87278 23214 87330
rect 23266 87278 23278 87330
rect 23874 87278 23886 87330
rect 23938 87278 23950 87330
rect 3390 87218 3442 87230
rect 3390 87154 3442 87166
rect 7870 87218 7922 87230
rect 19966 87218 20018 87230
rect 13570 87166 13582 87218
rect 13634 87166 13646 87218
rect 18834 87166 18846 87218
rect 18898 87166 18910 87218
rect 7870 87154 7922 87166
rect 19966 87154 20018 87166
rect 20750 87218 20802 87230
rect 20750 87154 20802 87166
rect 23550 87218 23602 87230
rect 30594 87166 30606 87218
rect 30658 87166 30670 87218
rect 23550 87154 23602 87166
rect 672 87050 31024 87084
rect 672 86998 4466 87050
rect 4518 86998 4570 87050
rect 4622 86998 4674 87050
rect 4726 86998 24466 87050
rect 24518 86998 24570 87050
rect 24622 86998 24674 87050
rect 24726 86998 31024 87050
rect 672 86964 31024 86998
rect 22878 86882 22930 86894
rect 6402 86830 6414 86882
rect 6466 86830 6478 86882
rect 9874 86830 9886 86882
rect 9938 86830 9950 86882
rect 22878 86818 22930 86830
rect 11454 86770 11506 86782
rect 12910 86770 12962 86782
rect 1586 86718 1598 86770
rect 1650 86718 1662 86770
rect 4162 86718 4174 86770
rect 4226 86718 4238 86770
rect 12450 86718 12462 86770
rect 12514 86718 12526 86770
rect 11454 86706 11506 86718
rect 12910 86706 12962 86718
rect 18846 86770 18898 86782
rect 23438 86770 23490 86782
rect 19842 86718 19854 86770
rect 19906 86718 19918 86770
rect 30594 86718 30606 86770
rect 30658 86718 30670 86770
rect 18846 86706 18898 86718
rect 23438 86706 23490 86718
rect 11006 86658 11058 86670
rect 20526 86658 20578 86670
rect 22766 86658 22818 86670
rect 23550 86658 23602 86670
rect 3714 86606 3726 86658
rect 3778 86606 3790 86658
rect 5954 86606 5966 86658
rect 6018 86606 6030 86658
rect 9426 86606 9438 86658
rect 9490 86606 9502 86658
rect 11778 86606 11790 86658
rect 11842 86606 11854 86658
rect 12338 86606 12350 86658
rect 12402 86606 12414 86658
rect 13458 86606 13470 86658
rect 13522 86606 13534 86658
rect 14578 86606 14590 86658
rect 14642 86606 14654 86658
rect 19282 86606 19294 86658
rect 19346 86606 19358 86658
rect 19618 86606 19630 86658
rect 19682 86606 19694 86658
rect 20850 86606 20862 86658
rect 20914 86606 20926 86658
rect 21858 86606 21870 86658
rect 21922 86606 21934 86658
rect 22978 86606 22990 86658
rect 23042 86606 23054 86658
rect 11006 86594 11058 86606
rect 20526 86594 20578 86606
rect 22766 86594 22818 86606
rect 23550 86594 23602 86606
rect 30270 86658 30322 86670
rect 30270 86594 30322 86606
rect 23998 86546 24050 86558
rect 1250 86494 1262 86546
rect 1314 86494 1326 86546
rect 23998 86482 24050 86494
rect 2830 86434 2882 86446
rect 2830 86370 2882 86382
rect 5294 86434 5346 86446
rect 5294 86370 5346 86382
rect 7534 86434 7586 86446
rect 7534 86370 7586 86382
rect 22542 86434 22594 86446
rect 22542 86370 22594 86382
rect 23438 86434 23490 86446
rect 23438 86370 23490 86382
rect 23886 86434 23938 86446
rect 23886 86370 23938 86382
rect 672 86266 31024 86300
rect 672 86214 3806 86266
rect 3858 86214 3910 86266
rect 3962 86214 4014 86266
rect 4066 86214 23806 86266
rect 23858 86214 23910 86266
rect 23962 86214 24014 86266
rect 24066 86214 31024 86266
rect 672 86180 31024 86214
rect 19966 86098 20018 86110
rect 19966 86034 20018 86046
rect 23326 86098 23378 86110
rect 23326 86034 23378 86046
rect 7982 85986 8034 85998
rect 15150 85986 15202 85998
rect 2706 85934 2718 85986
rect 2770 85934 2782 85986
rect 7074 85934 7086 85986
rect 7138 85934 7150 85986
rect 13010 85934 13022 85986
rect 13074 85934 13086 85986
rect 22306 85934 22318 85986
rect 22370 85934 22382 85986
rect 7982 85922 8034 85934
rect 15150 85922 15202 85934
rect 9438 85874 9490 85886
rect 19630 85874 19682 85886
rect 23550 85874 23602 85886
rect 1250 85822 1262 85874
rect 1314 85822 1326 85874
rect 8418 85822 8430 85874
rect 8482 85822 8494 85874
rect 8866 85822 8878 85874
rect 8930 85822 8942 85874
rect 10210 85822 10222 85874
rect 10274 85822 10286 85874
rect 10994 85822 11006 85874
rect 11058 85822 11070 85874
rect 15474 85822 15486 85874
rect 15538 85822 15550 85874
rect 16034 85822 16046 85874
rect 16098 85822 16110 85874
rect 17154 85822 17166 85874
rect 17218 85822 17230 85874
rect 18162 85822 18174 85874
rect 18226 85822 18238 85874
rect 22866 85822 22878 85874
rect 22930 85822 22942 85874
rect 23090 85822 23102 85874
rect 23154 85822 23166 85874
rect 9438 85810 9490 85822
rect 19630 85810 19682 85822
rect 23550 85810 23602 85822
rect 23774 85874 23826 85886
rect 23774 85810 23826 85822
rect 14590 85762 14642 85774
rect 16606 85762 16658 85774
rect 20750 85762 20802 85774
rect 1026 85710 1038 85762
rect 1090 85710 1102 85762
rect 6738 85710 6750 85762
rect 6802 85710 6814 85762
rect 8978 85710 8990 85762
rect 9042 85710 9054 85762
rect 13458 85710 13470 85762
rect 13522 85710 13534 85762
rect 16146 85710 16158 85762
rect 16210 85710 16222 85762
rect 19058 85710 19070 85762
rect 19122 85710 19134 85762
rect 19394 85710 19406 85762
rect 19458 85710 19470 85762
rect 14590 85698 14642 85710
rect 16606 85698 16658 85710
rect 20750 85698 20802 85710
rect 24110 85762 24162 85774
rect 24434 85710 24446 85762
rect 24498 85710 24510 85762
rect 24110 85698 24162 85710
rect 2158 85650 2210 85662
rect 4286 85650 4338 85662
rect 1810 85598 1822 85650
rect 1874 85598 1886 85650
rect 3154 85598 3166 85650
rect 3218 85598 3230 85650
rect 2158 85586 2210 85598
rect 4286 85586 4338 85598
rect 5518 85650 5570 85662
rect 23886 85650 23938 85662
rect 21858 85598 21870 85650
rect 21922 85598 21934 85650
rect 5518 85586 5570 85598
rect 23886 85586 23938 85598
rect 672 85482 31024 85516
rect 672 85430 4466 85482
rect 4518 85430 4570 85482
rect 4622 85430 4674 85482
rect 4726 85430 24466 85482
rect 24518 85430 24570 85482
rect 24622 85430 24674 85482
rect 24726 85430 31024 85482
rect 672 85396 31024 85430
rect 23102 85314 23154 85326
rect 17378 85262 17390 85314
rect 17442 85262 17454 85314
rect 20402 85262 20414 85314
rect 20466 85262 20478 85314
rect 23102 85250 23154 85262
rect 23550 85314 23602 85326
rect 23550 85250 23602 85262
rect 22990 85202 23042 85214
rect 30270 85202 30322 85214
rect 1026 85150 1038 85202
rect 1090 85150 1102 85202
rect 2818 85150 2830 85202
rect 2882 85150 2894 85202
rect 6738 85150 6750 85202
rect 6802 85150 6814 85202
rect 11218 85150 11230 85202
rect 11282 85150 11294 85202
rect 13906 85150 13918 85202
rect 13970 85150 13982 85202
rect 23874 85150 23886 85202
rect 23938 85150 23950 85202
rect 30594 85150 30606 85202
rect 30658 85150 30670 85202
rect 22990 85138 23042 85150
rect 30270 85138 30322 85150
rect 1374 85090 1426 85102
rect 3502 85090 3554 85102
rect 12462 85090 12514 85102
rect 14590 85090 14642 85102
rect 21086 85090 21138 85102
rect 2258 85038 2270 85090
rect 2322 85038 2334 85090
rect 2594 85038 2606 85090
rect 2658 85038 2670 85090
rect 3826 85038 3838 85090
rect 3890 85038 3902 85090
rect 4834 85038 4846 85090
rect 4898 85038 4910 85090
rect 7186 85038 7198 85090
rect 7250 85038 7262 85090
rect 10882 85038 10894 85090
rect 10946 85038 10958 85090
rect 13234 85038 13246 85090
rect 13298 85038 13310 85090
rect 13794 85038 13806 85090
rect 13858 85038 13870 85090
rect 14914 85038 14926 85090
rect 14978 85038 14990 85090
rect 16034 85038 16046 85090
rect 16098 85038 16110 85090
rect 16818 85038 16830 85090
rect 16882 85038 16894 85090
rect 19730 85038 19742 85090
rect 19794 85038 19806 85090
rect 20178 85038 20190 85090
rect 20242 85038 20254 85090
rect 21410 85038 21422 85090
rect 21474 85038 21486 85090
rect 22530 85038 22542 85090
rect 22594 85038 22606 85090
rect 1374 85026 1426 85038
rect 3502 85026 3554 85038
rect 12462 85026 12514 85038
rect 14590 85026 14642 85038
rect 21086 85026 21138 85038
rect 1822 84978 1874 84990
rect 1822 84914 1874 84926
rect 12910 84978 12962 84990
rect 12910 84914 12962 84926
rect 19406 84978 19458 84990
rect 19406 84914 19458 84926
rect 5518 84866 5570 84878
rect 5518 84802 5570 84814
rect 18510 84866 18562 84878
rect 18510 84802 18562 84814
rect 672 84698 31024 84732
rect 672 84646 3806 84698
rect 3858 84646 3910 84698
rect 3962 84646 4014 84698
rect 4066 84646 23806 84698
rect 23858 84646 23910 84698
rect 23962 84646 24014 84698
rect 24066 84646 31024 84698
rect 672 84612 31024 84646
rect 7422 84418 7474 84430
rect 7422 84354 7474 84366
rect 11342 84418 11394 84430
rect 11342 84354 11394 84366
rect 15038 84418 15090 84430
rect 15038 84354 15090 84366
rect 20638 84418 20690 84430
rect 20638 84354 20690 84366
rect 2830 84306 2882 84318
rect 8878 84306 8930 84318
rect 16494 84306 16546 84318
rect 19070 84306 19122 84318
rect 22094 84306 22146 84318
rect 1474 84254 1486 84306
rect 1538 84254 1550 84306
rect 2034 84254 2046 84306
rect 2098 84254 2110 84306
rect 3154 84254 3166 84306
rect 3218 84254 3230 84306
rect 3378 84254 3390 84306
rect 3442 84254 3454 84306
rect 4162 84254 4174 84306
rect 4226 84254 4238 84306
rect 5282 84254 5294 84306
rect 5346 84254 5358 84306
rect 7858 84254 7870 84306
rect 7922 84254 7934 84306
rect 8194 84254 8206 84306
rect 8258 84254 8270 84306
rect 9650 84254 9662 84306
rect 9714 84254 9726 84306
rect 10546 84254 10558 84306
rect 10610 84254 10622 84306
rect 15362 84254 15374 84306
rect 15426 84254 15438 84306
rect 15922 84254 15934 84306
rect 15986 84254 15998 84306
rect 17042 84254 17054 84306
rect 17106 84254 17118 84306
rect 17266 84254 17278 84306
rect 17330 84254 17342 84306
rect 18050 84254 18062 84306
rect 18114 84254 18126 84306
rect 20962 84254 20974 84306
rect 21026 84254 21038 84306
rect 21410 84254 21422 84306
rect 21474 84254 21486 84306
rect 22642 84254 22654 84306
rect 22706 84254 22718 84306
rect 23650 84254 23662 84306
rect 23714 84254 23726 84306
rect 2830 84242 2882 84254
rect 8878 84242 8930 84254
rect 16494 84242 16546 84254
rect 19070 84242 19122 84254
rect 22094 84242 22146 84254
rect 1150 84194 1202 84206
rect 13022 84194 13074 84206
rect 5842 84142 5854 84194
rect 5906 84142 5918 84194
rect 16034 84142 16046 84194
rect 16098 84142 16110 84194
rect 19282 84142 19294 84194
rect 19346 84142 19358 84194
rect 19618 84142 19630 84194
rect 19682 84142 19694 84194
rect 21634 84142 21646 84194
rect 21698 84142 21710 84194
rect 1150 84130 1202 84142
rect 13022 84130 13074 84142
rect 6974 84082 7026 84094
rect 12798 84082 12850 84094
rect 2146 84030 2158 84082
rect 2210 84030 2222 84082
rect 8418 84030 8430 84082
rect 8482 84030 8494 84082
rect 6974 84018 7026 84030
rect 12798 84018 12850 84030
rect 18734 84082 18786 84094
rect 18734 84018 18786 84030
rect 30270 84082 30322 84094
rect 30594 84030 30606 84082
rect 30658 84030 30670 84082
rect 30270 84018 30322 84030
rect 672 83914 31024 83948
rect 672 83862 4466 83914
rect 4518 83862 4570 83914
rect 4622 83862 4674 83914
rect 4726 83862 24466 83914
rect 24518 83862 24570 83914
rect 24622 83862 24674 83914
rect 24726 83862 31024 83914
rect 672 83828 31024 83862
rect 4286 83746 4338 83758
rect 22094 83746 22146 83758
rect 1362 83694 1374 83746
rect 1426 83694 1438 83746
rect 9874 83694 9886 83746
rect 9938 83694 9950 83746
rect 23650 83694 23662 83746
rect 23714 83694 23726 83746
rect 4286 83682 4338 83694
rect 22094 83682 22146 83694
rect 6526 83634 6578 83646
rect 2370 83582 2382 83634
rect 2434 83582 2446 83634
rect 3938 83582 3950 83634
rect 4002 83582 4014 83634
rect 6066 83582 6078 83634
rect 6130 83582 6142 83634
rect 6526 83570 6578 83582
rect 8878 83634 8930 83646
rect 16718 83634 16770 83646
rect 14914 83582 14926 83634
rect 14978 83582 14990 83634
rect 17714 83582 17726 83634
rect 17778 83582 17790 83634
rect 20850 83582 20862 83634
rect 20914 83582 20926 83634
rect 30594 83582 30606 83634
rect 30658 83582 30670 83634
rect 8878 83570 8930 83582
rect 16718 83570 16770 83582
rect 1038 83522 1090 83534
rect 10334 83522 10386 83534
rect 16046 83522 16098 83534
rect 18398 83522 18450 83534
rect 23326 83522 23378 83534
rect 1810 83470 1822 83522
rect 1874 83470 1886 83522
rect 5394 83470 5406 83522
rect 5458 83470 5470 83522
rect 5842 83470 5854 83522
rect 5906 83470 5918 83522
rect 7298 83470 7310 83522
rect 7362 83470 7374 83522
rect 8082 83470 8094 83522
rect 8146 83470 8158 83522
rect 9202 83470 9214 83522
rect 9266 83470 9278 83522
rect 9650 83470 9662 83522
rect 9714 83470 9726 83522
rect 11106 83470 11118 83522
rect 11170 83470 11182 83522
rect 12002 83470 12014 83522
rect 12066 83470 12078 83522
rect 13906 83470 13918 83522
rect 13970 83470 13982 83522
rect 17042 83470 17054 83522
rect 17106 83470 17118 83522
rect 17490 83470 17502 83522
rect 17554 83470 17566 83522
rect 18722 83470 18734 83522
rect 18786 83470 18798 83522
rect 19730 83470 19742 83522
rect 19794 83470 19806 83522
rect 20402 83470 20414 83522
rect 20466 83470 20478 83522
rect 1038 83458 1090 83470
rect 10334 83458 10386 83470
rect 16046 83458 16098 83470
rect 18398 83458 18450 83470
rect 23326 83458 23378 83470
rect 30270 83522 30322 83534
rect 30270 83458 30322 83470
rect 5070 83410 5122 83422
rect 14466 83358 14478 83410
rect 14530 83358 14542 83410
rect 5070 83346 5122 83358
rect 3502 83298 3554 83310
rect 3502 83234 3554 83246
rect 13358 83298 13410 83310
rect 13358 83234 13410 83246
rect 13470 83298 13522 83310
rect 13470 83234 13522 83246
rect 13694 83298 13746 83310
rect 13694 83234 13746 83246
rect 672 83130 31024 83164
rect 672 83078 3806 83130
rect 3858 83078 3910 83130
rect 3962 83078 4014 83130
rect 4066 83078 23806 83130
rect 23858 83078 23910 83130
rect 23962 83078 24014 83130
rect 24066 83078 31024 83130
rect 672 83044 31024 83078
rect 9886 82962 9938 82974
rect 9886 82898 9938 82910
rect 17726 82962 17778 82974
rect 17726 82898 17778 82910
rect 5842 82798 5854 82850
rect 5906 82798 5918 82850
rect 2830 82738 2882 82750
rect 1586 82686 1598 82738
rect 1650 82686 1662 82738
rect 1922 82686 1934 82738
rect 1986 82686 1998 82738
rect 3154 82686 3166 82738
rect 3218 82686 3230 82738
rect 4162 82686 4174 82738
rect 4226 82686 4238 82738
rect 8306 82686 8318 82738
rect 8370 82686 8382 82738
rect 10546 82686 10558 82738
rect 10610 82686 10622 82738
rect 14466 82686 14478 82738
rect 14530 82686 14542 82738
rect 16034 82686 16046 82738
rect 16098 82686 16110 82738
rect 18274 82686 18286 82738
rect 18338 82686 18350 82738
rect 2830 82674 2882 82686
rect 1150 82626 1202 82638
rect 6178 82574 6190 82626
rect 6242 82574 6254 82626
rect 8754 82574 8766 82626
rect 8818 82574 8830 82626
rect 10882 82574 10894 82626
rect 10946 82574 10958 82626
rect 14130 82574 14142 82626
rect 14194 82574 14206 82626
rect 16482 82574 16494 82626
rect 16546 82574 16558 82626
rect 22866 82574 22878 82626
rect 22930 82574 22942 82626
rect 1150 82562 1202 82574
rect 4958 82514 5010 82526
rect 7422 82514 7474 82526
rect 2146 82462 2158 82514
rect 2210 82462 2222 82514
rect 5282 82462 5294 82514
rect 5346 82462 5358 82514
rect 4958 82450 5010 82462
rect 7422 82450 7474 82462
rect 12126 82514 12178 82526
rect 12126 82450 12178 82462
rect 12910 82514 12962 82526
rect 22542 82514 22594 82526
rect 18498 82462 18510 82514
rect 18562 82462 18574 82514
rect 12910 82450 12962 82462
rect 22542 82450 22594 82462
rect 672 82346 31024 82380
rect 672 82294 4466 82346
rect 4518 82294 4570 82346
rect 4622 82294 4674 82346
rect 4726 82294 24466 82346
rect 24518 82294 24570 82346
rect 24622 82294 24674 82346
rect 24726 82294 31024 82346
rect 672 82260 31024 82294
rect 8318 82178 8370 82190
rect 8318 82114 8370 82126
rect 8990 82178 9042 82190
rect 8990 82114 9042 82126
rect 3726 82066 3778 82078
rect 5182 82066 5234 82078
rect 12014 82066 12066 82078
rect 13470 82066 13522 82078
rect 2146 82014 2158 82066
rect 2210 82014 2222 82066
rect 4722 82014 4734 82066
rect 4786 82014 4798 82066
rect 7298 82014 7310 82066
rect 7362 82014 7374 82066
rect 7970 82014 7982 82066
rect 8034 82014 8046 82066
rect 10210 82014 10222 82066
rect 10274 82014 10286 82066
rect 13010 82014 13022 82066
rect 13074 82014 13086 82066
rect 3726 82002 3778 82014
rect 5182 82002 5234 82014
rect 12014 82002 12066 82014
rect 13470 82002 13522 82014
rect 15710 82066 15762 82078
rect 30270 82066 30322 82078
rect 19954 82014 19966 82066
rect 20018 82014 20030 82066
rect 22754 82014 22766 82066
rect 22818 82014 22830 82066
rect 29810 82014 29822 82066
rect 29874 82014 29886 82066
rect 30594 82014 30606 82066
rect 30658 82014 30670 82066
rect 15710 82002 15762 82014
rect 30270 82002 30322 82014
rect 15486 81954 15538 81966
rect 4050 81902 4062 81954
rect 4114 81902 4126 81954
rect 4498 81902 4510 81954
rect 4562 81902 4574 81954
rect 5730 81902 5742 81954
rect 5794 81902 5806 81954
rect 6738 81902 6750 81954
rect 6802 81902 6814 81954
rect 7522 81902 7534 81954
rect 7586 81902 7598 81954
rect 10658 81902 10670 81954
rect 10722 81902 10734 81954
rect 12338 81902 12350 81954
rect 12402 81902 12414 81954
rect 12786 81902 12798 81954
rect 12850 81902 12862 81954
rect 14242 81902 14254 81954
rect 14306 81902 14318 81954
rect 15026 81902 15038 81954
rect 15090 81902 15102 81954
rect 15486 81890 15538 81902
rect 15822 81954 15874 81966
rect 29486 81954 29538 81966
rect 19394 81902 19406 81954
rect 19458 81902 19470 81954
rect 15822 81890 15874 81902
rect 29486 81890 29538 81902
rect 1698 81790 1710 81842
rect 1762 81790 1774 81842
rect 23202 81790 23214 81842
rect 23266 81790 23278 81842
rect 3278 81730 3330 81742
rect 3278 81666 3330 81678
rect 21086 81730 21138 81742
rect 21086 81666 21138 81678
rect 21646 81730 21698 81742
rect 21646 81666 21698 81678
rect 672 81562 31024 81596
rect 672 81510 3806 81562
rect 3858 81510 3910 81562
rect 3962 81510 4014 81562
rect 4066 81510 23806 81562
rect 23858 81510 23910 81562
rect 23962 81510 24014 81562
rect 24066 81510 31024 81562
rect 672 81476 31024 81510
rect 10882 81230 10894 81282
rect 10946 81230 10958 81282
rect 15698 81230 15710 81282
rect 15762 81230 15774 81282
rect 20850 81230 20862 81282
rect 20914 81230 20926 81282
rect 14590 81170 14642 81182
rect 1698 81118 1710 81170
rect 1762 81118 1774 81170
rect 6178 81118 6190 81170
rect 6242 81118 6254 81170
rect 8530 81118 8542 81170
rect 8594 81118 8606 81170
rect 12898 81118 12910 81170
rect 12962 81118 12974 81170
rect 14590 81106 14642 81118
rect 15038 81170 15090 81182
rect 15038 81106 15090 81118
rect 10558 81058 10610 81070
rect 2034 81006 2046 81058
rect 2098 81006 2110 81058
rect 6626 81006 6638 81058
rect 6690 81006 6702 81058
rect 8866 81006 8878 81058
rect 8930 81006 8942 81058
rect 16034 81006 16046 81058
rect 16098 81006 16110 81058
rect 21186 81006 21198 81058
rect 21250 81006 21262 81058
rect 10558 80994 10610 81006
rect 3278 80946 3330 80958
rect 4286 80946 4338 80958
rect 5294 80946 5346 80958
rect 3938 80894 3950 80946
rect 4002 80894 4014 80946
rect 4946 80894 4958 80946
rect 5010 80894 5022 80946
rect 3278 80882 3330 80894
rect 4286 80882 4338 80894
rect 5294 80882 5346 80894
rect 7870 80946 7922 80958
rect 7870 80882 7922 80894
rect 10110 80946 10162 80958
rect 10110 80882 10162 80894
rect 10782 80946 10834 80958
rect 15150 80946 15202 80958
rect 17278 80946 17330 80958
rect 13458 80894 13470 80946
rect 13522 80894 13534 80946
rect 16146 80894 16158 80946
rect 16210 80894 16222 80946
rect 10782 80882 10834 80894
rect 15150 80882 15202 80894
rect 17278 80882 17330 80894
rect 22430 80946 22482 80958
rect 22430 80882 22482 80894
rect 30270 80946 30322 80958
rect 30594 80894 30606 80946
rect 30658 80894 30670 80946
rect 30270 80882 30322 80894
rect 672 80778 31024 80812
rect 672 80726 4466 80778
rect 4518 80726 4570 80778
rect 4622 80726 4674 80778
rect 4726 80726 24466 80778
rect 24518 80726 24570 80778
rect 24622 80726 24674 80778
rect 24726 80726 31024 80778
rect 672 80692 31024 80726
rect 14030 80610 14082 80622
rect 12898 80558 12910 80610
rect 12962 80558 12974 80610
rect 14914 80558 14926 80610
rect 14978 80558 14990 80610
rect 18834 80558 18846 80610
rect 18898 80558 18910 80610
rect 21410 80558 21422 80610
rect 21474 80558 21486 80610
rect 29810 80558 29822 80610
rect 29874 80558 29886 80610
rect 14030 80546 14082 80558
rect 2942 80498 2994 80510
rect 2482 80446 2494 80498
rect 2546 80446 2558 80498
rect 2942 80434 2994 80446
rect 5070 80498 5122 80510
rect 6526 80498 6578 80510
rect 15262 80498 15314 80510
rect 6066 80446 6078 80498
rect 6130 80446 6142 80498
rect 9874 80446 9886 80498
rect 9938 80446 9950 80498
rect 15026 80446 15038 80498
rect 15090 80446 15102 80498
rect 5070 80434 5122 80446
rect 6526 80434 6578 80446
rect 15262 80434 15314 80446
rect 20414 80498 20466 80510
rect 20414 80434 20466 80446
rect 21870 80498 21922 80510
rect 21870 80434 21922 80446
rect 14814 80386 14866 80398
rect 29486 80386 29538 80398
rect 1922 80334 1934 80386
rect 1986 80334 1998 80386
rect 2370 80334 2382 80386
rect 2434 80334 2446 80386
rect 3602 80334 3614 80386
rect 3666 80334 3678 80386
rect 4498 80334 4510 80386
rect 4562 80334 4574 80386
rect 5506 80334 5518 80386
rect 5570 80334 5582 80386
rect 5842 80334 5854 80386
rect 5906 80334 5918 80386
rect 7074 80334 7086 80386
rect 7138 80334 7150 80386
rect 8082 80334 8094 80386
rect 8146 80334 8158 80386
rect 12338 80334 12350 80386
rect 12402 80334 12414 80386
rect 14466 80334 14478 80386
rect 14530 80334 14542 80386
rect 18386 80334 18398 80386
rect 18450 80334 18462 80386
rect 20850 80334 20862 80386
rect 20914 80334 20926 80386
rect 21186 80334 21198 80386
rect 21250 80334 21262 80386
rect 22642 80334 22654 80386
rect 22706 80334 22718 80386
rect 23538 80334 23550 80386
rect 23602 80334 23614 80386
rect 14814 80322 14866 80334
rect 29486 80322 29538 80334
rect 1486 80274 1538 80286
rect 9538 80222 9550 80274
rect 9602 80222 9614 80274
rect 1486 80210 1538 80222
rect 11118 80162 11170 80174
rect 11118 80098 11170 80110
rect 19966 80162 20018 80174
rect 19966 80098 20018 80110
rect 672 79994 31024 80028
rect 672 79942 3806 79994
rect 3858 79942 3910 79994
rect 3962 79942 4014 79994
rect 4066 79942 23806 79994
rect 23858 79942 23910 79994
rect 23962 79942 24014 79994
rect 24066 79942 31024 79994
rect 672 79908 31024 79942
rect 14366 79826 14418 79838
rect 14366 79762 14418 79774
rect 8430 79714 8482 79726
rect 8430 79650 8482 79662
rect 20638 79714 20690 79726
rect 20638 79650 20690 79662
rect 12238 79602 12290 79614
rect 15598 79602 15650 79614
rect 17278 79602 17330 79614
rect 22318 79602 22370 79614
rect 1250 79550 1262 79602
rect 1314 79550 1326 79602
rect 3378 79550 3390 79602
rect 3442 79550 3454 79602
rect 4274 79550 4286 79602
rect 4338 79550 4350 79602
rect 7186 79550 7198 79602
rect 7250 79550 7262 79602
rect 8754 79550 8766 79602
rect 8818 79550 8830 79602
rect 9202 79550 9214 79602
rect 9266 79550 9278 79602
rect 9986 79550 9998 79602
rect 10050 79550 10062 79602
rect 10658 79550 10670 79602
rect 10722 79550 10734 79602
rect 11442 79550 11454 79602
rect 11506 79550 11518 79602
rect 14354 79550 14366 79602
rect 14418 79550 14430 79602
rect 15922 79550 15934 79602
rect 15986 79550 15998 79602
rect 16370 79550 16382 79602
rect 16434 79550 16446 79602
rect 17826 79550 17838 79602
rect 17890 79550 17902 79602
rect 18610 79550 18622 79602
rect 18674 79550 18686 79602
rect 20962 79550 20974 79602
rect 21026 79550 21038 79602
rect 21410 79550 21422 79602
rect 21474 79550 21486 79602
rect 22642 79550 22654 79602
rect 22706 79550 22718 79602
rect 23762 79550 23774 79602
rect 23826 79550 23838 79602
rect 12238 79538 12290 79550
rect 15598 79538 15650 79550
rect 17278 79538 17330 79550
rect 22318 79538 22370 79550
rect 12126 79490 12178 79502
rect 6738 79438 6750 79490
rect 6802 79438 6814 79490
rect 12126 79426 12178 79438
rect 14030 79490 14082 79502
rect 22094 79490 22146 79502
rect 16594 79438 16606 79490
rect 16658 79438 16670 79490
rect 14030 79426 14082 79438
rect 22094 79426 22146 79438
rect 2830 79378 2882 79390
rect 5630 79378 5682 79390
rect 8094 79378 8146 79390
rect 11902 79378 11954 79390
rect 29486 79378 29538 79390
rect 30270 79378 30322 79390
rect 1698 79326 1710 79378
rect 1762 79326 1774 79378
rect 3602 79326 3614 79378
rect 3666 79326 3678 79378
rect 4050 79326 4062 79378
rect 4114 79326 4126 79378
rect 7746 79326 7758 79378
rect 7810 79326 7822 79378
rect 9426 79326 9438 79378
rect 9490 79326 9502 79378
rect 21634 79326 21646 79378
rect 21698 79326 21710 79378
rect 29810 79326 29822 79378
rect 29874 79326 29886 79378
rect 30594 79326 30606 79378
rect 30658 79326 30670 79378
rect 2830 79314 2882 79326
rect 5630 79314 5682 79326
rect 8094 79314 8146 79326
rect 11902 79314 11954 79326
rect 29486 79314 29538 79326
rect 30270 79314 30322 79326
rect 672 79210 31024 79244
rect 672 79158 4466 79210
rect 4518 79158 4570 79210
rect 4622 79158 4674 79210
rect 4726 79158 24466 79210
rect 24518 79158 24570 79210
rect 24622 79158 24674 79210
rect 24726 79158 31024 79210
rect 672 79124 31024 79158
rect 15934 79042 15986 79054
rect 11442 78990 11454 79042
rect 11506 78990 11518 79042
rect 17714 78990 17726 79042
rect 17778 78990 17790 79042
rect 15934 78978 15986 78990
rect 11902 78930 11954 78942
rect 16718 78930 16770 78942
rect 2370 78878 2382 78930
rect 2434 78878 2446 78930
rect 3938 78878 3950 78930
rect 4002 78878 4014 78930
rect 5506 78878 5518 78930
rect 5570 78878 5582 78930
rect 6850 78878 6862 78930
rect 6914 78878 6926 78930
rect 9538 78878 9550 78930
rect 9602 78878 9614 78930
rect 11666 78878 11678 78930
rect 11730 78878 11742 78930
rect 14802 78878 14814 78930
rect 14866 78878 14878 78930
rect 11902 78866 11954 78878
rect 16718 78866 16770 78878
rect 20302 78930 20354 78942
rect 21298 78878 21310 78930
rect 21362 78878 21374 78930
rect 30594 78878 30606 78930
rect 30658 78878 30670 78930
rect 20302 78866 20354 78878
rect 5854 78818 5906 78830
rect 12686 78818 12738 78830
rect 18174 78818 18226 78830
rect 21982 78818 22034 78830
rect 30270 78818 30322 78830
rect 2706 78766 2718 78818
rect 2770 78766 2782 78818
rect 6402 78766 6414 78818
rect 6466 78766 6478 78818
rect 11106 78766 11118 78818
rect 11170 78766 11182 78818
rect 14242 78766 14254 78818
rect 14306 78766 14318 78818
rect 17042 78766 17054 78818
rect 17106 78766 17118 78818
rect 17490 78766 17502 78818
rect 17554 78766 17566 78818
rect 18722 78766 18734 78818
rect 18786 78766 18798 78818
rect 19730 78766 19742 78818
rect 19794 78766 19806 78818
rect 20738 78766 20750 78818
rect 20802 78766 20814 78818
rect 21074 78766 21086 78818
rect 21138 78766 21150 78818
rect 22306 78766 22318 78818
rect 22370 78766 22382 78818
rect 23314 78766 23326 78818
rect 23378 78766 23390 78818
rect 5854 78754 5906 78766
rect 12686 78754 12738 78766
rect 18174 78754 18226 78766
rect 21982 78754 22034 78766
rect 30270 78754 30322 78766
rect 3490 78654 3502 78706
rect 3554 78654 3566 78706
rect 9090 78654 9102 78706
rect 9154 78654 9166 78706
rect 14354 78654 14366 78706
rect 14418 78654 14430 78706
rect 1150 78594 1202 78606
rect 1150 78530 1202 78542
rect 5070 78594 5122 78606
rect 5070 78530 5122 78542
rect 8094 78594 8146 78606
rect 8094 78530 8146 78542
rect 10670 78594 10722 78606
rect 10670 78530 10722 78542
rect 11454 78594 11506 78606
rect 11454 78530 11506 78542
rect 12238 78594 12290 78606
rect 12238 78530 12290 78542
rect 12350 78594 12402 78606
rect 12350 78530 12402 78542
rect 12574 78594 12626 78606
rect 12574 78530 12626 78542
rect 672 78426 31024 78460
rect 672 78374 3806 78426
rect 3858 78374 3910 78426
rect 3962 78374 4014 78426
rect 4066 78374 23806 78426
rect 23858 78374 23910 78426
rect 23962 78374 24014 78426
rect 24066 78374 31024 78426
rect 672 78340 31024 78374
rect 12126 78258 12178 78270
rect 12126 78194 12178 78206
rect 17614 78258 17666 78270
rect 17614 78194 17666 78206
rect 9438 78146 9490 78158
rect 12238 78146 12290 78158
rect 1250 78094 1262 78146
rect 1314 78094 1326 78146
rect 10098 78094 10110 78146
rect 10162 78094 10174 78146
rect 13010 78094 13022 78146
rect 13074 78094 13086 78146
rect 9438 78082 9490 78094
rect 12238 78082 12290 78094
rect 4162 77982 4174 78034
rect 4226 77982 4238 78034
rect 5618 77982 5630 78034
rect 5682 77982 5694 78034
rect 7858 77982 7870 78034
rect 7922 77982 7934 78034
rect 15474 77982 15486 78034
rect 15538 77982 15550 78034
rect 19170 77982 19182 78034
rect 19234 77982 19246 78034
rect 22418 77982 22430 78034
rect 22482 77982 22494 78034
rect 29486 77922 29538 77934
rect 1698 77870 1710 77922
rect 1762 77870 1774 77922
rect 6066 77870 6078 77922
rect 6130 77870 6142 77922
rect 8306 77870 8318 77922
rect 8370 77870 8382 77922
rect 13346 77870 13358 77922
rect 13410 77870 13422 77922
rect 15922 77870 15934 77922
rect 15986 77870 15998 77922
rect 21858 77870 21870 77922
rect 21922 77870 21934 77922
rect 29810 77870 29822 77922
rect 29874 77870 29886 77922
rect 29486 77858 29538 77870
rect 2830 77810 2882 77822
rect 2830 77746 2882 77758
rect 3278 77810 3330 77822
rect 7198 77810 7250 77822
rect 11678 77810 11730 77822
rect 3602 77758 3614 77810
rect 3666 77758 3678 77810
rect 3938 77758 3950 77810
rect 4002 77758 4014 77810
rect 10546 77758 10558 77810
rect 10610 77758 10622 77810
rect 3278 77746 3330 77758
rect 7198 77746 7250 77758
rect 11678 77746 11730 77758
rect 14590 77810 14642 77822
rect 14590 77746 14642 77758
rect 17054 77810 17106 77822
rect 20750 77810 20802 77822
rect 18722 77758 18734 77810
rect 18786 77758 18798 77810
rect 17054 77746 17106 77758
rect 20750 77746 20802 77758
rect 672 77642 31024 77676
rect 672 77590 4466 77642
rect 4518 77590 4570 77642
rect 4622 77590 4674 77642
rect 4726 77590 24466 77642
rect 24518 77590 24570 77642
rect 24622 77590 24674 77642
rect 24726 77590 31024 77642
rect 672 77556 31024 77590
rect 6626 77422 6638 77474
rect 6690 77422 6702 77474
rect 20178 77422 20190 77474
rect 20242 77422 20254 77474
rect 9886 77362 9938 77374
rect 1026 77310 1038 77362
rect 1090 77310 1102 77362
rect 1698 77310 1710 77362
rect 1762 77310 1774 77362
rect 3378 77310 3390 77362
rect 3442 77310 3454 77362
rect 9202 77310 9214 77362
rect 9266 77310 9278 77362
rect 10882 77310 10894 77362
rect 10946 77310 10958 77362
rect 13458 77310 13470 77362
rect 13522 77310 13534 77362
rect 14802 77310 14814 77362
rect 14866 77310 14878 77362
rect 17378 77310 17390 77362
rect 17442 77310 17454 77362
rect 21186 77310 21198 77362
rect 21250 77310 21262 77362
rect 21634 77310 21646 77362
rect 21698 77310 21710 77362
rect 9886 77298 9938 77310
rect 1374 77250 1426 77262
rect 1374 77186 1426 77198
rect 2046 77250 2098 77262
rect 2046 77186 2098 77198
rect 2382 77250 2434 77262
rect 3838 77250 3890 77262
rect 9550 77250 9602 77262
rect 11566 77250 11618 77262
rect 13806 77250 13858 77262
rect 16046 77250 16098 77262
rect 20638 77250 20690 77262
rect 2706 77198 2718 77250
rect 2770 77198 2782 77250
rect 3154 77198 3166 77250
rect 3218 77198 3230 77250
rect 4386 77198 4398 77250
rect 4450 77198 4462 77250
rect 5394 77198 5406 77250
rect 5458 77198 5470 77250
rect 10322 77198 10334 77250
rect 10386 77198 10398 77250
rect 10770 77198 10782 77250
rect 10834 77198 10846 77250
rect 11890 77198 11902 77250
rect 11954 77198 11966 77250
rect 12898 77198 12910 77250
rect 12962 77198 12974 77250
rect 14354 77198 14366 77250
rect 14418 77198 14430 77250
rect 16818 77198 16830 77250
rect 16882 77198 16894 77250
rect 19954 77198 19966 77250
rect 20018 77198 20030 77250
rect 2382 77186 2434 77198
rect 3838 77186 3890 77198
rect 9550 77186 9602 77198
rect 11566 77186 11618 77198
rect 13806 77186 13858 77198
rect 16046 77186 16098 77198
rect 20638 77186 20690 77198
rect 20974 77138 21026 77150
rect 6178 77086 6190 77138
rect 6242 77086 6254 77138
rect 20974 77074 21026 77086
rect 7758 77026 7810 77038
rect 7758 76962 7810 76974
rect 18510 77026 18562 77038
rect 18510 76962 18562 76974
rect 672 76858 31024 76892
rect 672 76806 3806 76858
rect 3858 76806 3910 76858
rect 3962 76806 4014 76858
rect 4066 76806 23806 76858
rect 23858 76806 23910 76858
rect 23962 76806 24014 76858
rect 24066 76806 31024 76858
rect 672 76772 31024 76806
rect 6638 76578 6690 76590
rect 1922 76526 1934 76578
rect 1986 76526 1998 76578
rect 6638 76514 6690 76526
rect 12910 76578 12962 76590
rect 12910 76514 12962 76526
rect 16494 76578 16546 76590
rect 16494 76514 16546 76526
rect 8094 76466 8146 76478
rect 12126 76466 12178 76478
rect 14590 76466 14642 76478
rect 18174 76466 18226 76478
rect 5058 76414 5070 76466
rect 5122 76414 5134 76466
rect 7074 76414 7086 76466
rect 7138 76414 7150 76466
rect 7410 76414 7422 76466
rect 7474 76414 7486 76466
rect 8866 76414 8878 76466
rect 8930 76414 8942 76466
rect 9762 76414 9774 76466
rect 9826 76414 9838 76466
rect 10434 76414 10446 76466
rect 10498 76414 10510 76466
rect 13234 76414 13246 76466
rect 13298 76414 13310 76466
rect 13682 76414 13694 76466
rect 13746 76414 13758 76466
rect 14914 76414 14926 76466
rect 14978 76414 14990 76466
rect 15922 76414 15934 76466
rect 15986 76414 15998 76466
rect 16930 76414 16942 76466
rect 16994 76414 17006 76466
rect 17266 76414 17278 76466
rect 17330 76414 17342 76466
rect 18610 76414 18622 76466
rect 18674 76414 18686 76466
rect 19506 76414 19518 76466
rect 19570 76414 19582 76466
rect 22306 76414 22318 76466
rect 22370 76414 22382 76466
rect 8094 76402 8146 76414
rect 12126 76402 12178 76414
rect 14590 76402 14642 76414
rect 18174 76402 18226 76414
rect 2370 76302 2382 76354
rect 2434 76302 2446 76354
rect 7634 76302 7646 76354
rect 7698 76302 7710 76354
rect 10882 76302 10894 76354
rect 10946 76302 10958 76354
rect 13906 76302 13918 76354
rect 13970 76302 13982 76354
rect 21858 76302 21870 76354
rect 21922 76302 21934 76354
rect 1374 76242 1426 76254
rect 1026 76190 1038 76242
rect 1090 76190 1102 76242
rect 1374 76178 1426 76190
rect 3502 76242 3554 76254
rect 3502 76178 3554 76190
rect 3950 76242 4002 76254
rect 5966 76242 6018 76254
rect 20750 76242 20802 76254
rect 4274 76190 4286 76242
rect 4338 76190 4350 76242
rect 5282 76190 5294 76242
rect 5346 76190 5358 76242
rect 5618 76190 5630 76242
rect 5682 76190 5694 76242
rect 17490 76190 17502 76242
rect 17554 76190 17566 76242
rect 3950 76178 4002 76190
rect 5966 76178 6018 76190
rect 20750 76178 20802 76190
rect 672 76074 31024 76108
rect 672 76022 4466 76074
rect 4518 76022 4570 76074
rect 4622 76022 4674 76074
rect 4726 76022 24466 76074
rect 24518 76022 24570 76074
rect 24622 76022 24674 76074
rect 24726 76022 31024 76074
rect 672 75988 31024 76022
rect 3154 75854 3166 75906
rect 3218 75854 3230 75906
rect 7074 75854 7086 75906
rect 7138 75854 7150 75906
rect 11666 75854 11678 75906
rect 11730 75854 11742 75906
rect 13010 75854 13022 75906
rect 13074 75854 13086 75906
rect 17490 75854 17502 75906
rect 17554 75854 17566 75906
rect 20066 75854 20078 75906
rect 20130 75854 20142 75906
rect 3614 75794 3666 75806
rect 1026 75742 1038 75794
rect 1090 75742 1102 75794
rect 3614 75730 3666 75742
rect 20414 75794 20466 75806
rect 20414 75730 20466 75742
rect 20750 75794 20802 75806
rect 21746 75742 21758 75794
rect 21810 75742 21822 75794
rect 20750 75730 20802 75742
rect 1374 75682 1426 75694
rect 1374 75618 1426 75630
rect 2158 75682 2210 75694
rect 8206 75682 8258 75694
rect 2594 75630 2606 75682
rect 2658 75630 2670 75682
rect 2930 75630 2942 75682
rect 2994 75630 3006 75682
rect 4162 75630 4174 75682
rect 4226 75630 4238 75682
rect 5170 75630 5182 75682
rect 5234 75630 5246 75682
rect 6626 75630 6638 75682
rect 6690 75630 6702 75682
rect 2158 75618 2210 75630
rect 8206 75618 8258 75630
rect 12014 75682 12066 75694
rect 12014 75618 12066 75630
rect 18622 75682 18674 75694
rect 22430 75682 22482 75694
rect 21074 75630 21086 75682
rect 21138 75630 21150 75682
rect 21522 75630 21534 75682
rect 21586 75630 21598 75682
rect 22978 75630 22990 75682
rect 23042 75630 23054 75682
rect 23762 75630 23774 75682
rect 23826 75630 23838 75682
rect 18622 75618 18674 75630
rect 22430 75618 22482 75630
rect 12562 75518 12574 75570
rect 12626 75518 12638 75570
rect 17042 75518 17054 75570
rect 17106 75518 17118 75570
rect 14142 75458 14194 75470
rect 14142 75394 14194 75406
rect 672 75290 31024 75324
rect 672 75238 3806 75290
rect 3858 75238 3910 75290
rect 3962 75238 4014 75290
rect 4066 75238 23806 75290
rect 23858 75238 23910 75290
rect 23962 75238 24014 75290
rect 24066 75238 31024 75290
rect 672 75204 31024 75238
rect 1810 74958 1822 75010
rect 1874 74958 1886 75010
rect 6066 74958 6078 75010
rect 6130 74958 6142 75010
rect 26898 74958 26910 75010
rect 26962 74958 26974 75010
rect 4398 74898 4450 74910
rect 12126 74898 12178 74910
rect 14254 74898 14306 74910
rect 18398 74898 18450 74910
rect 5394 74846 5406 74898
rect 5458 74846 5470 74898
rect 8306 74846 8318 74898
rect 8370 74846 8382 74898
rect 10546 74846 10558 74898
rect 10610 74846 10622 74898
rect 13122 74846 13134 74898
rect 13186 74846 13198 74898
rect 13570 74846 13582 74898
rect 13634 74846 13646 74898
rect 14914 74846 14926 74898
rect 14978 74846 14990 74898
rect 15810 74846 15822 74898
rect 15874 74846 15886 74898
rect 17042 74846 17054 74898
rect 17106 74846 17118 74898
rect 17602 74846 17614 74898
rect 17666 74846 17678 74898
rect 18834 74846 18846 74898
rect 18898 74846 18910 74898
rect 19730 74846 19742 74898
rect 19794 74846 19806 74898
rect 22866 74846 22878 74898
rect 22930 74846 22942 74898
rect 4398 74834 4450 74846
rect 12126 74834 12178 74846
rect 14254 74834 14306 74846
rect 18398 74834 18450 74846
rect 12798 74786 12850 74798
rect 16718 74786 16770 74798
rect 2258 74734 2270 74786
rect 2322 74734 2334 74786
rect 6514 74734 6526 74786
rect 6578 74734 6590 74786
rect 8082 74734 8094 74786
rect 8146 74734 8158 74786
rect 10994 74734 11006 74786
rect 11058 74734 11070 74786
rect 13794 74734 13806 74786
rect 13858 74734 13870 74786
rect 27682 74734 27694 74786
rect 27746 74734 27758 74786
rect 12798 74722 12850 74734
rect 16718 74722 16770 74734
rect 3390 74674 3442 74686
rect 7646 74674 7698 74686
rect 30270 74674 30322 74686
rect 4050 74622 4062 74674
rect 4114 74622 4126 74674
rect 5170 74622 5182 74674
rect 5234 74622 5246 74674
rect 17714 74622 17726 74674
rect 17778 74622 17790 74674
rect 30594 74622 30606 74674
rect 30658 74622 30670 74674
rect 3390 74610 3442 74622
rect 7646 74610 7698 74622
rect 30270 74610 30322 74622
rect 672 74506 31024 74540
rect 672 74454 4466 74506
rect 4518 74454 4570 74506
rect 4622 74454 4674 74506
rect 4726 74454 24466 74506
rect 24518 74454 24570 74506
rect 24622 74454 24674 74506
rect 24726 74454 31024 74506
rect 672 74420 31024 74454
rect 7534 74338 7586 74350
rect 3938 74286 3950 74338
rect 4002 74286 4014 74338
rect 7534 74274 7586 74286
rect 8206 74338 8258 74350
rect 8206 74274 8258 74286
rect 16046 74338 16098 74350
rect 17054 74338 17106 74350
rect 16706 74286 16718 74338
rect 16770 74286 16782 74338
rect 16046 74274 16098 74286
rect 17054 74274 17106 74286
rect 22990 74338 23042 74350
rect 22990 74274 23042 74286
rect 2942 74226 2994 74238
rect 1026 74174 1038 74226
rect 1090 74174 1102 74226
rect 2146 74174 2158 74226
rect 2210 74174 2222 74226
rect 6514 74174 6526 74226
rect 6578 74174 6590 74226
rect 7186 74174 7198 74226
rect 7250 74174 7262 74226
rect 9426 74174 9438 74226
rect 9490 74174 9502 74226
rect 11778 74174 11790 74226
rect 11842 74174 11854 74226
rect 14802 74174 14814 74226
rect 14866 74174 14878 74226
rect 18610 74174 18622 74226
rect 18674 74174 18686 74226
rect 21746 74174 21758 74226
rect 21810 74174 21822 74226
rect 30594 74174 30606 74226
rect 30658 74174 30670 74226
rect 2942 74162 2994 74174
rect 1374 74114 1426 74126
rect 4622 74114 4674 74126
rect 6862 74114 6914 74126
rect 1922 74062 1934 74114
rect 1986 74062 1998 74114
rect 3266 74062 3278 74114
rect 3330 74062 3342 74114
rect 3826 74062 3838 74114
rect 3890 74062 3902 74114
rect 5058 74062 5070 74114
rect 5122 74062 5134 74114
rect 5954 74062 5966 74114
rect 6018 74062 6030 74114
rect 1374 74050 1426 74062
rect 4622 74050 4674 74062
rect 6862 74050 6914 74062
rect 7982 74114 8034 74126
rect 7982 74050 8034 74062
rect 8318 74114 8370 74126
rect 19294 74114 19346 74126
rect 30270 74114 30322 74126
rect 8978 74062 8990 74114
rect 9042 74062 9054 74114
rect 14466 74062 14478 74114
rect 14530 74062 14542 74114
rect 18050 74062 18062 74114
rect 18114 74062 18126 74114
rect 18386 74062 18398 74114
rect 18450 74062 18462 74114
rect 19730 74062 19742 74114
rect 19794 74062 19806 74114
rect 20626 74062 20638 74114
rect 20690 74062 20702 74114
rect 21410 74062 21422 74114
rect 21474 74062 21486 74114
rect 8318 74050 8370 74062
rect 19294 74050 19346 74062
rect 30270 74050 30322 74062
rect 17614 74002 17666 74014
rect 11442 73950 11454 74002
rect 11506 73950 11518 74002
rect 17614 73938 17666 73950
rect 10670 73890 10722 73902
rect 10670 73826 10722 73838
rect 13022 73890 13074 73902
rect 13022 73826 13074 73838
rect 672 73722 31024 73756
rect 672 73670 3806 73722
rect 3858 73670 3910 73722
rect 3962 73670 4014 73722
rect 4066 73670 23806 73722
rect 23858 73670 23910 73722
rect 23962 73670 24014 73722
rect 24066 73670 31024 73722
rect 672 73636 31024 73670
rect 10558 73554 10610 73566
rect 10558 73490 10610 73502
rect 18398 73554 18450 73566
rect 18398 73490 18450 73502
rect 10222 73442 10274 73454
rect 10222 73378 10274 73390
rect 11342 73442 11394 73454
rect 11342 73378 11394 73390
rect 12798 73442 12850 73454
rect 12798 73378 12850 73390
rect 4174 73330 4226 73342
rect 8542 73330 8594 73342
rect 1810 73278 1822 73330
rect 1874 73278 1886 73330
rect 5842 73278 5854 73330
rect 5906 73278 5918 73330
rect 7186 73278 7198 73330
rect 7250 73278 7262 73330
rect 8082 73278 8094 73330
rect 8146 73278 8158 73330
rect 9314 73278 9326 73330
rect 9378 73278 9390 73330
rect 9762 73278 9774 73330
rect 9826 73278 9838 73330
rect 13122 73278 13134 73330
rect 13186 73278 13198 73330
rect 13682 73278 13694 73330
rect 13746 73278 13758 73330
rect 15026 73278 15038 73330
rect 15090 73278 15102 73330
rect 15810 73278 15822 73330
rect 15874 73278 15886 73330
rect 16818 73278 16830 73330
rect 16882 73278 16894 73330
rect 4174 73266 4226 73278
rect 8542 73266 8594 73278
rect 10782 73218 10834 73230
rect 2258 73166 2270 73218
rect 2322 73166 2334 73218
rect 3826 73166 3838 73218
rect 3890 73166 3902 73218
rect 4946 73166 4958 73218
rect 5010 73166 5022 73218
rect 10782 73154 10834 73166
rect 11230 73218 11282 73230
rect 14254 73218 14306 73230
rect 11890 73166 11902 73218
rect 11954 73166 11966 73218
rect 20626 73166 20638 73218
rect 20690 73166 20702 73218
rect 23314 73166 23326 73218
rect 23378 73166 23390 73218
rect 11230 73154 11282 73166
rect 14254 73154 14306 73166
rect 3390 73106 3442 73118
rect 3390 73042 3442 73054
rect 5294 73106 5346 73118
rect 6638 73106 6690 73118
rect 10670 73106 10722 73118
rect 5618 73054 5630 73106
rect 5682 73054 5694 73106
rect 6290 73054 6302 73106
rect 6354 73054 6366 73106
rect 9202 73054 9214 73106
rect 9266 73054 9278 73106
rect 5294 73042 5346 73054
rect 6638 73042 6690 73054
rect 10670 73042 10722 73054
rect 12238 73106 12290 73118
rect 20974 73106 21026 73118
rect 13794 73054 13806 73106
rect 13858 73054 13870 73106
rect 17266 73054 17278 73106
rect 17330 73054 17342 73106
rect 12238 73042 12290 73054
rect 20974 73042 21026 73054
rect 22990 73106 23042 73118
rect 22990 73042 23042 73054
rect 672 72938 31024 72972
rect 672 72886 4466 72938
rect 4518 72886 4570 72938
rect 4622 72886 4674 72938
rect 4726 72886 24466 72938
rect 24518 72886 24570 72938
rect 24622 72886 24674 72938
rect 24726 72886 31024 72938
rect 672 72852 31024 72886
rect 9438 72770 9490 72782
rect 12798 72770 12850 72782
rect 17726 72770 17778 72782
rect 3042 72718 3054 72770
rect 3106 72718 3118 72770
rect 10322 72718 10334 72770
rect 10386 72718 10398 72770
rect 17378 72718 17390 72770
rect 17442 72718 17454 72770
rect 21522 72718 21534 72770
rect 21586 72718 21598 72770
rect 9438 72706 9490 72718
rect 12798 72706 12850 72718
rect 17726 72706 17778 72718
rect 3502 72658 3554 72670
rect 9886 72658 9938 72670
rect 1026 72606 1038 72658
rect 1090 72606 1102 72658
rect 6290 72606 6302 72658
rect 6354 72606 6366 72658
rect 7858 72606 7870 72658
rect 7922 72606 7934 72658
rect 11666 72606 11678 72658
rect 11730 72606 11742 72658
rect 13906 72606 13918 72658
rect 13970 72606 13982 72658
rect 18834 72606 18846 72658
rect 18898 72606 18910 72658
rect 30594 72606 30606 72658
rect 30658 72606 30670 72658
rect 3502 72594 3554 72606
rect 9886 72594 9938 72606
rect 1374 72546 1426 72558
rect 8206 72546 8258 72558
rect 10334 72546 10386 72558
rect 20078 72546 20130 72558
rect 22206 72546 22258 72558
rect 30270 72546 30322 72558
rect 2370 72494 2382 72546
rect 2434 72494 2446 72546
rect 2930 72494 2942 72546
rect 2994 72494 3006 72546
rect 4274 72494 4286 72546
rect 4338 72494 4350 72546
rect 5058 72494 5070 72546
rect 5122 72494 5134 72546
rect 5842 72494 5854 72546
rect 5906 72494 5918 72546
rect 9538 72494 9550 72546
rect 9602 72494 9614 72546
rect 10098 72494 10110 72546
rect 10162 72494 10174 72546
rect 10658 72494 10670 72546
rect 10722 72494 10734 72546
rect 11218 72494 11230 72546
rect 11282 72494 11294 72546
rect 13458 72494 13470 72546
rect 13522 72494 13534 72546
rect 18386 72494 18398 72546
rect 18450 72494 18462 72546
rect 20850 72494 20862 72546
rect 20914 72494 20926 72546
rect 21298 72494 21310 72546
rect 21362 72494 21374 72546
rect 22642 72494 22654 72546
rect 22706 72494 22718 72546
rect 23650 72494 23662 72546
rect 23714 72494 23726 72546
rect 1374 72482 1426 72494
rect 8206 72482 8258 72494
rect 10334 72482 10386 72494
rect 20078 72482 20130 72494
rect 22206 72482 22258 72494
rect 30270 72482 30322 72494
rect 2046 72434 2098 72446
rect 2046 72370 2098 72382
rect 9326 72434 9378 72446
rect 9326 72370 9378 72382
rect 20526 72434 20578 72446
rect 20526 72370 20578 72382
rect 7422 72322 7474 72334
rect 7422 72258 7474 72270
rect 9102 72322 9154 72334
rect 9102 72258 9154 72270
rect 15038 72322 15090 72334
rect 15038 72258 15090 72270
rect 672 72154 31024 72188
rect 672 72102 3806 72154
rect 3858 72102 3910 72154
rect 3962 72102 4014 72154
rect 4066 72102 23806 72154
rect 23858 72102 23910 72154
rect 23962 72102 24014 72154
rect 24066 72102 31024 72154
rect 672 72068 31024 72102
rect 9774 71986 9826 71998
rect 9774 71922 9826 71934
rect 19966 71986 20018 71998
rect 19966 71922 20018 71934
rect 22654 71986 22706 71998
rect 22654 71922 22706 71934
rect 6078 71874 6130 71886
rect 14590 71874 14642 71886
rect 11330 71822 11342 71874
rect 11394 71822 11406 71874
rect 6078 71810 6130 71822
rect 14590 71810 14642 71822
rect 4286 71762 4338 71774
rect 1250 71710 1262 71762
rect 1314 71710 1326 71762
rect 2706 71710 2718 71762
rect 2770 71710 2782 71762
rect 6402 71710 6414 71762
rect 6466 71710 6478 71762
rect 6962 71710 6974 71762
rect 7026 71710 7038 71762
rect 7634 71710 7646 71762
rect 7698 71710 7710 71762
rect 8082 71710 8094 71762
rect 8146 71710 8158 71762
rect 9202 71710 9214 71762
rect 9266 71710 9278 71762
rect 15026 71710 15038 71762
rect 15090 71710 15102 71762
rect 15474 71710 15486 71762
rect 15538 71710 15550 71762
rect 16706 71710 16718 71762
rect 16770 71710 16782 71762
rect 17602 71710 17614 71762
rect 17666 71710 17678 71762
rect 18274 71710 18286 71762
rect 18338 71710 18350 71762
rect 21074 71710 21086 71762
rect 21138 71710 21150 71762
rect 23202 71710 23214 71762
rect 23266 71710 23278 71762
rect 30370 71710 30382 71762
rect 30434 71710 30446 71762
rect 4286 71698 4338 71710
rect 16046 71650 16098 71662
rect 3154 71598 3166 71650
rect 3218 71598 3230 71650
rect 10882 71598 10894 71650
rect 10946 71598 10958 71650
rect 13906 71598 13918 71650
rect 13970 71598 13982 71650
rect 21410 71598 21422 71650
rect 21474 71598 21486 71650
rect 23426 71598 23438 71650
rect 23490 71598 23502 71650
rect 16046 71586 16098 71598
rect 2046 71538 2098 71550
rect 5294 71538 5346 71550
rect 14254 71538 14306 71550
rect 1026 71486 1038 71538
rect 1090 71486 1102 71538
rect 1698 71486 1710 71538
rect 1762 71486 1774 71538
rect 4946 71486 4958 71538
rect 5010 71486 5022 71538
rect 7074 71486 7086 71538
rect 7138 71486 7150 71538
rect 15586 71486 15598 71538
rect 15650 71486 15662 71538
rect 18834 71486 18846 71538
rect 18898 71486 18910 71538
rect 30594 71486 30606 71538
rect 30658 71486 30670 71538
rect 2046 71474 2098 71486
rect 5294 71474 5346 71486
rect 14254 71474 14306 71486
rect 672 71370 31024 71404
rect 672 71318 4466 71370
rect 4518 71318 4570 71370
rect 4622 71318 4674 71370
rect 4726 71318 24466 71370
rect 24518 71318 24570 71370
rect 24622 71318 24674 71370
rect 24726 71318 31024 71370
rect 672 71284 31024 71318
rect 16046 71202 16098 71214
rect 6066 71150 6078 71202
rect 6130 71150 6142 71202
rect 29810 71150 29822 71202
rect 29874 71150 29886 71202
rect 16046 71138 16098 71150
rect 2482 71038 2494 71090
rect 2546 71038 2558 71090
rect 8866 71038 8878 71090
rect 8930 71038 8942 71090
rect 10994 71038 11006 71090
rect 11058 71038 11070 71090
rect 14802 71038 14814 71090
rect 14866 71038 14878 71090
rect 21522 71038 21534 71090
rect 21586 71038 21598 71090
rect 30594 71038 30606 71090
rect 30658 71038 30670 71090
rect 3166 70978 3218 70990
rect 29486 70978 29538 70990
rect 1810 70926 1822 70978
rect 1874 70926 1886 70978
rect 2258 70926 2270 70978
rect 2322 70926 2334 70978
rect 3490 70926 3502 70978
rect 3554 70926 3566 70978
rect 4498 70926 4510 70978
rect 4562 70926 4574 70978
rect 5506 70926 5518 70978
rect 5570 70926 5582 70978
rect 5842 70926 5854 70978
rect 5906 70926 5918 70978
rect 6626 70926 6638 70978
rect 6690 70926 6702 70978
rect 7298 70926 7310 70978
rect 7362 70926 7374 70978
rect 8082 70926 8094 70978
rect 8146 70926 8158 70978
rect 9090 70926 9102 70978
rect 9154 70926 9166 70978
rect 14354 70926 14366 70978
rect 14418 70926 14430 70978
rect 21074 70926 21086 70978
rect 21138 70926 21150 70978
rect 3166 70914 3218 70926
rect 29486 70914 29538 70926
rect 30270 70978 30322 70990
rect 30270 70914 30322 70926
rect 1486 70866 1538 70878
rect 1486 70802 1538 70814
rect 5070 70866 5122 70878
rect 18958 70866 19010 70878
rect 11330 70814 11342 70866
rect 11394 70814 11406 70866
rect 5070 70802 5122 70814
rect 18958 70802 19010 70814
rect 9774 70754 9826 70766
rect 9774 70690 9826 70702
rect 22766 70754 22818 70766
rect 22766 70690 22818 70702
rect 672 70586 31024 70620
rect 672 70534 3806 70586
rect 3858 70534 3910 70586
rect 3962 70534 4014 70586
rect 4066 70534 23806 70586
rect 23858 70534 23910 70586
rect 23962 70534 24014 70586
rect 24066 70534 31024 70586
rect 672 70500 31024 70534
rect 5630 70418 5682 70430
rect 5630 70354 5682 70366
rect 8990 70306 9042 70318
rect 7186 70254 7198 70306
rect 7250 70254 7262 70306
rect 15362 70254 15374 70306
rect 15426 70254 15438 70306
rect 8990 70242 9042 70254
rect 10446 70194 10498 70206
rect 1250 70142 1262 70194
rect 1314 70142 1326 70194
rect 3490 70142 3502 70194
rect 3554 70142 3566 70194
rect 4050 70142 4062 70194
rect 4114 70142 4126 70194
rect 7298 70142 7310 70194
rect 7362 70142 7374 70194
rect 9314 70142 9326 70194
rect 9378 70142 9390 70194
rect 9874 70142 9886 70194
rect 9938 70142 9950 70194
rect 11218 70142 11230 70194
rect 11282 70142 11294 70194
rect 12002 70142 12014 70194
rect 12066 70142 12078 70194
rect 17714 70142 17726 70194
rect 17778 70142 17790 70194
rect 21186 70142 21198 70194
rect 21250 70142 21262 70194
rect 10446 70130 10498 70142
rect 8094 70082 8146 70094
rect 3266 70030 3278 70082
rect 3330 70030 3342 70082
rect 4274 70030 4286 70082
rect 4338 70030 4350 70082
rect 7746 70030 7758 70082
rect 7810 70030 7822 70082
rect 14466 70030 14478 70082
rect 14530 70030 14542 70082
rect 18162 70030 18174 70082
rect 18226 70030 18238 70082
rect 19730 70030 19742 70082
rect 19794 70030 19806 70082
rect 8094 70018 8146 70030
rect 2830 69970 2882 69982
rect 14814 69970 14866 69982
rect 16942 69970 16994 69982
rect 1698 69918 1710 69970
rect 1762 69918 1774 69970
rect 6738 69918 6750 69970
rect 6802 69918 6814 69970
rect 9986 69918 9998 69970
rect 10050 69918 10062 69970
rect 15810 69918 15822 69970
rect 15874 69918 15886 69970
rect 2830 69906 2882 69918
rect 14814 69906 14866 69918
rect 16942 69906 16994 69918
rect 19294 69970 19346 69982
rect 19294 69906 19346 69918
rect 20078 69970 20130 69982
rect 22878 69970 22930 69982
rect 21746 69918 21758 69970
rect 21810 69918 21822 69970
rect 20078 69906 20130 69918
rect 22878 69906 22930 69918
rect 672 69802 31024 69836
rect 672 69750 4466 69802
rect 4518 69750 4570 69802
rect 4622 69750 4674 69802
rect 4726 69750 24466 69802
rect 24518 69750 24570 69802
rect 24622 69750 24674 69802
rect 24726 69750 31024 69802
rect 672 69716 31024 69750
rect 8318 69634 8370 69646
rect 8318 69570 8370 69582
rect 8990 69634 9042 69646
rect 10098 69582 10110 69634
rect 10162 69582 10174 69634
rect 11890 69582 11902 69634
rect 11954 69582 11966 69634
rect 22418 69582 22430 69634
rect 22482 69582 22494 69634
rect 8990 69570 9042 69582
rect 3390 69522 3442 69534
rect 1026 69470 1038 69522
rect 1090 69470 1102 69522
rect 2930 69470 2942 69522
rect 2994 69470 3006 69522
rect 6066 69470 6078 69522
rect 6130 69470 6142 69522
rect 7970 69470 7982 69522
rect 8034 69470 8046 69522
rect 14578 69470 14590 69522
rect 14642 69470 14654 69522
rect 17266 69470 17278 69522
rect 17330 69470 17342 69522
rect 19506 69470 19518 69522
rect 19570 69470 19582 69522
rect 30594 69470 30606 69522
rect 30658 69470 30670 69522
rect 3390 69458 3442 69470
rect 1374 69410 1426 69422
rect 12238 69410 12290 69422
rect 30270 69410 30322 69422
rect 2370 69358 2382 69410
rect 2434 69358 2446 69410
rect 2818 69358 2830 69410
rect 2882 69358 2894 69410
rect 3938 69358 3950 69410
rect 4002 69358 4014 69410
rect 4946 69358 4958 69410
rect 5010 69358 5022 69410
rect 16930 69358 16942 69410
rect 16994 69358 17006 69410
rect 19170 69358 19182 69410
rect 19234 69358 19246 69410
rect 22866 69358 22878 69410
rect 22930 69358 22942 69410
rect 23762 69358 23774 69410
rect 23826 69358 23838 69410
rect 1374 69346 1426 69358
rect 12238 69346 12290 69358
rect 30270 69346 30322 69358
rect 1934 69298 1986 69310
rect 5730 69246 5742 69298
rect 5794 69246 5806 69298
rect 10546 69246 10558 69298
rect 10610 69246 10622 69298
rect 14130 69246 14142 69298
rect 14194 69246 14206 69298
rect 1934 69234 1986 69246
rect 7310 69186 7362 69198
rect 7310 69122 7362 69134
rect 15710 69186 15762 69198
rect 15710 69122 15762 69134
rect 18510 69186 18562 69198
rect 18510 69122 18562 69134
rect 20750 69186 20802 69198
rect 20750 69122 20802 69134
rect 21310 69186 21362 69198
rect 21310 69122 21362 69134
rect 23438 69186 23490 69198
rect 23438 69122 23490 69134
rect 23774 69186 23826 69198
rect 23774 69122 23826 69134
rect 672 69018 31024 69052
rect 672 68966 3806 69018
rect 3858 68966 3910 69018
rect 3962 68966 4014 69018
rect 4066 68966 23806 69018
rect 23858 68966 23910 69018
rect 23962 68966 24014 69018
rect 24066 68966 31024 69018
rect 672 68932 31024 68966
rect 19966 68738 20018 68750
rect 5170 68686 5182 68738
rect 5234 68686 5246 68738
rect 10546 68686 10558 68738
rect 10610 68686 10622 68738
rect 14466 68686 14478 68738
rect 14530 68686 14542 68738
rect 19966 68674 20018 68686
rect 20638 68738 20690 68750
rect 20638 68674 20690 68686
rect 24334 68738 24386 68750
rect 24334 68674 24386 68686
rect 9774 68626 9826 68638
rect 1922 68574 1934 68626
rect 1986 68574 1998 68626
rect 4162 68574 4174 68626
rect 4226 68574 4238 68626
rect 7298 68574 7310 68626
rect 7362 68574 7374 68626
rect 9774 68562 9826 68574
rect 15262 68626 15314 68638
rect 19294 68626 19346 68638
rect 15698 68574 15710 68626
rect 15762 68574 15774 68626
rect 16146 68574 16158 68626
rect 16210 68574 16222 68626
rect 16818 68574 16830 68626
rect 16882 68574 16894 68626
rect 17266 68574 17278 68626
rect 17330 68574 17342 68626
rect 18386 68574 18398 68626
rect 18450 68574 18462 68626
rect 15262 68562 15314 68574
rect 19294 68562 19346 68574
rect 19630 68626 19682 68638
rect 19630 68562 19682 68574
rect 19742 68626 19794 68638
rect 19742 68562 19794 68574
rect 20078 68626 20130 68638
rect 22318 68626 22370 68638
rect 24222 68626 24274 68638
rect 21074 68574 21086 68626
rect 21138 68574 21150 68626
rect 21410 68574 21422 68626
rect 21474 68574 21486 68626
rect 22866 68574 22878 68626
rect 22930 68574 22942 68626
rect 23650 68574 23662 68626
rect 23714 68574 23726 68626
rect 20078 68562 20130 68574
rect 22318 68562 22370 68574
rect 24222 68562 24274 68574
rect 24670 68626 24722 68638
rect 24770 68574 24782 68626
rect 24834 68574 24846 68626
rect 24670 68562 24722 68574
rect 18958 68514 19010 68526
rect 2258 68462 2270 68514
rect 2322 68462 2334 68514
rect 5618 68462 5630 68514
rect 5682 68462 5694 68514
rect 7746 68462 7758 68514
rect 7810 68462 7822 68514
rect 10882 68462 10894 68514
rect 10946 68462 10958 68514
rect 14130 68462 14142 68514
rect 14194 68462 14206 68514
rect 16258 68462 16270 68514
rect 16322 68462 16334 68514
rect 18958 68450 19010 68462
rect 19070 68514 19122 68526
rect 21634 68462 21646 68514
rect 21698 68462 21710 68514
rect 24434 68462 24446 68514
rect 24498 68462 24510 68514
rect 29810 68462 29822 68514
rect 29874 68462 29886 68514
rect 19070 68450 19122 68462
rect 1374 68402 1426 68414
rect 1026 68350 1038 68402
rect 1090 68350 1102 68402
rect 1374 68338 1426 68350
rect 3502 68402 3554 68414
rect 6750 68402 6802 68414
rect 3938 68350 3950 68402
rect 4002 68350 4014 68402
rect 3502 68338 3554 68350
rect 6750 68338 6802 68350
rect 8990 68402 9042 68414
rect 12126 68402 12178 68414
rect 9426 68350 9438 68402
rect 9490 68350 9502 68402
rect 8990 68338 9042 68350
rect 12126 68338 12178 68350
rect 12910 68402 12962 68414
rect 12910 68338 12962 68350
rect 29486 68402 29538 68414
rect 29486 68338 29538 68350
rect 30270 68402 30322 68414
rect 30594 68350 30606 68402
rect 30658 68350 30670 68402
rect 30270 68338 30322 68350
rect 672 68234 31024 68268
rect 672 68182 4466 68234
rect 4518 68182 4570 68234
rect 4622 68182 4674 68234
rect 4726 68182 24466 68234
rect 24518 68182 24570 68234
rect 24622 68182 24674 68234
rect 24726 68182 31024 68234
rect 672 68148 31024 68182
rect 1810 68014 1822 68066
rect 1874 68014 1886 68066
rect 5954 68014 5966 68066
rect 6018 68014 6030 68066
rect 9986 68014 9998 68066
rect 10050 68014 10062 68066
rect 13122 68014 13134 68066
rect 13186 68014 13198 68066
rect 15810 68014 15822 68066
rect 15874 68014 15886 68066
rect 21410 68014 21422 68066
rect 21474 68014 21486 68066
rect 29810 68014 29822 68066
rect 29874 68014 29886 68066
rect 4958 67954 5010 67966
rect 1026 67902 1038 67954
rect 1090 67902 1102 67954
rect 3378 67902 3390 67954
rect 3442 67902 3454 67954
rect 4958 67890 5010 67902
rect 12126 67954 12178 67966
rect 12126 67890 12178 67902
rect 13582 67954 13634 67966
rect 13582 67890 13634 67902
rect 16158 67954 16210 67966
rect 16158 67890 16210 67902
rect 16830 67954 16882 67966
rect 21870 67954 21922 67966
rect 17826 67902 17838 67954
rect 17890 67902 17902 67954
rect 16830 67890 16882 67902
rect 21870 67890 21922 67902
rect 1374 67842 1426 67854
rect 1374 67778 1426 67790
rect 2158 67842 2210 67854
rect 2158 67778 2210 67790
rect 4510 67842 4562 67854
rect 6638 67842 6690 67854
rect 5282 67790 5294 67842
rect 5346 67790 5358 67842
rect 5842 67790 5854 67842
rect 5906 67790 5918 67842
rect 6962 67790 6974 67842
rect 7026 67790 7038 67842
rect 7186 67790 7198 67842
rect 7250 67790 7262 67842
rect 8082 67790 8094 67842
rect 8146 67790 8158 67842
rect 12450 67790 12462 67842
rect 12514 67790 12526 67842
rect 12898 67790 12910 67842
rect 12962 67790 12974 67842
rect 14130 67790 14142 67842
rect 14194 67790 14206 67842
rect 15250 67790 15262 67842
rect 15314 67790 15326 67842
rect 17266 67790 17278 67842
rect 17330 67790 17342 67842
rect 17602 67790 17614 67842
rect 17666 67790 17678 67842
rect 18386 67790 18398 67842
rect 18450 67790 18462 67842
rect 18834 67790 18846 67842
rect 18898 67790 18910 67842
rect 19954 67790 19966 67842
rect 20018 67790 20030 67842
rect 20738 67790 20750 67842
rect 20802 67790 20814 67842
rect 21186 67790 21198 67842
rect 21250 67790 21262 67842
rect 22418 67790 22430 67842
rect 22482 67790 22494 67842
rect 23426 67790 23438 67842
rect 23490 67790 23502 67842
rect 29586 67790 29598 67842
rect 29650 67790 29662 67842
rect 4510 67778 4562 67790
rect 6638 67778 6690 67790
rect 20414 67730 20466 67742
rect 2930 67678 2942 67730
rect 2994 67678 3006 67730
rect 9538 67678 9550 67730
rect 9602 67678 9614 67730
rect 20414 67666 20466 67678
rect 11118 67618 11170 67630
rect 11118 67554 11170 67566
rect 672 67450 31024 67484
rect 672 67398 3806 67450
rect 3858 67398 3910 67450
rect 3962 67398 4014 67450
rect 4066 67398 23806 67450
rect 23858 67398 23910 67450
rect 23962 67398 24014 67450
rect 24066 67398 31024 67450
rect 672 67364 31024 67398
rect 14142 67170 14194 67182
rect 22654 67170 22706 67182
rect 2706 67118 2718 67170
rect 2770 67118 2782 67170
rect 6962 67118 6974 67170
rect 7026 67118 7038 67170
rect 19394 67118 19406 67170
rect 19458 67118 19470 67170
rect 21074 67118 21086 67170
rect 21138 67118 21150 67170
rect 14142 67106 14194 67118
rect 22654 67106 22706 67118
rect 23102 67170 23154 67182
rect 23102 67106 23154 67118
rect 23214 67170 23266 67182
rect 23214 67106 23266 67118
rect 15822 67058 15874 67070
rect 9650 67006 9662 67058
rect 9714 67006 9726 67058
rect 14578 67006 14590 67058
rect 14642 67006 14654 67058
rect 14914 67006 14926 67058
rect 14978 67006 14990 67058
rect 16146 67006 16158 67058
rect 16210 67006 16222 67058
rect 17154 67006 17166 67058
rect 17218 67006 17230 67058
rect 30370 67006 30382 67058
rect 30434 67006 30446 67058
rect 15822 66994 15874 67006
rect 1474 66894 1486 66946
rect 1538 66894 1550 66946
rect 1810 66894 1822 66946
rect 1874 66894 1886 66946
rect 3042 66894 3054 66946
rect 3106 66894 3118 66946
rect 7298 66894 7310 66946
rect 7362 66894 7374 66946
rect 9986 66894 9998 66946
rect 10050 66894 10062 66946
rect 19058 66894 19070 66946
rect 19122 66894 19134 66946
rect 21410 66894 21422 66946
rect 21474 66894 21486 66946
rect 1150 66834 1202 66846
rect 1150 66770 1202 66782
rect 2158 66834 2210 66846
rect 2158 66770 2210 66782
rect 4286 66834 4338 66846
rect 4286 66770 4338 66782
rect 8542 66834 8594 66846
rect 8542 66770 8594 66782
rect 11230 66834 11282 66846
rect 13806 66834 13858 66846
rect 17838 66834 17890 66846
rect 13458 66782 13470 66834
rect 13522 66782 13534 66834
rect 15138 66782 15150 66834
rect 15202 66782 15214 66834
rect 30594 66782 30606 66834
rect 30658 66782 30670 66834
rect 11230 66770 11282 66782
rect 13806 66770 13858 66782
rect 17838 66770 17890 66782
rect 672 66666 31024 66700
rect 672 66614 4466 66666
rect 4518 66614 4570 66666
rect 4622 66614 4674 66666
rect 4726 66614 24466 66666
rect 24518 66614 24570 66666
rect 24622 66614 24674 66666
rect 24726 66614 31024 66666
rect 672 66580 31024 66614
rect 3278 66498 3330 66510
rect 15822 66498 15874 66510
rect 4274 66446 4286 66498
rect 4338 66446 4350 66498
rect 6066 66446 6078 66498
rect 6130 66446 6142 66498
rect 14690 66446 14702 66498
rect 14754 66446 14766 66498
rect 19170 66446 19182 66498
rect 19234 66446 19246 66498
rect 3278 66434 3330 66446
rect 15822 66434 15874 66446
rect 18174 66386 18226 66398
rect 1586 66334 1598 66386
rect 1650 66334 1662 66386
rect 3602 66334 3614 66386
rect 3666 66334 3678 66386
rect 10322 66334 10334 66386
rect 10386 66334 10398 66386
rect 30594 66334 30606 66386
rect 30658 66334 30670 66386
rect 18174 66322 18226 66334
rect 3950 66274 4002 66286
rect 11006 66274 11058 66286
rect 19854 66274 19906 66286
rect 30270 66274 30322 66286
rect 1250 66222 1262 66274
rect 1314 66222 1326 66274
rect 5394 66222 5406 66274
rect 5458 66222 5470 66274
rect 5842 66222 5854 66274
rect 5906 66222 5918 66274
rect 6626 66222 6638 66274
rect 6690 66222 6702 66274
rect 7298 66222 7310 66274
rect 7362 66222 7374 66274
rect 8082 66222 8094 66274
rect 8146 66222 8158 66274
rect 9650 66222 9662 66274
rect 9714 66222 9726 66274
rect 10098 66222 10110 66274
rect 10162 66222 10174 66274
rect 11330 66222 11342 66274
rect 11394 66222 11406 66274
rect 12338 66222 12350 66274
rect 12402 66222 12414 66274
rect 14242 66222 14254 66274
rect 14306 66222 14318 66274
rect 18498 66222 18510 66274
rect 18562 66222 18574 66274
rect 18946 66222 18958 66274
rect 19010 66222 19022 66274
rect 20178 66222 20190 66274
rect 20242 66222 20254 66274
rect 21186 66222 21198 66274
rect 21250 66222 21262 66274
rect 3950 66210 4002 66222
rect 11006 66210 11058 66222
rect 19854 66210 19906 66222
rect 30270 66210 30322 66222
rect 5070 66162 5122 66174
rect 5070 66098 5122 66110
rect 9326 66162 9378 66174
rect 9326 66098 9378 66110
rect 2830 66050 2882 66062
rect 2830 65986 2882 65998
rect 672 65882 31024 65916
rect 672 65830 3806 65882
rect 3858 65830 3910 65882
rect 3962 65830 4014 65882
rect 4066 65830 23806 65882
rect 23858 65830 23910 65882
rect 23962 65830 24014 65882
rect 24066 65830 31024 65882
rect 672 65796 31024 65830
rect 14590 65714 14642 65726
rect 14590 65650 14642 65662
rect 19854 65714 19906 65726
rect 19854 65650 19906 65662
rect 1922 65550 1934 65602
rect 1986 65550 1998 65602
rect 5842 65550 5854 65602
rect 5906 65550 5918 65602
rect 13010 65550 13022 65602
rect 13074 65550 13086 65602
rect 15810 65550 15822 65602
rect 15874 65550 15886 65602
rect 18274 65550 18286 65602
rect 18338 65550 18350 65602
rect 4398 65490 4450 65502
rect 10670 65490 10722 65502
rect 17390 65490 17442 65502
rect 1250 65438 1262 65490
rect 1314 65438 1326 65490
rect 9314 65438 9326 65490
rect 9378 65438 9390 65490
rect 9874 65438 9886 65490
rect 9938 65438 9950 65490
rect 10994 65438 11006 65490
rect 11058 65438 11070 65490
rect 11218 65438 11230 65490
rect 11282 65438 11294 65490
rect 12114 65438 12126 65490
rect 12178 65438 12190 65490
rect 4398 65426 4450 65438
rect 10670 65426 10722 65438
rect 17390 65426 17442 65438
rect 8990 65378 9042 65390
rect 2370 65326 2382 65378
rect 2434 65326 2446 65378
rect 13346 65326 13358 65378
rect 13410 65326 13422 65378
rect 16258 65326 16270 65378
rect 16322 65326 16334 65378
rect 20962 65326 20974 65378
rect 21026 65326 21038 65378
rect 8990 65314 9042 65326
rect 3502 65266 3554 65278
rect 5294 65266 5346 65278
rect 7422 65266 7474 65278
rect 20638 65266 20690 65278
rect 1026 65214 1038 65266
rect 1090 65214 1102 65266
rect 4050 65214 4062 65266
rect 4114 65214 4126 65266
rect 4946 65214 4958 65266
rect 5010 65214 5022 65266
rect 6290 65214 6302 65266
rect 6354 65214 6366 65266
rect 9986 65214 9998 65266
rect 10050 65214 10062 65266
rect 18722 65214 18734 65266
rect 18786 65214 18798 65266
rect 3502 65202 3554 65214
rect 5294 65202 5346 65214
rect 7422 65202 7474 65214
rect 20638 65202 20690 65214
rect 672 65098 31024 65132
rect 672 65046 4466 65098
rect 4518 65046 4570 65098
rect 4622 65046 4674 65098
rect 4726 65046 24466 65098
rect 24518 65046 24570 65098
rect 24622 65046 24674 65098
rect 24726 65046 31024 65098
rect 672 65012 31024 65046
rect 5966 64930 6018 64942
rect 3042 64878 3054 64930
rect 3106 64878 3118 64930
rect 13570 64878 13582 64930
rect 13634 64878 13646 64930
rect 5966 64866 6018 64878
rect 8990 64818 9042 64830
rect 1698 64766 1710 64818
rect 1762 64766 1774 64818
rect 5618 64766 5630 64818
rect 5682 64766 5694 64818
rect 6962 64766 6974 64818
rect 7026 64766 7038 64818
rect 9986 64766 9998 64818
rect 10050 64766 10062 64818
rect 19058 64766 19070 64818
rect 19122 64766 19134 64818
rect 20066 64766 20078 64818
rect 20130 64766 20142 64818
rect 30594 64766 30606 64818
rect 30658 64766 30670 64818
rect 8990 64754 9042 64766
rect 1374 64706 1426 64718
rect 8206 64706 8258 64718
rect 10446 64706 10498 64718
rect 30270 64706 30322 64718
rect 2370 64654 2382 64706
rect 2434 64654 2446 64706
rect 2818 64654 2830 64706
rect 2882 64654 2894 64706
rect 3602 64654 3614 64706
rect 3666 64654 3678 64706
rect 4274 64654 4286 64706
rect 4338 64654 4350 64706
rect 5058 64654 5070 64706
rect 5122 64654 5134 64706
rect 6514 64654 6526 64706
rect 6578 64654 6590 64706
rect 9314 64654 9326 64706
rect 9378 64654 9390 64706
rect 9874 64654 9886 64706
rect 9938 64654 9950 64706
rect 10994 64654 11006 64706
rect 11058 64654 11070 64706
rect 12114 64654 12126 64706
rect 12178 64654 12190 64706
rect 13122 64654 13134 64706
rect 13186 64654 13198 64706
rect 18834 64654 18846 64706
rect 18898 64654 18910 64706
rect 19618 64654 19630 64706
rect 19682 64654 19694 64706
rect 1374 64642 1426 64654
rect 8206 64642 8258 64654
rect 10446 64642 10498 64654
rect 30270 64642 30322 64654
rect 2046 64594 2098 64606
rect 2046 64530 2098 64542
rect 14702 64482 14754 64494
rect 14702 64418 14754 64430
rect 21310 64482 21362 64494
rect 21310 64418 21362 64430
rect 672 64314 31024 64348
rect 672 64262 3806 64314
rect 3858 64262 3910 64314
rect 3962 64262 4014 64314
rect 4066 64262 23806 64314
rect 23858 64262 23910 64314
rect 23962 64262 24014 64314
rect 24066 64262 31024 64314
rect 672 64228 31024 64262
rect 8206 64146 8258 64158
rect 8206 64082 8258 64094
rect 10782 64034 10834 64046
rect 8866 63982 8878 64034
rect 8930 63982 8942 64034
rect 14242 63982 14254 64034
rect 14306 63982 14318 64034
rect 20962 63982 20974 64034
rect 21026 63982 21038 64034
rect 10782 63970 10834 63982
rect 3502 63922 3554 63934
rect 1250 63870 1262 63922
rect 1314 63870 1326 63922
rect 1810 63870 1822 63922
rect 1874 63870 1886 63922
rect 4162 63870 4174 63922
rect 4226 63870 4238 63922
rect 5170 63870 5182 63922
rect 5234 63870 5246 63922
rect 6514 63870 6526 63922
rect 6578 63870 6590 63922
rect 18162 63870 18174 63922
rect 18226 63870 18238 63922
rect 3502 63858 3554 63870
rect 2370 63758 2382 63810
rect 2434 63758 2446 63810
rect 4946 63758 4958 63810
rect 5010 63758 5022 63810
rect 9314 63758 9326 63810
rect 9378 63758 9390 63810
rect 14690 63758 14702 63810
rect 14754 63758 14766 63810
rect 17378 63758 17390 63810
rect 17442 63758 17454 63810
rect 18722 63758 18734 63810
rect 18786 63758 18798 63810
rect 21298 63758 21310 63810
rect 21362 63758 21374 63810
rect 29810 63758 29822 63810
rect 29874 63758 29886 63810
rect 10446 63698 10498 63710
rect 1026 63646 1038 63698
rect 1090 63646 1102 63698
rect 3938 63646 3950 63698
rect 4002 63646 4014 63698
rect 7074 63646 7086 63698
rect 7138 63646 7150 63698
rect 10446 63634 10498 63646
rect 15822 63698 15874 63710
rect 15822 63634 15874 63646
rect 17726 63698 17778 63710
rect 17726 63634 17778 63646
rect 19854 63698 19906 63710
rect 19854 63634 19906 63646
rect 22542 63698 22594 63710
rect 22542 63634 22594 63646
rect 29486 63698 29538 63710
rect 29486 63634 29538 63646
rect 30270 63698 30322 63710
rect 30594 63646 30606 63698
rect 30658 63646 30670 63698
rect 30270 63634 30322 63646
rect 672 63530 31024 63564
rect 672 63478 4466 63530
rect 4518 63478 4570 63530
rect 4622 63478 4674 63530
rect 4726 63478 24466 63530
rect 24518 63478 24570 63530
rect 24622 63478 24674 63530
rect 24726 63478 31024 63530
rect 672 63444 31024 63478
rect 8318 63362 8370 63374
rect 9214 63362 9266 63374
rect 15150 63362 15202 63374
rect 1250 63310 1262 63362
rect 1314 63310 1326 63362
rect 2930 63310 2942 63362
rect 2994 63310 3006 63362
rect 6290 63310 6302 63362
rect 6354 63310 6366 63362
rect 7970 63310 7982 63362
rect 8034 63310 8046 63362
rect 8866 63310 8878 63362
rect 8930 63310 8942 63362
rect 11890 63310 11902 63362
rect 11954 63310 11966 63362
rect 17490 63310 17502 63362
rect 17554 63310 17566 63362
rect 20066 63310 20078 63362
rect 20130 63310 20142 63362
rect 29810 63310 29822 63362
rect 29874 63310 29886 63362
rect 8318 63298 8370 63310
rect 9214 63298 9266 63310
rect 15150 63298 15202 63310
rect 3390 63250 3442 63262
rect 3390 63186 3442 63198
rect 15934 63250 15986 63262
rect 15934 63186 15986 63198
rect 19070 63250 19122 63262
rect 30594 63198 30606 63250
rect 30658 63198 30670 63250
rect 19070 63186 19122 63198
rect 12350 63138 12402 63150
rect 14926 63138 14978 63150
rect 1474 63086 1486 63138
rect 1538 63086 1550 63138
rect 2370 63086 2382 63138
rect 2434 63086 2446 63138
rect 2706 63086 2718 63138
rect 2770 63086 2782 63138
rect 4162 63086 4174 63138
rect 4226 63086 4238 63138
rect 4946 63086 4958 63138
rect 5010 63086 5022 63138
rect 5730 63086 5742 63138
rect 5794 63086 5806 63138
rect 11218 63086 11230 63138
rect 11282 63086 11294 63138
rect 11666 63086 11678 63138
rect 11730 63086 11742 63138
rect 12898 63086 12910 63138
rect 12962 63086 12974 63138
rect 13906 63086 13918 63138
rect 13970 63086 13982 63138
rect 12350 63074 12402 63086
rect 14926 63074 14978 63086
rect 15262 63138 15314 63150
rect 20750 63138 20802 63150
rect 29486 63138 29538 63150
rect 16930 63086 16942 63138
rect 16994 63086 17006 63138
rect 19506 63086 19518 63138
rect 19570 63086 19582 63138
rect 19954 63086 19966 63138
rect 20018 63086 20030 63138
rect 21074 63086 21086 63138
rect 21138 63086 21150 63138
rect 22082 63086 22094 63138
rect 22146 63086 22158 63138
rect 15262 63074 15314 63086
rect 20750 63074 20802 63086
rect 29486 63074 29538 63086
rect 30270 63138 30322 63150
rect 30270 63074 30322 63086
rect 1934 63026 1986 63038
rect 1934 62962 1986 62974
rect 10894 63026 10946 63038
rect 10894 62962 10946 62974
rect 15710 63026 15762 63038
rect 15710 62962 15762 62974
rect 7422 62914 7474 62926
rect 7422 62850 7474 62862
rect 16046 62914 16098 62926
rect 16046 62850 16098 62862
rect 18622 62914 18674 62926
rect 18622 62850 18674 62862
rect 672 62746 31024 62780
rect 672 62694 3806 62746
rect 3858 62694 3910 62746
rect 3962 62694 4014 62746
rect 4066 62694 23806 62746
rect 23858 62694 23910 62746
rect 23962 62694 24014 62746
rect 24066 62694 31024 62746
rect 672 62660 31024 62694
rect 19630 62578 19682 62590
rect 19630 62514 19682 62526
rect 5630 62466 5682 62478
rect 5630 62402 5682 62414
rect 10894 62466 10946 62478
rect 10894 62402 10946 62414
rect 14254 62466 14306 62478
rect 18050 62414 18062 62466
rect 18114 62414 18126 62466
rect 14254 62402 14306 62414
rect 1150 62354 1202 62366
rect 2830 62354 2882 62366
rect 7310 62354 7362 62366
rect 9550 62354 9602 62366
rect 22318 62354 22370 62366
rect 1474 62302 1486 62354
rect 1538 62302 1550 62354
rect 2034 62302 2046 62354
rect 2098 62302 2110 62354
rect 3378 62302 3390 62354
rect 3442 62302 3454 62354
rect 4274 62302 4286 62354
rect 4338 62302 4350 62354
rect 5954 62302 5966 62354
rect 6018 62302 6030 62354
rect 6402 62302 6414 62354
rect 6466 62302 6478 62354
rect 7634 62302 7646 62354
rect 7698 62302 7710 62354
rect 8642 62302 8654 62354
rect 8706 62302 8718 62354
rect 14578 62302 14590 62354
rect 14642 62302 14654 62354
rect 15026 62302 15038 62354
rect 15090 62302 15102 62354
rect 15810 62302 15822 62354
rect 15874 62302 15886 62354
rect 16258 62302 16270 62354
rect 16322 62302 16334 62354
rect 17266 62302 17278 62354
rect 17330 62302 17342 62354
rect 21074 62302 21086 62354
rect 21138 62302 21150 62354
rect 21522 62302 21534 62354
rect 21586 62302 21598 62354
rect 22642 62302 22654 62354
rect 22706 62302 22718 62354
rect 23762 62302 23774 62354
rect 23826 62302 23838 62354
rect 1150 62290 1202 62302
rect 2830 62290 2882 62302
rect 7310 62290 7362 62302
rect 9550 62290 9602 62302
rect 22318 62290 22370 62302
rect 5294 62242 5346 62254
rect 20638 62242 20690 62254
rect 2146 62190 2158 62242
rect 2210 62190 2222 62242
rect 4946 62190 4958 62242
rect 5010 62190 5022 62242
rect 6626 62190 6638 62242
rect 6690 62190 6702 62242
rect 18386 62190 18398 62242
rect 18450 62190 18462 62242
rect 21634 62190 21646 62242
rect 21698 62190 21710 62242
rect 5294 62178 5346 62190
rect 20638 62178 20690 62190
rect 9202 62078 9214 62130
rect 9266 62078 9278 62130
rect 15250 62078 15262 62130
rect 15314 62078 15326 62130
rect 672 61962 31024 61996
rect 672 61910 4466 61962
rect 4518 61910 4570 61962
rect 4622 61910 4674 61962
rect 4726 61910 24466 61962
rect 24518 61910 24570 61962
rect 24622 61910 24674 61962
rect 24726 61910 31024 61962
rect 672 61876 31024 61910
rect 2158 61794 2210 61806
rect 17614 61794 17666 61806
rect 6066 61742 6078 61794
rect 6130 61742 6142 61794
rect 9986 61742 9998 61794
rect 10050 61742 10062 61794
rect 15698 61742 15710 61794
rect 15762 61742 15774 61794
rect 19170 61742 19182 61794
rect 19234 61742 19246 61794
rect 29810 61742 29822 61794
rect 29874 61742 29886 61794
rect 2158 61730 2210 61742
rect 17614 61730 17666 61742
rect 1374 61682 1426 61694
rect 5070 61682 5122 61694
rect 1026 61630 1038 61682
rect 1090 61630 1102 61682
rect 1810 61630 1822 61682
rect 1874 61630 1886 61682
rect 3490 61630 3502 61682
rect 3554 61630 3566 61682
rect 1374 61618 1426 61630
rect 5070 61618 5122 61630
rect 6526 61682 6578 61694
rect 6526 61618 6578 61630
rect 11566 61682 11618 61694
rect 15374 61682 15426 61694
rect 12562 61630 12574 61682
rect 12626 61630 12638 61682
rect 11566 61618 11618 61630
rect 15374 61618 15426 61630
rect 18174 61682 18226 61694
rect 30594 61630 30606 61682
rect 30658 61630 30670 61682
rect 18174 61618 18226 61630
rect 4622 61570 4674 61582
rect 11118 61570 11170 61582
rect 13022 61570 13074 61582
rect 16830 61570 16882 61582
rect 2930 61518 2942 61570
rect 2994 61518 3006 61570
rect 5394 61518 5406 61570
rect 5458 61518 5470 61570
rect 5954 61518 5966 61570
rect 6018 61518 6030 61570
rect 7298 61518 7310 61570
rect 7362 61518 7374 61570
rect 8194 61518 8206 61570
rect 8258 61518 8270 61570
rect 9426 61518 9438 61570
rect 9490 61518 9502 61570
rect 11890 61518 11902 61570
rect 11954 61518 11966 61570
rect 12450 61518 12462 61570
rect 12514 61518 12526 61570
rect 13570 61518 13582 61570
rect 13634 61518 13646 61570
rect 14578 61518 14590 61570
rect 14642 61518 14654 61570
rect 15586 61518 15598 61570
rect 15650 61518 15662 61570
rect 16034 61518 16046 61570
rect 16098 61518 16110 61570
rect 4622 61506 4674 61518
rect 11118 61506 11170 61518
rect 13022 61506 13074 61518
rect 16830 61506 16882 61518
rect 17054 61570 17106 61582
rect 30270 61570 30322 61582
rect 18610 61518 18622 61570
rect 18674 61518 18686 61570
rect 18946 61518 18958 61570
rect 19010 61518 19022 61570
rect 19730 61518 19742 61570
rect 19794 61518 19806 61570
rect 20402 61518 20414 61570
rect 20466 61518 20478 61570
rect 21186 61518 21198 61570
rect 21250 61518 21262 61570
rect 29586 61518 29598 61570
rect 29650 61518 29662 61570
rect 17054 61506 17106 61518
rect 30270 61506 30322 61518
rect 17726 61458 17778 61470
rect 17726 61394 17778 61406
rect 16718 61346 16770 61358
rect 15922 61294 15934 61346
rect 15986 61294 15998 61346
rect 16718 61282 16770 61294
rect 17166 61346 17218 61358
rect 17166 61282 17218 61294
rect 672 61178 31024 61212
rect 672 61126 3806 61178
rect 3858 61126 3910 61178
rect 3962 61126 4014 61178
rect 4066 61126 23806 61178
rect 23858 61126 23910 61178
rect 23962 61126 24014 61178
rect 24066 61126 31024 61178
rect 672 61092 31024 61126
rect 4286 61010 4338 61022
rect 4286 60946 4338 60958
rect 12126 61010 12178 61022
rect 12126 60946 12178 60958
rect 14814 61010 14866 61022
rect 14814 60946 14866 60958
rect 5630 60898 5682 60910
rect 20638 60898 20690 60910
rect 10546 60846 10558 60898
rect 10610 60846 10622 60898
rect 5630 60834 5682 60846
rect 20638 60834 20690 60846
rect 7310 60786 7362 60798
rect 19294 60786 19346 60798
rect 2594 60734 2606 60786
rect 2658 60734 2670 60786
rect 5954 60734 5966 60786
rect 6018 60734 6030 60786
rect 6402 60734 6414 60786
rect 6466 60734 6478 60786
rect 7634 60734 7646 60786
rect 7698 60734 7710 60786
rect 8642 60734 8654 60786
rect 8706 60734 8718 60786
rect 13122 60734 13134 60786
rect 13186 60734 13198 60786
rect 15362 60734 15374 60786
rect 15426 60734 15438 60786
rect 17602 60734 17614 60786
rect 17666 60734 17678 60786
rect 20962 60734 20974 60786
rect 21026 60734 21038 60786
rect 21410 60734 21422 60786
rect 21474 60734 21486 60786
rect 22642 60734 22654 60786
rect 22706 60734 22718 60786
rect 23650 60734 23662 60786
rect 23714 60734 23726 60786
rect 7310 60722 7362 60734
rect 19294 60722 19346 60734
rect 2158 60674 2210 60686
rect 22094 60674 22146 60686
rect 6626 60622 6638 60674
rect 6690 60622 6702 60674
rect 10994 60622 11006 60674
rect 11058 60622 11070 60674
rect 13682 60622 13694 60674
rect 13746 60622 13758 60674
rect 15922 60622 15934 60674
rect 15986 60622 15998 60674
rect 18162 60622 18174 60674
rect 18226 60622 18238 60674
rect 21634 60622 21646 60674
rect 21698 60622 21710 60674
rect 29810 60622 29822 60674
rect 29874 60622 29886 60674
rect 2158 60610 2210 60622
rect 22094 60610 22146 60622
rect 1374 60562 1426 60574
rect 17054 60562 17106 60574
rect 1026 60510 1038 60562
rect 1090 60510 1102 60562
rect 1810 60510 1822 60562
rect 1874 60510 1886 60562
rect 3154 60510 3166 60562
rect 3218 60510 3230 60562
rect 1374 60498 1426 60510
rect 17054 60498 17106 60510
rect 29486 60562 29538 60574
rect 29486 60498 29538 60510
rect 30270 60562 30322 60574
rect 30594 60510 30606 60562
rect 30658 60510 30670 60562
rect 30270 60498 30322 60510
rect 672 60394 31024 60428
rect 672 60342 4466 60394
rect 4518 60342 4570 60394
rect 4622 60342 4674 60394
rect 4726 60342 24466 60394
rect 24518 60342 24570 60394
rect 24622 60342 24674 60394
rect 24726 60342 31024 60394
rect 672 60308 31024 60342
rect 1150 60226 1202 60238
rect 5182 60226 5234 60238
rect 4050 60174 4062 60226
rect 4114 60174 4126 60226
rect 1150 60162 1202 60174
rect 5182 60162 5234 60174
rect 7422 60226 7474 60238
rect 7422 60162 7474 60174
rect 11118 60226 11170 60238
rect 11118 60162 11170 60174
rect 11902 60226 11954 60238
rect 15934 60226 15986 60238
rect 14802 60174 14814 60226
rect 14866 60174 14878 60226
rect 11902 60162 11954 60174
rect 15934 60162 15986 60174
rect 20638 60226 20690 60238
rect 29810 60174 29822 60226
rect 29874 60174 29886 60226
rect 20638 60162 20690 60174
rect 16942 60114 16994 60126
rect 2370 60062 2382 60114
rect 2434 60062 2446 60114
rect 6290 60062 6302 60114
rect 6354 60062 6366 60114
rect 9874 60062 9886 60114
rect 9938 60062 9950 60114
rect 11554 60062 11566 60114
rect 11618 60062 11630 60114
rect 17938 60062 17950 60114
rect 18002 60062 18014 60114
rect 21858 60062 21870 60114
rect 21922 60062 21934 60114
rect 16942 60050 16994 60062
rect 16606 60002 16658 60014
rect 29486 60002 29538 60014
rect 9538 59950 9550 60002
rect 9602 59950 9614 60002
rect 14242 59950 14254 60002
rect 14306 59950 14318 60002
rect 17266 59950 17278 60002
rect 17330 59950 17342 60002
rect 17826 59950 17838 60002
rect 17890 59950 17902 60002
rect 18498 59950 18510 60002
rect 18562 59950 18574 60002
rect 18946 59950 18958 60002
rect 19010 59950 19022 60002
rect 20066 59950 20078 60002
rect 20130 59950 20142 60002
rect 16606 59938 16658 59950
rect 29486 59938 29538 59950
rect 2706 59838 2718 59890
rect 2770 59838 2782 59890
rect 3602 59838 3614 59890
rect 3666 59838 3678 59890
rect 5842 59838 5854 59890
rect 5906 59838 5918 59890
rect 22194 59838 22206 59890
rect 22258 59838 22270 59890
rect 672 59610 31024 59644
rect 672 59558 3806 59610
rect 3858 59558 3910 59610
rect 3962 59558 4014 59610
rect 4066 59558 23806 59610
rect 23858 59558 23910 59610
rect 23962 59558 24014 59610
rect 24066 59558 31024 59610
rect 672 59524 31024 59558
rect 18510 59442 18562 59454
rect 18510 59378 18562 59390
rect 18958 59330 19010 59342
rect 18958 59266 19010 59278
rect 2158 59218 2210 59230
rect 8306 59166 8318 59218
rect 8370 59166 8382 59218
rect 14690 59166 14702 59218
rect 14754 59166 14766 59218
rect 16818 59166 16830 59218
rect 16882 59166 16894 59218
rect 2158 59154 2210 59166
rect 2830 59106 2882 59118
rect 2482 59054 2494 59106
rect 2546 59054 2558 59106
rect 8754 59054 8766 59106
rect 8818 59054 8830 59106
rect 15026 59054 15038 59106
rect 15090 59054 15102 59106
rect 17378 59054 17390 59106
rect 17442 59054 17454 59106
rect 2830 59042 2882 59054
rect 1374 58994 1426 59006
rect 9886 58994 9938 59006
rect 1026 58942 1038 58994
rect 1090 58942 1102 58994
rect 1810 58942 1822 58994
rect 1874 58942 1886 58994
rect 1374 58930 1426 58942
rect 9886 58930 9938 58942
rect 16270 58994 16322 59006
rect 16270 58930 16322 58942
rect 30270 58994 30322 59006
rect 30594 58942 30606 58994
rect 30658 58942 30670 58994
rect 30270 58930 30322 58942
rect 672 58826 31024 58860
rect 672 58774 4466 58826
rect 4518 58774 4570 58826
rect 4622 58774 4674 58826
rect 4726 58774 24466 58826
rect 24518 58774 24570 58826
rect 24622 58774 24674 58826
rect 24726 58774 31024 58826
rect 672 58740 31024 58774
rect 1374 58658 1426 58670
rect 17054 58658 17106 58670
rect 16706 58606 16718 58658
rect 16770 58606 16782 58658
rect 1374 58594 1426 58606
rect 17054 58594 17106 58606
rect 20638 58658 20690 58670
rect 29810 58606 29822 58658
rect 29874 58606 29886 58658
rect 20638 58594 20690 58606
rect 1026 58494 1038 58546
rect 1090 58494 1102 58546
rect 1698 58494 1710 58546
rect 1762 58494 1774 58546
rect 9986 58494 9998 58546
rect 10050 58494 10062 58546
rect 14018 58494 14030 58546
rect 14082 58494 14094 58546
rect 19394 58494 19406 58546
rect 19458 58494 19470 58546
rect 30594 58494 30606 58546
rect 30658 58494 30670 58546
rect 2046 58434 2098 58446
rect 29486 58434 29538 58446
rect 9650 58382 9662 58434
rect 9714 58382 9726 58434
rect 13682 58382 13694 58434
rect 13746 58382 13758 58434
rect 19058 58382 19070 58434
rect 19122 58382 19134 58434
rect 2046 58370 2098 58382
rect 29486 58370 29538 58382
rect 30270 58434 30322 58446
rect 30270 58370 30322 58382
rect 11230 58210 11282 58222
rect 11230 58146 11282 58158
rect 15262 58210 15314 58222
rect 15262 58146 15314 58158
rect 672 58042 31024 58076
rect 672 57990 3806 58042
rect 3858 57990 3910 58042
rect 3962 57990 4014 58042
rect 4066 57990 23806 58042
rect 23858 57990 23910 58042
rect 23962 57990 24014 58042
rect 24066 57990 31024 58042
rect 672 57956 31024 57990
rect 14590 57762 14642 57774
rect 8082 57710 8094 57762
rect 8146 57710 8158 57762
rect 10322 57710 10334 57762
rect 10386 57710 10398 57762
rect 14590 57698 14642 57710
rect 18958 57762 19010 57774
rect 18958 57698 19010 57710
rect 1374 57650 1426 57662
rect 16270 57650 16322 57662
rect 15026 57598 15038 57650
rect 15090 57598 15102 57650
rect 15362 57598 15374 57650
rect 15426 57598 15438 57650
rect 16706 57598 16718 57650
rect 16770 57598 16782 57650
rect 17714 57598 17726 57650
rect 17778 57598 17790 57650
rect 1374 57586 1426 57598
rect 16270 57586 16322 57598
rect 1026 57486 1038 57538
rect 1090 57486 1102 57538
rect 8530 57486 8542 57538
rect 8594 57486 8606 57538
rect 10770 57486 10782 57538
rect 10834 57486 10846 57538
rect 13570 57486 13582 57538
rect 13634 57486 13646 57538
rect 13906 57486 13918 57538
rect 13970 57486 13982 57538
rect 29810 57486 29822 57538
rect 29874 57486 29886 57538
rect 9662 57426 9714 57438
rect 9662 57362 9714 57374
rect 11902 57426 11954 57438
rect 11902 57362 11954 57374
rect 13246 57426 13298 57438
rect 13246 57362 13298 57374
rect 14254 57426 14306 57438
rect 29486 57426 29538 57438
rect 15586 57374 15598 57426
rect 15650 57374 15662 57426
rect 14254 57362 14306 57374
rect 29486 57362 29538 57374
rect 672 57258 31024 57292
rect 672 57206 4466 57258
rect 4518 57206 4570 57258
rect 4622 57206 4674 57258
rect 4726 57206 24466 57258
rect 24518 57206 24570 57258
rect 24622 57206 24674 57258
rect 24726 57206 31024 57258
rect 672 57172 31024 57206
rect 18958 57090 19010 57102
rect 18958 57026 19010 57038
rect 10110 56978 10162 56990
rect 4834 56926 4846 56978
rect 4898 56926 4910 56978
rect 7074 56926 7086 56978
rect 7138 56926 7150 56978
rect 11106 56926 11118 56978
rect 11170 56926 11182 56978
rect 30594 56926 30606 56978
rect 30658 56926 30670 56978
rect 10110 56914 10162 56926
rect 6626 56814 6638 56866
rect 6690 56814 6702 56866
rect 10434 56814 10446 56866
rect 10498 56814 10510 56866
rect 10994 56814 11006 56866
rect 11058 56814 11070 56866
rect 11666 56814 11678 56866
rect 11730 56814 11742 56866
rect 12338 56814 12350 56866
rect 12402 56814 12414 56866
rect 13122 56814 13134 56866
rect 13186 56814 13198 56866
rect 30370 56814 30382 56866
rect 30434 56814 30446 56866
rect 4386 56702 4398 56754
rect 4450 56702 4462 56754
rect 5966 56642 6018 56654
rect 5966 56578 6018 56590
rect 8206 56642 8258 56654
rect 8206 56578 8258 56590
rect 672 56474 31024 56508
rect 672 56422 3806 56474
rect 3858 56422 3910 56474
rect 3962 56422 4014 56474
rect 4066 56422 23806 56474
rect 23858 56422 23910 56474
rect 23962 56422 24014 56474
rect 24066 56422 31024 56474
rect 672 56388 31024 56422
rect 8990 56194 9042 56206
rect 18958 56194 19010 56206
rect 5842 56142 5854 56194
rect 5906 56142 5918 56194
rect 14466 56142 14478 56194
rect 14530 56142 14542 56194
rect 8990 56130 9042 56142
rect 18958 56130 19010 56142
rect 10670 56082 10722 56094
rect 9426 56030 9438 56082
rect 9490 56030 9502 56082
rect 9874 56030 9886 56082
rect 9938 56030 9950 56082
rect 11218 56030 11230 56082
rect 11282 56030 11294 56082
rect 12114 56030 12126 56082
rect 12178 56030 12190 56082
rect 10670 56018 10722 56030
rect 14018 55918 14030 55970
rect 14082 55918 14094 55970
rect 21298 55918 21310 55970
rect 21362 55918 21374 55970
rect 7422 55858 7474 55870
rect 12910 55858 12962 55870
rect 6290 55806 6302 55858
rect 6354 55806 6366 55858
rect 9986 55806 9998 55858
rect 10050 55806 10062 55858
rect 7422 55794 7474 55806
rect 12910 55794 12962 55806
rect 20974 55858 21026 55870
rect 20974 55794 21026 55806
rect 30270 55858 30322 55870
rect 30594 55806 30606 55858
rect 30658 55806 30670 55858
rect 30270 55794 30322 55806
rect 672 55690 31024 55724
rect 672 55638 4466 55690
rect 4518 55638 4570 55690
rect 4622 55638 4674 55690
rect 4726 55638 24466 55690
rect 24518 55638 24570 55690
rect 24622 55638 24674 55690
rect 24726 55638 31024 55690
rect 672 55604 31024 55638
rect 18958 55522 19010 55534
rect 30482 55470 30494 55522
rect 30546 55470 30558 55522
rect 18958 55458 19010 55470
rect 5070 55410 5122 55422
rect 3490 55358 3502 55410
rect 3554 55358 3566 55410
rect 6066 55358 6078 55410
rect 6130 55358 6142 55410
rect 9762 55358 9774 55410
rect 9826 55358 9838 55410
rect 14130 55358 14142 55410
rect 14194 55358 14206 55410
rect 5070 55346 5122 55358
rect 4622 55298 4674 55310
rect 6526 55298 6578 55310
rect 30158 55298 30210 55310
rect 2930 55246 2942 55298
rect 2994 55246 3006 55298
rect 5394 55246 5406 55298
rect 5458 55246 5470 55298
rect 5842 55246 5854 55298
rect 5906 55246 5918 55298
rect 7298 55246 7310 55298
rect 7362 55246 7374 55298
rect 8082 55246 8094 55298
rect 8146 55246 8158 55298
rect 9314 55246 9326 55298
rect 9378 55246 9390 55298
rect 28354 55246 28366 55298
rect 28418 55246 28430 55298
rect 4622 55234 4674 55246
rect 6526 55234 6578 55246
rect 30158 55234 30210 55246
rect 13682 55134 13694 55186
rect 13746 55134 13758 55186
rect 24770 55134 24782 55186
rect 24834 55134 24846 55186
rect 11006 55074 11058 55086
rect 11006 55010 11058 55022
rect 15262 55074 15314 55086
rect 15262 55010 15314 55022
rect 672 54906 31024 54940
rect 672 54854 3806 54906
rect 3858 54854 3910 54906
rect 3962 54854 4014 54906
rect 4066 54854 23806 54906
rect 23858 54854 23910 54906
rect 23962 54854 24014 54906
rect 24066 54854 31024 54906
rect 672 54820 31024 54854
rect 3726 54738 3778 54750
rect 3726 54674 3778 54686
rect 5742 54626 5794 54638
rect 2146 54574 2158 54626
rect 2210 54574 2222 54626
rect 5742 54562 5794 54574
rect 14142 54626 14194 54638
rect 14142 54562 14194 54574
rect 7422 54514 7474 54526
rect 15822 54514 15874 54526
rect 6066 54462 6078 54514
rect 6130 54462 6142 54514
rect 6514 54462 6526 54514
rect 6578 54462 6590 54514
rect 7746 54462 7758 54514
rect 7810 54462 7822 54514
rect 8754 54462 8766 54514
rect 8818 54462 8830 54514
rect 10434 54462 10446 54514
rect 10498 54462 10510 54514
rect 14578 54462 14590 54514
rect 14642 54462 14654 54514
rect 14914 54462 14926 54514
rect 14978 54462 14990 54514
rect 16146 54462 16158 54514
rect 16210 54462 16222 54514
rect 17154 54462 17166 54514
rect 17218 54462 17230 54514
rect 7422 54450 7474 54462
rect 15822 54450 15874 54462
rect 2482 54350 2494 54402
rect 2546 54350 2558 54402
rect 10882 54350 10894 54402
rect 10946 54350 10958 54402
rect 30594 54350 30606 54402
rect 30658 54350 30670 54402
rect 12126 54290 12178 54302
rect 30270 54290 30322 54302
rect 6738 54238 6750 54290
rect 6802 54238 6814 54290
rect 15138 54238 15150 54290
rect 15202 54238 15214 54290
rect 12126 54226 12178 54238
rect 30270 54226 30322 54238
rect 672 54122 31024 54156
rect 672 54070 4466 54122
rect 4518 54070 4570 54122
rect 4622 54070 4674 54122
rect 4726 54070 24466 54122
rect 24518 54070 24570 54122
rect 24622 54070 24674 54122
rect 24726 54070 31024 54122
rect 672 54036 31024 54070
rect 3490 53790 3502 53842
rect 3554 53790 3566 53842
rect 10546 53790 10558 53842
rect 10610 53790 10622 53842
rect 15586 53790 15598 53842
rect 15650 53790 15662 53842
rect 21746 53790 21758 53842
rect 21810 53790 21822 53842
rect 30594 53790 30606 53842
rect 30658 53790 30670 53842
rect 6750 53730 6802 53742
rect 2930 53678 2942 53730
rect 2994 53678 3006 53730
rect 6750 53666 6802 53678
rect 9550 53730 9602 53742
rect 15262 53730 15314 53742
rect 9874 53678 9886 53730
rect 9938 53678 9950 53730
rect 10322 53678 10334 53730
rect 10386 53678 10398 53730
rect 11106 53678 11118 53730
rect 11170 53678 11182 53730
rect 11666 53678 11678 53730
rect 11730 53678 11742 53730
rect 12562 53678 12574 53730
rect 12626 53678 12638 53730
rect 9550 53666 9602 53678
rect 15262 53666 15314 53678
rect 21422 53730 21474 53742
rect 30370 53678 30382 53730
rect 30434 53678 30446 53730
rect 21422 53666 21474 53678
rect 14030 53618 14082 53630
rect 14030 53554 14082 53566
rect 4622 53506 4674 53518
rect 4622 53442 4674 53454
rect 672 53338 31024 53372
rect 672 53286 3806 53338
rect 3858 53286 3910 53338
rect 3962 53286 4014 53338
rect 4066 53286 23806 53338
rect 23858 53286 23910 53338
rect 23962 53286 24014 53338
rect 24066 53286 31024 53338
rect 672 53252 31024 53286
rect 10894 53170 10946 53182
rect 10894 53106 10946 53118
rect 16046 53170 16098 53182
rect 16046 53106 16098 53118
rect 8430 52946 8482 52958
rect 11230 52946 11282 52958
rect 16494 52946 16546 52958
rect 2594 52894 2606 52946
rect 2658 52894 2670 52946
rect 6962 52894 6974 52946
rect 7026 52894 7038 52946
rect 8082 52894 8094 52946
rect 8146 52894 8158 52946
rect 9202 52894 9214 52946
rect 9266 52894 9278 52946
rect 9650 52894 9662 52946
rect 9714 52894 9726 52946
rect 12002 52894 12014 52946
rect 12066 52894 12078 52946
rect 14466 52894 14478 52946
rect 14530 52894 14542 52946
rect 8430 52882 8482 52894
rect 11230 52882 11282 52894
rect 16494 52882 16546 52894
rect 10110 52834 10162 52846
rect 3042 52782 3054 52834
rect 3106 52782 3118 52834
rect 11778 52782 11790 52834
rect 11842 52782 11854 52834
rect 14914 52782 14926 52834
rect 14978 52782 14990 52834
rect 10110 52770 10162 52782
rect 4286 52722 4338 52734
rect 30270 52722 30322 52734
rect 9090 52670 9102 52722
rect 9154 52670 9166 52722
rect 16818 52670 16830 52722
rect 16882 52670 16894 52722
rect 30594 52670 30606 52722
rect 30658 52670 30670 52722
rect 4286 52658 4338 52670
rect 30270 52658 30322 52670
rect 672 52554 31024 52588
rect 672 52502 4466 52554
rect 4518 52502 4570 52554
rect 4622 52502 4674 52554
rect 4726 52502 24466 52554
rect 24518 52502 24570 52554
rect 24622 52502 24674 52554
rect 24726 52502 31024 52554
rect 672 52468 31024 52502
rect 4510 52386 4562 52398
rect 11106 52334 11118 52386
rect 11170 52334 11182 52386
rect 14914 52334 14926 52386
rect 14978 52334 14990 52386
rect 4510 52322 4562 52334
rect 10110 52274 10162 52286
rect 3266 52222 3278 52274
rect 3330 52222 3342 52274
rect 17042 52222 17054 52274
rect 17106 52222 17118 52274
rect 10110 52210 10162 52222
rect 6862 52162 6914 52174
rect 11566 52162 11618 52174
rect 10434 52110 10446 52162
rect 10498 52110 10510 52162
rect 10882 52110 10894 52162
rect 10946 52110 10958 52162
rect 12114 52110 12126 52162
rect 12178 52110 12190 52162
rect 13122 52110 13134 52162
rect 13186 52110 13198 52162
rect 16818 52110 16830 52162
rect 16882 52110 16894 52162
rect 6862 52098 6914 52110
rect 11566 52098 11618 52110
rect 2930 51998 2942 52050
rect 2994 51998 3006 52050
rect 15362 51998 15374 52050
rect 15426 51998 15438 52050
rect 13806 51938 13858 51950
rect 13806 51874 13858 51886
rect 672 51770 31024 51804
rect 672 51718 3806 51770
rect 3858 51718 3910 51770
rect 3962 51718 4014 51770
rect 4066 51718 23806 51770
rect 23858 51718 23910 51770
rect 23962 51718 24014 51770
rect 24066 51718 31024 51770
rect 672 51684 31024 51718
rect 4958 51490 5010 51502
rect 4958 51426 5010 51438
rect 6414 51378 6466 51390
rect 10670 51378 10722 51390
rect 14254 51378 14306 51390
rect 2706 51326 2718 51378
rect 2770 51326 2782 51378
rect 5282 51326 5294 51378
rect 5346 51326 5358 51378
rect 5842 51326 5854 51378
rect 5906 51326 5918 51378
rect 7074 51326 7086 51378
rect 7138 51326 7150 51378
rect 7970 51326 7982 51378
rect 8034 51326 8046 51378
rect 9314 51326 9326 51378
rect 9378 51326 9390 51378
rect 9874 51326 9886 51378
rect 9938 51326 9950 51378
rect 11218 51326 11230 51378
rect 11282 51326 11294 51378
rect 12002 51326 12014 51378
rect 12066 51326 12078 51378
rect 13122 51326 13134 51378
rect 13186 51326 13198 51378
rect 13682 51326 13694 51378
rect 13746 51326 13758 51378
rect 14802 51326 14814 51378
rect 14866 51326 14878 51378
rect 15810 51326 15822 51378
rect 15874 51326 15886 51378
rect 6414 51314 6466 51326
rect 10670 51314 10722 51326
rect 14254 51314 14306 51326
rect 8990 51266 9042 51278
rect 12798 51266 12850 51278
rect 3042 51214 3054 51266
rect 3106 51214 3118 51266
rect 9986 51214 9998 51266
rect 10050 51214 10062 51266
rect 8990 51202 9042 51214
rect 12798 51202 12850 51214
rect 4286 51154 4338 51166
rect 16942 51154 16994 51166
rect 30270 51154 30322 51166
rect 5954 51102 5966 51154
rect 6018 51102 6030 51154
rect 13794 51102 13806 51154
rect 13858 51102 13870 51154
rect 17266 51102 17278 51154
rect 17330 51102 17342 51154
rect 30594 51102 30606 51154
rect 30658 51102 30670 51154
rect 4286 51090 4338 51102
rect 16942 51090 16994 51102
rect 30270 51090 30322 51102
rect 672 50986 31024 51020
rect 672 50934 4466 50986
rect 4518 50934 4570 50986
rect 4622 50934 4674 50986
rect 4726 50934 24466 50986
rect 24518 50934 24570 50986
rect 24622 50934 24674 50986
rect 24726 50934 31024 50986
rect 672 50900 31024 50934
rect 1150 50818 1202 50830
rect 2482 50766 2494 50818
rect 2546 50766 2558 50818
rect 5058 50766 5070 50818
rect 5122 50766 5134 50818
rect 10770 50766 10782 50818
rect 10834 50766 10846 50818
rect 17938 50766 17950 50818
rect 18002 50766 18014 50818
rect 1150 50754 1202 50766
rect 3614 50706 3666 50718
rect 1474 50654 1486 50706
rect 1538 50654 1550 50706
rect 3614 50642 3666 50654
rect 5518 50706 5570 50718
rect 12786 50654 12798 50706
rect 12850 50654 12862 50706
rect 30594 50654 30606 50706
rect 30658 50654 30670 50706
rect 5518 50642 5570 50654
rect 13246 50594 13298 50606
rect 2034 50542 2046 50594
rect 2098 50542 2110 50594
rect 4386 50542 4398 50594
rect 4450 50542 4462 50594
rect 4946 50542 4958 50594
rect 5010 50542 5022 50594
rect 6066 50542 6078 50594
rect 6130 50542 6142 50594
rect 7074 50542 7086 50594
rect 7138 50542 7150 50594
rect 11218 50542 11230 50594
rect 11282 50542 11294 50594
rect 12114 50542 12126 50594
rect 12178 50542 12190 50594
rect 12562 50542 12574 50594
rect 12626 50542 12638 50594
rect 13794 50542 13806 50594
rect 13858 50542 13870 50594
rect 14018 50542 14030 50594
rect 14082 50542 14094 50594
rect 14802 50542 14814 50594
rect 14866 50542 14878 50594
rect 30370 50542 30382 50594
rect 30434 50542 30446 50594
rect 13246 50530 13298 50542
rect 4062 50482 4114 50494
rect 4062 50418 4114 50430
rect 11790 50482 11842 50494
rect 11790 50418 11842 50430
rect 15262 50482 15314 50494
rect 18386 50430 18398 50482
rect 18450 50430 18462 50482
rect 15262 50418 15314 50430
rect 9662 50370 9714 50382
rect 9662 50306 9714 50318
rect 16830 50370 16882 50382
rect 16830 50306 16882 50318
rect 672 50202 31024 50236
rect 672 50150 3806 50202
rect 3858 50150 3910 50202
rect 3962 50150 4014 50202
rect 4066 50150 23806 50202
rect 23858 50150 23910 50202
rect 23962 50150 24014 50202
rect 24066 50150 31024 50202
rect 672 50116 31024 50150
rect 8542 50034 8594 50046
rect 8542 49970 8594 49982
rect 12126 50034 12178 50046
rect 12126 49970 12178 49982
rect 13246 50034 13298 50046
rect 13246 49970 13298 49982
rect 9886 49810 9938 49822
rect 16830 49810 16882 49822
rect 1474 49758 1486 49810
rect 1538 49758 1550 49810
rect 6962 49758 6974 49810
rect 7026 49758 7038 49810
rect 10546 49758 10558 49810
rect 10610 49758 10622 49810
rect 14802 49758 14814 49810
rect 14866 49758 14878 49810
rect 15810 49758 15822 49810
rect 15874 49758 15886 49810
rect 16146 49758 16158 49810
rect 16210 49758 16222 49810
rect 17378 49758 17390 49810
rect 17442 49758 17454 49810
rect 18386 49758 18398 49810
rect 18450 49758 18462 49810
rect 9886 49746 9938 49758
rect 16830 49746 16882 49758
rect 15374 49698 15426 49710
rect 1922 49646 1934 49698
rect 1986 49646 1998 49698
rect 10994 49646 11006 49698
rect 11058 49646 11070 49698
rect 14466 49646 14478 49698
rect 14530 49646 14542 49698
rect 15374 49634 15426 49646
rect 3166 49586 3218 49598
rect 9998 49586 10050 49598
rect 7410 49534 7422 49586
rect 7474 49534 7486 49586
rect 16370 49534 16382 49586
rect 16434 49534 16446 49586
rect 3166 49522 3218 49534
rect 9998 49522 10050 49534
rect 672 49418 31024 49452
rect 672 49366 4466 49418
rect 4518 49366 4570 49418
rect 4622 49366 4674 49418
rect 4726 49366 24466 49418
rect 24518 49366 24570 49418
rect 24622 49366 24674 49418
rect 24726 49366 31024 49418
rect 672 49332 31024 49366
rect 2270 49250 2322 49262
rect 2270 49186 2322 49198
rect 8206 49250 8258 49262
rect 11566 49250 11618 49262
rect 10434 49198 10446 49250
rect 10498 49198 10510 49250
rect 12674 49198 12686 49250
rect 12738 49198 12750 49250
rect 8206 49186 8258 49198
rect 11566 49186 11618 49198
rect 1362 49086 1374 49138
rect 1426 49086 1438 49138
rect 1586 49086 1598 49138
rect 1650 49086 1662 49138
rect 3714 49086 3726 49138
rect 3778 49086 3790 49138
rect 7074 49086 7086 49138
rect 7138 49086 7150 49138
rect 19730 49086 19742 49138
rect 19794 49086 19806 49138
rect 30594 49086 30606 49138
rect 30658 49086 30670 49138
rect 1934 49026 1986 49038
rect 4174 49026 4226 49038
rect 19406 49026 19458 49038
rect 3042 48974 3054 49026
rect 3106 48974 3118 49026
rect 3602 48974 3614 49026
rect 3666 48974 3678 49026
rect 4834 48974 4846 49026
rect 4898 48974 4910 49026
rect 5842 48974 5854 49026
rect 5906 48974 5918 49026
rect 6626 48974 6638 49026
rect 6690 48974 6702 49026
rect 12114 48974 12126 49026
rect 12178 48974 12190 49026
rect 1934 48962 1986 48974
rect 4174 48962 4226 48974
rect 19406 48962 19458 48974
rect 30270 49026 30322 49038
rect 30270 48962 30322 48974
rect 2718 48914 2770 48926
rect 15262 48914 15314 48926
rect 9986 48862 9998 48914
rect 10050 48862 10062 48914
rect 2718 48850 2770 48862
rect 15262 48850 15314 48862
rect 13806 48802 13858 48814
rect 13806 48738 13858 48750
rect 672 48634 31024 48668
rect 672 48582 3806 48634
rect 3858 48582 3910 48634
rect 3962 48582 4014 48634
rect 4066 48582 23806 48634
rect 23858 48582 23910 48634
rect 23962 48582 24014 48634
rect 24066 48582 31024 48634
rect 672 48548 31024 48582
rect 2158 48466 2210 48478
rect 2158 48402 2210 48414
rect 15934 48466 15986 48478
rect 15934 48402 15986 48414
rect 12226 48302 12238 48354
rect 12290 48302 12302 48354
rect 16594 48302 16606 48354
rect 16658 48302 16670 48354
rect 11902 48242 11954 48254
rect 3714 48190 3726 48242
rect 3778 48190 3790 48242
rect 6626 48190 6638 48242
rect 6690 48190 6702 48242
rect 10770 48190 10782 48242
rect 10834 48190 10846 48242
rect 11902 48178 11954 48190
rect 13358 48242 13410 48254
rect 13358 48178 13410 48190
rect 13470 48242 13522 48254
rect 13570 48190 13582 48242
rect 13634 48190 13646 48242
rect 14354 48190 14366 48242
rect 14418 48190 14430 48242
rect 13470 48178 13522 48190
rect 11342 48130 11394 48142
rect 3378 48078 3390 48130
rect 3442 48078 3454 48130
rect 7074 48078 7086 48130
rect 7138 48078 7150 48130
rect 11342 48066 11394 48078
rect 11454 48130 11506 48142
rect 11454 48066 11506 48078
rect 11678 48130 11730 48142
rect 11678 48066 11730 48078
rect 13022 48130 13074 48142
rect 13234 48078 13246 48130
rect 13298 48078 13310 48130
rect 16930 48078 16942 48130
rect 16994 48078 17006 48130
rect 18946 48078 18958 48130
rect 19010 48078 19022 48130
rect 13022 48066 13074 48078
rect 8318 48018 8370 48030
rect 8318 47954 8370 47966
rect 9102 48018 9154 48030
rect 12126 48018 12178 48030
rect 10210 47966 10222 48018
rect 10274 47966 10286 48018
rect 9102 47954 9154 47966
rect 12126 47954 12178 47966
rect 13806 48018 13858 48030
rect 18174 48018 18226 48030
rect 14802 47966 14814 48018
rect 14866 47966 14878 48018
rect 13806 47954 13858 47966
rect 18174 47954 18226 47966
rect 18622 48018 18674 48030
rect 18622 47954 18674 47966
rect 30270 48018 30322 48030
rect 30594 47966 30606 48018
rect 30658 47966 30670 48018
rect 30270 47954 30322 47966
rect 672 47850 31024 47884
rect 672 47798 4466 47850
rect 4518 47798 4570 47850
rect 4622 47798 4674 47850
rect 4726 47798 24466 47850
rect 24518 47798 24570 47850
rect 24622 47798 24674 47850
rect 24726 47798 31024 47850
rect 672 47764 31024 47798
rect 3266 47630 3278 47682
rect 3330 47630 3342 47682
rect 10210 47630 10222 47682
rect 10274 47630 10286 47682
rect 14802 47630 14814 47682
rect 14866 47630 14878 47682
rect 3726 47570 3778 47582
rect 9214 47570 9266 47582
rect 1922 47518 1934 47570
rect 1986 47518 1998 47570
rect 6514 47518 6526 47570
rect 6578 47518 6590 47570
rect 3726 47506 3778 47518
rect 9214 47506 9266 47518
rect 10670 47570 10722 47582
rect 10670 47506 10722 47518
rect 13470 47570 13522 47582
rect 18174 47570 18226 47582
rect 17714 47518 17726 47570
rect 17778 47518 17790 47570
rect 30594 47518 30606 47570
rect 30658 47518 30670 47570
rect 13470 47506 13522 47518
rect 18174 47506 18226 47518
rect 13022 47458 13074 47470
rect 1698 47406 1710 47458
rect 1762 47406 1774 47458
rect 2706 47406 2718 47458
rect 2770 47406 2782 47458
rect 3042 47406 3054 47458
rect 3106 47406 3118 47458
rect 4274 47406 4286 47458
rect 4338 47406 4350 47458
rect 5394 47406 5406 47458
rect 5458 47406 5470 47458
rect 9538 47406 9550 47458
rect 9602 47406 9614 47458
rect 9986 47406 9998 47458
rect 10050 47406 10062 47458
rect 11218 47406 11230 47458
rect 11282 47406 11294 47458
rect 12226 47406 12238 47458
rect 12290 47406 12302 47458
rect 13022 47394 13074 47406
rect 15934 47458 15986 47470
rect 30270 47458 30322 47470
rect 17042 47406 17054 47458
rect 17106 47406 17118 47458
rect 17490 47406 17502 47458
rect 17554 47406 17566 47458
rect 18722 47406 18734 47458
rect 18786 47406 18798 47458
rect 19730 47406 19742 47458
rect 19794 47406 19806 47458
rect 15934 47394 15986 47406
rect 30270 47394 30322 47406
rect 2270 47346 2322 47358
rect 8206 47346 8258 47358
rect 16718 47346 16770 47358
rect 6066 47294 6078 47346
rect 6130 47294 6142 47346
rect 14354 47294 14366 47346
rect 14418 47294 14430 47346
rect 2270 47282 2322 47294
rect 8206 47282 8258 47294
rect 16718 47282 16770 47294
rect 7646 47234 7698 47246
rect 7646 47170 7698 47182
rect 8094 47234 8146 47246
rect 8094 47170 8146 47182
rect 13134 47234 13186 47246
rect 13134 47170 13186 47182
rect 13358 47234 13410 47246
rect 13358 47170 13410 47182
rect 672 47066 31024 47100
rect 672 47014 3806 47066
rect 3858 47014 3910 47066
rect 3962 47014 4014 47066
rect 4066 47014 23806 47066
rect 23858 47014 23910 47066
rect 23962 47014 24014 47066
rect 24066 47014 31024 47066
rect 672 46980 31024 47014
rect 3166 46898 3218 46910
rect 3166 46834 3218 46846
rect 12910 46898 12962 46910
rect 12910 46834 12962 46846
rect 5854 46674 5906 46686
rect 1474 46622 1486 46674
rect 1538 46622 1550 46674
rect 5170 46622 5182 46674
rect 5234 46622 5246 46674
rect 7186 46622 7198 46674
rect 7250 46622 7262 46674
rect 7522 46622 7534 46674
rect 7586 46622 7598 46674
rect 8306 46622 8318 46674
rect 8370 46622 8382 46674
rect 8978 46622 8990 46674
rect 9042 46622 9054 46674
rect 9874 46622 9886 46674
rect 9938 46622 9950 46674
rect 12002 46622 12014 46674
rect 12066 46622 12078 46674
rect 14466 46622 14478 46674
rect 14530 46622 14542 46674
rect 5854 46610 5906 46622
rect 6750 46562 6802 46574
rect 1922 46510 1934 46562
rect 1986 46510 1998 46562
rect 5058 46510 5070 46562
rect 5122 46510 5134 46562
rect 7746 46510 7758 46562
rect 7810 46510 7822 46562
rect 16370 46510 16382 46562
rect 16434 46510 16446 46562
rect 23538 46510 23550 46562
rect 23602 46510 23614 46562
rect 6750 46498 6802 46510
rect 6190 46450 6242 46462
rect 6190 46386 6242 46398
rect 10446 46450 10498 46462
rect 16046 46450 16098 46462
rect 11554 46398 11566 46450
rect 11618 46398 11630 46450
rect 14018 46398 14030 46450
rect 14082 46398 14094 46450
rect 10446 46386 10498 46398
rect 16046 46386 16098 46398
rect 16606 46450 16658 46462
rect 16606 46386 16658 46398
rect 23214 46450 23266 46462
rect 23214 46386 23266 46398
rect 672 46282 31024 46316
rect 672 46230 4466 46282
rect 4518 46230 4570 46282
rect 4622 46230 4674 46282
rect 4726 46230 24466 46282
rect 24518 46230 24570 46282
rect 24622 46230 24674 46282
rect 24726 46230 31024 46282
rect 672 46196 31024 46230
rect 9662 46114 9714 46126
rect 9662 46050 9714 46062
rect 17838 46114 17890 46126
rect 22642 46062 22654 46114
rect 22706 46062 22718 46114
rect 17838 46050 17890 46062
rect 1586 45950 1598 46002
rect 1650 45950 1662 46002
rect 4834 45950 4846 46002
rect 4898 45950 4910 46002
rect 7074 45950 7086 46002
rect 7138 45950 7150 46002
rect 11330 45950 11342 46002
rect 11394 45950 11406 46002
rect 18834 45950 18846 46002
rect 18898 45950 18910 46002
rect 20066 45950 20078 46002
rect 20130 45950 20142 46002
rect 30594 45950 30606 46002
rect 30658 45950 30670 46002
rect 8206 45890 8258 45902
rect 6514 45838 6526 45890
rect 6578 45838 6590 45890
rect 8206 45826 8258 45838
rect 8878 45890 8930 45902
rect 12014 45890 12066 45902
rect 22318 45890 22370 45902
rect 9090 45838 9102 45890
rect 9154 45838 9166 45890
rect 9650 45838 9662 45890
rect 9714 45838 9726 45890
rect 10658 45838 10670 45890
rect 10722 45838 10734 45890
rect 11106 45838 11118 45890
rect 11170 45838 11182 45890
rect 12338 45838 12350 45890
rect 12402 45838 12414 45890
rect 13346 45838 13358 45890
rect 13410 45838 13422 45890
rect 18946 45838 18958 45890
rect 19010 45838 19022 45890
rect 8878 45826 8930 45838
rect 12014 45826 12066 45838
rect 22318 45826 22370 45838
rect 30270 45890 30322 45902
rect 30270 45826 30322 45838
rect 10334 45778 10386 45790
rect 1250 45726 1262 45778
rect 1314 45726 1326 45778
rect 4386 45726 4398 45778
rect 4450 45726 4462 45778
rect 6626 45726 6638 45778
rect 6690 45726 6702 45778
rect 19730 45726 19742 45778
rect 19794 45726 19806 45778
rect 10334 45714 10386 45726
rect 2830 45666 2882 45678
rect 2830 45602 2882 45614
rect 5966 45666 6018 45678
rect 18174 45666 18226 45678
rect 9426 45614 9438 45666
rect 9490 45614 9502 45666
rect 5966 45602 6018 45614
rect 18174 45602 18226 45614
rect 21310 45666 21362 45678
rect 21310 45602 21362 45614
rect 672 45498 31024 45532
rect 672 45446 3806 45498
rect 3858 45446 3910 45498
rect 3962 45446 4014 45498
rect 4066 45446 23806 45498
rect 23858 45446 23910 45498
rect 23962 45446 24014 45498
rect 24066 45446 31024 45498
rect 672 45412 31024 45446
rect 12126 45330 12178 45342
rect 12126 45266 12178 45278
rect 18958 45330 19010 45342
rect 18958 45266 19010 45278
rect 9774 45218 9826 45230
rect 13458 45166 13470 45218
rect 13522 45166 13534 45218
rect 9774 45154 9826 45166
rect 5854 45106 5906 45118
rect 7534 45106 7586 45118
rect 1250 45054 1262 45106
rect 1314 45054 1326 45106
rect 6514 45054 6526 45106
rect 6578 45054 6590 45106
rect 6850 45054 6862 45106
rect 6914 45054 6926 45106
rect 8194 45054 8206 45106
rect 8258 45054 8270 45106
rect 9202 45054 9214 45106
rect 9266 45054 9278 45106
rect 10434 45054 10446 45106
rect 10498 45054 10510 45106
rect 17378 45054 17390 45106
rect 17442 45054 17454 45106
rect 5854 45042 5906 45054
rect 7534 45042 7586 45054
rect 5518 44994 5570 45006
rect 5518 44930 5570 44942
rect 6078 44994 6130 45006
rect 9662 44994 9714 45006
rect 7074 44942 7086 44994
rect 7138 44942 7150 44994
rect 13794 44942 13806 44994
rect 13858 44942 13870 44994
rect 17826 44942 17838 44994
rect 17890 44942 17902 44994
rect 29810 44942 29822 44994
rect 29874 44942 29886 44994
rect 6078 44930 6130 44942
rect 9662 44930 9714 44942
rect 2830 44882 2882 44894
rect 1698 44830 1710 44882
rect 1762 44830 1774 44882
rect 2830 44818 2882 44830
rect 5630 44882 5682 44894
rect 5630 44818 5682 44830
rect 9886 44882 9938 44894
rect 15038 44882 15090 44894
rect 10994 44830 11006 44882
rect 11058 44830 11070 44882
rect 9886 44818 9938 44830
rect 15038 44818 15090 44830
rect 29486 44882 29538 44894
rect 29486 44818 29538 44830
rect 30270 44882 30322 44894
rect 30594 44830 30606 44882
rect 30658 44830 30670 44882
rect 30270 44818 30322 44830
rect 672 44714 31024 44748
rect 672 44662 4466 44714
rect 4518 44662 4570 44714
rect 4622 44662 4674 44714
rect 4726 44662 24466 44714
rect 24518 44662 24570 44714
rect 24622 44662 24674 44714
rect 24726 44662 31024 44714
rect 672 44628 31024 44662
rect 8206 44546 8258 44558
rect 2930 44494 2942 44546
rect 2994 44494 3006 44546
rect 10882 44494 10894 44546
rect 10946 44494 10958 44546
rect 14802 44494 14814 44546
rect 14866 44494 14878 44546
rect 19842 44494 19854 44546
rect 19906 44494 19918 44546
rect 22642 44494 22654 44546
rect 22706 44494 22718 44546
rect 29810 44494 29822 44546
rect 29874 44494 29886 44546
rect 8206 44482 8258 44494
rect 3390 44434 3442 44446
rect 9438 44434 9490 44446
rect 7074 44382 7086 44434
rect 7138 44382 7150 44434
rect 3390 44370 3442 44382
rect 9438 44370 9490 44382
rect 9886 44434 9938 44446
rect 17266 44382 17278 44434
rect 17330 44382 17342 44434
rect 9886 44370 9938 44382
rect 8990 44322 9042 44334
rect 2370 44270 2382 44322
rect 2434 44270 2446 44322
rect 2818 44270 2830 44322
rect 2882 44270 2894 44322
rect 4162 44270 4174 44322
rect 4226 44270 4238 44322
rect 4946 44270 4958 44322
rect 5010 44270 5022 44322
rect 6626 44270 6638 44322
rect 6690 44270 6702 44322
rect 8990 44258 9042 44270
rect 9102 44322 9154 44334
rect 11566 44322 11618 44334
rect 10210 44270 10222 44322
rect 10274 44270 10286 44322
rect 10770 44270 10782 44322
rect 10834 44270 10846 44322
rect 11890 44270 11902 44322
rect 11954 44270 11966 44322
rect 13010 44270 13022 44322
rect 13074 44270 13086 44322
rect 14354 44270 14366 44322
rect 14418 44270 14430 44322
rect 16818 44270 16830 44322
rect 16882 44270 16894 44322
rect 19282 44270 19294 44322
rect 19346 44270 19358 44322
rect 29586 44270 29598 44322
rect 29650 44270 29662 44322
rect 9102 44258 9154 44270
rect 11566 44258 11618 44270
rect 1934 44210 1986 44222
rect 19394 44158 19406 44210
rect 19458 44158 19470 44210
rect 23090 44158 23102 44210
rect 23154 44158 23166 44210
rect 1934 44146 1986 44158
rect 9326 44098 9378 44110
rect 9326 44034 9378 44046
rect 15934 44098 15986 44110
rect 15934 44034 15986 44046
rect 18510 44098 18562 44110
rect 18510 44034 18562 44046
rect 20974 44098 21026 44110
rect 20974 44034 21026 44046
rect 21534 44098 21586 44110
rect 21534 44034 21586 44046
rect 672 43930 31024 43964
rect 672 43878 3806 43930
rect 3858 43878 3910 43930
rect 3962 43878 4014 43930
rect 4066 43878 23806 43930
rect 23858 43878 23910 43930
rect 23962 43878 24014 43930
rect 24066 43878 31024 43930
rect 672 43844 31024 43878
rect 11566 43762 11618 43774
rect 11566 43698 11618 43710
rect 6862 43650 6914 43662
rect 5282 43598 5294 43650
rect 5346 43598 5358 43650
rect 6862 43586 6914 43598
rect 9326 43650 9378 43662
rect 9326 43586 9378 43598
rect 2606 43538 2658 43550
rect 15710 43538 15762 43550
rect 22094 43538 22146 43550
rect 1586 43486 1598 43538
rect 1650 43486 1662 43538
rect 2034 43486 2046 43538
rect 2098 43486 2110 43538
rect 3154 43486 3166 43538
rect 3218 43486 3230 43538
rect 4162 43486 4174 43538
rect 4226 43486 4238 43538
rect 7746 43486 7758 43538
rect 7810 43486 7822 43538
rect 9986 43486 9998 43538
rect 10050 43486 10062 43538
rect 14466 43486 14478 43538
rect 14530 43486 14542 43538
rect 14802 43486 14814 43538
rect 14866 43486 14878 43538
rect 16034 43486 16046 43538
rect 16098 43486 16110 43538
rect 17154 43486 17166 43538
rect 17218 43486 17230 43538
rect 17714 43486 17726 43538
rect 17778 43486 17790 43538
rect 20962 43486 20974 43538
rect 21026 43486 21038 43538
rect 21410 43486 21422 43538
rect 21474 43486 21486 43538
rect 22642 43486 22654 43538
rect 22706 43486 22718 43538
rect 23650 43486 23662 43538
rect 23714 43486 23726 43538
rect 2606 43474 2658 43486
rect 15710 43474 15762 43486
rect 22094 43474 22146 43486
rect 1150 43426 1202 43438
rect 14030 43426 14082 43438
rect 20638 43426 20690 43438
rect 2146 43374 2158 43426
rect 2210 43374 2222 43426
rect 8194 43374 8206 43426
rect 8258 43374 8270 43426
rect 10322 43374 10334 43426
rect 10386 43374 10398 43426
rect 18274 43374 18286 43426
rect 18338 43374 18350 43426
rect 21634 43374 21646 43426
rect 21698 43374 21710 43426
rect 1150 43362 1202 43374
rect 14030 43362 14082 43374
rect 20638 43362 20690 43374
rect 19406 43314 19458 43326
rect 5730 43262 5742 43314
rect 5794 43262 5806 43314
rect 15026 43262 15038 43314
rect 15090 43262 15102 43314
rect 19406 43250 19458 43262
rect 29486 43314 29538 43326
rect 30270 43314 30322 43326
rect 29810 43262 29822 43314
rect 29874 43262 29886 43314
rect 30594 43262 30606 43314
rect 30658 43262 30670 43314
rect 29486 43250 29538 43262
rect 30270 43250 30322 43262
rect 672 43146 31024 43180
rect 672 43094 4466 43146
rect 4518 43094 4570 43146
rect 4622 43094 4674 43146
rect 4726 43094 24466 43146
rect 24518 43094 24570 43146
rect 24622 43094 24674 43146
rect 24726 43094 31024 43146
rect 672 43060 31024 43094
rect 6178 42926 6190 42978
rect 6242 42926 6254 42978
rect 15138 42926 15150 42978
rect 15202 42926 15214 42978
rect 18834 42926 18846 42978
rect 18898 42926 18910 42978
rect 9326 42866 9378 42878
rect 2930 42814 2942 42866
rect 2994 42814 3006 42866
rect 10322 42814 10334 42866
rect 10386 42814 10398 42866
rect 22754 42814 22766 42866
rect 22818 42814 22830 42866
rect 30594 42814 30606 42866
rect 30658 42814 30670 42866
rect 9326 42802 9378 42814
rect 3390 42754 3442 42766
rect 10782 42754 10834 42766
rect 14478 42754 14530 42766
rect 30270 42754 30322 42766
rect 2370 42702 2382 42754
rect 2434 42702 2446 42754
rect 2818 42702 2830 42754
rect 2882 42702 2894 42754
rect 4050 42702 4062 42754
rect 4114 42702 4126 42754
rect 4946 42702 4958 42754
rect 5010 42702 5022 42754
rect 5730 42702 5742 42754
rect 5794 42702 5806 42754
rect 9650 42702 9662 42754
rect 9714 42702 9726 42754
rect 10098 42702 10110 42754
rect 10162 42702 10174 42754
rect 11442 42702 11454 42754
rect 11506 42702 11518 42754
rect 12338 42702 12350 42754
rect 12402 42702 12414 42754
rect 13122 42702 13134 42754
rect 13186 42702 13198 42754
rect 13906 42702 13918 42754
rect 13970 42702 13982 42754
rect 15250 42702 15262 42754
rect 15314 42702 15326 42754
rect 15698 42702 15710 42754
rect 15762 42702 15774 42754
rect 18274 42702 18286 42754
rect 18338 42702 18350 42754
rect 18610 42702 18622 42754
rect 18674 42702 18686 42754
rect 19394 42702 19406 42754
rect 19458 42702 19470 42754
rect 19842 42702 19854 42754
rect 19906 42702 19918 42754
rect 20850 42702 20862 42754
rect 20914 42702 20926 42754
rect 23202 42702 23214 42754
rect 23266 42702 23278 42754
rect 3390 42690 3442 42702
rect 10782 42690 10834 42702
rect 14478 42690 14530 42702
rect 30270 42690 30322 42702
rect 1934 42642 1986 42654
rect 1934 42578 1986 42590
rect 16158 42642 16210 42654
rect 16158 42578 16210 42590
rect 17838 42642 17890 42654
rect 17838 42578 17890 42590
rect 7310 42530 7362 42542
rect 7310 42466 7362 42478
rect 21534 42530 21586 42542
rect 21534 42466 21586 42478
rect 672 42362 31024 42396
rect 672 42310 3806 42362
rect 3858 42310 3910 42362
rect 3962 42310 4014 42362
rect 4066 42310 23806 42362
rect 23858 42310 23910 42362
rect 23962 42310 24014 42362
rect 24066 42310 31024 42362
rect 672 42276 31024 42310
rect 10334 42194 10386 42206
rect 10334 42130 10386 42142
rect 13806 42194 13858 42206
rect 13806 42130 13858 42142
rect 8990 42082 9042 42094
rect 11890 42030 11902 42082
rect 11954 42030 11966 42082
rect 15362 42030 15374 42082
rect 15426 42030 15438 42082
rect 16482 42030 16494 42082
rect 16546 42030 16558 42082
rect 8990 42018 9042 42030
rect 4958 41970 5010 41982
rect 8654 41970 8706 41982
rect 1586 41918 1598 41970
rect 1650 41918 1662 41970
rect 1922 41918 1934 41970
rect 1986 41918 1998 41970
rect 2706 41918 2718 41970
rect 2770 41918 2782 41970
rect 3154 41918 3166 41970
rect 3218 41918 3230 41970
rect 4162 41918 4174 41970
rect 4226 41918 4238 41970
rect 5282 41918 5294 41970
rect 5346 41918 5358 41970
rect 5730 41918 5742 41970
rect 5794 41918 5806 41970
rect 6514 41918 6526 41970
rect 6578 41918 6590 41970
rect 7186 41918 7198 41970
rect 7250 41918 7262 41970
rect 7970 41918 7982 41970
rect 8034 41918 8046 41970
rect 4958 41906 5010 41918
rect 8654 41906 8706 41918
rect 19630 41970 19682 41982
rect 19630 41906 19682 41918
rect 20638 41970 20690 41982
rect 20962 41918 20974 41970
rect 21026 41918 21038 41970
rect 21410 41918 21422 41970
rect 21474 41918 21486 41970
rect 22642 41918 22654 41970
rect 22706 41918 22718 41970
rect 23650 41918 23662 41970
rect 23714 41918 23726 41970
rect 20638 41906 20690 41918
rect 1150 41858 1202 41870
rect 22094 41858 22146 41870
rect 9202 41806 9214 41858
rect 9266 41806 9278 41858
rect 9538 41806 9550 41858
rect 9602 41806 9614 41858
rect 11442 41806 11454 41858
rect 11506 41806 11518 41858
rect 15026 41806 15038 41858
rect 15090 41806 15102 41858
rect 16930 41806 16942 41858
rect 16994 41806 17006 41858
rect 18946 41806 18958 41858
rect 19010 41806 19022 41858
rect 19282 41806 19294 41858
rect 19346 41806 19358 41858
rect 21634 41806 21646 41858
rect 21698 41806 21710 41858
rect 29810 41806 29822 41858
rect 29874 41806 29886 41858
rect 1150 41794 1202 41806
rect 22094 41794 22146 41806
rect 18062 41746 18114 41758
rect 2146 41694 2158 41746
rect 2210 41694 2222 41746
rect 5954 41694 5966 41746
rect 6018 41694 6030 41746
rect 18062 41682 18114 41694
rect 19966 41746 20018 41758
rect 19966 41682 20018 41694
rect 29486 41746 29538 41758
rect 29486 41682 29538 41694
rect 672 41578 31024 41612
rect 672 41526 4466 41578
rect 4518 41526 4570 41578
rect 4622 41526 4674 41578
rect 4726 41526 24466 41578
rect 24518 41526 24570 41578
rect 24622 41526 24674 41578
rect 24726 41526 31024 41578
rect 672 41492 31024 41526
rect 4398 41410 4450 41422
rect 21758 41410 21810 41422
rect 3266 41358 3278 41410
rect 3330 41358 3342 41410
rect 5842 41358 5854 41410
rect 5906 41358 5918 41410
rect 10994 41358 11006 41410
rect 11058 41358 11070 41410
rect 19058 41358 19070 41410
rect 19122 41358 19134 41410
rect 22866 41358 22878 41410
rect 22930 41358 22942 41410
rect 4398 41346 4450 41358
rect 21758 41346 21810 41358
rect 19518 41298 19570 41310
rect 30270 41298 30322 41310
rect 14802 41246 14814 41298
rect 14866 41246 14878 41298
rect 29810 41246 29822 41298
rect 29874 41246 29886 41298
rect 30594 41246 30606 41298
rect 30658 41246 30670 41298
rect 19518 41234 19570 41246
rect 30270 41234 30322 41246
rect 4846 41186 4898 41198
rect 6526 41186 6578 41198
rect 11454 41186 11506 41198
rect 29486 41186 29538 41198
rect 5282 41134 5294 41186
rect 5346 41134 5358 41186
rect 5618 41134 5630 41186
rect 5682 41134 5694 41186
rect 7074 41134 7086 41186
rect 7138 41134 7150 41186
rect 7858 41134 7870 41186
rect 7922 41134 7934 41186
rect 10322 41134 10334 41186
rect 10386 41134 10398 41186
rect 10770 41134 10782 41186
rect 10834 41134 10846 41186
rect 12002 41134 12014 41186
rect 12066 41134 12078 41186
rect 12226 41134 12238 41186
rect 12290 41134 12302 41186
rect 13010 41134 13022 41186
rect 13074 41134 13086 41186
rect 14466 41134 14478 41186
rect 14530 41134 14542 41186
rect 18498 41134 18510 41186
rect 18562 41134 18574 41186
rect 18834 41134 18846 41186
rect 18898 41134 18910 41186
rect 20178 41134 20190 41186
rect 20242 41134 20254 41186
rect 21074 41134 21086 41186
rect 21138 41134 21150 41186
rect 23314 41134 23326 41186
rect 23378 41134 23390 41186
rect 4846 41122 4898 41134
rect 6526 41122 6578 41134
rect 11454 41122 11506 41134
rect 29486 41122 29538 41134
rect 9998 41074 10050 41086
rect 2818 41022 2830 41074
rect 2882 41022 2894 41074
rect 9998 41010 10050 41022
rect 18062 41074 18114 41086
rect 18062 41010 18114 41022
rect 16046 40962 16098 40974
rect 16046 40898 16098 40910
rect 672 40794 31024 40828
rect 672 40742 3806 40794
rect 3858 40742 3910 40794
rect 3962 40742 4014 40794
rect 4066 40742 23806 40794
rect 23858 40742 23910 40794
rect 23962 40742 24014 40794
rect 24066 40742 31024 40794
rect 672 40708 31024 40742
rect 5854 40626 5906 40638
rect 5854 40562 5906 40574
rect 8430 40626 8482 40638
rect 8430 40562 8482 40574
rect 8990 40626 9042 40638
rect 8990 40562 9042 40574
rect 14590 40626 14642 40638
rect 14590 40562 14642 40574
rect 20638 40514 20690 40526
rect 1698 40462 1710 40514
rect 1762 40462 1774 40514
rect 6850 40462 6862 40514
rect 6914 40462 6926 40514
rect 10546 40462 10558 40514
rect 10610 40462 10622 40514
rect 13010 40462 13022 40514
rect 13074 40462 13086 40514
rect 20638 40450 20690 40462
rect 3278 40402 3330 40414
rect 17838 40402 17890 40414
rect 30270 40402 30322 40414
rect 5170 40350 5182 40402
rect 5234 40350 5246 40402
rect 16482 40350 16494 40402
rect 16546 40350 16558 40402
rect 16930 40350 16942 40402
rect 16994 40350 17006 40402
rect 18162 40350 18174 40402
rect 18226 40350 18238 40402
rect 19170 40350 19182 40402
rect 19234 40350 19246 40402
rect 20962 40350 20974 40402
rect 21026 40350 21038 40402
rect 21522 40350 21534 40402
rect 21586 40350 21598 40402
rect 22194 40350 22206 40402
rect 22258 40350 22270 40402
rect 22754 40350 22766 40402
rect 22818 40350 22830 40402
rect 23650 40350 23662 40402
rect 23714 40350 23726 40402
rect 3278 40338 3330 40350
rect 17838 40338 17890 40350
rect 30270 40338 30322 40350
rect 16158 40290 16210 40302
rect 2034 40238 2046 40290
rect 2098 40238 2110 40290
rect 5058 40238 5070 40290
rect 5122 40238 5134 40290
rect 10098 40238 10110 40290
rect 10162 40238 10174 40290
rect 13458 40238 13470 40290
rect 13522 40238 13534 40290
rect 17154 40238 17166 40290
rect 17218 40238 17230 40290
rect 21634 40238 21646 40290
rect 21698 40238 21710 40290
rect 29810 40238 29822 40290
rect 29874 40238 29886 40290
rect 16158 40226 16210 40238
rect 6190 40178 6242 40190
rect 29486 40178 29538 40190
rect 7298 40126 7310 40178
rect 7362 40126 7374 40178
rect 30594 40126 30606 40178
rect 30658 40126 30670 40178
rect 6190 40114 6242 40126
rect 29486 40114 29538 40126
rect 672 40010 31024 40044
rect 672 39958 4466 40010
rect 4518 39958 4570 40010
rect 4622 39958 4674 40010
rect 4726 39958 24466 40010
rect 24518 39958 24570 40010
rect 24622 39958 24674 40010
rect 24726 39958 31024 40010
rect 672 39924 31024 39958
rect 2830 39842 2882 39854
rect 2830 39778 2882 39790
rect 6526 39842 6578 39854
rect 6526 39778 6578 39790
rect 10894 39730 10946 39742
rect 1586 39678 1598 39730
rect 1650 39678 1662 39730
rect 5394 39678 5406 39730
rect 5458 39678 5470 39730
rect 7074 39678 7086 39730
rect 7138 39678 7150 39730
rect 7634 39678 7646 39730
rect 7698 39678 7710 39730
rect 11890 39678 11902 39730
rect 11954 39678 11966 39730
rect 10894 39666 10946 39678
rect 12350 39618 12402 39630
rect 4946 39566 4958 39618
rect 5010 39566 5022 39618
rect 11218 39566 11230 39618
rect 11282 39566 11294 39618
rect 11666 39566 11678 39618
rect 11730 39566 11742 39618
rect 12898 39566 12910 39618
rect 12962 39566 12974 39618
rect 13906 39566 13918 39618
rect 13970 39566 13982 39618
rect 12350 39554 12402 39566
rect 1250 39454 1262 39506
rect 1314 39454 1326 39506
rect 7870 39394 7922 39406
rect 7870 39330 7922 39342
rect 8206 39394 8258 39406
rect 8206 39330 8258 39342
rect 672 39226 31024 39260
rect 672 39174 3806 39226
rect 3858 39174 3910 39226
rect 3962 39174 4014 39226
rect 4066 39174 23806 39226
rect 23858 39174 23910 39226
rect 23962 39174 24014 39226
rect 24066 39174 31024 39226
rect 672 39140 31024 39174
rect 2830 39058 2882 39070
rect 2830 38994 2882 39006
rect 9886 39058 9938 39070
rect 9886 38994 9938 39006
rect 12126 39058 12178 39070
rect 12126 38994 12178 39006
rect 1250 38894 1262 38946
rect 1314 38894 1326 38946
rect 8306 38894 8318 38946
rect 8370 38894 8382 38946
rect 10546 38894 10558 38946
rect 10610 38894 10622 38946
rect 15374 38834 15426 38846
rect 5506 38782 5518 38834
rect 5570 38782 5582 38834
rect 14018 38782 14030 38834
rect 14082 38782 14094 38834
rect 14466 38782 14478 38834
rect 14530 38782 14542 38834
rect 15698 38782 15710 38834
rect 15762 38782 15774 38834
rect 16706 38782 16718 38834
rect 16770 38782 16782 38834
rect 20850 38782 20862 38834
rect 20914 38782 20926 38834
rect 15374 38770 15426 38782
rect 13694 38722 13746 38734
rect 1586 38670 1598 38722
rect 1650 38670 1662 38722
rect 6066 38670 6078 38722
rect 6130 38670 6142 38722
rect 8754 38670 8766 38722
rect 8818 38670 8830 38722
rect 10882 38670 10894 38722
rect 10946 38670 10958 38722
rect 14690 38670 14702 38722
rect 14754 38670 14766 38722
rect 21410 38670 21422 38722
rect 21474 38670 21486 38722
rect 13694 38658 13746 38670
rect 7198 38610 7250 38622
rect 7198 38546 7250 38558
rect 22542 38610 22594 38622
rect 22542 38546 22594 38558
rect 672 38442 31024 38476
rect 672 38390 4466 38442
rect 4518 38390 4570 38442
rect 4622 38390 4674 38442
rect 4726 38390 24466 38442
rect 24518 38390 24570 38442
rect 24622 38390 24674 38442
rect 24726 38390 31024 38442
rect 672 38356 31024 38390
rect 11006 38274 11058 38286
rect 13246 38274 13298 38286
rect 6066 38222 6078 38274
rect 6130 38222 6142 38274
rect 9874 38222 9886 38274
rect 9938 38222 9950 38274
rect 12114 38222 12126 38274
rect 12178 38222 12190 38274
rect 11006 38210 11058 38222
rect 13246 38210 13298 38222
rect 15486 38274 15538 38286
rect 15486 38210 15538 38222
rect 18622 38274 18674 38286
rect 18622 38210 18674 38222
rect 20078 38162 20130 38174
rect 1922 38110 1934 38162
rect 1986 38110 1998 38162
rect 14242 38110 14254 38162
rect 14306 38110 14318 38162
rect 21298 38110 21310 38162
rect 21362 38110 21374 38162
rect 20078 38098 20130 38110
rect 18734 38050 18786 38062
rect 1362 37998 1374 38050
rect 1426 37998 1438 38050
rect 18734 37986 18786 37998
rect 19518 38050 19570 38062
rect 19842 37998 19854 38050
rect 19906 37998 19918 38050
rect 19518 37986 19570 37998
rect 19182 37938 19234 37950
rect 1474 37886 1486 37938
rect 1538 37886 1550 37938
rect 5618 37886 5630 37938
rect 5682 37886 5694 37938
rect 9426 37886 9438 37938
rect 9490 37886 9502 37938
rect 11666 37886 11678 37938
rect 11730 37886 11742 37938
rect 13906 37886 13918 37938
rect 13970 37886 13982 37938
rect 20066 37886 20078 37938
rect 20130 37886 20142 37938
rect 20850 37886 20862 37938
rect 20914 37886 20926 37938
rect 19182 37874 19234 37886
rect 3054 37826 3106 37838
rect 3054 37762 3106 37774
rect 7198 37826 7250 37838
rect 7198 37762 7250 37774
rect 18622 37826 18674 37838
rect 18622 37762 18674 37774
rect 19070 37826 19122 37838
rect 19070 37762 19122 37774
rect 22430 37826 22482 37838
rect 22430 37762 22482 37774
rect 672 37658 31024 37692
rect 672 37606 3806 37658
rect 3858 37606 3910 37658
rect 3962 37606 4014 37658
rect 4066 37606 23806 37658
rect 23858 37606 23910 37658
rect 23962 37606 24014 37658
rect 24066 37606 31024 37658
rect 672 37572 31024 37606
rect 2706 37326 2718 37378
rect 2770 37326 2782 37378
rect 15934 37266 15986 37278
rect 1922 37214 1934 37266
rect 1986 37214 1998 37266
rect 6850 37214 6862 37266
rect 6914 37214 6926 37266
rect 7186 37214 7198 37266
rect 7250 37214 7262 37266
rect 8642 37214 8654 37266
rect 8706 37214 8718 37266
rect 9426 37214 9438 37266
rect 9490 37214 9502 37266
rect 10098 37214 10110 37266
rect 10162 37214 10174 37266
rect 14690 37214 14702 37266
rect 14754 37214 14766 37266
rect 15026 37214 15038 37266
rect 15090 37214 15102 37266
rect 16258 37214 16270 37266
rect 16322 37214 16334 37266
rect 17266 37214 17278 37266
rect 17330 37214 17342 37266
rect 18050 37214 18062 37266
rect 18114 37214 18126 37266
rect 20850 37214 20862 37266
rect 20914 37214 20926 37266
rect 15934 37202 15986 37214
rect 6414 37154 6466 37166
rect 7870 37154 7922 37166
rect 7410 37102 7422 37154
rect 7474 37102 7486 37154
rect 6414 37090 6466 37102
rect 7870 37090 7922 37102
rect 14254 37154 14306 37166
rect 18386 37102 18398 37154
rect 18450 37102 18462 37154
rect 14254 37090 14306 37102
rect 4286 37042 4338 37054
rect 11790 37042 11842 37054
rect 19630 37042 19682 37054
rect 22542 37042 22594 37054
rect 2146 36990 2158 37042
rect 2210 36990 2222 37042
rect 3154 36990 3166 37042
rect 3218 36990 3230 37042
rect 10658 36990 10670 37042
rect 10722 36990 10734 37042
rect 15250 36990 15262 37042
rect 15314 36990 15326 37042
rect 21410 36990 21422 37042
rect 21474 36990 21486 37042
rect 4286 36978 4338 36990
rect 11790 36978 11842 36990
rect 19630 36978 19682 36990
rect 22542 36978 22594 36990
rect 672 36874 31024 36908
rect 672 36822 4466 36874
rect 4518 36822 4570 36874
rect 4622 36822 4674 36874
rect 4726 36822 24466 36874
rect 24518 36822 24570 36874
rect 24622 36822 24674 36874
rect 24726 36822 31024 36874
rect 672 36788 31024 36822
rect 16046 36706 16098 36718
rect 23662 36706 23714 36718
rect 2482 36654 2494 36706
rect 2546 36654 2558 36706
rect 17938 36654 17950 36706
rect 18002 36654 18014 36706
rect 16046 36642 16098 36654
rect 23662 36642 23714 36654
rect 11790 36594 11842 36606
rect 7298 36542 7310 36594
rect 7362 36542 7374 36594
rect 11330 36542 11342 36594
rect 11394 36542 11406 36594
rect 14802 36542 14814 36594
rect 14866 36542 14878 36594
rect 19618 36542 19630 36594
rect 19682 36542 19694 36594
rect 19954 36542 19966 36594
rect 20018 36542 20030 36594
rect 21298 36542 21310 36594
rect 21362 36542 21374 36594
rect 23986 36542 23998 36594
rect 24050 36542 24062 36594
rect 11790 36530 11842 36542
rect 1486 36482 1538 36494
rect 2942 36482 2994 36494
rect 8318 36482 8370 36494
rect 1810 36430 1822 36482
rect 1874 36430 1886 36482
rect 2258 36430 2270 36482
rect 2322 36430 2334 36482
rect 3490 36430 3502 36482
rect 3554 36430 3566 36482
rect 3714 36430 3726 36482
rect 3778 36430 3790 36482
rect 4498 36430 4510 36482
rect 4562 36430 4574 36482
rect 5170 36430 5182 36482
rect 5234 36430 5246 36482
rect 6066 36430 6078 36482
rect 6130 36430 6142 36482
rect 6738 36430 6750 36482
rect 6802 36430 6814 36482
rect 7522 36430 7534 36482
rect 7586 36430 7598 36482
rect 7858 36430 7870 36482
rect 7922 36430 7934 36482
rect 1486 36418 1538 36430
rect 2942 36418 2994 36430
rect 8318 36418 8370 36430
rect 10334 36482 10386 36494
rect 10658 36430 10670 36482
rect 10722 36430 10734 36482
rect 11106 36430 11118 36482
rect 11170 36430 11182 36482
rect 12338 36430 12350 36482
rect 12402 36430 12414 36482
rect 13346 36430 13358 36482
rect 13410 36430 13422 36482
rect 14354 36430 14366 36482
rect 14418 36430 14430 36482
rect 20850 36430 20862 36482
rect 20914 36430 20926 36482
rect 10334 36418 10386 36430
rect 18386 36318 18398 36370
rect 18450 36318 18462 36370
rect 16830 36258 16882 36270
rect 16830 36194 16882 36206
rect 19070 36258 19122 36270
rect 19070 36194 19122 36206
rect 19406 36258 19458 36270
rect 19406 36194 19458 36206
rect 22542 36258 22594 36270
rect 22542 36194 22594 36206
rect 672 36090 31024 36124
rect 672 36038 3806 36090
rect 3858 36038 3910 36090
rect 3962 36038 4014 36090
rect 4066 36038 23806 36090
rect 23858 36038 23910 36090
rect 23962 36038 24014 36090
rect 24066 36038 31024 36090
rect 672 36004 31024 36038
rect 15038 35922 15090 35934
rect 19294 35922 19346 35934
rect 16930 35870 16942 35922
rect 16994 35870 17006 35922
rect 15038 35858 15090 35870
rect 19294 35858 19346 35870
rect 1150 35810 1202 35822
rect 1150 35746 1202 35758
rect 12238 35810 12290 35822
rect 12238 35746 12290 35758
rect 20974 35810 21026 35822
rect 20974 35746 21026 35758
rect 6862 35698 6914 35710
rect 10558 35698 10610 35710
rect 16382 35698 16434 35710
rect 30270 35698 30322 35710
rect 1474 35646 1486 35698
rect 1538 35646 1550 35698
rect 2034 35646 2046 35698
rect 2098 35646 2110 35698
rect 2706 35646 2718 35698
rect 2770 35646 2782 35698
rect 3266 35646 3278 35698
rect 3330 35646 3342 35698
rect 4162 35646 4174 35698
rect 4226 35646 4238 35698
rect 5730 35646 5742 35698
rect 5794 35646 5806 35698
rect 6178 35646 6190 35698
rect 6242 35646 6254 35698
rect 7410 35646 7422 35698
rect 7474 35646 7486 35698
rect 8418 35646 8430 35698
rect 8482 35646 8494 35698
rect 9202 35646 9214 35698
rect 9266 35646 9278 35698
rect 10210 35646 10222 35698
rect 10274 35646 10286 35698
rect 11330 35646 11342 35698
rect 11394 35646 11406 35698
rect 11778 35646 11790 35698
rect 11842 35646 11854 35698
rect 13458 35646 13470 35698
rect 13522 35646 13534 35698
rect 17154 35646 17166 35698
rect 17218 35646 17230 35698
rect 17714 35646 17726 35698
rect 17778 35646 17790 35698
rect 21410 35646 21422 35698
rect 21474 35646 21486 35698
rect 21746 35646 21758 35698
rect 21810 35646 21822 35698
rect 22530 35646 22542 35698
rect 22594 35646 22606 35698
rect 22978 35646 22990 35698
rect 23042 35646 23054 35698
rect 24098 35646 24110 35698
rect 24162 35646 24174 35698
rect 6862 35634 6914 35646
rect 10558 35634 10610 35646
rect 16382 35634 16434 35646
rect 30270 35634 30322 35646
rect 5406 35586 5458 35598
rect 16046 35586 16098 35598
rect 19742 35586 19794 35598
rect 6402 35534 6414 35586
rect 6466 35534 6478 35586
rect 16594 35534 16606 35586
rect 16658 35534 16670 35586
rect 18050 35534 18062 35586
rect 18114 35534 18126 35586
rect 5406 35522 5458 35534
rect 16046 35522 16098 35534
rect 19742 35522 19794 35534
rect 15710 35474 15762 35486
rect 2146 35422 2158 35474
rect 2210 35422 2222 35474
rect 11218 35422 11230 35474
rect 11282 35422 11294 35474
rect 13906 35422 13918 35474
rect 13970 35422 13982 35474
rect 15710 35410 15762 35422
rect 15934 35474 15986 35486
rect 15934 35410 15986 35422
rect 17166 35474 17218 35486
rect 17166 35410 17218 35422
rect 19854 35474 19906 35486
rect 19854 35410 19906 35422
rect 19966 35474 20018 35486
rect 21970 35422 21982 35474
rect 22034 35422 22046 35474
rect 30594 35422 30606 35474
rect 30658 35422 30670 35474
rect 19966 35410 20018 35422
rect 672 35306 31024 35340
rect 672 35254 4466 35306
rect 4518 35254 4570 35306
rect 4622 35254 4674 35306
rect 4726 35254 24466 35306
rect 24518 35254 24570 35306
rect 24622 35254 24674 35306
rect 24726 35254 31024 35306
rect 672 35220 31024 35254
rect 20302 35138 20354 35150
rect 30270 35138 30322 35150
rect 3714 35086 3726 35138
rect 3778 35086 3790 35138
rect 13906 35086 13918 35138
rect 13970 35086 13982 35138
rect 21746 35086 21758 35138
rect 21810 35086 21822 35138
rect 20302 35074 20354 35086
rect 30270 35074 30322 35086
rect 6526 35026 6578 35038
rect 12462 35026 12514 35038
rect 6066 34974 6078 35026
rect 6130 34974 6142 35026
rect 9090 34974 9102 35026
rect 9154 34974 9166 35026
rect 11330 34974 11342 35026
rect 11394 34974 11406 35026
rect 6526 34962 6578 34974
rect 12462 34962 12514 34974
rect 17502 35026 17554 35038
rect 20750 35026 20802 35038
rect 17826 34974 17838 35026
rect 17890 34974 17902 35026
rect 19170 34974 19182 35026
rect 19234 34974 19246 35026
rect 24770 34974 24782 35026
rect 24834 34974 24846 35026
rect 30594 34974 30606 35026
rect 30658 34974 30670 35026
rect 17502 34962 17554 34974
rect 20750 34962 20802 34974
rect 3278 34914 3330 34926
rect 4734 34914 4786 34926
rect 9774 34914 9826 34926
rect 14366 34914 14418 34926
rect 17166 34914 17218 34926
rect 1698 34862 1710 34914
rect 1762 34862 1774 34914
rect 2706 34862 2718 34914
rect 2770 34862 2782 34914
rect 3278 34850 3330 34862
rect 3826 34850 3838 34902
rect 3890 34850 3902 34902
rect 4274 34862 4286 34914
rect 4338 34862 4350 34914
rect 5506 34862 5518 34914
rect 5570 34862 5582 34914
rect 5842 34862 5854 34914
rect 5906 34862 5918 34914
rect 7074 34862 7086 34914
rect 7138 34862 7150 34914
rect 7298 34862 7310 34914
rect 7362 34862 7374 34914
rect 8082 34862 8094 34914
rect 8146 34862 8158 34914
rect 9202 34862 9214 34914
rect 9266 34862 9278 34914
rect 13234 34862 13246 34914
rect 13298 34862 13310 34914
rect 13794 34862 13806 34914
rect 13858 34862 13870 34914
rect 14914 34862 14926 34914
rect 14978 34862 14990 34914
rect 15922 34862 15934 34914
rect 15986 34862 15998 34914
rect 4734 34850 4786 34862
rect 9774 34850 9826 34862
rect 14366 34850 14418 34862
rect 17166 34850 17218 34862
rect 17278 34914 17330 34926
rect 17278 34850 17330 34862
rect 18062 34914 18114 34926
rect 22430 34914 22482 34926
rect 25454 34914 25506 34926
rect 21186 34862 21198 34914
rect 21250 34862 21262 34914
rect 21522 34862 21534 34914
rect 21586 34862 21598 34914
rect 22754 34862 22766 34914
rect 22818 34862 22830 34914
rect 23762 34862 23774 34914
rect 23826 34862 23838 34914
rect 24658 34862 24670 34914
rect 24722 34862 24734 34914
rect 18062 34850 18114 34862
rect 22430 34850 22482 34862
rect 25454 34850 25506 34862
rect 5070 34802 5122 34814
rect 12910 34802 12962 34814
rect 10882 34750 10894 34802
rect 10946 34750 10958 34802
rect 5070 34738 5122 34750
rect 12910 34738 12962 34750
rect 16718 34802 16770 34814
rect 18162 34750 18174 34802
rect 18226 34750 18238 34802
rect 18722 34750 18734 34802
rect 18786 34750 18798 34802
rect 16718 34738 16770 34750
rect 10110 34690 10162 34702
rect 10110 34626 10162 34638
rect 16830 34690 16882 34702
rect 16830 34626 16882 34638
rect 25790 34690 25842 34702
rect 25790 34626 25842 34638
rect 672 34522 31024 34556
rect 672 34470 3806 34522
rect 3858 34470 3910 34522
rect 3962 34470 4014 34522
rect 4066 34470 23806 34522
rect 23858 34470 23910 34522
rect 23962 34470 24014 34522
rect 24066 34470 31024 34522
rect 672 34436 31024 34470
rect 7870 34354 7922 34366
rect 7870 34290 7922 34302
rect 2382 34242 2434 34254
rect 16830 34242 16882 34254
rect 6290 34190 6302 34242
rect 6354 34190 6366 34242
rect 2382 34178 2434 34190
rect 16830 34178 16882 34190
rect 20974 34242 21026 34254
rect 20974 34178 21026 34190
rect 10446 34130 10498 34142
rect 22654 34130 22706 34142
rect 25454 34130 25506 34142
rect 3938 34078 3950 34130
rect 4002 34078 4014 34130
rect 9090 34078 9102 34130
rect 9154 34078 9166 34130
rect 9650 34078 9662 34130
rect 9714 34078 9726 34130
rect 10770 34078 10782 34130
rect 10834 34078 10846 34130
rect 11890 34078 11902 34130
rect 11954 34078 11966 34130
rect 14690 34078 14702 34130
rect 14754 34078 14766 34130
rect 17266 34078 17278 34130
rect 17330 34078 17342 34130
rect 17602 34078 17614 34130
rect 17666 34078 17678 34130
rect 18834 34078 18846 34130
rect 18898 34078 18910 34130
rect 19842 34078 19854 34130
rect 19906 34078 19918 34130
rect 21410 34078 21422 34130
rect 21474 34078 21486 34130
rect 21746 34078 21758 34130
rect 21810 34078 21822 34130
rect 22978 34078 22990 34130
rect 23042 34078 23054 34130
rect 23986 34078 23998 34130
rect 24050 34078 24062 34130
rect 24882 34078 24894 34130
rect 24946 34078 24958 34130
rect 10446 34066 10498 34078
rect 22654 34066 22706 34078
rect 25454 34066 25506 34078
rect 30270 34130 30322 34142
rect 30270 34066 30322 34078
rect 8766 34018 8818 34030
rect 18286 34018 18338 34030
rect 3490 33966 3502 34018
rect 3554 33966 3566 34018
rect 6626 33966 6638 34018
rect 6690 33966 6702 34018
rect 9762 33966 9774 34018
rect 9826 33966 9838 34018
rect 17826 33966 17838 34018
rect 17890 33966 17902 34018
rect 21970 33966 21982 34018
rect 22034 33966 22046 34018
rect 24658 33966 24670 34018
rect 24722 33966 24734 34018
rect 8766 33954 8818 33966
rect 18286 33954 18338 33966
rect 12798 33906 12850 33918
rect 16382 33906 16434 33918
rect 15250 33854 15262 33906
rect 15314 33854 15326 33906
rect 12798 33842 12850 33854
rect 16382 33842 16434 33854
rect 25790 33906 25842 33918
rect 30594 33854 30606 33906
rect 30658 33854 30670 33906
rect 25790 33842 25842 33854
rect 672 33738 31024 33772
rect 672 33686 4466 33738
rect 4518 33686 4570 33738
rect 4622 33686 4674 33738
rect 4726 33686 24466 33738
rect 24518 33686 24570 33738
rect 24622 33686 24674 33738
rect 24726 33686 31024 33738
rect 672 33652 31024 33686
rect 6302 33570 6354 33582
rect 6302 33506 6354 33518
rect 17726 33570 17778 33582
rect 17726 33506 17778 33518
rect 19070 33570 19122 33582
rect 21746 33518 21758 33570
rect 21810 33518 21822 33570
rect 19070 33506 19122 33518
rect 2158 33458 2210 33470
rect 1810 33406 1822 33458
rect 1874 33406 1886 33458
rect 2158 33394 2210 33406
rect 2606 33458 2658 33470
rect 19294 33458 19346 33470
rect 3602 33406 3614 33458
rect 3666 33406 3678 33458
rect 7410 33406 7422 33458
rect 7474 33406 7486 33458
rect 11666 33406 11678 33458
rect 11730 33406 11742 33458
rect 14690 33406 14702 33458
rect 14754 33406 14766 33458
rect 18274 33406 18286 33458
rect 18338 33406 18350 33458
rect 2606 33394 2658 33406
rect 19294 33394 19346 33406
rect 19630 33458 19682 33470
rect 19630 33394 19682 33406
rect 20750 33458 20802 33470
rect 30594 33406 30606 33458
rect 30658 33406 30670 33458
rect 20750 33394 20802 33406
rect 4286 33346 4338 33358
rect 17054 33346 17106 33358
rect 2930 33294 2942 33346
rect 2994 33294 3006 33346
rect 3378 33294 3390 33346
rect 3442 33294 3454 33346
rect 4610 33294 4622 33346
rect 4674 33294 4686 33346
rect 4834 33294 4846 33346
rect 4898 33294 4910 33346
rect 5618 33294 5630 33346
rect 5682 33294 5694 33346
rect 14130 33294 14142 33346
rect 14194 33294 14206 33346
rect 4286 33282 4338 33294
rect 17054 33282 17106 33294
rect 17502 33346 17554 33358
rect 18510 33346 18562 33358
rect 18050 33294 18062 33346
rect 18114 33294 18126 33346
rect 17502 33282 17554 33294
rect 18510 33282 18562 33294
rect 18958 33346 19010 33358
rect 18958 33282 19010 33294
rect 19518 33346 19570 33358
rect 21074 33294 21086 33346
rect 21138 33294 21150 33346
rect 21522 33294 21534 33346
rect 21586 33294 21598 33346
rect 22306 33294 22318 33346
rect 22370 33294 22382 33346
rect 22754 33294 22766 33346
rect 22818 33294 22830 33346
rect 23762 33294 23774 33346
rect 23826 33294 23838 33346
rect 30370 33294 30382 33346
rect 30434 33294 30446 33346
rect 19518 33282 19570 33294
rect 16718 33234 16770 33246
rect 7858 33182 7870 33234
rect 7922 33182 7934 33234
rect 11218 33182 11230 33234
rect 11282 33182 11294 33234
rect 16718 33170 16770 33182
rect 16830 33234 16882 33246
rect 16830 33170 16882 33182
rect 17614 33234 17666 33246
rect 17614 33170 17666 33182
rect 18734 33234 18786 33246
rect 18734 33170 18786 33182
rect 19854 33234 19906 33246
rect 19854 33170 19906 33182
rect 29598 33234 29650 33246
rect 29598 33170 29650 33182
rect 12798 33122 12850 33134
rect 12798 33058 12850 33070
rect 15822 33122 15874 33134
rect 15822 33058 15874 33070
rect 20078 33122 20130 33134
rect 20078 33058 20130 33070
rect 29710 33122 29762 33134
rect 29710 33058 29762 33070
rect 672 32954 31024 32988
rect 672 32902 3806 32954
rect 3858 32902 3910 32954
rect 3962 32902 4014 32954
rect 4066 32902 23806 32954
rect 23858 32902 23910 32954
rect 23962 32902 24014 32954
rect 24066 32902 31024 32954
rect 672 32868 31024 32902
rect 1150 32786 1202 32798
rect 1150 32722 1202 32734
rect 7982 32786 8034 32798
rect 7982 32722 8034 32734
rect 9886 32786 9938 32798
rect 9886 32722 9938 32734
rect 13694 32786 13746 32798
rect 23438 32786 23490 32798
rect 19282 32734 19294 32786
rect 19346 32734 19358 32786
rect 13694 32722 13746 32734
rect 23438 32722 23490 32734
rect 15150 32674 15202 32686
rect 6402 32622 6414 32674
rect 6466 32622 6478 32674
rect 15150 32610 15202 32622
rect 21086 32674 21138 32686
rect 21086 32610 21138 32622
rect 16606 32562 16658 32574
rect 18734 32562 18786 32574
rect 20526 32562 20578 32574
rect 2818 32510 2830 32562
rect 2882 32510 2894 32562
rect 11442 32510 11454 32562
rect 11506 32510 11518 32562
rect 13010 32510 13022 32562
rect 13074 32510 13086 32562
rect 15586 32510 15598 32562
rect 15650 32510 15662 32562
rect 15922 32510 15934 32562
rect 15986 32510 15998 32562
rect 17266 32510 17278 32562
rect 17330 32510 17342 32562
rect 18162 32510 18174 32562
rect 18226 32510 18238 32562
rect 18946 32510 18958 32562
rect 19010 32510 19022 32562
rect 19394 32510 19406 32562
rect 19458 32510 19470 32562
rect 16606 32498 16658 32510
rect 18734 32498 18786 32510
rect 20526 32498 20578 32510
rect 20974 32562 21026 32574
rect 20974 32498 21026 32510
rect 21198 32562 21250 32574
rect 21858 32510 21870 32562
rect 21922 32510 21934 32562
rect 21198 32498 21250 32510
rect 2370 32398 2382 32450
rect 2434 32398 2446 32450
rect 10994 32398 11006 32450
rect 11058 32398 11070 32450
rect 12898 32398 12910 32450
rect 12962 32398 12974 32450
rect 16146 32398 16158 32450
rect 16210 32398 16222 32450
rect 14030 32338 14082 32350
rect 6850 32286 6862 32338
rect 6914 32286 6926 32338
rect 14030 32274 14082 32286
rect 19518 32338 19570 32350
rect 22306 32286 22318 32338
rect 22370 32286 22382 32338
rect 19518 32274 19570 32286
rect 672 32170 31024 32204
rect 672 32118 4466 32170
rect 4518 32118 4570 32170
rect 4622 32118 4674 32170
rect 4726 32118 24466 32170
rect 24518 32118 24570 32170
rect 24622 32118 24674 32170
rect 24726 32118 31024 32170
rect 672 32084 31024 32118
rect 13806 32002 13858 32014
rect 13806 31938 13858 31950
rect 18062 32002 18114 32014
rect 18062 31938 18114 31950
rect 18286 32002 18338 32014
rect 30270 32002 30322 32014
rect 22082 31950 22094 32002
rect 22146 31950 22158 32002
rect 18286 31938 18338 31950
rect 30270 31938 30322 31950
rect 5630 31890 5682 31902
rect 10670 31890 10722 31902
rect 16046 31890 16098 31902
rect 2930 31838 2942 31890
rect 2994 31838 3006 31890
rect 6738 31838 6750 31890
rect 6802 31838 6814 31890
rect 9538 31838 9550 31890
rect 9602 31838 9614 31890
rect 11890 31838 11902 31890
rect 11954 31838 11966 31890
rect 14914 31838 14926 31890
rect 14978 31838 14990 31890
rect 5630 31826 5682 31838
rect 10670 31826 10722 31838
rect 16046 31826 16098 31838
rect 17390 31890 17442 31902
rect 17390 31826 17442 31838
rect 19070 31890 19122 31902
rect 19070 31826 19122 31838
rect 23214 31890 23266 31902
rect 30594 31838 30606 31890
rect 30658 31838 30670 31890
rect 23214 31826 23266 31838
rect 3614 31778 3666 31790
rect 16158 31778 16210 31790
rect 17614 31778 17666 31790
rect 19518 31778 19570 31790
rect 2370 31726 2382 31778
rect 2434 31726 2446 31778
rect 2706 31726 2718 31778
rect 2770 31726 2782 31778
rect 4162 31726 4174 31778
rect 4226 31726 4238 31778
rect 4946 31726 4958 31778
rect 5010 31726 5022 31778
rect 17042 31726 17054 31778
rect 17106 31726 17118 31778
rect 19282 31726 19294 31778
rect 19346 31726 19358 31778
rect 21522 31726 21534 31778
rect 21586 31726 21598 31778
rect 3614 31714 3666 31726
rect 16158 31714 16210 31726
rect 17614 31714 17666 31726
rect 19518 31714 19570 31726
rect 1934 31666 1986 31678
rect 18174 31666 18226 31678
rect 7186 31614 7198 31666
rect 7250 31614 7262 31666
rect 9090 31614 9102 31666
rect 9154 31614 9166 31666
rect 11554 31614 11566 31666
rect 11618 31614 11630 31666
rect 15362 31614 15374 31666
rect 15426 31614 15438 31666
rect 19618 31614 19630 31666
rect 19682 31614 19694 31666
rect 1934 31602 1986 31614
rect 18174 31602 18226 31614
rect 13134 31554 13186 31566
rect 13134 31490 13186 31502
rect 17054 31554 17106 31566
rect 17054 31490 17106 31502
rect 18622 31554 18674 31566
rect 18622 31490 18674 31502
rect 18734 31554 18786 31566
rect 18734 31490 18786 31502
rect 672 31386 31024 31420
rect 672 31334 3806 31386
rect 3858 31334 3910 31386
rect 3962 31334 4014 31386
rect 4066 31334 23806 31386
rect 23858 31334 23910 31386
rect 23962 31334 24014 31386
rect 24066 31334 31024 31386
rect 672 31300 31024 31334
rect 3166 31218 3218 31230
rect 3166 31154 3218 31166
rect 5070 31218 5122 31230
rect 5070 31154 5122 31166
rect 8990 31218 9042 31230
rect 8990 31154 9042 31166
rect 15150 31218 15202 31230
rect 15150 31154 15202 31166
rect 18510 31218 18562 31230
rect 18510 31154 18562 31166
rect 17166 31106 17218 31118
rect 7410 31054 7422 31106
rect 7474 31054 7486 31106
rect 17166 31042 17218 31054
rect 15486 30994 15538 31006
rect 1586 30942 1598 30994
rect 1650 30942 1662 30994
rect 6738 30942 6750 30994
rect 6802 30942 6814 30994
rect 10434 30942 10446 30994
rect 10498 30942 10510 30994
rect 13010 30942 13022 30994
rect 13074 30942 13086 30994
rect 15486 30930 15538 30942
rect 16606 30994 16658 31006
rect 16606 30930 16658 30942
rect 17054 30994 17106 31006
rect 17054 30930 17106 30942
rect 17278 30994 17330 31006
rect 19742 30994 19794 31006
rect 18050 30942 18062 30994
rect 18114 30942 18126 30994
rect 20066 30942 20078 30994
rect 20130 30942 20142 30994
rect 30370 30942 30382 30994
rect 30434 30942 30446 30994
rect 17278 30930 17330 30942
rect 19742 30930 19794 30942
rect 19294 30882 19346 30894
rect 2034 30830 2046 30882
rect 2098 30830 2110 30882
rect 6178 30830 6190 30882
rect 6242 30830 6254 30882
rect 10994 30830 11006 30882
rect 11058 30830 11070 30882
rect 13346 30830 13358 30882
rect 13410 30830 13422 30882
rect 15698 30830 15710 30882
rect 15762 30830 15774 30882
rect 16034 30830 16046 30882
rect 16098 30830 16110 30882
rect 17714 30830 17726 30882
rect 17778 30830 17790 30882
rect 19506 30830 19518 30882
rect 19570 30830 19582 30882
rect 19294 30818 19346 30830
rect 12126 30770 12178 30782
rect 7858 30718 7870 30770
rect 7922 30718 7934 30770
rect 12126 30706 12178 30718
rect 14590 30770 14642 30782
rect 14590 30706 14642 30718
rect 18846 30770 18898 30782
rect 18846 30706 18898 30718
rect 20078 30770 20130 30782
rect 30594 30718 30606 30770
rect 30658 30718 30670 30770
rect 20078 30706 20130 30718
rect 672 30602 31024 30636
rect 672 30550 4466 30602
rect 4518 30550 4570 30602
rect 4622 30550 4674 30602
rect 4726 30550 24466 30602
rect 24518 30550 24570 30602
rect 24622 30550 24674 30602
rect 24726 30550 31024 30602
rect 672 30516 31024 30550
rect 16270 30434 16322 30446
rect 7074 30382 7086 30434
rect 7138 30382 7150 30434
rect 10210 30382 10222 30434
rect 10274 30382 10286 30434
rect 12786 30382 12798 30434
rect 12850 30382 12862 30434
rect 16270 30370 16322 30382
rect 17838 30434 17890 30446
rect 20750 30434 20802 30446
rect 18834 30382 18846 30434
rect 18898 30382 18910 30434
rect 17838 30370 17890 30382
rect 20750 30370 20802 30382
rect 2718 30322 2770 30334
rect 15934 30322 15986 30334
rect 3714 30270 3726 30322
rect 3778 30270 3790 30322
rect 2718 30258 2770 30270
rect 15934 30258 15986 30270
rect 16046 30322 16098 30334
rect 16046 30258 16098 30270
rect 17054 30322 17106 30334
rect 17054 30258 17106 30270
rect 21310 30322 21362 30334
rect 21310 30258 21362 30270
rect 21422 30322 21474 30334
rect 30594 30270 30606 30322
rect 30658 30270 30670 30322
rect 21422 30258 21474 30270
rect 11790 30210 11842 30222
rect 13470 30210 13522 30222
rect 20302 30210 20354 30222
rect 3042 30158 3054 30210
rect 3106 30158 3118 30210
rect 3490 30158 3502 30210
rect 3554 30158 3566 30210
rect 4274 30158 4286 30210
rect 4338 30158 4350 30210
rect 4834 30158 4846 30210
rect 4898 30158 4910 30210
rect 5730 30158 5742 30210
rect 5794 30158 5806 30210
rect 6626 30158 6638 30210
rect 6690 30158 6702 30210
rect 9762 30158 9774 30210
rect 9826 30158 9838 30210
rect 12226 30158 12238 30210
rect 12290 30158 12302 30210
rect 12562 30158 12574 30210
rect 12626 30158 12638 30210
rect 13794 30158 13806 30210
rect 13858 30158 13870 30210
rect 14802 30158 14814 30210
rect 14866 30158 14878 30210
rect 17266 30158 17278 30210
rect 17330 30158 17342 30210
rect 17826 30158 17838 30210
rect 17890 30158 17902 30210
rect 11790 30146 11842 30158
rect 13470 30146 13522 30158
rect 20302 30146 20354 30158
rect 20862 30210 20914 30222
rect 20862 30146 20914 30158
rect 20974 30210 21026 30222
rect 20974 30146 21026 30158
rect 21646 30210 21698 30222
rect 21646 30146 21698 30158
rect 30270 30210 30322 30222
rect 30270 30146 30322 30158
rect 18386 30046 18398 30098
rect 18450 30046 18462 30098
rect 8206 29986 8258 29998
rect 8206 29922 8258 29934
rect 11342 29986 11394 29998
rect 19966 29986 20018 29998
rect 17602 29934 17614 29986
rect 17666 29934 17678 29986
rect 11342 29922 11394 29934
rect 19966 29922 20018 29934
rect 672 29818 31024 29852
rect 672 29766 3806 29818
rect 3858 29766 3910 29818
rect 3962 29766 4014 29818
rect 4066 29766 23806 29818
rect 23858 29766 23910 29818
rect 23962 29766 24014 29818
rect 24066 29766 31024 29818
rect 672 29732 31024 29766
rect 1150 29650 1202 29662
rect 1150 29586 1202 29598
rect 5070 29650 5122 29662
rect 5070 29586 5122 29598
rect 20750 29650 20802 29662
rect 20750 29586 20802 29598
rect 16830 29538 16882 29550
rect 2706 29486 2718 29538
rect 2770 29486 2782 29538
rect 6626 29486 6638 29538
rect 6690 29486 6702 29538
rect 7522 29486 7534 29538
rect 7586 29486 7598 29538
rect 16830 29474 16882 29486
rect 18286 29426 18338 29438
rect 20638 29426 20690 29438
rect 21870 29426 21922 29438
rect 10546 29374 10558 29426
rect 10610 29374 10622 29426
rect 14354 29374 14366 29426
rect 14418 29374 14430 29426
rect 17154 29374 17166 29426
rect 17218 29374 17230 29426
rect 17602 29374 17614 29426
rect 17666 29374 17678 29426
rect 18834 29374 18846 29426
rect 18898 29374 18910 29426
rect 19842 29374 19854 29426
rect 19906 29374 19918 29426
rect 21298 29374 21310 29426
rect 21362 29374 21374 29426
rect 18286 29362 18338 29374
rect 20638 29362 20690 29374
rect 21870 29362 21922 29374
rect 22206 29426 22258 29438
rect 22206 29362 22258 29374
rect 30270 29426 30322 29438
rect 30270 29362 30322 29374
rect 20974 29314 21026 29326
rect 2258 29262 2270 29314
rect 2322 29262 2334 29314
rect 6178 29262 6190 29314
rect 6242 29262 6254 29314
rect 7970 29262 7982 29314
rect 8034 29262 8046 29314
rect 10994 29262 11006 29314
rect 11058 29262 11070 29314
rect 14802 29262 14814 29314
rect 14866 29262 14878 29314
rect 17826 29262 17838 29314
rect 17890 29262 17902 29314
rect 20974 29250 21026 29262
rect 21534 29314 21586 29326
rect 21534 29250 21586 29262
rect 22542 29314 22594 29326
rect 22542 29250 22594 29262
rect 9102 29202 9154 29214
rect 9102 29138 9154 29150
rect 12126 29202 12178 29214
rect 12126 29138 12178 29150
rect 15934 29202 15986 29214
rect 15934 29138 15986 29150
rect 21422 29202 21474 29214
rect 21422 29138 21474 29150
rect 22094 29202 22146 29214
rect 30594 29150 30606 29202
rect 30658 29150 30670 29202
rect 22094 29138 22146 29150
rect 672 29034 31024 29068
rect 672 28982 4466 29034
rect 4518 28982 4570 29034
rect 4622 28982 4674 29034
rect 4726 28982 24466 29034
rect 24518 28982 24570 29034
rect 24622 28982 24674 29034
rect 24726 28982 31024 29034
rect 672 28948 31024 28982
rect 3278 28866 3330 28878
rect 17502 28866 17554 28878
rect 2146 28814 2158 28866
rect 2210 28814 2222 28866
rect 7298 28814 7310 28866
rect 7362 28814 7374 28866
rect 18610 28814 18622 28866
rect 18674 28814 18686 28866
rect 21298 28814 21310 28866
rect 21362 28814 21374 28866
rect 3278 28802 3330 28814
rect 17502 28802 17554 28814
rect 8318 28754 8370 28766
rect 19630 28754 19682 28766
rect 9874 28702 9886 28754
rect 9938 28702 9950 28754
rect 13906 28702 13918 28754
rect 13970 28702 13982 28754
rect 8318 28690 8370 28702
rect 19630 28690 19682 28702
rect 30270 28754 30322 28766
rect 30594 28702 30606 28754
rect 30658 28702 30670 28754
rect 30270 28690 30322 28702
rect 6862 28642 6914 28654
rect 11790 28647 11842 28659
rect 1698 28590 1710 28642
rect 1762 28590 1774 28642
rect 5170 28590 5182 28642
rect 5234 28590 5246 28642
rect 6066 28590 6078 28642
rect 6130 28590 6142 28642
rect 7522 28590 7534 28642
rect 7586 28590 7598 28642
rect 7970 28590 7982 28642
rect 8034 28590 8046 28642
rect 9202 28590 9214 28642
rect 9266 28590 9278 28642
rect 9762 28590 9774 28642
rect 9826 28590 9838 28642
rect 10434 28590 10446 28642
rect 10498 28590 10510 28642
rect 10882 28590 10894 28642
rect 10946 28590 10958 28642
rect 11106 28590 11118 28642
rect 11170 28590 11182 28642
rect 14590 28642 14642 28654
rect 19966 28642 20018 28654
rect 6862 28578 6914 28590
rect 11790 28583 11842 28595
rect 13234 28590 13246 28642
rect 13298 28590 13310 28642
rect 13794 28590 13806 28642
rect 13858 28590 13870 28642
rect 15026 28590 15038 28642
rect 15090 28590 15102 28642
rect 15922 28590 15934 28642
rect 15986 28590 15998 28642
rect 14590 28578 14642 28590
rect 19966 28578 20018 28590
rect 8878 28530 8930 28542
rect 8878 28466 8930 28478
rect 12910 28530 12962 28542
rect 19742 28530 19794 28542
rect 19058 28478 19070 28530
rect 19122 28478 19134 28530
rect 20850 28478 20862 28530
rect 20914 28478 20926 28530
rect 12910 28466 12962 28478
rect 19742 28466 19794 28478
rect 20078 28418 20130 28430
rect 20078 28354 20130 28366
rect 22430 28418 22482 28430
rect 22430 28354 22482 28366
rect 672 28250 31024 28284
rect 672 28198 3806 28250
rect 3858 28198 3910 28250
rect 3962 28198 4014 28250
rect 4066 28198 23806 28250
rect 23858 28198 23910 28250
rect 23962 28198 24014 28250
rect 24066 28198 31024 28250
rect 672 28164 31024 28198
rect 19966 28082 20018 28094
rect 19966 28018 20018 28030
rect 21870 28082 21922 28094
rect 21870 28018 21922 28030
rect 1150 27970 1202 27982
rect 8318 27970 8370 27982
rect 6290 27918 6302 27970
rect 6354 27918 6366 27970
rect 1150 27906 1202 27918
rect 8318 27906 8370 27918
rect 20862 27970 20914 27982
rect 20862 27906 20914 27918
rect 21982 27970 22034 27982
rect 21982 27906 22034 27918
rect 15822 27858 15874 27870
rect 20638 27858 20690 27870
rect 1586 27806 1598 27858
rect 1650 27806 1662 27858
rect 2034 27806 2046 27858
rect 2098 27806 2110 27858
rect 2706 27806 2718 27858
rect 2770 27806 2782 27858
rect 3266 27806 3278 27858
rect 3330 27806 3342 27858
rect 4162 27806 4174 27858
rect 4226 27806 4238 27858
rect 8642 27806 8654 27858
rect 8706 27806 8718 27858
rect 9090 27806 9102 27858
rect 9154 27806 9166 27858
rect 10546 27806 10558 27858
rect 10610 27806 10622 27858
rect 11442 27806 11454 27858
rect 11506 27806 11518 27858
rect 14466 27806 14478 27858
rect 14530 27806 14542 27858
rect 14914 27806 14926 27858
rect 14978 27806 14990 27858
rect 16146 27806 16158 27858
rect 16210 27806 16222 27858
rect 17154 27806 17166 27858
rect 17218 27806 17230 27858
rect 18386 27806 18398 27858
rect 18450 27806 18462 27858
rect 15822 27794 15874 27806
rect 20638 27794 20690 27806
rect 21086 27858 21138 27870
rect 21646 27858 21698 27870
rect 21298 27806 21310 27858
rect 21362 27806 21374 27858
rect 21086 27794 21138 27806
rect 21646 27794 21698 27806
rect 29598 27858 29650 27870
rect 29598 27794 29650 27806
rect 30270 27858 30322 27870
rect 30270 27794 30322 27806
rect 9774 27746 9826 27758
rect 6626 27694 6638 27746
rect 6690 27694 6702 27746
rect 9774 27682 9826 27694
rect 14142 27746 14194 27758
rect 29710 27746 29762 27758
rect 18722 27694 18734 27746
rect 18786 27694 18798 27746
rect 14142 27682 14194 27694
rect 29710 27682 29762 27694
rect 7870 27634 7922 27646
rect 20750 27634 20802 27646
rect 2146 27582 2158 27634
rect 2210 27582 2222 27634
rect 9314 27582 9326 27634
rect 9378 27582 9390 27634
rect 15138 27582 15150 27634
rect 15202 27582 15214 27634
rect 30594 27582 30606 27634
rect 30658 27582 30670 27634
rect 7870 27570 7922 27582
rect 20750 27570 20802 27582
rect 672 27466 31024 27500
rect 672 27414 4466 27466
rect 4518 27414 4570 27466
rect 4622 27414 4674 27466
rect 4726 27414 24466 27466
rect 24518 27414 24570 27466
rect 24622 27414 24674 27466
rect 24726 27414 31024 27466
rect 672 27380 31024 27414
rect 18622 27298 18674 27310
rect 18622 27234 18674 27246
rect 19182 27298 19234 27310
rect 19182 27234 19234 27246
rect 21086 27298 21138 27310
rect 21086 27234 21138 27246
rect 30270 27298 30322 27310
rect 30270 27234 30322 27246
rect 1486 27186 1538 27198
rect 8318 27186 8370 27198
rect 10334 27186 10386 27198
rect 2482 27134 2494 27186
rect 2546 27134 2558 27186
rect 7298 27134 7310 27186
rect 7362 27134 7374 27186
rect 9874 27134 9886 27186
rect 9938 27134 9950 27186
rect 1486 27122 1538 27134
rect 8318 27122 8370 27134
rect 10334 27122 10386 27134
rect 14702 27186 14754 27198
rect 16158 27186 16210 27198
rect 18510 27186 18562 27198
rect 15138 27134 15150 27186
rect 15202 27134 15214 27186
rect 16930 27134 16942 27186
rect 16994 27134 17006 27186
rect 14702 27122 14754 27134
rect 16158 27122 16210 27134
rect 18510 27122 18562 27134
rect 19294 27186 19346 27198
rect 19294 27122 19346 27134
rect 19630 27186 19682 27198
rect 19630 27122 19682 27134
rect 19742 27186 19794 27198
rect 30594 27134 30606 27186
rect 30658 27134 30670 27186
rect 19742 27122 19794 27134
rect 3166 27074 3218 27086
rect 17614 27074 17666 27086
rect 1810 27022 1822 27074
rect 1874 27022 1886 27074
rect 2370 27022 2382 27074
rect 2434 27022 2446 27074
rect 3714 27022 3726 27074
rect 3778 27022 3790 27074
rect 4498 27022 4510 27074
rect 4562 27022 4574 27074
rect 5170 27022 5182 27074
rect 5234 27022 5246 27074
rect 6066 27022 6078 27074
rect 6130 27022 6142 27074
rect 6738 27022 6750 27074
rect 6802 27022 6814 27074
rect 7522 27022 7534 27074
rect 7586 27022 7598 27074
rect 7858 27022 7870 27074
rect 7922 27022 7934 27074
rect 9202 27022 9214 27074
rect 9266 27022 9278 27074
rect 9762 27022 9774 27074
rect 9826 27022 9838 27074
rect 10882 27022 10894 27074
rect 10946 27022 10958 27074
rect 11890 27022 11902 27074
rect 11954 27022 11966 27074
rect 13010 27022 13022 27074
rect 13074 27022 13086 27074
rect 13906 27022 13918 27074
rect 13970 27022 13982 27074
rect 15250 27022 15262 27074
rect 15314 27022 15326 27074
rect 15698 27022 15710 27074
rect 15762 27022 15774 27074
rect 16818 27022 16830 27074
rect 16882 27022 16894 27074
rect 3166 27010 3218 27022
rect 17614 27010 17666 27022
rect 8878 26962 8930 26974
rect 8878 26898 8930 26910
rect 21198 26962 21250 26974
rect 21198 26898 21250 26910
rect 21310 26962 21362 26974
rect 21310 26898 21362 26910
rect 21646 26962 21698 26974
rect 21646 26898 21698 26910
rect 21758 26962 21810 26974
rect 21758 26898 21810 26910
rect 17950 26850 18002 26862
rect 17950 26786 18002 26798
rect 18622 26850 18674 26862
rect 18622 26786 18674 26798
rect 19182 26850 19234 26862
rect 19182 26786 19234 26798
rect 672 26682 31024 26716
rect 672 26630 3806 26682
rect 3858 26630 3910 26682
rect 3962 26630 4014 26682
rect 4066 26630 23806 26682
rect 23858 26630 23910 26682
rect 23962 26630 24014 26682
rect 24066 26630 31024 26682
rect 672 26596 31024 26630
rect 2830 26514 2882 26526
rect 2830 26450 2882 26462
rect 16158 26514 16210 26526
rect 16158 26450 16210 26462
rect 20750 26514 20802 26526
rect 20750 26450 20802 26462
rect 8766 26402 8818 26414
rect 1250 26350 1262 26402
rect 1314 26350 1326 26402
rect 8766 26338 8818 26350
rect 13918 26402 13970 26414
rect 13918 26338 13970 26350
rect 8318 26290 8370 26302
rect 6626 26238 6638 26290
rect 6690 26238 6702 26290
rect 9090 26238 9102 26290
rect 9154 26238 9166 26290
rect 9538 26238 9550 26290
rect 9602 26238 9614 26290
rect 10322 26238 10334 26290
rect 10386 26238 10398 26290
rect 10882 26238 10894 26290
rect 10946 26238 10958 26290
rect 11890 26238 11902 26290
rect 11954 26238 11966 26290
rect 14466 26238 14478 26290
rect 14530 26238 14542 26290
rect 17154 26238 17166 26290
rect 17218 26238 17230 26290
rect 22306 26238 22318 26290
rect 22370 26238 22382 26290
rect 8318 26226 8370 26238
rect 1586 26126 1598 26178
rect 1650 26126 1662 26178
rect 14030 26066 14082 26078
rect 16606 26066 16658 26078
rect 7186 26014 7198 26066
rect 7250 26014 7262 26066
rect 9762 26014 9774 26066
rect 9826 26014 9838 26066
rect 15026 26014 15038 26066
rect 15090 26014 15102 26066
rect 14030 26002 14082 26014
rect 16606 26002 16658 26014
rect 16718 26066 16770 26078
rect 16718 26002 16770 26014
rect 16830 26066 16882 26078
rect 21858 26014 21870 26066
rect 21922 26014 21934 26066
rect 16830 26002 16882 26014
rect 672 25898 31024 25932
rect 672 25846 4466 25898
rect 4518 25846 4570 25898
rect 4622 25846 4674 25898
rect 4726 25846 24466 25898
rect 24518 25846 24570 25898
rect 24622 25846 24674 25898
rect 24726 25846 31024 25898
rect 672 25812 31024 25846
rect 7310 25730 7362 25742
rect 4162 25678 4174 25730
rect 4226 25678 4238 25730
rect 6178 25678 6190 25730
rect 6242 25678 6254 25730
rect 7310 25666 7362 25678
rect 15598 25730 15650 25742
rect 15598 25666 15650 25678
rect 17278 25730 17330 25742
rect 17278 25666 17330 25678
rect 17726 25730 17778 25742
rect 17726 25666 17778 25678
rect 17950 25730 18002 25742
rect 22318 25730 22370 25742
rect 20738 25678 20750 25730
rect 20802 25678 20814 25730
rect 17950 25666 18002 25678
rect 22318 25666 22370 25678
rect 30270 25730 30322 25742
rect 30270 25666 30322 25678
rect 3726 25618 3778 25630
rect 3726 25554 3778 25566
rect 5182 25618 5234 25630
rect 16046 25618 16098 25630
rect 9538 25566 9550 25618
rect 9602 25566 9614 25618
rect 12898 25566 12910 25618
rect 12962 25566 12974 25618
rect 5182 25554 5234 25566
rect 16046 25554 16098 25566
rect 18062 25618 18114 25630
rect 30594 25566 30606 25618
rect 30658 25566 30670 25618
rect 18062 25554 18114 25566
rect 15710 25506 15762 25518
rect 2146 25454 2158 25506
rect 2210 25454 2222 25506
rect 2930 25454 2942 25506
rect 2994 25454 3006 25506
rect 3154 25454 3166 25506
rect 3218 25454 3230 25506
rect 4274 25454 4286 25506
rect 4338 25454 4350 25506
rect 4834 25454 4846 25506
rect 4898 25454 4910 25506
rect 5730 25454 5742 25506
rect 5794 25454 5806 25506
rect 9090 25454 9102 25506
rect 9154 25454 9166 25506
rect 12226 25454 12238 25506
rect 12290 25454 12302 25506
rect 12786 25454 12798 25506
rect 12850 25454 12862 25506
rect 13458 25454 13470 25506
rect 13522 25454 13534 25506
rect 13906 25454 13918 25506
rect 13970 25454 13982 25506
rect 14914 25454 14926 25506
rect 14978 25454 14990 25506
rect 15710 25442 15762 25454
rect 15822 25506 15874 25518
rect 15822 25442 15874 25454
rect 16270 25506 16322 25518
rect 16270 25442 16322 25454
rect 16718 25506 16770 25518
rect 16718 25442 16770 25454
rect 16942 25506 16994 25518
rect 16942 25442 16994 25454
rect 17166 25506 17218 25518
rect 17166 25442 17218 25454
rect 17390 25506 17442 25518
rect 17390 25442 17442 25454
rect 21870 25506 21922 25518
rect 22530 25454 22542 25506
rect 22594 25454 22606 25506
rect 22754 25454 22766 25506
rect 22818 25454 22830 25506
rect 21870 25442 21922 25454
rect 11902 25394 11954 25406
rect 20290 25342 20302 25394
rect 20354 25342 20366 25394
rect 11902 25330 11954 25342
rect 10670 25282 10722 25294
rect 10670 25218 10722 25230
rect 22206 25282 22258 25294
rect 22206 25218 22258 25230
rect 672 25114 31024 25148
rect 672 25062 3806 25114
rect 3858 25062 3910 25114
rect 3962 25062 4014 25114
rect 4066 25062 23806 25114
rect 23858 25062 23910 25114
rect 23962 25062 24014 25114
rect 24066 25062 31024 25114
rect 672 25028 31024 25062
rect 2830 24946 2882 24958
rect 2830 24882 2882 24894
rect 6750 24946 6802 24958
rect 6750 24882 6802 24894
rect 8094 24946 8146 24958
rect 8094 24882 8146 24894
rect 14590 24946 14642 24958
rect 14590 24882 14642 24894
rect 15598 24946 15650 24958
rect 15598 24882 15650 24894
rect 21422 24946 21474 24958
rect 21422 24882 21474 24894
rect 22206 24946 22258 24958
rect 22206 24882 22258 24894
rect 20862 24834 20914 24846
rect 5170 24782 5182 24834
rect 5234 24782 5246 24834
rect 10546 24782 10558 24834
rect 10610 24782 10622 24834
rect 13010 24782 13022 24834
rect 13074 24782 13086 24834
rect 20862 24770 20914 24782
rect 21646 24834 21698 24846
rect 21646 24770 21698 24782
rect 22094 24722 22146 24734
rect 1250 24670 1262 24722
rect 1314 24670 1326 24722
rect 7298 24670 7310 24722
rect 7362 24670 7374 24722
rect 17266 24670 17278 24722
rect 17330 24670 17342 24722
rect 20626 24670 20638 24722
rect 20690 24670 20702 24722
rect 22094 24658 22146 24670
rect 30270 24722 30322 24734
rect 30270 24658 30322 24670
rect 8990 24610 9042 24622
rect 20974 24610 21026 24622
rect 1586 24558 1598 24610
rect 1650 24558 1662 24610
rect 5506 24558 5518 24610
rect 5570 24558 5582 24610
rect 7522 24558 7534 24610
rect 7586 24558 7598 24610
rect 13346 24558 13358 24610
rect 13410 24558 13422 24610
rect 16706 24558 16718 24610
rect 16770 24558 16782 24610
rect 8990 24546 9042 24558
rect 20974 24546 21026 24558
rect 21870 24610 21922 24622
rect 21870 24546 21922 24558
rect 8430 24498 8482 24510
rect 10098 24446 10110 24498
rect 10162 24446 10174 24498
rect 30594 24446 30606 24498
rect 30658 24446 30670 24498
rect 8430 24434 8482 24446
rect 672 24330 31024 24364
rect 672 24278 4466 24330
rect 4518 24278 4570 24330
rect 4622 24278 4674 24330
rect 4726 24278 24466 24330
rect 24518 24278 24570 24330
rect 24622 24278 24674 24330
rect 24726 24278 31024 24330
rect 672 24244 31024 24278
rect 1374 24162 1426 24174
rect 1374 24098 1426 24110
rect 7422 24162 7474 24174
rect 7422 24098 7474 24110
rect 3390 24050 3442 24062
rect 19854 24050 19906 24062
rect 1026 23998 1038 24050
rect 1090 23998 1102 24050
rect 2930 23998 2942 24050
rect 2994 23998 3006 24050
rect 6178 23998 6190 24050
rect 6242 23998 6254 24050
rect 10770 23998 10782 24050
rect 10834 23998 10846 24050
rect 14802 23998 14814 24050
rect 14866 23998 14878 24050
rect 3390 23986 3442 23998
rect 19854 23986 19906 23998
rect 20302 24050 20354 24062
rect 30270 24050 30322 24062
rect 21634 23998 21646 24050
rect 21698 23998 21710 24050
rect 30594 23998 30606 24050
rect 30658 23998 30670 24050
rect 20302 23986 20354 23998
rect 30270 23986 30322 23998
rect 2370 23886 2382 23938
rect 2434 23886 2446 23938
rect 2706 23886 2718 23938
rect 2770 23886 2782 23938
rect 4050 23886 4062 23938
rect 4114 23886 4126 23938
rect 4946 23886 4958 23938
rect 5010 23886 5022 23938
rect 14466 23886 14478 23938
rect 14530 23886 14542 23938
rect 19394 23886 19406 23938
rect 19458 23886 19470 23938
rect 19618 23886 19630 23938
rect 19682 23886 19694 23938
rect 23538 23886 23550 23938
rect 23602 23886 23614 23938
rect 1934 23826 1986 23838
rect 20414 23826 20466 23838
rect 23326 23826 23378 23838
rect 5842 23774 5854 23826
rect 5906 23774 5918 23826
rect 10434 23774 10446 23826
rect 10498 23774 10510 23826
rect 21186 23774 21198 23826
rect 21250 23774 21262 23826
rect 1934 23762 1986 23774
rect 20414 23762 20466 23774
rect 23326 23762 23378 23774
rect 12014 23714 12066 23726
rect 12014 23650 12066 23662
rect 16046 23714 16098 23726
rect 16046 23650 16098 23662
rect 19518 23714 19570 23726
rect 19518 23650 19570 23662
rect 20526 23714 20578 23726
rect 20526 23650 20578 23662
rect 22766 23714 22818 23726
rect 22766 23650 22818 23662
rect 23214 23714 23266 23726
rect 23214 23650 23266 23662
rect 672 23546 31024 23580
rect 672 23494 3806 23546
rect 3858 23494 3910 23546
rect 3962 23494 4014 23546
rect 4066 23494 23806 23546
rect 23858 23494 23910 23546
rect 23962 23494 24014 23546
rect 24066 23494 31024 23546
rect 672 23460 31024 23494
rect 4286 23378 4338 23390
rect 4286 23314 4338 23326
rect 6750 23378 6802 23390
rect 6750 23314 6802 23326
rect 11678 23378 11730 23390
rect 16034 23326 16046 23378
rect 16098 23326 16110 23378
rect 11678 23314 11730 23326
rect 5170 23214 5182 23266
rect 5234 23214 5246 23266
rect 14018 23214 14030 23266
rect 14082 23214 14094 23266
rect 15486 23154 15538 23166
rect 1250 23102 1262 23154
rect 1314 23102 1326 23154
rect 2706 23102 2718 23154
rect 2770 23102 2782 23154
rect 7634 23102 7646 23154
rect 7698 23102 7710 23154
rect 8082 23102 8094 23154
rect 8146 23102 8158 23154
rect 9426 23102 9438 23154
rect 9490 23102 9502 23154
rect 10210 23102 10222 23154
rect 10274 23102 10286 23154
rect 10994 23102 11006 23154
rect 11058 23102 11070 23154
rect 14578 23102 14590 23154
rect 14642 23102 14654 23154
rect 15250 23102 15262 23154
rect 15314 23102 15326 23154
rect 15486 23090 15538 23102
rect 16830 23154 16882 23166
rect 16830 23090 16882 23102
rect 17278 23154 17330 23166
rect 17278 23090 17330 23102
rect 17502 23154 17554 23166
rect 23214 23154 23266 23166
rect 18386 23102 18398 23154
rect 18450 23102 18462 23154
rect 22418 23102 22430 23154
rect 22482 23102 22494 23154
rect 23090 23102 23102 23154
rect 23154 23102 23166 23154
rect 17502 23090 17554 23102
rect 23214 23090 23266 23102
rect 23326 23154 23378 23166
rect 23326 23090 23378 23102
rect 23662 23154 23714 23166
rect 23662 23090 23714 23102
rect 23886 23154 23938 23166
rect 23886 23090 23938 23102
rect 30270 23154 30322 23166
rect 30270 23090 30322 23102
rect 7198 23042 7250 23054
rect 7198 22978 7250 22990
rect 8654 23042 8706 23054
rect 12014 23042 12066 23054
rect 10882 22990 10894 23042
rect 10946 22990 10958 23042
rect 8654 22978 8706 22990
rect 12014 22978 12066 22990
rect 13134 23042 13186 23054
rect 13134 22978 13186 22990
rect 13246 23042 13298 23054
rect 13246 22978 13298 22990
rect 13694 23042 13746 23054
rect 13694 22978 13746 22990
rect 14366 23042 14418 23054
rect 14366 22978 14418 22990
rect 14926 23042 14978 23054
rect 14926 22978 14978 22990
rect 15598 23042 15650 23054
rect 15598 22978 15650 22990
rect 16718 23042 16770 23054
rect 24222 23042 24274 23054
rect 18834 22990 18846 23042
rect 18898 22990 18910 23042
rect 21858 22990 21870 23042
rect 21922 22990 21934 23042
rect 16718 22978 16770 22990
rect 24222 22978 24274 22990
rect 2046 22930 2098 22942
rect 13470 22930 13522 22942
rect 1026 22878 1038 22930
rect 1090 22878 1102 22930
rect 1698 22878 1710 22930
rect 1762 22878 1774 22930
rect 3154 22878 3166 22930
rect 3218 22878 3230 22930
rect 5618 22878 5630 22930
rect 5682 22878 5694 22930
rect 8194 22878 8206 22930
rect 8258 22878 8270 22930
rect 2046 22866 2098 22878
rect 13470 22866 13522 22878
rect 13918 22930 13970 22942
rect 13918 22866 13970 22878
rect 14814 22930 14866 22942
rect 14814 22866 14866 22878
rect 17614 22930 17666 22942
rect 17614 22866 17666 22878
rect 19966 22930 20018 22942
rect 19966 22866 20018 22878
rect 20750 22930 20802 22942
rect 24110 22930 24162 22942
rect 23202 22878 23214 22930
rect 23266 22878 23278 22930
rect 30594 22878 30606 22930
rect 30658 22878 30670 22930
rect 20750 22866 20802 22878
rect 24110 22866 24162 22878
rect 672 22762 31024 22796
rect 672 22710 4466 22762
rect 4518 22710 4570 22762
rect 4622 22710 4674 22762
rect 4726 22710 24466 22762
rect 24518 22710 24570 22762
rect 24622 22710 24674 22762
rect 24726 22710 31024 22762
rect 672 22676 31024 22710
rect 3726 22594 3778 22606
rect 3726 22530 3778 22542
rect 4286 22594 4338 22606
rect 4286 22530 4338 22542
rect 14926 22594 14978 22606
rect 14926 22530 14978 22542
rect 16942 22594 16994 22606
rect 23438 22594 23490 22606
rect 18050 22542 18062 22594
rect 18114 22542 18126 22594
rect 16942 22530 16994 22542
rect 23438 22530 23490 22542
rect 30270 22594 30322 22606
rect 30270 22530 30322 22542
rect 16158 22482 16210 22494
rect 21198 22482 21250 22494
rect 2594 22430 2606 22482
rect 2658 22430 2670 22482
rect 5394 22430 5406 22482
rect 5458 22430 5470 22482
rect 7074 22430 7086 22482
rect 7138 22430 7150 22482
rect 10434 22430 10446 22482
rect 10498 22430 10510 22482
rect 12786 22430 12798 22482
rect 12850 22430 12862 22482
rect 20738 22430 20750 22482
rect 20802 22430 20814 22482
rect 30594 22430 30606 22482
rect 30658 22430 30670 22482
rect 16158 22418 16210 22430
rect 21198 22418 21250 22430
rect 14366 22370 14418 22382
rect 14366 22306 14418 22318
rect 14814 22370 14866 22382
rect 14814 22306 14866 22318
rect 15038 22370 15090 22382
rect 15038 22306 15090 22318
rect 15598 22370 15650 22382
rect 23550 22370 23602 22382
rect 15922 22318 15934 22370
rect 15986 22318 15998 22370
rect 20066 22318 20078 22370
rect 20130 22318 20142 22370
rect 20514 22318 20526 22370
rect 20578 22318 20590 22370
rect 21970 22318 21982 22370
rect 22034 22318 22046 22370
rect 22754 22318 22766 22370
rect 22818 22318 22830 22370
rect 23314 22318 23326 22370
rect 23378 22318 23390 22370
rect 15598 22306 15650 22318
rect 23550 22306 23602 22318
rect 19742 22258 19794 22270
rect 2146 22206 2158 22258
rect 2210 22206 2222 22258
rect 5842 22206 5854 22258
rect 5906 22206 5918 22258
rect 6626 22206 6638 22258
rect 6690 22206 6702 22258
rect 10098 22206 10110 22258
rect 10162 22206 10174 22258
rect 12338 22206 12350 22258
rect 12402 22206 12414 22258
rect 16146 22206 16158 22258
rect 16210 22206 16222 22258
rect 17042 22206 17054 22258
rect 17106 22206 17118 22258
rect 17602 22206 17614 22258
rect 17666 22206 17678 22258
rect 19742 22194 19794 22206
rect 23774 22258 23826 22270
rect 23774 22194 23826 22206
rect 8206 22146 8258 22158
rect 8206 22082 8258 22094
rect 11678 22146 11730 22158
rect 11678 22082 11730 22094
rect 13918 22146 13970 22158
rect 13918 22082 13970 22094
rect 16718 22146 16770 22158
rect 16718 22082 16770 22094
rect 19182 22146 19234 22158
rect 19182 22082 19234 22094
rect 672 21978 31024 22012
rect 672 21926 3806 21978
rect 3858 21926 3910 21978
rect 3962 21926 4014 21978
rect 4066 21926 23806 21978
rect 23858 21926 23910 21978
rect 23962 21926 24014 21978
rect 24066 21926 31024 21978
rect 672 21892 31024 21926
rect 2942 21810 2994 21822
rect 2942 21746 2994 21758
rect 5742 21810 5794 21822
rect 5742 21746 5794 21758
rect 22542 21810 22594 21822
rect 22542 21746 22594 21758
rect 23102 21810 23154 21822
rect 23102 21746 23154 21758
rect 16830 21698 16882 21710
rect 1362 21646 1374 21698
rect 1426 21646 1438 21698
rect 20962 21646 20974 21698
rect 21026 21646 21038 21698
rect 16830 21634 16882 21646
rect 14254 21586 14306 21598
rect 22990 21586 23042 21598
rect 7298 21534 7310 21586
rect 7362 21534 7374 21586
rect 8082 21534 8094 21586
rect 8146 21534 8158 21586
rect 13122 21534 13134 21586
rect 13186 21534 13198 21586
rect 13570 21534 13582 21586
rect 13634 21534 13646 21586
rect 14802 21534 14814 21586
rect 14866 21534 14878 21586
rect 15810 21534 15822 21586
rect 15874 21534 15886 21586
rect 17154 21534 17166 21586
rect 17218 21534 17230 21586
rect 17714 21534 17726 21586
rect 17778 21534 17790 21586
rect 18386 21534 18398 21586
rect 18450 21534 18462 21586
rect 19058 21534 19070 21586
rect 19122 21534 19134 21586
rect 19842 21534 19854 21586
rect 19906 21534 19918 21586
rect 20850 21534 20862 21586
rect 20914 21534 20926 21586
rect 14254 21522 14306 21534
rect 22990 21522 23042 21534
rect 12798 21474 12850 21486
rect 1810 21422 1822 21474
rect 1874 21422 1886 21474
rect 6850 21422 6862 21474
rect 6914 21422 6926 21474
rect 7858 21422 7870 21474
rect 7922 21422 7934 21474
rect 12798 21410 12850 21422
rect 16494 21474 16546 21486
rect 21410 21422 21422 21474
rect 21474 21422 21486 21474
rect 16494 21410 16546 21422
rect 4062 21362 4114 21374
rect 3714 21310 3726 21362
rect 3778 21310 3790 21362
rect 4062 21298 4114 21310
rect 8542 21362 8594 21374
rect 16382 21362 16434 21374
rect 30270 21362 30322 21374
rect 13794 21310 13806 21362
rect 13858 21310 13870 21362
rect 17826 21310 17838 21362
rect 17890 21310 17902 21362
rect 30594 21310 30606 21362
rect 30658 21310 30670 21362
rect 8542 21298 8594 21310
rect 16382 21298 16434 21310
rect 30270 21298 30322 21310
rect 672 21194 31024 21228
rect 672 21142 4466 21194
rect 4518 21142 4570 21194
rect 4622 21142 4674 21194
rect 4726 21142 24466 21194
rect 24518 21142 24570 21194
rect 24622 21142 24674 21194
rect 24726 21142 31024 21194
rect 672 21108 31024 21142
rect 16830 21026 16882 21038
rect 16830 20962 16882 20974
rect 20750 21026 20802 21038
rect 20750 20962 20802 20974
rect 11678 20914 11730 20926
rect 16158 20914 16210 20926
rect 21198 20914 21250 20926
rect 3714 20862 3726 20914
rect 3778 20862 3790 20914
rect 6066 20862 6078 20914
rect 6130 20862 6142 20914
rect 9986 20862 9998 20914
rect 10050 20862 10062 20914
rect 12674 20862 12686 20914
rect 12738 20862 12750 20914
rect 18050 20862 18062 20914
rect 18114 20862 18126 20914
rect 19506 20862 19518 20914
rect 19570 20862 19582 20914
rect 30594 20862 30606 20914
rect 30658 20862 30670 20914
rect 11678 20850 11730 20862
rect 16158 20850 16210 20862
rect 21198 20850 21250 20862
rect 3054 20802 3106 20814
rect 6526 20802 6578 20814
rect 11230 20802 11282 20814
rect 13134 20802 13186 20814
rect 15934 20802 15986 20814
rect 21310 20802 21362 20814
rect 1698 20750 1710 20802
rect 1762 20750 1774 20802
rect 2594 20750 2606 20802
rect 2658 20750 2670 20802
rect 3826 20750 3838 20802
rect 3890 20750 3902 20802
rect 4274 20750 4286 20802
rect 4338 20750 4350 20802
rect 5506 20750 5518 20802
rect 5570 20750 5582 20802
rect 5954 20750 5966 20802
rect 6018 20750 6030 20802
rect 7298 20750 7310 20802
rect 7362 20750 7374 20802
rect 8082 20750 8094 20802
rect 8146 20750 8158 20802
rect 12114 20750 12126 20802
rect 12178 20750 12190 20802
rect 12450 20750 12462 20802
rect 12514 20750 12526 20802
rect 13906 20750 13918 20802
rect 13970 20750 13982 20802
rect 14690 20750 14702 20802
rect 14754 20750 14766 20802
rect 18386 20750 18398 20802
rect 18450 20750 18462 20802
rect 3054 20738 3106 20750
rect 6526 20738 6578 20750
rect 11230 20738 11282 20750
rect 13134 20738 13186 20750
rect 15934 20738 15986 20750
rect 21310 20738 21362 20750
rect 21534 20802 21586 20814
rect 21534 20738 21586 20750
rect 21758 20802 21810 20814
rect 21758 20738 21810 20750
rect 30270 20802 30322 20814
rect 30270 20738 30322 20750
rect 4734 20690 4786 20702
rect 4734 20626 4786 20638
rect 5070 20690 5122 20702
rect 9650 20638 9662 20690
rect 9714 20638 9726 20690
rect 19170 20638 19182 20690
rect 19234 20638 19246 20690
rect 5070 20626 5122 20638
rect 15374 20578 15426 20590
rect 15374 20514 15426 20526
rect 15598 20578 15650 20590
rect 15598 20514 15650 20526
rect 16046 20578 16098 20590
rect 16046 20514 16098 20526
rect 21982 20578 22034 20590
rect 21982 20514 22034 20526
rect 672 20410 31024 20444
rect 672 20358 3806 20410
rect 3858 20358 3910 20410
rect 3962 20358 4014 20410
rect 4066 20358 23806 20410
rect 23858 20358 23910 20410
rect 23962 20358 24014 20410
rect 24066 20358 31024 20410
rect 672 20324 31024 20358
rect 14814 20242 14866 20254
rect 14814 20178 14866 20190
rect 20638 20242 20690 20254
rect 20638 20178 20690 20190
rect 1150 20130 1202 20142
rect 1150 20066 1202 20078
rect 17166 20130 17218 20142
rect 17166 20066 17218 20078
rect 17614 20130 17666 20142
rect 17614 20066 17666 20078
rect 20750 20130 20802 20142
rect 20750 20066 20802 20078
rect 6750 20018 6802 20030
rect 10110 20018 10162 20030
rect 1474 19966 1486 20018
rect 1538 19966 1550 20018
rect 2034 19966 2046 20018
rect 2098 19966 2110 20018
rect 3154 19966 3166 20018
rect 3218 19966 3230 20018
rect 3378 19966 3390 20018
rect 3442 19966 3454 20018
rect 4162 19966 4174 20018
rect 4226 19966 4238 20018
rect 5394 19966 5406 20018
rect 5458 19966 5470 20018
rect 5842 19966 5854 20018
rect 5906 19966 5918 20018
rect 7298 19966 7310 20018
rect 7362 19966 7374 20018
rect 8082 19966 8094 20018
rect 8146 19966 8158 20018
rect 8978 19966 8990 20018
rect 9042 19966 9054 20018
rect 9426 19966 9438 20018
rect 9490 19966 9502 20018
rect 10658 19966 10670 20018
rect 10722 19966 10734 20018
rect 11666 19966 11678 20018
rect 11730 19966 11742 20018
rect 13122 19966 13134 20018
rect 13186 19966 13198 20018
rect 15586 19966 15598 20018
rect 15650 19966 15662 20018
rect 18386 19966 18398 20018
rect 18450 19966 18462 20018
rect 6750 19954 6802 19966
rect 10110 19954 10162 19966
rect 2606 19906 2658 19918
rect 2606 19842 2658 19854
rect 5070 19906 5122 19918
rect 5070 19842 5122 19854
rect 8654 19906 8706 19918
rect 17726 19906 17778 19918
rect 13682 19854 13694 19906
rect 13746 19854 13758 19906
rect 16034 19854 16046 19906
rect 16098 19854 16110 19906
rect 8654 19842 8706 19854
rect 17726 19842 17778 19854
rect 19966 19906 20018 19918
rect 19966 19842 20018 19854
rect 2146 19742 2158 19794
rect 2210 19742 2222 19794
rect 6066 19742 6078 19794
rect 6130 19742 6142 19794
rect 9650 19742 9662 19794
rect 9714 19742 9726 19794
rect 18834 19742 18846 19794
rect 18898 19742 18910 19794
rect 672 19626 31024 19660
rect 672 19574 4466 19626
rect 4518 19574 4570 19626
rect 4622 19574 4674 19626
rect 4726 19574 24466 19626
rect 24518 19574 24570 19626
rect 24622 19574 24674 19626
rect 24726 19574 31024 19626
rect 672 19540 31024 19574
rect 8206 19458 8258 19470
rect 8206 19394 8258 19406
rect 15150 19458 15202 19470
rect 15150 19394 15202 19406
rect 16270 19458 16322 19470
rect 18510 19458 18562 19470
rect 17378 19406 17390 19458
rect 17442 19406 17454 19458
rect 16270 19394 16322 19406
rect 18510 19394 18562 19406
rect 19854 19458 19906 19470
rect 19854 19394 19906 19406
rect 19966 19458 20018 19470
rect 19966 19394 20018 19406
rect 30270 19458 30322 19470
rect 30270 19394 30322 19406
rect 1262 19346 1314 19358
rect 1934 19346 1986 19358
rect 11566 19346 11618 19358
rect 15710 19346 15762 19358
rect 1586 19294 1598 19346
rect 1650 19294 1662 19346
rect 2930 19294 2942 19346
rect 2994 19294 3006 19346
rect 5506 19294 5518 19346
rect 5570 19294 5582 19346
rect 7074 19294 7086 19346
rect 7138 19294 7150 19346
rect 9986 19294 9998 19346
rect 10050 19294 10062 19346
rect 12562 19294 12574 19346
rect 12626 19294 12638 19346
rect 1262 19282 1314 19294
rect 1934 19282 1986 19294
rect 11566 19282 11618 19294
rect 15710 19282 15762 19294
rect 15934 19346 15986 19358
rect 15934 19282 15986 19294
rect 16158 19346 16210 19358
rect 16158 19282 16210 19294
rect 20078 19346 20130 19358
rect 30594 19294 30606 19346
rect 30658 19294 30670 19346
rect 20078 19282 20130 19294
rect 11118 19234 11170 19246
rect 2370 19182 2382 19234
rect 2434 19182 2446 19234
rect 2706 19182 2718 19234
rect 2770 19182 2782 19234
rect 3490 19182 3502 19234
rect 3554 19182 3566 19234
rect 3938 19182 3950 19234
rect 4002 19182 4014 19234
rect 4946 19182 4958 19234
rect 5010 19182 5022 19234
rect 5730 19182 5742 19234
rect 5794 19182 5806 19234
rect 9538 19182 9550 19234
rect 9602 19182 9614 19234
rect 11890 19182 11902 19234
rect 11954 19182 11966 19234
rect 12338 19182 12350 19234
rect 12402 19182 12414 19234
rect 13122 19182 13134 19234
rect 13186 19182 13198 19234
rect 13570 19182 13582 19234
rect 13634 19182 13646 19234
rect 14578 19182 14590 19234
rect 14642 19182 14654 19234
rect 16930 19182 16942 19234
rect 16994 19182 17006 19234
rect 11118 19170 11170 19182
rect 15262 19122 15314 19134
rect 6626 19070 6638 19122
rect 6690 19070 6702 19122
rect 15262 19058 15314 19070
rect 672 18842 31024 18876
rect 672 18790 3806 18842
rect 3858 18790 3910 18842
rect 3962 18790 4014 18842
rect 4066 18790 23806 18842
rect 23858 18790 23910 18842
rect 23962 18790 24014 18842
rect 24066 18790 31024 18842
rect 672 18756 31024 18790
rect 16830 18674 16882 18686
rect 16830 18610 16882 18622
rect 17278 18674 17330 18686
rect 17278 18610 17330 18622
rect 18286 18674 18338 18686
rect 18286 18610 18338 18622
rect 8654 18562 8706 18574
rect 6626 18510 6638 18562
rect 6690 18510 6702 18562
rect 13010 18510 13022 18562
rect 13074 18510 13086 18562
rect 15250 18510 15262 18562
rect 15314 18510 15326 18562
rect 17490 18510 17502 18562
rect 17554 18510 17566 18562
rect 18050 18510 18062 18562
rect 18114 18510 18126 18562
rect 8654 18498 8706 18510
rect 3278 18450 3330 18462
rect 8206 18450 8258 18462
rect 1698 18398 1710 18450
rect 1762 18398 1774 18450
rect 4162 18398 4174 18450
rect 4226 18398 4238 18450
rect 3278 18386 3330 18398
rect 8206 18386 8258 18398
rect 8990 18450 9042 18462
rect 10670 18450 10722 18462
rect 14590 18450 14642 18462
rect 30270 18450 30322 18462
rect 9426 18398 9438 18450
rect 9490 18398 9502 18450
rect 9874 18398 9886 18450
rect 9938 18398 9950 18450
rect 10994 18398 11006 18450
rect 11058 18398 11070 18450
rect 12002 18398 12014 18450
rect 12066 18398 12078 18450
rect 17938 18398 17950 18450
rect 18002 18398 18014 18450
rect 8990 18386 9042 18398
rect 10670 18386 10722 18398
rect 14590 18386 14642 18398
rect 30270 18386 30322 18398
rect 17502 18338 17554 18350
rect 2146 18286 2158 18338
rect 2210 18286 2222 18338
rect 3938 18286 3950 18338
rect 4002 18286 4014 18338
rect 6962 18286 6974 18338
rect 7026 18286 7038 18338
rect 13458 18286 13470 18338
rect 13522 18286 13534 18338
rect 15586 18286 15598 18338
rect 15650 18286 15662 18338
rect 17502 18274 17554 18286
rect 5294 18226 5346 18238
rect 5966 18226 6018 18238
rect 4946 18174 4958 18226
rect 5010 18174 5022 18226
rect 5618 18174 5630 18226
rect 5682 18174 5694 18226
rect 9986 18174 9998 18226
rect 10050 18174 10062 18226
rect 30594 18174 30606 18226
rect 30658 18174 30670 18226
rect 5294 18162 5346 18174
rect 5966 18162 6018 18174
rect 672 18058 31024 18092
rect 672 18006 4466 18058
rect 4518 18006 4570 18058
rect 4622 18006 4674 18058
rect 4726 18006 24466 18058
rect 24518 18006 24570 18058
rect 24622 18006 24674 18058
rect 24726 18006 31024 18058
rect 672 17972 31024 18006
rect 1150 17890 1202 17902
rect 5518 17890 5570 17902
rect 2258 17838 2270 17890
rect 2322 17838 2334 17890
rect 1150 17826 1202 17838
rect 5518 17826 5570 17838
rect 7758 17890 7810 17902
rect 10670 17890 10722 17902
rect 13022 17890 13074 17902
rect 9538 17838 9550 17890
rect 9602 17838 9614 17890
rect 11890 17838 11902 17890
rect 11954 17838 11966 17890
rect 7758 17826 7810 17838
rect 10670 17826 10722 17838
rect 13022 17826 13074 17838
rect 13806 17890 13858 17902
rect 13806 17826 13858 17838
rect 16046 17890 16098 17902
rect 16046 17826 16098 17838
rect 16942 17890 16994 17902
rect 16942 17826 16994 17838
rect 30270 17890 30322 17902
rect 30270 17826 30322 17838
rect 13694 17778 13746 17790
rect 4274 17726 4286 17778
rect 4338 17726 4350 17778
rect 6626 17726 6638 17778
rect 6690 17726 6702 17778
rect 13694 17714 13746 17726
rect 13918 17778 13970 17790
rect 17054 17778 17106 17790
rect 18622 17778 18674 17790
rect 14914 17726 14926 17778
rect 14978 17726 14990 17778
rect 18274 17726 18286 17778
rect 18338 17726 18350 17778
rect 13918 17714 13970 17726
rect 17054 17714 17106 17726
rect 18622 17714 18674 17726
rect 18958 17778 19010 17790
rect 19954 17726 19966 17778
rect 20018 17726 20030 17778
rect 30594 17726 30606 17778
rect 30658 17726 30670 17778
rect 18958 17714 19010 17726
rect 20638 17666 20690 17678
rect 2706 17614 2718 17666
rect 2770 17614 2782 17666
rect 6178 17614 6190 17666
rect 6242 17614 6254 17666
rect 9090 17614 9102 17666
rect 9154 17614 9166 17666
rect 11330 17614 11342 17666
rect 11394 17614 11406 17666
rect 14466 17614 14478 17666
rect 14530 17614 14542 17666
rect 16706 17614 16718 17666
rect 16770 17614 16782 17666
rect 19394 17614 19406 17666
rect 19458 17614 19470 17666
rect 19730 17614 19742 17666
rect 19794 17614 19806 17666
rect 21186 17614 21198 17666
rect 21250 17614 21262 17666
rect 21970 17614 21982 17666
rect 22034 17614 22046 17666
rect 20638 17602 20690 17614
rect 3938 17502 3950 17554
rect 4002 17502 4014 17554
rect 672 17274 31024 17308
rect 672 17222 3806 17274
rect 3858 17222 3910 17274
rect 3962 17222 4014 17274
rect 4066 17222 23806 17274
rect 23858 17222 23910 17274
rect 23962 17222 24014 17274
rect 24066 17222 31024 17274
rect 672 17188 31024 17222
rect 1150 17106 1202 17118
rect 1150 17042 1202 17054
rect 6974 17106 7026 17118
rect 6974 17042 7026 17054
rect 9438 17106 9490 17118
rect 9438 17042 9490 17054
rect 12910 17106 12962 17118
rect 12910 17042 12962 17054
rect 19742 17106 19794 17118
rect 19742 17042 19794 17054
rect 2706 16942 2718 16994
rect 2770 16942 2782 16994
rect 5394 16942 5406 16994
rect 5458 16942 5470 16994
rect 7858 16942 7870 16994
rect 7922 16942 7934 16994
rect 11554 16942 11566 16994
rect 11618 16942 11630 16994
rect 4286 16882 4338 16894
rect 4286 16818 4338 16830
rect 9998 16882 10050 16894
rect 14578 16830 14590 16882
rect 14642 16830 14654 16882
rect 18050 16830 18062 16882
rect 18114 16830 18126 16882
rect 9998 16818 10050 16830
rect 2258 16718 2270 16770
rect 2322 16718 2334 16770
rect 3266 16718 3278 16770
rect 3330 16718 3342 16770
rect 3938 16718 3950 16770
rect 4002 16718 4014 16770
rect 5730 16718 5742 16770
rect 5794 16718 5806 16770
rect 8194 16718 8206 16770
rect 8258 16718 8270 16770
rect 14130 16718 14142 16770
rect 14194 16718 14206 16770
rect 18498 16718 18510 16770
rect 18562 16718 18574 16770
rect 3614 16658 3666 16670
rect 30270 16658 30322 16670
rect 11106 16606 11118 16658
rect 11170 16606 11182 16658
rect 30594 16606 30606 16658
rect 30658 16606 30670 16658
rect 3614 16594 3666 16606
rect 30270 16594 30322 16606
rect 672 16490 31024 16524
rect 672 16438 4466 16490
rect 4518 16438 4570 16490
rect 4622 16438 4674 16490
rect 4726 16438 24466 16490
rect 24518 16438 24570 16490
rect 24622 16438 24674 16490
rect 24726 16438 31024 16490
rect 672 16404 31024 16438
rect 3278 16322 3330 16334
rect 4958 16322 5010 16334
rect 7086 16322 7138 16334
rect 20974 16322 21026 16334
rect 2146 16270 2158 16322
rect 2210 16270 2222 16322
rect 4610 16270 4622 16322
rect 4674 16270 4686 16322
rect 5954 16270 5966 16322
rect 6018 16270 6030 16322
rect 7970 16270 7982 16322
rect 8034 16270 8046 16322
rect 9538 16270 9550 16322
rect 9602 16270 9614 16322
rect 16706 16270 16718 16322
rect 16770 16270 16782 16322
rect 19842 16270 19854 16322
rect 19906 16270 19918 16322
rect 3278 16258 3330 16270
rect 4958 16258 5010 16270
rect 7086 16258 7138 16270
rect 20974 16258 21026 16270
rect 30270 16322 30322 16334
rect 30270 16258 30322 16270
rect 11566 16210 11618 16222
rect 3938 16158 3950 16210
rect 4002 16158 4014 16210
rect 11218 16158 11230 16210
rect 11282 16158 11294 16210
rect 12898 16158 12910 16210
rect 12962 16158 12974 16210
rect 17378 16158 17390 16210
rect 17442 16158 17454 16210
rect 22642 16158 22654 16210
rect 22706 16158 22718 16210
rect 30594 16158 30606 16210
rect 30658 16158 30670 16210
rect 11566 16146 11618 16158
rect 4286 16098 4338 16110
rect 8318 16098 8370 16110
rect 17054 16098 17106 16110
rect 1698 16046 1710 16098
rect 1762 16046 1774 16098
rect 5506 16046 5518 16098
rect 5570 16046 5582 16098
rect 8978 16046 8990 16098
rect 9042 16046 9054 16098
rect 12226 16046 12238 16098
rect 12290 16046 12302 16098
rect 12786 16046 12798 16098
rect 12850 16046 12862 16098
rect 13458 16046 13470 16098
rect 13522 16046 13534 16098
rect 14018 16046 14030 16098
rect 14082 16046 14094 16098
rect 14914 16046 14926 16098
rect 14978 16046 14990 16098
rect 4286 16034 4338 16046
rect 8318 16034 8370 16046
rect 17054 16034 17106 16046
rect 17726 16098 17778 16110
rect 23090 16046 23102 16098
rect 23154 16046 23166 16098
rect 17726 16034 17778 16046
rect 11902 15986 11954 15998
rect 19394 15934 19406 15986
rect 19458 15934 19470 15986
rect 11902 15922 11954 15934
rect 10670 15874 10722 15886
rect 10670 15810 10722 15822
rect 21534 15874 21586 15886
rect 21534 15810 21586 15822
rect 672 15706 31024 15740
rect 672 15654 3806 15706
rect 3858 15654 3910 15706
rect 3962 15654 4014 15706
rect 4066 15654 23806 15706
rect 23858 15654 23910 15706
rect 23962 15654 24014 15706
rect 24066 15654 31024 15706
rect 672 15620 31024 15654
rect 2830 15538 2882 15550
rect 2830 15474 2882 15486
rect 5070 15538 5122 15550
rect 5070 15474 5122 15486
rect 1250 15374 1262 15426
rect 1314 15374 1326 15426
rect 6626 15374 6638 15426
rect 6690 15374 6702 15426
rect 14466 15374 14478 15426
rect 14530 15374 14542 15426
rect 21186 15374 21198 15426
rect 21250 15374 21262 15426
rect 3614 15314 3666 15326
rect 10110 15314 10162 15326
rect 8754 15262 8766 15314
rect 8818 15262 8830 15314
rect 9314 15262 9326 15314
rect 9378 15262 9390 15314
rect 10658 15262 10670 15314
rect 10722 15262 10734 15314
rect 11554 15262 11566 15314
rect 11618 15262 11630 15314
rect 15922 15262 15934 15314
rect 15986 15262 15998 15314
rect 18050 15262 18062 15314
rect 18114 15262 18126 15314
rect 30370 15262 30382 15314
rect 30434 15262 30446 15314
rect 3614 15250 3666 15262
rect 10110 15250 10162 15262
rect 4398 15202 4450 15214
rect 1586 15150 1598 15202
rect 1650 15150 1662 15202
rect 3266 15150 3278 15202
rect 3330 15150 3342 15202
rect 4050 15150 4062 15202
rect 4114 15150 4126 15202
rect 4398 15138 4450 15150
rect 8430 15202 8482 15214
rect 12910 15202 12962 15214
rect 9426 15150 9438 15202
rect 9490 15150 9502 15202
rect 14018 15150 14030 15202
rect 14082 15150 14094 15202
rect 15026 15150 15038 15202
rect 15090 15150 15102 15202
rect 16258 15150 16270 15202
rect 16322 15150 16334 15202
rect 18610 15150 18622 15202
rect 18674 15150 18686 15202
rect 21634 15150 21646 15202
rect 21698 15150 21710 15202
rect 8430 15138 8482 15150
rect 12910 15138 12962 15150
rect 8094 15090 8146 15102
rect 6178 15038 6190 15090
rect 6242 15038 6254 15090
rect 7746 15038 7758 15090
rect 7810 15038 7822 15090
rect 8094 15026 8146 15038
rect 15374 15090 15426 15102
rect 15374 15026 15426 15038
rect 17502 15090 17554 15102
rect 17502 15026 17554 15038
rect 19742 15090 19794 15102
rect 19742 15026 19794 15038
rect 22766 15090 22818 15102
rect 30594 15038 30606 15090
rect 30658 15038 30670 15090
rect 22766 15026 22818 15038
rect 672 14922 31024 14956
rect 672 14870 4466 14922
rect 4518 14870 4570 14922
rect 4622 14870 4674 14922
rect 4726 14870 24466 14922
rect 24518 14870 24570 14922
rect 24622 14870 24674 14922
rect 24726 14870 31024 14922
rect 672 14836 31024 14870
rect 12462 14754 12514 14766
rect 30270 14754 30322 14766
rect 6066 14702 6078 14754
rect 6130 14702 6142 14754
rect 13906 14702 13918 14754
rect 13970 14702 13982 14754
rect 17714 14702 17726 14754
rect 17778 14702 17790 14754
rect 12462 14690 12514 14702
rect 30270 14690 30322 14702
rect 5070 14642 5122 14654
rect 3714 14590 3726 14642
rect 3778 14590 3790 14642
rect 8866 14590 8878 14642
rect 8930 14590 8942 14642
rect 9538 14590 9550 14642
rect 9602 14590 9614 14642
rect 11330 14590 11342 14642
rect 11394 14590 11406 14642
rect 21746 14590 21758 14642
rect 21810 14590 21822 14642
rect 30594 14590 30606 14642
rect 30658 14590 30670 14642
rect 5070 14578 5122 14590
rect 3278 14530 3330 14542
rect 9886 14530 9938 14542
rect 14590 14530 14642 14542
rect 18174 14530 18226 14542
rect 22430 14530 22482 14542
rect 1698 14478 1710 14530
rect 1762 14478 1774 14530
rect 2706 14478 2718 14530
rect 2770 14478 2782 14530
rect 3826 14478 3838 14530
rect 3890 14478 3902 14530
rect 4386 14478 4398 14530
rect 4450 14478 4462 14530
rect 5506 14478 5518 14530
rect 5570 14478 5582 14530
rect 5842 14478 5854 14530
rect 5906 14478 5918 14530
rect 6626 14478 6638 14530
rect 6690 14478 6702 14530
rect 7298 14478 7310 14530
rect 7362 14478 7374 14530
rect 8082 14478 8094 14530
rect 8146 14478 8158 14530
rect 9090 14478 9102 14530
rect 9154 14478 9166 14530
rect 13346 14478 13358 14530
rect 13410 14478 13422 14530
rect 13682 14478 13694 14530
rect 13746 14478 13758 14530
rect 15026 14478 15038 14530
rect 15090 14478 15102 14530
rect 15922 14478 15934 14530
rect 15986 14478 15998 14530
rect 17154 14478 17166 14530
rect 17218 14478 17230 14530
rect 17490 14478 17502 14530
rect 17554 14478 17566 14530
rect 18722 14478 18734 14530
rect 18786 14478 18798 14530
rect 19730 14478 19742 14530
rect 19794 14478 19806 14530
rect 21074 14478 21086 14530
rect 21138 14478 21150 14530
rect 21522 14478 21534 14530
rect 21586 14478 21598 14530
rect 22754 14478 22766 14530
rect 22818 14478 22830 14530
rect 23762 14478 23774 14530
rect 23826 14478 23838 14530
rect 3278 14466 3330 14478
rect 9886 14466 9938 14478
rect 14590 14466 14642 14478
rect 18174 14466 18226 14478
rect 22430 14466 22482 14478
rect 4734 14418 4786 14430
rect 12910 14418 12962 14430
rect 10882 14366 10894 14418
rect 10946 14366 10958 14418
rect 4734 14354 4786 14366
rect 12910 14354 12962 14366
rect 16718 14418 16770 14430
rect 16718 14354 16770 14366
rect 20750 14418 20802 14430
rect 20750 14354 20802 14366
rect 672 14138 31024 14172
rect 672 14086 3806 14138
rect 3858 14086 3910 14138
rect 3962 14086 4014 14138
rect 4066 14086 23806 14138
rect 23858 14086 23910 14138
rect 23962 14086 24014 14138
rect 24066 14086 31024 14138
rect 672 14052 31024 14086
rect 7870 13970 7922 13982
rect 7870 13906 7922 13918
rect 15038 13970 15090 13982
rect 15038 13906 15090 13918
rect 18174 13970 18226 13982
rect 18174 13906 18226 13918
rect 8318 13858 8370 13870
rect 8318 13794 8370 13806
rect 30158 13858 30210 13870
rect 30158 13794 30210 13806
rect 5294 13746 5346 13758
rect 9998 13746 10050 13758
rect 22206 13746 22258 13758
rect 1250 13694 1262 13746
rect 1314 13694 1326 13746
rect 2258 13694 2270 13746
rect 2322 13694 2334 13746
rect 3490 13694 3502 13746
rect 3554 13694 3566 13746
rect 4050 13694 4062 13746
rect 4114 13694 4126 13746
rect 6290 13694 6302 13746
rect 6354 13694 6366 13746
rect 8642 13694 8654 13746
rect 8706 13694 8718 13746
rect 9090 13694 9102 13746
rect 9154 13694 9166 13746
rect 10322 13694 10334 13746
rect 10386 13694 10398 13746
rect 11330 13694 11342 13746
rect 11394 13694 11406 13746
rect 13458 13694 13470 13746
rect 13522 13694 13534 13746
rect 16594 13694 16606 13746
rect 16658 13694 16670 13746
rect 21186 13694 21198 13746
rect 21250 13694 21262 13746
rect 21522 13694 21534 13746
rect 21586 13694 21598 13746
rect 22754 13694 22766 13746
rect 22818 13694 22830 13746
rect 23762 13694 23774 13746
rect 23826 13694 23838 13746
rect 5294 13682 5346 13694
rect 9998 13682 10050 13694
rect 22206 13682 22258 13694
rect 2942 13634 2994 13646
rect 2942 13570 2994 13582
rect 4398 13634 4450 13646
rect 12238 13634 12290 13646
rect 20750 13634 20802 13646
rect 4946 13582 4958 13634
rect 5010 13582 5022 13634
rect 6738 13582 6750 13634
rect 6802 13582 6814 13634
rect 9314 13582 9326 13634
rect 9378 13582 9390 13634
rect 11890 13582 11902 13634
rect 11954 13582 11966 13634
rect 13906 13582 13918 13634
rect 13970 13582 13982 13634
rect 16930 13582 16942 13634
rect 16994 13582 17006 13634
rect 21746 13582 21758 13634
rect 21810 13582 21822 13634
rect 4398 13570 4450 13582
rect 12238 13570 12290 13582
rect 20750 13570 20802 13582
rect 3378 13470 3390 13522
rect 3442 13470 3454 13522
rect 672 13354 31024 13388
rect 672 13302 4466 13354
rect 4518 13302 4570 13354
rect 4622 13302 4674 13354
rect 4726 13302 24466 13354
rect 24518 13302 24570 13354
rect 24622 13302 24674 13354
rect 24726 13302 31024 13354
rect 672 13268 31024 13302
rect 8878 13186 8930 13198
rect 8878 13122 8930 13134
rect 11902 13186 11954 13198
rect 14142 13186 14194 13198
rect 21422 13186 21474 13198
rect 13010 13134 13022 13186
rect 13074 13134 13086 13186
rect 18722 13134 18734 13186
rect 18786 13134 18798 13186
rect 11902 13122 11954 13134
rect 14142 13122 14194 13134
rect 21422 13122 21474 13134
rect 30270 13186 30322 13198
rect 30270 13122 30322 13134
rect 5070 13074 5122 13086
rect 17726 13074 17778 13086
rect 3714 13022 3726 13074
rect 3778 13022 3790 13074
rect 6066 13022 6078 13074
rect 6130 13022 6142 13074
rect 9202 13022 9214 13074
rect 9266 13022 9278 13074
rect 10770 13022 10782 13074
rect 10834 13022 10846 13074
rect 17042 13022 17054 13074
rect 17106 13022 17118 13074
rect 22530 13022 22542 13074
rect 22594 13022 22606 13074
rect 30594 13022 30606 13074
rect 30658 13022 30670 13074
rect 5070 13010 5122 13022
rect 17726 13010 17778 13022
rect 3054 12962 3106 12974
rect 6750 12962 6802 12974
rect 17390 12962 17442 12974
rect 19406 12962 19458 12974
rect 1698 12910 1710 12962
rect 1762 12910 1774 12962
rect 2482 12910 2494 12962
rect 2546 12910 2558 12962
rect 3938 12910 3950 12962
rect 4002 12910 4014 12962
rect 4386 12910 4398 12962
rect 4450 12910 4462 12962
rect 5394 12910 5406 12962
rect 5458 12910 5470 12962
rect 5842 12910 5854 12962
rect 5906 12910 5918 12962
rect 7074 12910 7086 12962
rect 7138 12910 7150 12962
rect 8082 12910 8094 12962
rect 8146 12910 8158 12962
rect 18162 12910 18174 12962
rect 18226 12910 18238 12962
rect 18610 12910 18622 12962
rect 18674 12910 18686 12962
rect 19954 12910 19966 12962
rect 20018 12910 20030 12962
rect 20738 12910 20750 12962
rect 20802 12910 20814 12962
rect 3054 12898 3106 12910
rect 6750 12898 6802 12910
rect 17390 12898 17442 12910
rect 19406 12898 19458 12910
rect 4734 12850 4786 12862
rect 10322 12798 10334 12850
rect 10386 12798 10398 12850
rect 12562 12798 12574 12850
rect 12626 12798 12638 12850
rect 22978 12798 22990 12850
rect 23042 12798 23054 12850
rect 4734 12786 4786 12798
rect 672 12570 31024 12604
rect 672 12518 3806 12570
rect 3858 12518 3910 12570
rect 3962 12518 4014 12570
rect 4066 12518 23806 12570
rect 23858 12518 23910 12570
rect 23962 12518 24014 12570
rect 24066 12518 31024 12570
rect 672 12484 31024 12518
rect 3390 12402 3442 12414
rect 3390 12338 3442 12350
rect 7870 12402 7922 12414
rect 7870 12338 7922 12350
rect 10110 12402 10162 12414
rect 10110 12338 10162 12350
rect 18286 12402 18338 12414
rect 18286 12338 18338 12350
rect 20750 12402 20802 12414
rect 20750 12338 20802 12350
rect 14466 12238 14478 12290
rect 14530 12238 14542 12290
rect 11230 12178 11282 12190
rect 1810 12126 1822 12178
rect 1874 12126 1886 12178
rect 6290 12126 6302 12178
rect 6354 12126 6366 12178
rect 8418 12126 8430 12178
rect 8482 12126 8494 12178
rect 12114 12126 12126 12178
rect 12178 12126 12190 12178
rect 16706 12126 16718 12178
rect 16770 12126 16782 12178
rect 22418 12126 22430 12178
rect 22482 12126 22494 12178
rect 30370 12126 30382 12178
rect 30434 12126 30446 12178
rect 11230 12114 11282 12126
rect 10894 12066 10946 12078
rect 2258 12014 2270 12066
rect 2322 12014 2334 12066
rect 4946 12014 4958 12066
rect 5010 12014 5022 12066
rect 14018 12014 14030 12066
rect 14082 12014 14094 12066
rect 10894 12002 10946 12014
rect 4174 11954 4226 11966
rect 3826 11902 3838 11954
rect 3890 11902 3902 11954
rect 4174 11890 4226 11902
rect 5294 11954 5346 11966
rect 12910 11954 12962 11966
rect 6738 11902 6750 11954
rect 6802 11902 6814 11954
rect 8978 11902 8990 11954
rect 9042 11902 9054 11954
rect 10546 11902 10558 11954
rect 10610 11902 10622 11954
rect 11554 11902 11566 11954
rect 11618 11902 11630 11954
rect 11890 11902 11902 11954
rect 11954 11902 11966 11954
rect 17154 11902 17166 11954
rect 17218 11902 17230 11954
rect 21858 11902 21870 11954
rect 21922 11902 21934 11954
rect 30594 11902 30606 11954
rect 30658 11902 30670 11954
rect 5294 11890 5346 11902
rect 12910 11890 12962 11902
rect 672 11786 31024 11820
rect 672 11734 4466 11786
rect 4518 11734 4570 11786
rect 4622 11734 4674 11786
rect 4726 11734 24466 11786
rect 24518 11734 24570 11786
rect 24622 11734 24674 11786
rect 24726 11734 31024 11786
rect 672 11700 31024 11734
rect 2830 11618 2882 11630
rect 2830 11554 2882 11566
rect 3390 11618 3442 11630
rect 3390 11554 3442 11566
rect 7310 11618 7362 11630
rect 30270 11618 30322 11630
rect 11442 11566 11454 11618
rect 11506 11566 11518 11618
rect 19170 11566 19182 11618
rect 19234 11566 19246 11618
rect 7310 11554 7362 11566
rect 30270 11554 30322 11566
rect 18174 11506 18226 11518
rect 1586 11454 1598 11506
rect 1650 11454 1662 11506
rect 4610 11454 4622 11506
rect 4674 11454 4686 11506
rect 6066 11454 6078 11506
rect 6130 11454 6142 11506
rect 7746 11454 7758 11506
rect 7810 11454 7822 11506
rect 8866 11454 8878 11506
rect 8930 11454 8942 11506
rect 10098 11454 10110 11506
rect 10162 11454 10174 11506
rect 13906 11454 13918 11506
rect 13970 11454 13982 11506
rect 30594 11454 30606 11506
rect 30658 11454 30670 11506
rect 18174 11442 18226 11454
rect 8094 11394 8146 11406
rect 10446 11394 10498 11406
rect 4946 11342 4958 11394
rect 5010 11342 5022 11394
rect 9090 11342 9102 11394
rect 9154 11342 9166 11394
rect 10994 11342 11006 11394
rect 11058 11342 11070 11394
rect 13458 11342 13470 11394
rect 13522 11342 13534 11394
rect 18498 11342 18510 11394
rect 18562 11342 18574 11394
rect 18946 11342 18958 11394
rect 19010 11342 19022 11394
rect 19730 11342 19742 11394
rect 19794 11342 19806 11394
rect 20402 11342 20414 11394
rect 20466 11342 20478 11394
rect 21186 11342 21198 11394
rect 21250 11342 21262 11394
rect 8094 11330 8146 11342
rect 10446 11330 10498 11342
rect 1250 11230 1262 11282
rect 1314 11230 1326 11282
rect 5730 11230 5742 11282
rect 5794 11230 5806 11282
rect 12574 11170 12626 11182
rect 12574 11106 12626 11118
rect 15038 11170 15090 11182
rect 15038 11106 15090 11118
rect 672 11002 31024 11036
rect 672 10950 3806 11002
rect 3858 10950 3910 11002
rect 3962 10950 4014 11002
rect 4066 10950 23806 11002
rect 23858 10950 23910 11002
rect 23962 10950 24014 11002
rect 24066 10950 31024 11002
rect 672 10916 31024 10950
rect 2830 10834 2882 10846
rect 2830 10770 2882 10782
rect 7198 10834 7250 10846
rect 7198 10770 7250 10782
rect 18510 10834 18562 10846
rect 18510 10770 18562 10782
rect 1250 10670 1262 10722
rect 1314 10670 1326 10722
rect 3490 10558 3502 10610
rect 3554 10558 3566 10610
rect 4162 10558 4174 10610
rect 4226 10558 4238 10610
rect 5618 10558 5630 10610
rect 5682 10558 5694 10610
rect 8754 10558 8766 10610
rect 8818 10558 8830 10610
rect 9650 10558 9662 10610
rect 9714 10558 9726 10610
rect 10994 10558 11006 10610
rect 11058 10558 11070 10610
rect 11554 10558 11566 10610
rect 11618 10558 11630 10610
rect 13010 10558 13022 10610
rect 13074 10558 13086 10610
rect 13682 10558 13694 10610
rect 13746 10558 13758 10610
rect 16930 10558 16942 10610
rect 16994 10558 17006 10610
rect 22306 10558 22318 10610
rect 22370 10558 22382 10610
rect 10446 10498 10498 10510
rect 11902 10498 11954 10510
rect 20750 10498 20802 10510
rect 1586 10446 1598 10498
rect 1650 10446 1662 10498
rect 3938 10446 3950 10498
rect 4002 10446 4014 10498
rect 5954 10446 5966 10498
rect 6018 10446 6030 10498
rect 7634 10446 7646 10498
rect 7698 10446 7710 10498
rect 10882 10446 10894 10498
rect 10946 10446 10958 10498
rect 12786 10446 12798 10498
rect 12850 10446 12862 10498
rect 14130 10446 14142 10498
rect 14194 10446 14206 10498
rect 15698 10446 15710 10498
rect 15762 10446 15774 10498
rect 17266 10446 17278 10498
rect 17330 10446 17342 10498
rect 21858 10446 21870 10498
rect 21922 10446 21934 10498
rect 10446 10434 10498 10446
rect 11902 10434 11954 10446
rect 20750 10434 20802 10446
rect 7982 10386 8034 10398
rect 3266 10334 3278 10386
rect 3330 10334 3342 10386
rect 7982 10322 8034 10334
rect 15262 10386 15314 10398
rect 15262 10322 15314 10334
rect 16046 10386 16098 10398
rect 17378 10334 17390 10386
rect 17442 10334 17454 10386
rect 16046 10322 16098 10334
rect 672 10218 31024 10252
rect 672 10166 4466 10218
rect 4518 10166 4570 10218
rect 4622 10166 4674 10218
rect 4726 10166 24466 10218
rect 24518 10166 24570 10218
rect 24622 10166 24674 10218
rect 24726 10166 31024 10218
rect 672 10132 31024 10166
rect 1150 10050 1202 10062
rect 5966 10050 6018 10062
rect 14926 10050 14978 10062
rect 19742 10050 19794 10062
rect 2258 9998 2270 10050
rect 2322 9998 2334 10050
rect 10322 9998 10334 10050
rect 10386 9998 10398 10050
rect 12002 9998 12014 10050
rect 12066 9998 12078 10050
rect 16706 9998 16718 10050
rect 16770 9998 16782 10050
rect 21186 9998 21198 10050
rect 21250 9998 21262 10050
rect 1150 9986 1202 9998
rect 5966 9986 6018 9998
rect 14926 9986 14978 9998
rect 19742 9986 19794 9998
rect 4722 9886 4734 9938
rect 4786 9886 4798 9938
rect 7074 9886 7086 9938
rect 7138 9886 7150 9938
rect 8866 9886 8878 9938
rect 8930 9886 8942 9938
rect 9538 9886 9550 9938
rect 9602 9886 9614 9938
rect 14578 9886 14590 9938
rect 14642 9886 14654 9938
rect 15250 9886 15262 9938
rect 15314 9886 15326 9938
rect 18498 9886 18510 9938
rect 18562 9886 18574 9938
rect 10670 9826 10722 9838
rect 17054 9826 17106 9838
rect 21870 9826 21922 9838
rect 6514 9774 6526 9826
rect 6578 9774 6590 9826
rect 9090 9774 9102 9826
rect 9154 9774 9166 9826
rect 9762 9774 9774 9826
rect 9826 9774 9838 9826
rect 11330 9774 11342 9826
rect 11394 9774 11406 9826
rect 11778 9774 11790 9826
rect 11842 9774 11854 9826
rect 12562 9774 12574 9826
rect 12626 9774 12638 9826
rect 13010 9774 13022 9826
rect 13074 9774 13086 9826
rect 14018 9774 14030 9826
rect 14082 9774 14094 9826
rect 15474 9774 15486 9826
rect 15538 9774 15550 9826
rect 18050 9774 18062 9826
rect 18114 9774 18126 9826
rect 20626 9774 20638 9826
rect 20690 9774 20702 9826
rect 10670 9762 10722 9774
rect 17054 9762 17106 9774
rect 21074 9762 21086 9814
rect 21138 9762 21150 9814
rect 22194 9774 22206 9826
rect 22258 9774 22270 9826
rect 22418 9774 22430 9826
rect 22482 9774 22494 9826
rect 23314 9774 23326 9826
rect 23378 9774 23390 9826
rect 21870 9762 21922 9774
rect 11006 9714 11058 9726
rect 2706 9662 2718 9714
rect 2770 9662 2782 9714
rect 4386 9662 4398 9714
rect 4450 9662 4462 9714
rect 11006 9650 11058 9662
rect 20190 9714 20242 9726
rect 20190 9650 20242 9662
rect 8206 9602 8258 9614
rect 8206 9538 8258 9550
rect 672 9434 31024 9468
rect 672 9382 3806 9434
rect 3858 9382 3910 9434
rect 3962 9382 4014 9434
rect 4066 9382 23806 9434
rect 23858 9382 23910 9434
rect 23962 9382 24014 9434
rect 24066 9382 31024 9434
rect 672 9348 31024 9382
rect 4286 9266 4338 9278
rect 4286 9202 4338 9214
rect 22430 9266 22482 9278
rect 22430 9202 22482 9214
rect 13582 9154 13634 9166
rect 13582 9090 13634 9102
rect 17278 9154 17330 9166
rect 18834 9102 18846 9154
rect 18898 9102 18910 9154
rect 24546 9102 24558 9154
rect 24610 9102 24622 9154
rect 17278 9090 17330 9102
rect 1374 9042 1426 9054
rect 1374 8978 1426 8990
rect 2046 9042 2098 9054
rect 5294 9042 5346 9054
rect 2706 8990 2718 9042
rect 2770 8990 2782 9042
rect 2046 8978 2098 8990
rect 5294 8978 5346 8990
rect 5966 9042 6018 9054
rect 12126 9042 12178 9054
rect 6850 8990 6862 9042
rect 6914 8990 6926 9042
rect 7298 8990 7310 9042
rect 7362 8990 7374 9042
rect 8418 8990 8430 9042
rect 8482 8990 8494 9042
rect 9426 8990 9438 9042
rect 9490 8990 9502 9042
rect 10546 8990 10558 9042
rect 10610 8990 10622 9042
rect 13906 8990 13918 9042
rect 13970 8990 13982 9042
rect 14354 8990 14366 9042
rect 14418 8990 14430 9042
rect 15138 8990 15150 9042
rect 15202 8990 15214 9042
rect 15586 8990 15598 9042
rect 15650 8990 15662 9042
rect 16594 8990 16606 9042
rect 16658 8990 16670 9042
rect 20850 8990 20862 9042
rect 20914 8990 20926 9042
rect 5966 8978 6018 8990
rect 12126 8978 12178 8990
rect 6414 8930 6466 8942
rect 1026 8878 1038 8930
rect 1090 8878 1102 8930
rect 1698 8878 1710 8930
rect 1762 8878 1774 8930
rect 3154 8878 3166 8930
rect 3218 8878 3230 8930
rect 6414 8866 6466 8878
rect 7870 8930 7922 8942
rect 14578 8878 14590 8930
rect 14642 8878 14654 8930
rect 18498 8878 18510 8930
rect 18562 8878 18574 8930
rect 21186 8878 21198 8930
rect 21250 8878 21262 8930
rect 24098 8878 24110 8930
rect 24162 8878 24174 8930
rect 7870 8866 7922 8878
rect 12798 8818 12850 8830
rect 20078 8818 20130 8830
rect 4946 8766 4958 8818
rect 5010 8766 5022 8818
rect 5618 8766 5630 8818
rect 5682 8766 5694 8818
rect 7410 8766 7422 8818
rect 7474 8766 7486 8818
rect 10994 8766 11006 8818
rect 11058 8766 11070 8818
rect 13122 8766 13134 8818
rect 13186 8766 13198 8818
rect 19730 8766 19742 8818
rect 19794 8766 19806 8818
rect 12798 8754 12850 8766
rect 20078 8754 20130 8766
rect 22990 8818 23042 8830
rect 22990 8754 23042 8766
rect 672 8650 31024 8684
rect 672 8598 4466 8650
rect 4518 8598 4570 8650
rect 4622 8598 4674 8650
rect 4726 8598 24466 8650
rect 24518 8598 24570 8650
rect 24622 8598 24674 8650
rect 24726 8598 31024 8650
rect 672 8564 31024 8598
rect 11118 8482 11170 8494
rect 11118 8418 11170 8430
rect 20750 8482 20802 8494
rect 20750 8418 20802 8430
rect 7646 8370 7698 8382
rect 13022 8370 13074 8382
rect 15486 8370 15538 8382
rect 1026 8318 1038 8370
rect 1090 8318 1102 8370
rect 1810 8318 1822 8370
rect 1874 8318 1886 8370
rect 4050 8318 4062 8370
rect 4114 8318 4126 8370
rect 6626 8318 6638 8370
rect 6690 8318 6702 8370
rect 7298 8318 7310 8370
rect 7362 8318 7374 8370
rect 7970 8318 7982 8370
rect 8034 8318 8046 8370
rect 9986 8318 9998 8370
rect 10050 8318 10062 8370
rect 12562 8318 12574 8370
rect 12626 8318 12638 8370
rect 15138 8318 15150 8370
rect 15202 8318 15214 8370
rect 15810 8318 15822 8370
rect 15874 8318 15886 8370
rect 17938 8318 17950 8370
rect 18002 8318 18014 8370
rect 19506 8318 19518 8370
rect 19570 8318 19582 8370
rect 21746 8318 21758 8370
rect 21810 8318 21822 8370
rect 7646 8306 7698 8318
rect 13022 8306 13074 8318
rect 15486 8306 15538 8318
rect 1374 8258 1426 8270
rect 1374 8194 1426 8206
rect 2158 8258 2210 8270
rect 4734 8258 4786 8270
rect 6974 8258 7026 8270
rect 16158 8258 16210 8270
rect 3490 8206 3502 8258
rect 3554 8206 3566 8258
rect 3938 8206 3950 8258
rect 4002 8206 4014 8258
rect 5058 8206 5070 8258
rect 5122 8206 5134 8258
rect 6066 8206 6078 8258
rect 6130 8206 6142 8258
rect 8194 8206 8206 8258
rect 8258 8206 8270 8258
rect 11890 8206 11902 8258
rect 11954 8206 11966 8258
rect 12338 8206 12350 8258
rect 12402 8206 12414 8258
rect 13570 8206 13582 8258
rect 13634 8206 13646 8258
rect 14578 8206 14590 8258
rect 14642 8206 14654 8258
rect 18386 8206 18398 8258
rect 18450 8206 18462 8258
rect 19170 8206 19182 8258
rect 19234 8206 19246 8258
rect 2158 8194 2210 8206
rect 4734 8194 4786 8206
rect 6974 8194 7026 8206
rect 16158 8194 16210 8206
rect 3054 8146 3106 8158
rect 11566 8146 11618 8158
rect 9538 8094 9550 8146
rect 9602 8094 9614 8146
rect 21410 8094 21422 8146
rect 21474 8094 21486 8146
rect 3054 8082 3106 8094
rect 11566 8082 11618 8094
rect 16830 8034 16882 8046
rect 16830 7970 16882 7982
rect 22990 8034 23042 8046
rect 22990 7970 23042 7982
rect 672 7866 31024 7900
rect 672 7814 3806 7866
rect 3858 7814 3910 7866
rect 3962 7814 4014 7866
rect 4066 7814 23806 7866
rect 23858 7814 23910 7866
rect 23962 7814 24014 7866
rect 24066 7814 31024 7866
rect 672 7780 31024 7814
rect 3390 7698 3442 7710
rect 3390 7634 3442 7646
rect 12126 7698 12178 7710
rect 12126 7634 12178 7646
rect 6750 7586 6802 7598
rect 14590 7586 14642 7598
rect 19966 7586 20018 7598
rect 10546 7534 10558 7586
rect 10610 7534 10622 7586
rect 18386 7534 18398 7586
rect 18450 7534 18462 7586
rect 6750 7522 6802 7534
rect 14590 7522 14642 7534
rect 19966 7522 20018 7534
rect 20638 7586 20690 7598
rect 20638 7522 20690 7534
rect 5294 7474 5346 7486
rect 1810 7422 1822 7474
rect 1874 7422 1886 7474
rect 5730 7422 5742 7474
rect 5794 7422 5806 7474
rect 7186 7422 7198 7474
rect 7250 7422 7262 7474
rect 7634 7425 7646 7477
rect 7698 7425 7710 7477
rect 16270 7474 16322 7486
rect 22318 7474 22370 7486
rect 8754 7422 8766 7474
rect 8818 7422 8830 7474
rect 9762 7422 9774 7474
rect 9826 7422 9838 7474
rect 15026 7422 15038 7474
rect 15090 7422 15102 7474
rect 15362 7422 15374 7474
rect 15426 7422 15438 7474
rect 16706 7422 16718 7474
rect 16770 7422 16782 7474
rect 17602 7422 17614 7474
rect 17666 7422 17678 7474
rect 20962 7422 20974 7474
rect 21026 7422 21038 7474
rect 21410 7422 21422 7474
rect 21474 7422 21486 7474
rect 22866 7422 22878 7474
rect 22930 7422 22942 7474
rect 23650 7422 23662 7474
rect 23714 7422 23726 7474
rect 5294 7410 5346 7422
rect 16270 7410 16322 7422
rect 22318 7410 22370 7422
rect 8206 7362 8258 7374
rect 2258 7310 2270 7362
rect 2322 7310 2334 7362
rect 4946 7310 4958 7362
rect 5010 7310 5022 7362
rect 5954 7310 5966 7362
rect 6018 7310 6030 7362
rect 8206 7298 8258 7310
rect 13246 7362 13298 7374
rect 15586 7310 15598 7362
rect 15650 7310 15662 7362
rect 18834 7310 18846 7362
rect 18898 7310 18910 7362
rect 21634 7310 21646 7362
rect 21698 7310 21710 7362
rect 13246 7298 13298 7310
rect 13918 7250 13970 7262
rect 7746 7198 7758 7250
rect 7810 7198 7822 7250
rect 10994 7198 11006 7250
rect 11058 7198 11070 7250
rect 13570 7198 13582 7250
rect 13634 7198 13646 7250
rect 14242 7198 14254 7250
rect 14306 7198 14318 7250
rect 13918 7186 13970 7198
rect 672 7082 31024 7116
rect 672 7030 4466 7082
rect 4518 7030 4570 7082
rect 4622 7030 4674 7082
rect 4726 7030 24466 7082
rect 24518 7030 24570 7082
rect 24622 7030 24674 7082
rect 24726 7030 31024 7082
rect 672 6996 31024 7030
rect 6626 6862 6638 6914
rect 6690 6862 6702 6914
rect 8306 6862 8318 6914
rect 8370 6862 8382 6914
rect 11330 6862 11342 6914
rect 11394 6862 11406 6914
rect 13906 6862 13918 6914
rect 13970 6862 13982 6914
rect 3054 6802 3106 6814
rect 20078 6802 20130 6814
rect 1698 6750 1710 6802
rect 1762 6750 1774 6802
rect 2370 6750 2382 6802
rect 2434 6750 2446 6802
rect 4050 6750 4062 6802
rect 4114 6750 4126 6802
rect 7298 6750 7310 6802
rect 7362 6750 7374 6802
rect 8866 6750 8878 6802
rect 8930 6750 8942 6802
rect 10322 6750 10334 6802
rect 10386 6750 10398 6802
rect 19058 6750 19070 6802
rect 19122 6750 19134 6802
rect 21410 6750 21422 6802
rect 21474 6750 21486 6802
rect 3054 6738 3106 6750
rect 20078 6738 20130 6750
rect 1374 6690 1426 6702
rect 4734 6690 4786 6702
rect 6974 6690 7026 6702
rect 2146 6638 2158 6690
rect 2210 6638 2222 6690
rect 3378 6638 3390 6690
rect 3442 6638 3454 6690
rect 3938 6638 3950 6690
rect 4002 6638 4014 6690
rect 5058 6638 5070 6690
rect 5122 6638 5134 6690
rect 6066 6638 6078 6690
rect 6130 6638 6142 6690
rect 1374 6626 1426 6638
rect 4734 6626 4786 6638
rect 6974 6626 7026 6638
rect 7646 6690 7698 6702
rect 7646 6626 7698 6638
rect 7982 6690 8034 6702
rect 12462 6690 12514 6702
rect 14366 6690 14418 6702
rect 18622 6690 18674 6702
rect 22094 6690 22146 6702
rect 9090 6638 9102 6690
rect 9154 6638 9166 6690
rect 10098 6638 10110 6690
rect 10162 6638 10174 6690
rect 13346 6638 13358 6690
rect 13410 6638 13422 6690
rect 13682 6638 13694 6690
rect 13746 6638 13758 6690
rect 14914 6638 14926 6690
rect 14978 6638 14990 6690
rect 15922 6638 15934 6690
rect 15986 6638 15998 6690
rect 16930 6638 16942 6690
rect 16994 6638 17006 6690
rect 18050 6638 18062 6690
rect 18114 6638 18126 6690
rect 19170 6638 19182 6690
rect 19234 6638 19246 6690
rect 19730 6638 19742 6690
rect 19794 6638 19806 6690
rect 20738 6638 20750 6690
rect 20802 6638 20814 6690
rect 21298 6638 21310 6690
rect 21362 6638 21374 6690
rect 22418 6638 22430 6690
rect 22482 6638 22494 6690
rect 23426 6638 23438 6690
rect 23490 6638 23502 6690
rect 7982 6626 8034 6638
rect 12462 6626 12514 6638
rect 14366 6626 14418 6638
rect 18622 6626 18674 6638
rect 22094 6626 22146 6638
rect 12910 6578 12962 6590
rect 10882 6526 10894 6578
rect 10946 6526 10958 6578
rect 12910 6514 12962 6526
rect 20414 6578 20466 6590
rect 20414 6514 20466 6526
rect 672 6298 31024 6332
rect 672 6246 3806 6298
rect 3858 6246 3910 6298
rect 3962 6246 4014 6298
rect 4066 6246 23806 6298
rect 23858 6246 23910 6298
rect 23962 6246 24014 6298
rect 24066 6246 31024 6298
rect 672 6212 31024 6246
rect 20750 6130 20802 6142
rect 20750 6066 20802 6078
rect 22990 6130 23042 6142
rect 22990 6066 23042 6078
rect 10110 6018 10162 6030
rect 10110 5954 10162 5966
rect 14814 6018 14866 6030
rect 14814 5954 14866 5966
rect 3838 5906 3890 5918
rect 8430 5906 8482 5918
rect 1250 5854 1262 5906
rect 1314 5854 1326 5906
rect 2258 5854 2270 5906
rect 2322 5854 2334 5906
rect 5058 5854 5070 5906
rect 5122 5854 5134 5906
rect 6962 5854 6974 5906
rect 7026 5854 7038 5906
rect 7858 5854 7870 5906
rect 7922 5854 7934 5906
rect 9202 5854 9214 5906
rect 9266 5854 9278 5906
rect 9650 5854 9662 5906
rect 9714 5854 9726 5906
rect 12002 5854 12014 5906
rect 12066 5854 12078 5906
rect 13458 5854 13470 5906
rect 13522 5854 13534 5906
rect 14130 5854 14142 5906
rect 14194 5854 14206 5906
rect 15250 5854 15262 5906
rect 15314 5854 15326 5906
rect 15586 5854 15598 5906
rect 15650 5854 15662 5906
rect 16818 5854 16830 5906
rect 16882 5854 16894 5906
rect 17826 5854 17838 5906
rect 17890 5854 17902 5906
rect 18610 5854 18622 5906
rect 18674 5854 18686 5906
rect 19618 5854 19630 5906
rect 19682 5854 19694 5906
rect 22306 5854 22318 5906
rect 22370 5854 22382 5906
rect 24546 5854 24558 5906
rect 24610 5854 24622 5906
rect 25330 5854 25342 5906
rect 25394 5854 25406 5906
rect 3838 5842 3890 5854
rect 8430 5842 8482 5854
rect 16270 5794 16322 5806
rect 26910 5794 26962 5806
rect 1026 5742 1038 5794
rect 1090 5742 1102 5794
rect 5954 5742 5966 5794
rect 6018 5742 6030 5794
rect 9090 5742 9102 5794
rect 9154 5742 9166 5794
rect 12226 5742 12238 5794
rect 12290 5742 12302 5794
rect 15810 5742 15822 5794
rect 15874 5742 15886 5794
rect 19394 5742 19406 5794
rect 19458 5742 19470 5794
rect 21858 5742 21870 5794
rect 21922 5742 21934 5794
rect 24098 5742 24110 5794
rect 24162 5742 24174 5794
rect 25778 5742 25790 5794
rect 25842 5742 25854 5794
rect 16270 5730 16322 5742
rect 26910 5730 26962 5742
rect 5630 5682 5682 5694
rect 2706 5630 2718 5682
rect 2770 5630 2782 5682
rect 5282 5630 5294 5682
rect 5346 5630 5358 5682
rect 5630 5618 5682 5630
rect 10558 5682 10610 5694
rect 11230 5682 11282 5694
rect 10882 5630 10894 5682
rect 10946 5630 10958 5682
rect 11554 5630 11566 5682
rect 11618 5630 11630 5682
rect 13234 5630 13246 5682
rect 13298 5630 13310 5682
rect 13906 5630 13918 5682
rect 13970 5630 13982 5682
rect 18386 5630 18398 5682
rect 18450 5630 18462 5682
rect 10558 5618 10610 5630
rect 11230 5618 11282 5630
rect 672 5514 31024 5548
rect 672 5462 4466 5514
rect 4518 5462 4570 5514
rect 4622 5462 4674 5514
rect 4726 5462 24466 5514
rect 24518 5462 24570 5514
rect 24622 5462 24674 5514
rect 24726 5462 31024 5514
rect 672 5428 31024 5462
rect 1374 5346 1426 5358
rect 1026 5294 1038 5346
rect 1090 5294 1102 5346
rect 1374 5282 1426 5294
rect 2046 5346 2098 5358
rect 2046 5282 2098 5294
rect 2382 5346 2434 5358
rect 7086 5346 7138 5358
rect 2706 5294 2718 5346
rect 2770 5294 2782 5346
rect 5394 5294 5406 5346
rect 5458 5294 5470 5346
rect 2382 5282 2434 5294
rect 7086 5282 7138 5294
rect 7982 5346 8034 5358
rect 7982 5282 8034 5294
rect 10670 5346 10722 5358
rect 10670 5282 10722 5294
rect 15374 5346 15426 5358
rect 15374 5282 15426 5294
rect 18734 5346 18786 5358
rect 18734 5282 18786 5294
rect 23326 5346 23378 5358
rect 23326 5282 23378 5294
rect 23998 5346 24050 5358
rect 23998 5282 24050 5294
rect 24446 5346 24498 5358
rect 24446 5282 24498 5294
rect 26350 5346 26402 5358
rect 26350 5282 26402 5294
rect 4958 5234 5010 5246
rect 1698 5182 1710 5234
rect 1762 5182 1774 5234
rect 4958 5170 5010 5182
rect 6414 5234 6466 5246
rect 19406 5234 19458 5246
rect 25118 5234 25170 5246
rect 6738 5182 6750 5234
rect 6802 5182 6814 5234
rect 8306 5182 8318 5234
rect 8370 5182 8382 5234
rect 9538 5182 9550 5234
rect 9602 5182 9614 5234
rect 12226 5182 12238 5234
rect 12290 5182 12302 5234
rect 15026 5182 15038 5234
rect 15090 5182 15102 5234
rect 16146 5182 16158 5234
rect 16210 5182 16222 5234
rect 17490 5182 17502 5234
rect 17554 5182 17566 5234
rect 20402 5182 20414 5234
rect 20466 5182 20478 5234
rect 22978 5182 22990 5234
rect 23042 5182 23054 5234
rect 23650 5182 23662 5234
rect 23714 5182 23726 5234
rect 6414 5170 6466 5182
rect 19406 5170 19458 5182
rect 25118 5170 25170 5182
rect 11230 5122 11282 5134
rect 12686 5122 12738 5134
rect 15822 5122 15874 5134
rect 21086 5122 21138 5134
rect 3378 5070 3390 5122
rect 3442 5070 3454 5122
rect 4162 5070 4174 5122
rect 4226 5070 4238 5122
rect 5618 5070 5630 5122
rect 5682 5070 5694 5122
rect 6066 5070 6078 5122
rect 6130 5070 6142 5122
rect 11554 5070 11566 5122
rect 11618 5070 11630 5122
rect 12114 5070 12126 5122
rect 12178 5070 12190 5122
rect 13234 5070 13246 5122
rect 13298 5070 13310 5122
rect 14242 5070 14254 5122
rect 14306 5070 14318 5122
rect 19730 5070 19742 5122
rect 19794 5070 19806 5122
rect 20290 5070 20302 5122
rect 20354 5070 20366 5122
rect 21522 5070 21534 5122
rect 21586 5070 21598 5122
rect 22418 5070 22430 5122
rect 22482 5070 22494 5122
rect 11230 5058 11282 5070
rect 12686 5058 12738 5070
rect 15822 5058 15874 5070
rect 21086 5058 21138 5070
rect 9090 4958 9102 5010
rect 9154 4958 9166 5010
rect 17154 4958 17166 5010
rect 17218 4958 17230 5010
rect 672 4730 31024 4764
rect 672 4678 3806 4730
rect 3858 4678 3910 4730
rect 3962 4678 4014 4730
rect 4066 4678 23806 4730
rect 23858 4678 23910 4730
rect 23962 4678 24014 4730
rect 24066 4678 31024 4730
rect 672 4644 31024 4678
rect 4286 4562 4338 4574
rect 4286 4498 4338 4510
rect 15598 4562 15650 4574
rect 15598 4498 15650 4510
rect 17838 4562 17890 4574
rect 17838 4498 17890 4510
rect 22430 4562 22482 4574
rect 22430 4498 22482 4510
rect 22990 4562 23042 4574
rect 22990 4498 23042 4510
rect 10110 4450 10162 4462
rect 10110 4386 10162 4398
rect 1374 4338 1426 4350
rect 1374 4274 1426 4286
rect 2046 4338 2098 4350
rect 10558 4338 10610 4350
rect 2706 4286 2718 4338
rect 2770 4286 2782 4338
rect 5170 4286 5182 4338
rect 5234 4286 5246 4338
rect 6962 4286 6974 4338
rect 7026 4286 7038 4338
rect 7858 4286 7870 4338
rect 7922 4286 7934 4338
rect 9202 4286 9214 4338
rect 9266 4286 9278 4338
rect 9762 4286 9774 4338
rect 9826 4286 9838 4338
rect 2046 4274 2098 4286
rect 10558 4274 10610 4286
rect 11566 4338 11618 4350
rect 11566 4274 11618 4286
rect 12238 4338 12290 4350
rect 18286 4338 18338 4350
rect 13346 4286 13358 4338
rect 13410 4286 13422 4338
rect 14018 4286 14030 4338
rect 14082 4286 14094 4338
rect 16258 4286 16270 4338
rect 16322 4286 16334 4338
rect 12238 4274 12290 4286
rect 18286 4274 18338 4286
rect 19294 4338 19346 4350
rect 19294 4274 19346 4286
rect 19630 4338 19682 4350
rect 20850 4286 20862 4338
rect 20914 4286 20926 4338
rect 24658 4286 24670 4338
rect 24722 4286 24734 4338
rect 19630 4274 19682 4286
rect 8654 4226 8706 4238
rect 26350 4226 26402 4238
rect 1026 4174 1038 4226
rect 1090 4174 1102 4226
rect 1698 4174 1710 4226
rect 1762 4174 1774 4226
rect 3154 4174 3166 4226
rect 3218 4174 3230 4226
rect 5394 4174 5406 4226
rect 5458 4174 5470 4226
rect 6066 4174 6078 4226
rect 6130 4174 6142 4226
rect 9090 4174 9102 4226
rect 9154 4174 9166 4226
rect 10882 4174 10894 4226
rect 10946 4174 10958 4226
rect 11890 4174 11902 4226
rect 11954 4174 11966 4226
rect 16594 4174 16606 4226
rect 16658 4174 16670 4226
rect 18946 4174 18958 4226
rect 19010 4174 19022 4226
rect 19954 4174 19966 4226
rect 20018 4174 20030 4226
rect 21186 4174 21198 4226
rect 21250 4174 21262 4226
rect 24098 4174 24110 4226
rect 24162 4174 24174 4226
rect 25106 4174 25118 4226
rect 25170 4174 25182 4226
rect 8654 4162 8706 4174
rect 26350 4162 26402 4174
rect 5742 4114 5794 4126
rect 25454 4114 25506 4126
rect 11218 4062 11230 4114
rect 11282 4062 11294 4114
rect 13122 4062 13134 4114
rect 13186 4062 13198 4114
rect 14466 4062 14478 4114
rect 14530 4062 14542 4114
rect 18610 4062 18622 4114
rect 18674 4062 18686 4114
rect 5742 4050 5794 4062
rect 25454 4050 25506 4062
rect 672 3946 31024 3980
rect 672 3894 4466 3946
rect 4518 3894 4570 3946
rect 4622 3894 4674 3946
rect 4726 3894 24466 3946
rect 24518 3894 24570 3946
rect 24622 3894 24674 3946
rect 24726 3894 31024 3946
rect 672 3860 31024 3894
rect 1374 3778 1426 3790
rect 2046 3778 2098 3790
rect 1026 3726 1038 3778
rect 1090 3726 1102 3778
rect 1698 3726 1710 3778
rect 1762 3726 1774 3778
rect 1374 3714 1426 3726
rect 2046 3714 2098 3726
rect 2718 3778 2770 3790
rect 7310 3778 7362 3790
rect 10894 3778 10946 3790
rect 21422 3778 21474 3790
rect 23550 3778 23602 3790
rect 5394 3726 5406 3778
rect 5458 3726 5470 3778
rect 7634 3726 7646 3778
rect 7698 3726 7710 3778
rect 9762 3726 9774 3778
rect 9826 3726 9838 3778
rect 13570 3726 13582 3778
rect 13634 3726 13646 3778
rect 15810 3726 15822 3778
rect 15874 3726 15886 3778
rect 17042 3726 17054 3778
rect 17106 3726 17118 3778
rect 18722 3726 18734 3778
rect 18786 3726 18798 3778
rect 22530 3726 22542 3778
rect 22594 3726 22606 3778
rect 2718 3714 2770 3726
rect 7310 3714 7362 3726
rect 10894 3714 10946 3726
rect 21422 3714 21474 3726
rect 23550 3714 23602 3726
rect 24558 3778 24610 3790
rect 25566 3778 25618 3790
rect 24882 3726 24894 3778
rect 24946 3726 24958 3778
rect 24558 3714 24610 3726
rect 4958 3666 5010 3678
rect 2370 3614 2382 3666
rect 2434 3614 2446 3666
rect 4958 3602 5010 3614
rect 6414 3666 6466 3678
rect 17726 3666 17778 3678
rect 25218 3670 25230 3722
rect 25282 3670 25294 3722
rect 25566 3714 25618 3726
rect 26238 3778 26290 3790
rect 26562 3726 26574 3778
rect 26626 3726 26638 3778
rect 26238 3714 26290 3726
rect 8306 3614 8318 3666
rect 8370 3614 8382 3666
rect 15474 3614 15486 3666
rect 15538 3614 15550 3666
rect 23874 3614 23886 3666
rect 23938 3614 23950 3666
rect 25890 3614 25902 3666
rect 25954 3614 25966 3666
rect 6414 3602 6466 3614
rect 17726 3602 17778 3614
rect 3378 3502 3390 3554
rect 3442 3502 3454 3554
rect 4162 3502 4174 3554
rect 4226 3502 4238 3554
rect 5618 3502 5630 3554
rect 5682 3502 5694 3554
rect 6066 3502 6078 3554
rect 6130 3502 6142 3554
rect 8082 3502 8094 3554
rect 8146 3502 8158 3554
rect 11442 3507 11454 3559
rect 11506 3507 11518 3559
rect 12910 3554 12962 3566
rect 14590 3554 14642 3566
rect 12338 3502 12350 3554
rect 12402 3502 12414 3554
rect 13682 3502 13694 3554
rect 13746 3502 13758 3554
rect 14242 3502 14254 3554
rect 14306 3502 14318 3554
rect 12910 3490 12962 3502
rect 14590 3490 14642 3502
rect 15150 3554 15202 3566
rect 19182 3554 19234 3566
rect 16034 3502 16046 3554
rect 16098 3502 16110 3554
rect 16818 3502 16830 3554
rect 16882 3502 16894 3554
rect 18162 3502 18174 3554
rect 18226 3502 18238 3554
rect 18498 3502 18510 3554
rect 18562 3502 18574 3554
rect 19954 3502 19966 3554
rect 20018 3502 20030 3554
rect 20738 3502 20750 3554
rect 20802 3502 20814 3554
rect 26786 3502 26798 3554
rect 26850 3502 26862 3554
rect 15150 3490 15202 3502
rect 19182 3490 19234 3502
rect 9314 3390 9326 3442
rect 9378 3390 9390 3442
rect 22978 3390 22990 3442
rect 23042 3390 23054 3442
rect 672 3162 31024 3196
rect 672 3110 3806 3162
rect 3858 3110 3910 3162
rect 3962 3110 4014 3162
rect 4066 3110 23806 3162
rect 23858 3110 23910 3162
rect 23962 3110 24014 3162
rect 24066 3110 31024 3162
rect 672 3076 31024 3110
rect 3390 2994 3442 3006
rect 3390 2930 3442 2942
rect 6862 2994 6914 3006
rect 6862 2930 6914 2942
rect 15262 2994 15314 3006
rect 15262 2930 15314 2942
rect 18174 2994 18226 3006
rect 18174 2930 18226 2942
rect 20750 2994 20802 3006
rect 20750 2930 20802 2942
rect 22990 2994 23042 3006
rect 22990 2930 23042 2942
rect 10894 2882 10946 2894
rect 10894 2818 10946 2830
rect 11230 2882 11282 2894
rect 13682 2830 13694 2882
rect 13746 2830 13758 2882
rect 16594 2830 16606 2882
rect 16658 2830 16670 2882
rect 24546 2830 24558 2882
rect 24610 2830 24622 2882
rect 11230 2818 11282 2830
rect 3838 2770 3890 2782
rect 9438 2770 9490 2782
rect 15710 2770 15762 2782
rect 1698 2718 1710 2770
rect 1762 2718 1774 2770
rect 5282 2718 5294 2770
rect 5346 2718 5358 2770
rect 7746 2718 7758 2770
rect 7810 2718 7822 2770
rect 8642 2718 8654 2770
rect 8706 2718 8718 2770
rect 10098 2718 10110 2770
rect 10162 2718 10174 2770
rect 10546 2718 10558 2770
rect 10610 2718 10622 2770
rect 12002 2718 12014 2770
rect 12066 2718 12078 2770
rect 13010 2718 13022 2770
rect 13074 2718 13086 2770
rect 3838 2706 3890 2718
rect 9438 2706 9490 2718
rect 15710 2706 15762 2718
rect 18622 2770 18674 2782
rect 18622 2706 18674 2718
rect 19630 2770 19682 2782
rect 25454 2770 25506 2782
rect 22306 2718 22318 2770
rect 22370 2718 22382 2770
rect 19630 2706 19682 2718
rect 25454 2706 25506 2718
rect 26126 2770 26178 2782
rect 26674 2718 26686 2770
rect 26738 2718 26750 2770
rect 27346 2718 27358 2770
rect 27410 2718 27422 2770
rect 26126 2706 26178 2718
rect 2146 2606 2158 2658
rect 2210 2606 2222 2658
rect 4162 2606 4174 2658
rect 4226 2606 4238 2658
rect 5730 2606 5742 2658
rect 5794 2606 5806 2658
rect 9874 2606 9886 2658
rect 9938 2606 9950 2658
rect 12786 2606 12798 2658
rect 12850 2606 12862 2658
rect 14018 2606 14030 2658
rect 14082 2606 14094 2658
rect 16034 2606 16046 2658
rect 16098 2606 16110 2658
rect 17042 2606 17054 2658
rect 17106 2606 17118 2658
rect 18946 2606 18958 2658
rect 19010 2606 19022 2658
rect 11566 2546 11618 2558
rect 12226 2494 12238 2546
rect 12290 2494 12302 2546
rect 19282 2494 19294 2546
rect 19346 2494 19358 2546
rect 21858 2494 21870 2546
rect 21922 2494 21934 2546
rect 24098 2494 24110 2546
rect 24162 2494 24174 2546
rect 25106 2494 25118 2546
rect 25170 2494 25182 2546
rect 25778 2494 25790 2546
rect 25842 2494 25854 2546
rect 26450 2494 26462 2546
rect 26514 2494 26526 2546
rect 27122 2494 27134 2546
rect 27186 2494 27198 2546
rect 11566 2482 11618 2494
rect 672 2378 31024 2412
rect 672 2326 4466 2378
rect 4518 2326 4570 2378
rect 4622 2326 4674 2378
rect 4726 2326 24466 2378
rect 24518 2326 24570 2378
rect 24622 2326 24674 2378
rect 24726 2326 31024 2378
rect 672 2292 31024 2326
rect 1150 2210 1202 2222
rect 1822 2210 1874 2222
rect 4958 2210 5010 2222
rect 7198 2210 7250 2222
rect 1474 2158 1486 2210
rect 1538 2158 1550 2210
rect 2482 2158 2494 2210
rect 2546 2158 2558 2210
rect 6066 2158 6078 2210
rect 6130 2158 6142 2210
rect 1150 2146 1202 2158
rect 1822 2146 1874 2158
rect 4958 2146 5010 2158
rect 7198 2146 7250 2158
rect 7982 2210 8034 2222
rect 9214 2210 9266 2222
rect 8306 2158 8318 2210
rect 8370 2158 8382 2210
rect 7982 2146 8034 2158
rect 9214 2146 9266 2158
rect 11678 2210 11730 2222
rect 11678 2146 11730 2158
rect 13918 2210 13970 2222
rect 15374 2210 15426 2222
rect 15026 2158 15038 2210
rect 15090 2158 15102 2210
rect 13918 2146 13970 2158
rect 15374 2146 15426 2158
rect 15710 2210 15762 2222
rect 19294 2210 19346 2222
rect 21534 2210 21586 2222
rect 18162 2158 18174 2210
rect 18226 2158 18238 2210
rect 20402 2158 20414 2210
rect 20466 2158 20478 2210
rect 15710 2146 15762 2158
rect 19294 2146 19346 2158
rect 21534 2146 21586 2158
rect 22094 2210 22146 2222
rect 22094 2146 22146 2158
rect 24670 2210 24722 2222
rect 24670 2146 24722 2158
rect 27806 2210 27858 2222
rect 27806 2146 27858 2158
rect 28478 2210 28530 2222
rect 28478 2146 28530 2158
rect 7646 2098 7698 2110
rect 17166 2098 17218 2110
rect 2146 2046 2158 2098
rect 2210 2046 2222 2098
rect 3826 2046 3838 2098
rect 3890 2046 3902 2098
rect 9538 2046 9550 2098
rect 9602 2046 9614 2098
rect 10434 2046 10446 2098
rect 10498 2046 10510 2098
rect 12786 2046 12798 2098
rect 12850 2046 12862 2098
rect 14690 2046 14702 2098
rect 14754 2046 14766 2098
rect 16034 2046 16046 2098
rect 16098 2046 16110 2098
rect 16818 2046 16830 2098
rect 16882 2046 16894 2098
rect 23202 2046 23214 2098
rect 23266 2046 23278 2098
rect 25890 2046 25902 2098
rect 25954 2046 25966 2098
rect 26786 2046 26798 2098
rect 26850 2046 26862 2098
rect 27458 2046 27470 2098
rect 27522 2046 27534 2098
rect 28130 2046 28142 2098
rect 28194 2046 28206 2098
rect 7646 2034 7698 2046
rect 17166 2034 17218 2046
rect 14366 1986 14418 1998
rect 2706 1934 2718 1986
rect 2770 1934 2782 1986
rect 3378 1934 3390 1986
rect 3442 1934 3454 1986
rect 5618 1934 5630 1986
rect 5682 1934 5694 1986
rect 12338 1934 12350 1986
rect 12402 1934 12414 1986
rect 17602 1934 17614 1986
rect 17666 1934 17678 1986
rect 19842 1934 19854 1986
rect 19906 1934 19918 1986
rect 23650 1934 23662 1986
rect 23714 1934 23726 1986
rect 27010 1934 27022 1986
rect 27074 1934 27086 1986
rect 14366 1922 14418 1934
rect 10098 1822 10110 1874
rect 10162 1822 10174 1874
rect 26226 1822 26238 1874
rect 26290 1822 26302 1874
rect 672 1594 31024 1628
rect 672 1542 3806 1594
rect 3858 1542 3910 1594
rect 3962 1542 4014 1594
rect 4066 1542 23806 1594
rect 23858 1542 23910 1594
rect 23962 1542 24014 1594
rect 24066 1542 31024 1594
rect 672 1508 31024 1542
rect 3390 1426 3442 1438
rect 3390 1362 3442 1374
rect 7982 1426 8034 1438
rect 7982 1362 8034 1374
rect 11790 1426 11842 1438
rect 11790 1362 11842 1374
rect 14254 1426 14306 1438
rect 14254 1362 14306 1374
rect 19406 1426 19458 1438
rect 19406 1362 19458 1374
rect 20190 1426 20242 1438
rect 20190 1362 20242 1374
rect 23998 1426 24050 1438
rect 23998 1362 24050 1374
rect 1810 1262 1822 1314
rect 1874 1262 1886 1314
rect 6402 1262 6414 1314
rect 6466 1262 6478 1314
rect 17826 1262 17838 1314
rect 17890 1262 17902 1314
rect 25554 1262 25566 1314
rect 25618 1262 25630 1314
rect 3838 1202 3890 1214
rect 23326 1202 23378 1214
rect 28030 1202 28082 1214
rect 5618 1150 5630 1202
rect 5682 1150 5694 1202
rect 9314 1150 9326 1202
rect 9378 1150 9390 1202
rect 10210 1150 10222 1202
rect 10274 1150 10286 1202
rect 12674 1150 12686 1202
rect 12738 1150 12750 1202
rect 14802 1150 14814 1202
rect 14866 1150 14878 1202
rect 15474 1150 15486 1202
rect 15538 1150 15550 1202
rect 21746 1150 21758 1202
rect 21810 1150 21822 1202
rect 22530 1150 22542 1202
rect 22594 1150 22606 1202
rect 26338 1150 26350 1202
rect 26402 1150 26414 1202
rect 28578 1150 28590 1202
rect 28642 1150 28654 1202
rect 29250 1150 29262 1202
rect 29314 1150 29326 1202
rect 3838 1138 3890 1150
rect 23326 1138 23378 1150
rect 28030 1138 28082 1150
rect 4846 1090 4898 1102
rect 2258 1038 2270 1090
rect 2322 1038 2334 1090
rect 4162 1038 4174 1090
rect 4226 1038 4238 1090
rect 6850 1038 6862 1090
rect 6914 1038 6926 1090
rect 10658 1038 10670 1090
rect 10722 1038 10734 1090
rect 18162 1038 18174 1090
rect 18226 1038 18238 1090
rect 21410 1038 21422 1090
rect 21474 1038 21486 1090
rect 25218 1038 25230 1090
rect 25282 1038 25294 1090
rect 26114 1038 26126 1090
rect 26178 1038 26190 1090
rect 27682 1038 27694 1090
rect 27746 1038 27758 1090
rect 28354 1038 28366 1090
rect 28418 1038 28430 1090
rect 4846 1026 4898 1038
rect 16942 978 16994 990
rect 27134 978 27186 990
rect 5170 926 5182 978
rect 5234 926 5246 978
rect 5842 926 5854 978
rect 5906 926 5918 978
rect 9538 926 9550 978
rect 9602 926 9614 978
rect 13122 926 13134 978
rect 13186 926 13198 978
rect 15026 926 15038 978
rect 15090 926 15102 978
rect 15698 926 15710 978
rect 15762 926 15774 978
rect 16594 926 16606 978
rect 16658 926 16670 978
rect 22306 926 22318 978
rect 22370 926 22382 978
rect 22978 926 22990 978
rect 23042 926 23054 978
rect 26786 926 26798 978
rect 26850 926 26862 978
rect 29026 926 29038 978
rect 29090 926 29102 978
rect 16942 914 16994 926
rect 27134 914 27186 926
rect 672 810 31024 844
rect 672 758 4466 810
rect 4518 758 4570 810
rect 4622 758 4674 810
rect 4726 758 24466 810
rect 24518 758 24570 810
rect 24622 758 24674 810
rect 24726 758 31024 810
rect 672 724 31024 758
<< via1 >>
rect 4466 113654 4518 113706
rect 4570 113654 4622 113706
rect 4674 113654 4726 113706
rect 24466 113654 24518 113706
rect 24570 113654 24622 113706
rect 24674 113654 24726 113706
rect 1486 113486 1538 113538
rect 4846 113486 4898 113538
rect 5182 113486 5234 113538
rect 14702 113486 14754 113538
rect 15374 113486 15426 113538
rect 18510 113486 18562 113538
rect 19182 113486 19234 113538
rect 22318 113486 22370 113538
rect 22990 113486 23042 113538
rect 24558 113486 24610 113538
rect 25454 113486 25506 113538
rect 26126 113486 26178 113538
rect 26798 113486 26850 113538
rect 27694 113486 27746 113538
rect 28366 113486 28418 113538
rect 29038 113486 29090 113538
rect 29822 113486 29874 113538
rect 2942 113374 2994 113426
rect 5518 113374 5570 113426
rect 5854 113374 5906 113426
rect 6862 113374 6914 113426
rect 9662 113374 9714 113426
rect 11566 113374 11618 113426
rect 12574 113374 12626 113426
rect 13694 113374 13746 113426
rect 17614 113374 17666 113426
rect 21310 113374 21362 113426
rect 23886 113374 23938 113426
rect 1262 113262 1314 113314
rect 6302 113262 6354 113314
rect 11790 113262 11842 113314
rect 15038 113262 15090 113314
rect 15598 113262 15650 113314
rect 18846 113262 18898 113314
rect 19518 113262 19570 113314
rect 22542 113262 22594 113314
rect 23214 113262 23266 113314
rect 24222 113262 24274 113314
rect 24782 113262 24834 113314
rect 25790 113262 25842 113314
rect 26350 113262 26402 113314
rect 27022 113262 27074 113314
rect 27918 113262 27970 113314
rect 28590 113262 28642 113314
rect 29262 113262 29314 113314
rect 30046 113262 30098 113314
rect 2606 113150 2658 113202
rect 9214 113150 9266 113202
rect 11230 113150 11282 113202
rect 14142 113150 14194 113202
rect 17950 113150 18002 113202
rect 21758 113150 21810 113202
rect 25230 113150 25282 113202
rect 4174 113038 4226 113090
rect 7982 113038 8034 113090
rect 10782 113038 10834 113090
rect 16382 113038 16434 113090
rect 20190 113038 20242 113090
rect 3806 112870 3858 112922
rect 3910 112870 3962 112922
rect 4014 112870 4066 112922
rect 23806 112870 23858 112922
rect 23910 112870 23962 112922
rect 24014 112870 24066 112922
rect 16718 112590 16770 112642
rect 18958 112590 19010 112642
rect 2718 112478 2770 112530
rect 8430 112478 8482 112530
rect 10782 112478 10834 112530
rect 14478 112478 14530 112530
rect 15150 112478 15202 112530
rect 23550 112478 23602 112530
rect 24222 112478 24274 112530
rect 25790 112478 25842 112530
rect 1486 112366 1538 112418
rect 6078 112366 6130 112418
rect 10222 112366 10274 112418
rect 11566 112366 11618 112418
rect 12238 112366 12290 112418
rect 16382 112366 16434 112418
rect 18622 112366 18674 112418
rect 19518 112366 19570 112418
rect 20638 112366 20690 112418
rect 21310 112366 21362 112418
rect 21982 112366 22034 112418
rect 23326 112366 23378 112418
rect 23998 112366 24050 112418
rect 24670 112366 24722 112418
rect 25566 112366 25618 112418
rect 26462 112366 26514 112418
rect 27134 112366 27186 112418
rect 27470 112366 27522 112418
rect 28478 112366 28530 112418
rect 29150 112366 29202 112418
rect 29822 112366 29874 112418
rect 1150 112254 1202 112306
rect 1822 112254 1874 112306
rect 2158 112254 2210 112306
rect 3166 112254 3218 112306
rect 4286 112254 4338 112306
rect 5070 112254 5122 112306
rect 5406 112254 5458 112306
rect 5742 112254 5794 112306
rect 6862 112254 6914 112306
rect 7982 112254 8034 112306
rect 9102 112254 9154 112306
rect 11230 112254 11282 112306
rect 11902 112254 11954 112306
rect 12910 112254 12962 112306
rect 14030 112254 14082 112306
rect 17390 112254 17442 112306
rect 19854 112254 19906 112306
rect 20974 112254 21026 112306
rect 21646 112254 21698 112306
rect 22318 112254 22370 112306
rect 22654 112254 22706 112306
rect 22990 112254 23042 112306
rect 25006 112254 25058 112306
rect 25342 112254 25394 112306
rect 26238 112254 26290 112306
rect 26798 112254 26850 112306
rect 28814 112254 28866 112306
rect 29486 112254 29538 112306
rect 30158 112254 30210 112306
rect 4466 112086 4518 112138
rect 4570 112086 4622 112138
rect 4674 112086 4726 112138
rect 24466 112086 24518 112138
rect 24570 112086 24622 112138
rect 24674 112086 24726 112138
rect 8094 111918 8146 111970
rect 9214 111918 9266 111970
rect 10894 111918 10946 111970
rect 21198 111918 21250 111970
rect 21870 111918 21922 111970
rect 22878 111918 22930 111970
rect 24894 111918 24946 111970
rect 26574 111918 26626 111970
rect 27246 111918 27298 111970
rect 27582 111918 27634 111970
rect 28254 111918 28306 111970
rect 28926 111918 28978 111970
rect 29934 111918 29986 111970
rect 1598 111806 1650 111858
rect 3838 111806 3890 111858
rect 5070 111806 5122 111858
rect 6190 111806 6242 111858
rect 12462 111806 12514 111858
rect 14926 111806 14978 111858
rect 17950 111806 18002 111858
rect 20190 111806 20242 111858
rect 21534 111806 21586 111858
rect 22206 111806 22258 111858
rect 23662 111806 23714 111858
rect 25566 111806 25618 111858
rect 29262 111806 29314 111858
rect 30606 111806 30658 111858
rect 5630 111694 5682 111746
rect 7758 111694 7810 111746
rect 8990 111694 9042 111746
rect 10558 111694 10610 111746
rect 12014 111694 12066 111746
rect 14366 111694 14418 111746
rect 20750 111694 20802 111746
rect 22542 111694 22594 111746
rect 23326 111694 23378 111746
rect 24558 111694 24610 111746
rect 25230 111694 25282 111746
rect 26014 111694 26066 111746
rect 26238 111694 26290 111746
rect 27022 111694 27074 111746
rect 27806 111694 27858 111746
rect 28478 111694 28530 111746
rect 29598 111694 29650 111746
rect 30270 111694 30322 111746
rect 1262 111582 1314 111634
rect 3502 111582 3554 111634
rect 9662 111582 9714 111634
rect 9998 111582 10050 111634
rect 11230 111582 11282 111634
rect 11566 111582 11618 111634
rect 18398 111582 18450 111634
rect 2830 111470 2882 111522
rect 7310 111470 7362 111522
rect 13582 111470 13634 111522
rect 16046 111470 16098 111522
rect 16830 111470 16882 111522
rect 19070 111470 19122 111522
rect 3806 111302 3858 111354
rect 3910 111302 3962 111354
rect 4014 111302 4066 111354
rect 23806 111302 23858 111354
rect 23910 111302 23962 111354
rect 24014 111302 24066 111354
rect 9662 111022 9714 111074
rect 11566 111022 11618 111074
rect 19518 111022 19570 111074
rect 1262 110910 1314 110962
rect 5518 110910 5570 110962
rect 6414 110910 6466 110962
rect 6862 110910 6914 110962
rect 7534 110910 7586 110962
rect 8094 110910 8146 110962
rect 9102 110910 9154 110962
rect 9998 110910 10050 110962
rect 10558 110910 10610 110962
rect 10894 110910 10946 110962
rect 12014 110910 12066 110962
rect 13582 110910 13634 110962
rect 15150 110910 15202 110962
rect 15822 110910 15874 110962
rect 17950 110910 18002 110962
rect 20862 110910 20914 110962
rect 21310 110910 21362 110962
rect 21982 110910 22034 110962
rect 22766 110910 22818 110962
rect 23326 110910 23378 110962
rect 23998 110910 24050 110962
rect 24670 110910 24722 110962
rect 26126 110910 26178 110962
rect 30270 110910 30322 110962
rect 1598 110798 1650 110850
rect 3726 110798 3778 110850
rect 4398 110798 4450 110850
rect 6078 110798 6130 110850
rect 10222 110798 10274 110850
rect 19070 110798 19122 110850
rect 20638 110798 20690 110850
rect 22318 110798 22370 110850
rect 22990 110798 23042 110850
rect 23662 110798 23714 110850
rect 24334 110798 24386 110850
rect 25006 110798 25058 110850
rect 25678 110798 25730 110850
rect 26798 110798 26850 110850
rect 27470 110798 27522 110850
rect 29822 110798 29874 110850
rect 2830 110686 2882 110738
rect 3390 110686 3442 110738
rect 4062 110686 4114 110738
rect 5742 110686 5794 110738
rect 7086 110686 7138 110738
rect 11230 110686 11282 110738
rect 12238 110686 12290 110738
rect 14030 110686 14082 110738
rect 16270 110686 16322 110738
rect 17390 110686 17442 110738
rect 21646 110686 21698 110738
rect 25342 110686 25394 110738
rect 26462 110686 26514 110738
rect 27134 110686 27186 110738
rect 29486 110686 29538 110738
rect 30606 110686 30658 110738
rect 4466 110518 4518 110570
rect 4570 110518 4622 110570
rect 4674 110518 4726 110570
rect 24466 110518 24518 110570
rect 24570 110518 24622 110570
rect 24674 110518 24726 110570
rect 1710 110350 1762 110402
rect 9998 110350 10050 110402
rect 13918 110350 13970 110402
rect 18958 110350 19010 110402
rect 19966 110350 20018 110402
rect 20302 110350 20354 110402
rect 21646 110350 21698 110402
rect 21982 110350 22034 110402
rect 22654 110350 22706 110402
rect 23886 110350 23938 110402
rect 24894 110350 24946 110402
rect 25566 110350 25618 110402
rect 27022 110350 27074 110402
rect 27358 110350 27410 110402
rect 2718 110238 2770 110290
rect 4622 110238 4674 110290
rect 4958 110238 5010 110290
rect 6638 110238 6690 110290
rect 9214 110238 9266 110290
rect 11342 110238 11394 110290
rect 17950 110238 18002 110290
rect 19630 110238 19682 110290
rect 20638 110238 20690 110290
rect 20974 110238 21026 110290
rect 25230 110238 25282 110290
rect 26574 110238 26626 110290
rect 27694 110238 27746 110290
rect 30606 110238 30658 110290
rect 1374 110126 1426 110178
rect 8878 110126 8930 110178
rect 10334 110126 10386 110178
rect 10894 110126 10946 110178
rect 13358 110126 13410 110178
rect 13694 110126 13746 110178
rect 14590 110126 14642 110178
rect 15038 110126 15090 110178
rect 15934 110126 15986 110178
rect 19294 110126 19346 110178
rect 21198 110126 21250 110178
rect 22318 110126 22370 110178
rect 23550 110126 23602 110178
rect 24670 110126 24722 110178
rect 26350 110126 26402 110178
rect 30270 110126 30322 110178
rect 2270 110014 2322 110066
rect 5630 110014 5682 110066
rect 6302 110014 6354 110066
rect 9550 110014 9602 110066
rect 12910 110014 12962 110066
rect 18398 110014 18450 110066
rect 25902 110014 25954 110066
rect 26798 110014 26850 110066
rect 3838 109902 3890 109954
rect 5294 109902 5346 109954
rect 7870 109902 7922 109954
rect 12462 109902 12514 109954
rect 16830 109902 16882 109954
rect 3806 109734 3858 109786
rect 3910 109734 3962 109786
rect 4014 109734 4066 109786
rect 23806 109734 23858 109786
rect 23910 109734 23962 109786
rect 24014 109734 24066 109786
rect 1262 109454 1314 109506
rect 6078 109454 6130 109506
rect 13470 109454 13522 109506
rect 4174 109342 4226 109394
rect 6526 109342 6578 109394
rect 6862 109342 6914 109394
rect 7646 109342 7698 109394
rect 8094 109342 8146 109394
rect 9102 109342 9154 109394
rect 9886 109342 9938 109394
rect 11118 109342 11170 109394
rect 15934 109342 15986 109394
rect 16382 109342 16434 109394
rect 17166 109342 17218 109394
rect 17502 109342 17554 109394
rect 18622 109342 18674 109394
rect 19070 109342 19122 109394
rect 19854 109342 19906 109394
rect 22990 109342 23042 109394
rect 29486 109342 29538 109394
rect 1598 109230 1650 109282
rect 3390 109230 3442 109282
rect 3726 109230 3778 109282
rect 4398 109230 4450 109282
rect 5406 109230 5458 109282
rect 5742 109230 5794 109282
rect 7086 109230 7138 109282
rect 11454 109230 11506 109282
rect 11790 109230 11842 109282
rect 12126 109230 12178 109282
rect 13918 109230 13970 109282
rect 15038 109230 15090 109282
rect 15486 109230 15538 109282
rect 19406 109230 19458 109282
rect 23214 109230 23266 109282
rect 26798 109230 26850 109282
rect 29822 109230 29874 109282
rect 2830 109118 2882 109170
rect 9662 109118 9714 109170
rect 10782 109118 10834 109170
rect 16494 109118 16546 109170
rect 20078 109118 20130 109170
rect 23550 109118 23602 109170
rect 25230 109118 25282 109170
rect 26126 109118 26178 109170
rect 27022 109118 27074 109170
rect 4466 108950 4518 109002
rect 4570 108950 4622 109002
rect 4674 108950 4726 109002
rect 24466 108950 24518 109002
rect 24570 108950 24622 109002
rect 24674 108950 24726 109002
rect 3390 108782 3442 108834
rect 9214 108782 9266 108834
rect 9550 108782 9602 108834
rect 10222 108782 10274 108834
rect 10558 108782 10610 108834
rect 14814 108782 14866 108834
rect 5742 108670 5794 108722
rect 6190 108670 6242 108722
rect 11902 108670 11954 108722
rect 16158 108670 16210 108722
rect 17950 108670 18002 108722
rect 23438 108670 23490 108722
rect 29822 108670 29874 108722
rect 30270 108670 30322 108722
rect 30606 108670 30658 108722
rect 1262 108558 1314 108610
rect 2270 108558 2322 108610
rect 2942 108558 2994 108610
rect 3502 108558 3554 108610
rect 3950 108558 4002 108610
rect 5070 108558 5122 108610
rect 5630 108558 5682 108610
rect 6750 108558 6802 108610
rect 7870 108558 7922 108610
rect 8878 108558 8930 108610
rect 9886 108558 9938 108610
rect 11230 108558 11282 108610
rect 11678 108558 11730 108610
rect 12462 108558 12514 108610
rect 12910 108558 12962 108610
rect 13918 108558 13970 108610
rect 15038 108558 15090 108610
rect 15822 108558 15874 108610
rect 18510 108558 18562 108610
rect 29598 108558 29650 108610
rect 4398 108446 4450 108498
rect 4734 108446 4786 108498
rect 8318 108446 8370 108498
rect 10894 108446 10946 108498
rect 15374 108446 15426 108498
rect 25118 108446 25170 108498
rect 26126 108446 26178 108498
rect 16830 108334 16882 108386
rect 3806 108166 3858 108218
rect 3910 108166 3962 108218
rect 4014 108166 4066 108218
rect 23806 108166 23858 108218
rect 23910 108166 23962 108218
rect 24014 108166 24066 108218
rect 6302 107886 6354 107938
rect 25118 107886 25170 107938
rect 1262 107774 1314 107826
rect 2382 107774 2434 107826
rect 2942 107774 2994 107826
rect 3614 107774 3666 107826
rect 4062 107774 4114 107826
rect 5182 107774 5234 107826
rect 9326 107774 9378 107826
rect 9774 107774 9826 107826
rect 11006 107774 11058 107826
rect 12014 107774 12066 107826
rect 13470 107774 13522 107826
rect 14254 107774 14306 107826
rect 15150 107774 15202 107826
rect 15598 107774 15650 107826
rect 16830 107774 16882 107826
rect 17726 107774 17778 107826
rect 30382 107774 30434 107826
rect 3390 107662 3442 107714
rect 4398 107662 4450 107714
rect 5406 107662 5458 107714
rect 7870 107662 7922 107714
rect 8654 107662 8706 107714
rect 8990 107662 9042 107714
rect 10446 107662 10498 107714
rect 13694 107662 13746 107714
rect 14030 107662 14082 107714
rect 14702 107662 14754 107714
rect 15710 107662 15762 107714
rect 16158 107662 16210 107714
rect 6750 107550 6802 107602
rect 8318 107550 8370 107602
rect 9998 107550 10050 107602
rect 30606 107550 30658 107602
rect 4466 107382 4518 107434
rect 4570 107382 4622 107434
rect 4674 107382 4726 107434
rect 24466 107382 24518 107434
rect 24570 107382 24622 107434
rect 24674 107382 24726 107434
rect 1150 107214 1202 107266
rect 7310 107214 7362 107266
rect 10110 107214 10162 107266
rect 12686 107214 12738 107266
rect 14030 107214 14082 107266
rect 25118 107214 25170 107266
rect 4062 107102 4114 107154
rect 5406 107102 5458 107154
rect 17950 107102 18002 107154
rect 30606 107102 30658 107154
rect 1486 106990 1538 107042
rect 1934 106990 1986 107042
rect 2830 106990 2882 107042
rect 3390 106990 3442 107042
rect 4174 106990 4226 107042
rect 4734 106990 4786 107042
rect 5742 106990 5794 107042
rect 9886 106990 9938 107042
rect 13806 106990 13858 107042
rect 16830 106990 16882 107042
rect 30270 106990 30322 107042
rect 5070 106878 5122 106930
rect 7758 106878 7810 106930
rect 8318 106878 8370 106930
rect 8878 106878 8930 106930
rect 9550 106878 9602 106930
rect 10782 106878 10834 106930
rect 13134 106878 13186 106930
rect 14590 106878 14642 106930
rect 18398 106878 18450 106930
rect 6190 106766 6242 106818
rect 11566 106766 11618 106818
rect 3806 106598 3858 106650
rect 3910 106598 3962 106650
rect 4014 106598 4066 106650
rect 23806 106598 23858 106650
rect 23910 106598 23962 106650
rect 24014 106598 24066 106650
rect 5406 106318 5458 106370
rect 15150 106318 15202 106370
rect 1262 106206 1314 106258
rect 2158 106206 2210 106258
rect 2942 106206 2994 106258
rect 3614 106206 3666 106258
rect 4062 106206 4114 106258
rect 7646 106206 7698 106258
rect 13022 106206 13074 106258
rect 16718 106206 16770 106258
rect 4398 106094 4450 106146
rect 9998 106094 10050 106146
rect 13358 106094 13410 106146
rect 29822 106094 29874 106146
rect 3390 105982 3442 106034
rect 5854 105982 5906 106034
rect 6974 105982 7026 106034
rect 8094 105982 8146 106034
rect 9214 105982 9266 106034
rect 9662 105982 9714 106034
rect 10334 105982 10386 106034
rect 10670 105982 10722 106034
rect 11118 105982 11170 106034
rect 14590 105982 14642 106034
rect 16270 105982 16322 106034
rect 29486 105982 29538 106034
rect 4466 105814 4518 105866
rect 4570 105814 4622 105866
rect 4674 105814 4726 105866
rect 24466 105814 24518 105866
rect 24570 105814 24622 105866
rect 24674 105814 24726 105866
rect 9214 105646 9266 105698
rect 11118 105646 11170 105698
rect 16046 105646 16098 105698
rect 22094 105646 22146 105698
rect 1598 105534 1650 105586
rect 2606 105534 2658 105586
rect 4734 105534 4786 105586
rect 6974 105534 7026 105586
rect 13358 105534 13410 105586
rect 14926 105534 14978 105586
rect 19070 105534 19122 105586
rect 19406 105534 19458 105586
rect 30270 105534 30322 105586
rect 30606 105534 30658 105586
rect 1262 105422 1314 105474
rect 8990 105422 9042 105474
rect 11342 105422 11394 105474
rect 14366 105422 14418 105474
rect 21870 105422 21922 105474
rect 2158 105310 2210 105362
rect 4398 105310 4450 105362
rect 6638 105310 6690 105362
rect 9662 105310 9714 105362
rect 13694 105310 13746 105362
rect 3726 105198 3778 105250
rect 5966 105198 6018 105250
rect 8206 105198 8258 105250
rect 12126 105198 12178 105250
rect 3806 105030 3858 105082
rect 3910 105030 3962 105082
rect 4014 105030 4066 105082
rect 23806 105030 23858 105082
rect 23910 105030 23962 105082
rect 24014 105030 24066 105082
rect 11678 104862 11730 104914
rect 1262 104750 1314 104802
rect 6078 104750 6130 104802
rect 12798 104750 12850 104802
rect 16606 104750 16658 104802
rect 3502 104638 3554 104690
rect 4286 104638 4338 104690
rect 5070 104638 5122 104690
rect 6414 104638 6466 104690
rect 6974 104638 7026 104690
rect 7534 104638 7586 104690
rect 8094 104638 8146 104690
rect 9214 104638 9266 104690
rect 11566 104638 11618 104690
rect 13134 104638 13186 104690
rect 13582 104638 13634 104690
rect 14478 104638 14530 104690
rect 15038 104638 15090 104690
rect 15822 104638 15874 104690
rect 1710 104526 1762 104578
rect 3726 104526 3778 104578
rect 4062 104526 4114 104578
rect 5294 104526 5346 104578
rect 7086 104526 7138 104578
rect 12014 104526 12066 104578
rect 12238 104526 12290 104578
rect 16942 104526 16994 104578
rect 2830 104414 2882 104466
rect 9662 104414 9714 104466
rect 11118 104414 11170 104466
rect 11454 104414 11506 104466
rect 13806 104414 13858 104466
rect 18174 104414 18226 104466
rect 30270 104414 30322 104466
rect 30606 104414 30658 104466
rect 4466 104246 4518 104298
rect 4570 104246 4622 104298
rect 4674 104246 4726 104298
rect 24466 104246 24518 104298
rect 24570 104246 24622 104298
rect 24674 104246 24726 104298
rect 12350 104078 12402 104130
rect 14254 104078 14306 104130
rect 20526 104078 20578 104130
rect 20862 104078 20914 104130
rect 1598 103966 1650 104018
rect 2606 103966 2658 104018
rect 4734 103966 4786 104018
rect 7086 103966 7138 104018
rect 11454 103966 11506 104018
rect 12574 103966 12626 104018
rect 12686 103966 12738 104018
rect 15262 103966 15314 104018
rect 18958 103966 19010 104018
rect 1374 103854 1426 103906
rect 15598 103854 15650 103906
rect 15822 103854 15874 103906
rect 16830 103854 16882 103906
rect 17726 103854 17778 103906
rect 18510 103854 18562 103906
rect 19070 103854 19122 103906
rect 19518 103854 19570 103906
rect 2158 103742 2210 103794
rect 4398 103742 4450 103794
rect 6638 103742 6690 103794
rect 11902 103742 11954 103794
rect 14702 103742 14754 103794
rect 19966 103742 20018 103794
rect 3726 103630 3778 103682
rect 5966 103630 6018 103682
rect 8206 103630 8258 103682
rect 10334 103630 10386 103682
rect 13134 103630 13186 103682
rect 15374 103630 15426 103682
rect 3806 103462 3858 103514
rect 3910 103462 3962 103514
rect 4014 103462 4066 103514
rect 23806 103462 23858 103514
rect 23910 103462 23962 103514
rect 24014 103462 24066 103514
rect 11678 103294 11730 103346
rect 12238 103294 12290 103346
rect 12798 103294 12850 103346
rect 18734 103294 18786 103346
rect 1262 103182 1314 103234
rect 6302 103182 6354 103234
rect 10110 103182 10162 103234
rect 12126 103182 12178 103234
rect 12910 103182 12962 103234
rect 3390 103070 3442 103122
rect 5070 103070 5122 103122
rect 6750 103070 6802 103122
rect 7198 103070 7250 103122
rect 7982 103070 8034 103122
rect 8542 103070 8594 103122
rect 9326 103070 9378 103122
rect 13134 103070 13186 103122
rect 13694 103070 13746 103122
rect 17054 103070 17106 103122
rect 19182 103070 19234 103122
rect 1598 102958 1650 103010
rect 3726 102958 3778 103010
rect 4398 102958 4450 103010
rect 5966 102958 6018 103010
rect 7310 102958 7362 103010
rect 17614 102958 17666 103010
rect 2830 102846 2882 102898
rect 4062 102846 4114 102898
rect 5294 102846 5346 102898
rect 5630 102846 5682 102898
rect 10558 102846 10610 102898
rect 14142 102846 14194 102898
rect 15262 102846 15314 102898
rect 16606 102846 16658 102898
rect 19518 102846 19570 102898
rect 30270 102846 30322 102898
rect 30606 102846 30658 102898
rect 4466 102678 4518 102730
rect 4570 102678 4622 102730
rect 4674 102678 4726 102730
rect 24466 102678 24518 102730
rect 24570 102678 24622 102730
rect 24674 102678 24726 102730
rect 1710 102398 1762 102450
rect 6078 102398 6130 102450
rect 7086 102398 7138 102450
rect 7982 102398 8034 102450
rect 8318 102398 8370 102450
rect 9102 102398 9154 102450
rect 10110 102398 10162 102450
rect 11342 102398 11394 102450
rect 12910 102398 12962 102450
rect 13918 102398 13970 102450
rect 17614 102398 17666 102450
rect 30270 102398 30322 102450
rect 30606 102398 30658 102450
rect 1262 102286 1314 102338
rect 3950 102286 4002 102338
rect 4846 102286 4898 102338
rect 5406 102286 5458 102338
rect 6190 102286 6242 102338
rect 6638 102286 6690 102338
rect 10222 102286 10274 102338
rect 13246 102286 13298 102338
rect 13694 102286 13746 102338
rect 14590 102286 14642 102338
rect 15150 102286 15202 102338
rect 16046 102286 16098 102338
rect 17278 102286 17330 102338
rect 10894 102174 10946 102226
rect 2942 102062 2994 102114
rect 9438 102062 9490 102114
rect 12462 102062 12514 102114
rect 3806 101894 3858 101946
rect 3910 101894 3962 101946
rect 4014 101894 4066 101946
rect 23806 101894 23858 101946
rect 23910 101894 23962 101946
rect 24014 101894 24066 101946
rect 13246 101614 13298 101666
rect 1374 101502 1426 101554
rect 2158 101502 2210 101554
rect 2942 101502 2994 101554
rect 3502 101502 3554 101554
rect 4062 101502 4114 101554
rect 5182 101502 5234 101554
rect 5854 101502 5906 101554
rect 8990 101502 9042 101554
rect 9550 101502 9602 101554
rect 10670 101502 10722 101554
rect 11678 101502 11730 101554
rect 13582 101502 13634 101554
rect 14030 101502 14082 101554
rect 14926 101502 14978 101554
rect 15262 101502 15314 101554
rect 16270 101502 16322 101554
rect 3390 101390 3442 101442
rect 4398 101390 4450 101442
rect 5406 101390 5458 101442
rect 8654 101390 8706 101442
rect 9662 101390 9714 101442
rect 10110 101390 10162 101442
rect 6414 101278 6466 101330
rect 7534 101278 7586 101330
rect 14254 101278 14306 101330
rect 4466 101110 4518 101162
rect 4570 101110 4622 101162
rect 4674 101110 4726 101162
rect 24466 101110 24518 101162
rect 24570 101110 24622 101162
rect 24674 101110 24726 101162
rect 2382 100942 2434 100994
rect 5966 100830 6018 100882
rect 6974 100830 7026 100882
rect 7310 100830 7362 100882
rect 10558 100830 10610 100882
rect 14254 100830 14306 100882
rect 17614 100830 17666 100882
rect 29822 100830 29874 100882
rect 30606 100830 30658 100882
rect 2830 100718 2882 100770
rect 3838 100718 3890 100770
rect 4734 100718 4786 100770
rect 5294 100718 5346 100770
rect 6190 100718 6242 100770
rect 6638 100718 6690 100770
rect 7646 100718 7698 100770
rect 9886 100718 9938 100770
rect 10334 100718 10386 100770
rect 11230 100718 11282 100770
rect 11566 100718 11618 100770
rect 12574 100718 12626 100770
rect 13918 100718 13970 100770
rect 15486 100718 15538 100770
rect 17278 100718 17330 100770
rect 29486 100718 29538 100770
rect 30270 100718 30322 100770
rect 9550 100606 9602 100658
rect 1262 100494 1314 100546
rect 3806 100326 3858 100378
rect 3910 100326 3962 100378
rect 4014 100326 4066 100378
rect 23806 100326 23858 100378
rect 23910 100326 23962 100378
rect 24014 100326 24066 100378
rect 12910 100158 12962 100210
rect 5182 100046 5234 100098
rect 8990 100046 9042 100098
rect 14478 100046 14530 100098
rect 1262 99934 1314 99986
rect 2158 99934 2210 99986
rect 2942 99934 2994 99986
rect 3614 99934 3666 99986
rect 4062 99934 4114 99986
rect 9326 99934 9378 99986
rect 9886 99934 9938 99986
rect 10670 99934 10722 99986
rect 11230 99934 11282 99986
rect 12126 99934 12178 99986
rect 17166 99934 17218 99986
rect 4398 99822 4450 99874
rect 5630 99822 5682 99874
rect 9998 99822 10050 99874
rect 17726 99822 17778 99874
rect 22542 99822 22594 99874
rect 3390 99710 3442 99762
rect 6750 99710 6802 99762
rect 14030 99710 14082 99762
rect 18846 99710 18898 99762
rect 22206 99710 22258 99762
rect 30270 99710 30322 99762
rect 30606 99710 30658 99762
rect 4466 99542 4518 99594
rect 4570 99542 4622 99594
rect 4674 99542 4726 99594
rect 24466 99542 24518 99594
rect 24570 99542 24622 99594
rect 24674 99542 24726 99594
rect 14814 99374 14866 99426
rect 18958 99374 19010 99426
rect 1934 99262 1986 99314
rect 4398 99262 4450 99314
rect 6638 99262 6690 99314
rect 10894 99262 10946 99314
rect 17390 99262 17442 99314
rect 19294 99262 19346 99314
rect 30270 99262 30322 99314
rect 30606 99262 30658 99314
rect 3166 99150 3218 99202
rect 3838 99150 3890 99202
rect 8318 99150 8370 99202
rect 10222 99156 10274 99208
rect 10782 99150 10834 99202
rect 11454 99150 11506 99202
rect 11902 99150 11954 99202
rect 12910 99150 12962 99202
rect 16942 99150 16994 99202
rect 1598 99038 1650 99090
rect 6190 99038 6242 99090
rect 7758 99038 7810 99090
rect 9886 99038 9938 99090
rect 14366 99038 14418 99090
rect 5518 98926 5570 98978
rect 8206 98926 8258 98978
rect 15934 98926 15986 98978
rect 18510 98926 18562 98978
rect 3806 98758 3858 98810
rect 3910 98758 3962 98810
rect 4014 98758 4066 98810
rect 23806 98758 23858 98810
rect 23910 98758 23962 98810
rect 24014 98758 24066 98810
rect 11342 98590 11394 98642
rect 1822 98478 1874 98530
rect 5294 98478 5346 98530
rect 9774 98478 9826 98530
rect 18846 98478 18898 98530
rect 19966 98478 20018 98530
rect 7422 98366 7474 98418
rect 13022 98366 13074 98418
rect 15598 98366 15650 98418
rect 16046 98366 16098 98418
rect 16830 98366 16882 98418
rect 17166 98366 17218 98418
rect 18174 98366 18226 98418
rect 18958 98366 19010 98418
rect 19182 98366 19234 98418
rect 19294 98366 19346 98418
rect 4174 98254 4226 98306
rect 4286 98254 4338 98306
rect 5742 98254 5794 98306
rect 7982 98254 8034 98306
rect 10110 98254 10162 98306
rect 13582 98254 13634 98306
rect 15150 98254 15202 98306
rect 16158 98254 16210 98306
rect 18734 98254 18786 98306
rect 2270 98142 2322 98194
rect 3390 98142 3442 98194
rect 4510 98142 4562 98194
rect 6862 98142 6914 98194
rect 9102 98142 9154 98194
rect 14702 98142 14754 98194
rect 19854 98142 19906 98194
rect 4466 97974 4518 98026
rect 4570 97974 4622 98026
rect 4674 97974 4726 98026
rect 24466 97974 24518 98026
rect 24570 97974 24622 98026
rect 24674 97974 24726 98026
rect 1710 97806 1762 97858
rect 8094 97806 8146 97858
rect 11790 97806 11842 97858
rect 14926 97806 14978 97858
rect 16830 97806 16882 97858
rect 19070 97806 19122 97858
rect 21982 97806 22034 97858
rect 4062 97694 4114 97746
rect 5070 97694 5122 97746
rect 10222 97694 10274 97746
rect 18062 97694 18114 97746
rect 29822 97694 29874 97746
rect 30270 97694 30322 97746
rect 30606 97694 30658 97746
rect 1150 97582 1202 97634
rect 4398 97582 4450 97634
rect 4846 97582 4898 97634
rect 5630 97582 5682 97634
rect 6190 97582 6242 97634
rect 7086 97582 7138 97634
rect 7758 97582 7810 97634
rect 7982 97582 8034 97634
rect 8206 97582 8258 97634
rect 10558 97582 10610 97634
rect 11342 97582 11394 97634
rect 18398 97582 18450 97634
rect 19182 97582 19234 97634
rect 21758 97582 21810 97634
rect 29486 97582 29538 97634
rect 8990 97470 9042 97522
rect 14478 97470 14530 97522
rect 2830 97358 2882 97410
rect 12910 97358 12962 97410
rect 16046 97358 16098 97410
rect 19070 97358 19122 97410
rect 19406 97358 19458 97410
rect 3806 97190 3858 97242
rect 3910 97190 3962 97242
rect 4014 97190 4066 97242
rect 23806 97190 23858 97242
rect 23910 97190 23962 97242
rect 24014 97190 24066 97242
rect 18286 97022 18338 97074
rect 18622 97022 18674 97074
rect 5518 96910 5570 96962
rect 7758 96910 7810 96962
rect 9998 96910 10050 96962
rect 14702 96910 14754 96962
rect 2718 96798 2770 96850
rect 11566 96798 11618 96850
rect 13022 96798 13074 96850
rect 13694 96798 13746 96850
rect 15038 96798 15090 96850
rect 15486 96798 15538 96850
rect 16158 96798 16210 96850
rect 16942 96798 16994 96850
rect 17726 96798 17778 96850
rect 18622 96798 18674 96850
rect 19518 96798 19570 96850
rect 22318 96798 22370 96850
rect 8206 96686 8258 96738
rect 12910 96686 12962 96738
rect 3166 96574 3218 96626
rect 4286 96574 4338 96626
rect 5966 96574 6018 96626
rect 7086 96574 7138 96626
rect 9326 96574 9378 96626
rect 10446 96574 10498 96626
rect 14030 96574 14082 96626
rect 15710 96574 15762 96626
rect 19854 96574 19906 96626
rect 20750 96574 20802 96626
rect 21870 96574 21922 96626
rect 30270 96574 30322 96626
rect 30606 96574 30658 96626
rect 4466 96406 4518 96458
rect 4570 96406 4622 96458
rect 4674 96406 4726 96458
rect 24466 96406 24518 96458
rect 24570 96406 24622 96458
rect 24674 96406 24726 96458
rect 8094 96238 8146 96290
rect 11454 96238 11506 96290
rect 16830 96238 16882 96290
rect 19966 96238 20018 96290
rect 22206 96238 22258 96290
rect 29486 96238 29538 96290
rect 29822 96238 29874 96290
rect 1710 96126 1762 96178
rect 4734 96126 4786 96178
rect 7310 96126 7362 96178
rect 17054 96126 17106 96178
rect 17166 96126 17218 96178
rect 18958 96126 19010 96178
rect 4174 96014 4226 96066
rect 4622 96014 4674 96066
rect 5406 96014 5458 96066
rect 5742 96014 5794 96066
rect 6750 96014 6802 96066
rect 7646 96014 7698 96066
rect 7758 96014 7810 96066
rect 7870 96014 7922 96066
rect 10894 96014 10946 96066
rect 11230 96014 11282 96066
rect 12126 96014 12178 96066
rect 12462 96014 12514 96066
rect 13470 96014 13522 96066
rect 18622 96014 18674 96066
rect 1374 95902 1426 95954
rect 3726 95902 3778 95954
rect 10446 95902 10498 95954
rect 19518 95902 19570 95954
rect 21758 95902 21810 95954
rect 2942 95790 2994 95842
rect 21086 95790 21138 95842
rect 23326 95790 23378 95842
rect 3806 95622 3858 95674
rect 3910 95622 3962 95674
rect 4014 95622 4066 95674
rect 23806 95622 23858 95674
rect 23910 95622 23962 95674
rect 24014 95622 24066 95674
rect 12910 95454 12962 95506
rect 7086 95342 7138 95394
rect 14478 95342 14530 95394
rect 1486 95230 1538 95282
rect 1934 95230 1986 95282
rect 2494 95230 2546 95282
rect 3054 95230 3106 95282
rect 4174 95230 4226 95282
rect 8542 95230 8594 95282
rect 8878 95230 8930 95282
rect 9550 95230 9602 95282
rect 10334 95230 10386 95282
rect 11118 95230 11170 95282
rect 18398 95230 18450 95282
rect 21086 95230 21138 95282
rect 21422 95230 21474 95282
rect 22206 95230 22258 95282
rect 22878 95230 22930 95282
rect 23774 95230 23826 95282
rect 1038 95118 1090 95170
rect 6638 95118 6690 95170
rect 8094 95118 8146 95170
rect 14142 95118 14194 95170
rect 20638 95118 20690 95170
rect 2046 95006 2098 95058
rect 5518 95006 5570 95058
rect 9102 95006 9154 95058
rect 18846 95006 18898 95058
rect 19966 95006 20018 95058
rect 21646 95006 21698 95058
rect 30270 95006 30322 95058
rect 30606 95006 30658 95058
rect 4466 94838 4518 94890
rect 4570 94838 4622 94890
rect 4674 94838 4726 94890
rect 24466 94838 24518 94890
rect 24570 94838 24622 94890
rect 24674 94838 24726 94890
rect 6638 94670 6690 94722
rect 12014 94670 12066 94722
rect 16830 94670 16882 94722
rect 18174 94670 18226 94722
rect 23662 94670 23714 94722
rect 1822 94558 1874 94610
rect 2830 94558 2882 94610
rect 9214 94558 9266 94610
rect 9662 94558 9714 94610
rect 14814 94558 14866 94610
rect 17166 94558 17218 94610
rect 20750 94558 20802 94610
rect 23326 94558 23378 94610
rect 30606 94558 30658 94610
rect 2270 94446 2322 94498
rect 2718 94446 2770 94498
rect 3390 94446 3442 94498
rect 4062 94446 4114 94498
rect 4846 94446 4898 94498
rect 7086 94446 7138 94498
rect 11454 94446 11506 94498
rect 11902 94446 11954 94498
rect 12686 94446 12738 94498
rect 13022 94446 13074 94498
rect 13246 94446 13298 94498
rect 14142 94446 14194 94498
rect 14702 94446 14754 94498
rect 20190 94446 20242 94498
rect 20526 94446 20578 94498
rect 21310 94446 21362 94498
rect 21870 94446 21922 94498
rect 22766 94446 22818 94498
rect 30382 94446 30434 94498
rect 11006 94334 11058 94386
rect 15822 94334 15874 94386
rect 17726 94334 17778 94386
rect 19742 94334 19794 94386
rect 5518 94222 5570 94274
rect 9886 94222 9938 94274
rect 10222 94222 10274 94274
rect 15486 94222 15538 94274
rect 19294 94222 19346 94274
rect 3806 94054 3858 94106
rect 3910 94054 3962 94106
rect 4014 94054 4066 94106
rect 23806 94054 23858 94106
rect 23910 94054 23962 94106
rect 24014 94054 24066 94106
rect 4398 93774 4450 93826
rect 8542 93774 8594 93826
rect 22766 93774 22818 93826
rect 1262 93662 1314 93714
rect 2158 93662 2210 93714
rect 2942 93662 2994 93714
rect 3502 93662 3554 93714
rect 3950 93662 4002 93714
rect 5742 93662 5794 93714
rect 8990 93662 9042 93714
rect 9326 93662 9378 93714
rect 10222 93662 10274 93714
rect 10782 93662 10834 93714
rect 11566 93662 11618 93714
rect 13582 93662 13634 93714
rect 15150 93662 15202 93714
rect 16046 93662 16098 93714
rect 16382 93662 16434 93714
rect 17054 93662 17106 93714
rect 17838 93662 17890 93714
rect 18622 93662 18674 93714
rect 26910 93662 26962 93714
rect 6078 93550 6130 93602
rect 9550 93550 9602 93602
rect 15598 93550 15650 93602
rect 3390 93438 3442 93490
rect 7310 93438 7362 93490
rect 14030 93438 14082 93490
rect 16606 93438 16658 93490
rect 19182 93438 19234 93490
rect 19518 93438 19570 93490
rect 4466 93270 4518 93322
rect 4570 93270 4622 93322
rect 4674 93270 4726 93322
rect 24466 93270 24518 93322
rect 24570 93270 24622 93322
rect 24674 93270 24726 93322
rect 7086 93102 7138 93154
rect 8206 93102 8258 93154
rect 9886 93102 9938 93154
rect 13806 93102 13858 93154
rect 17614 93102 17666 93154
rect 30270 93102 30322 93154
rect 1038 92990 1090 93042
rect 2046 92990 2098 93042
rect 2494 92990 2546 93042
rect 4958 92990 5010 93042
rect 5294 92990 5346 93042
rect 8878 92990 8930 93042
rect 12910 92990 12962 93042
rect 14814 92990 14866 93042
rect 17502 92990 17554 93042
rect 19742 92990 19794 93042
rect 20750 92990 20802 93042
rect 21198 92990 21250 93042
rect 24670 92990 24722 93042
rect 30606 92990 30658 93042
rect 1486 92878 1538 92930
rect 1934 92878 1986 92930
rect 3054 92878 3106 92930
rect 4174 92878 4226 92930
rect 5630 92878 5682 92930
rect 6638 92878 6690 92930
rect 9326 92878 9378 92930
rect 9662 92878 9714 92930
rect 10446 92878 10498 92930
rect 10894 92878 10946 92930
rect 11902 92878 11954 92930
rect 12686 92878 12738 92930
rect 14478 92878 14530 92930
rect 17054 92878 17106 92930
rect 20190 92878 20242 92930
rect 20526 92878 20578 92930
rect 21870 92878 21922 92930
rect 22766 92878 22818 92930
rect 24894 92878 24946 92930
rect 5966 92766 6018 92818
rect 13470 92654 13522 92706
rect 16046 92654 16098 92706
rect 18734 92654 18786 92706
rect 25454 92654 25506 92706
rect 25790 92654 25842 92706
rect 3806 92486 3858 92538
rect 3910 92486 3962 92538
rect 4014 92486 4066 92538
rect 23806 92486 23858 92538
rect 23910 92486 23962 92538
rect 24014 92486 24066 92538
rect 5070 92318 5122 92370
rect 5406 92206 5458 92258
rect 8206 92206 8258 92258
rect 15598 92206 15650 92258
rect 2718 92094 2770 92146
rect 6190 92094 6242 92146
rect 8542 92094 8594 92146
rect 8990 92094 9042 92146
rect 9662 92094 9714 92146
rect 10222 92094 10274 92146
rect 10446 92094 10498 92146
rect 11230 92094 11282 92146
rect 13582 92094 13634 92146
rect 15934 92094 15986 92146
rect 16382 92094 16434 92146
rect 17054 92094 17106 92146
rect 17838 92094 17890 92146
rect 18622 92094 18674 92146
rect 21086 92094 21138 92146
rect 21422 92094 21474 92146
rect 22094 92094 22146 92146
rect 22654 92094 22706 92146
rect 22878 92094 22930 92146
rect 23662 92094 23714 92146
rect 2270 91982 2322 92034
rect 6638 91982 6690 92034
rect 9214 91982 9266 92034
rect 14030 91982 14082 92034
rect 20638 91982 20690 92034
rect 21646 91982 21698 92034
rect 1150 91870 1202 91922
rect 5294 91870 5346 91922
rect 7758 91870 7810 91922
rect 15150 91870 15202 91922
rect 16606 91870 16658 91922
rect 19182 91870 19234 91922
rect 19518 91870 19570 91922
rect 30270 91870 30322 91922
rect 30606 91870 30658 91922
rect 4466 91702 4518 91754
rect 4570 91702 4622 91754
rect 4674 91702 4726 91754
rect 24466 91702 24518 91754
rect 24570 91702 24622 91754
rect 24674 91702 24726 91754
rect 7086 91534 7138 91586
rect 8206 91534 8258 91586
rect 13918 91534 13970 91586
rect 1710 91422 1762 91474
rect 4622 91422 4674 91474
rect 10894 91422 10946 91474
rect 12910 91422 12962 91474
rect 17726 91422 17778 91474
rect 21534 91422 21586 91474
rect 30606 91422 30658 91474
rect 6526 91310 6578 91362
rect 12126 91310 12178 91362
rect 13358 91310 13410 91362
rect 13806 91310 13858 91362
rect 14366 91310 14418 91362
rect 14926 91310 14978 91362
rect 15934 91310 15986 91362
rect 17054 91310 17106 91362
rect 17502 91310 17554 91362
rect 18174 91310 18226 91362
rect 18734 91310 18786 91362
rect 19742 91310 19794 91362
rect 21086 91310 21138 91362
rect 30270 91310 30322 91362
rect 1262 91198 1314 91250
rect 4958 91198 5010 91250
rect 10558 91198 10610 91250
rect 16718 91198 16770 91250
rect 2830 91086 2882 91138
rect 3390 91086 3442 91138
rect 22766 91086 22818 91138
rect 3806 90918 3858 90970
rect 3910 90918 3962 90970
rect 4014 90918 4066 90970
rect 23806 90918 23858 90970
rect 23910 90918 23962 90970
rect 24014 90918 24066 90970
rect 9998 90750 10050 90802
rect 15262 90750 15314 90802
rect 2718 90638 2770 90690
rect 6078 90638 6130 90690
rect 22318 90638 22370 90690
rect 6526 90526 6578 90578
rect 6862 90526 6914 90578
rect 7534 90526 7586 90578
rect 8094 90526 8146 90578
rect 9214 90526 9266 90578
rect 11678 90526 11730 90578
rect 13582 90526 13634 90578
rect 16046 90526 16098 90578
rect 16494 90526 16546 90578
rect 17166 90526 17218 90578
rect 17726 90526 17778 90578
rect 18846 90526 18898 90578
rect 7086 90414 7138 90466
rect 12798 90414 12850 90466
rect 13134 90414 13186 90466
rect 15710 90414 15762 90466
rect 21534 90414 21586 90466
rect 22094 90414 22146 90466
rect 1150 90302 1202 90354
rect 2270 90302 2322 90354
rect 11118 90302 11170 90354
rect 14142 90302 14194 90354
rect 16718 90302 16770 90354
rect 22654 90302 22706 90354
rect 4466 90134 4518 90186
rect 4570 90134 4622 90186
rect 4674 90134 4726 90186
rect 24466 90134 24518 90186
rect 24570 90134 24622 90186
rect 24674 90134 24726 90186
rect 4062 89966 4114 90018
rect 12238 89966 12290 90018
rect 13918 89966 13970 90018
rect 1598 89854 1650 89906
rect 4510 89854 4562 89906
rect 6750 89854 6802 89906
rect 7198 89854 7250 89906
rect 10110 89854 10162 89906
rect 12574 89854 12626 89906
rect 14366 89854 14418 89906
rect 18286 89854 18338 89906
rect 19518 89854 19570 89906
rect 30270 89854 30322 89906
rect 30606 89854 30658 89906
rect 1486 89742 1538 89794
rect 2270 89742 2322 89794
rect 3502 89742 3554 89794
rect 3838 89742 3890 89794
rect 5294 89742 5346 89794
rect 6190 89742 6242 89794
rect 13246 89742 13298 89794
rect 13806 89742 13858 89794
rect 14590 89742 14642 89794
rect 15038 89742 15090 89794
rect 16046 89742 16098 89794
rect 18734 89742 18786 89794
rect 19406 89742 19458 89794
rect 20190 89742 20242 89794
rect 3054 89630 3106 89682
rect 7534 89630 7586 89682
rect 9662 89630 9714 89682
rect 12910 89630 12962 89682
rect 2606 89518 2658 89570
rect 7870 89518 7922 89570
rect 11230 89518 11282 89570
rect 17166 89518 17218 89570
rect 20526 89518 20578 89570
rect 3806 89350 3858 89402
rect 3910 89350 3962 89402
rect 4014 89350 4066 89402
rect 23806 89350 23858 89402
rect 23910 89350 23962 89402
rect 24014 89350 24066 89402
rect 14590 89182 14642 89234
rect 18174 89182 18226 89234
rect 5854 89070 5906 89122
rect 9662 89070 9714 89122
rect 13022 89070 13074 89122
rect 2606 88958 2658 89010
rect 6190 88958 6242 89010
rect 6638 88958 6690 89010
rect 7310 88958 7362 89010
rect 8094 88958 8146 89010
rect 8990 88958 9042 89010
rect 17502 88958 17554 89010
rect 21422 88958 21474 89010
rect 3166 88846 3218 88898
rect 6862 88846 6914 88898
rect 9998 88846 10050 88898
rect 13358 88846 13410 88898
rect 17390 88846 17442 88898
rect 21982 88846 22034 88898
rect 4286 88734 4338 88786
rect 11230 88734 11282 88786
rect 18510 88734 18562 88786
rect 23102 88734 23154 88786
rect 30270 88734 30322 88786
rect 30606 88734 30658 88786
rect 4466 88566 4518 88618
rect 4570 88566 4622 88618
rect 4674 88566 4726 88618
rect 24466 88566 24518 88618
rect 24570 88566 24622 88618
rect 24674 88566 24726 88618
rect 1710 88398 1762 88450
rect 21758 88398 21810 88450
rect 29822 88398 29874 88450
rect 4286 88286 4338 88338
rect 11454 88286 11506 88338
rect 13694 88286 13746 88338
rect 18398 88286 18450 88338
rect 3614 88174 3666 88226
rect 4062 88174 4114 88226
rect 4846 88174 4898 88226
rect 5294 88174 5346 88226
rect 6414 88174 6466 88226
rect 13246 88174 13298 88226
rect 21198 88174 21250 88226
rect 29486 88174 29538 88226
rect 1262 88062 1314 88114
rect 3278 88062 3330 88114
rect 7310 88062 7362 88114
rect 11006 88062 11058 88114
rect 18062 88062 18114 88114
rect 2830 87950 2882 88002
rect 12574 87950 12626 88002
rect 14814 87950 14866 88002
rect 19630 87950 19682 88002
rect 22878 87950 22930 88002
rect 3806 87782 3858 87834
rect 3910 87782 3962 87834
rect 4014 87782 4066 87834
rect 23806 87782 23858 87834
rect 23910 87782 23962 87834
rect 24014 87782 24066 87834
rect 1822 87502 1874 87554
rect 6302 87502 6354 87554
rect 12238 87502 12290 87554
rect 13134 87502 13186 87554
rect 22318 87502 22370 87554
rect 9102 87390 9154 87442
rect 10110 87390 10162 87442
rect 10782 87390 10834 87442
rect 11454 87390 11506 87442
rect 11790 87390 11842 87442
rect 14702 87390 14754 87442
rect 18286 87390 18338 87442
rect 22878 87390 22930 87442
rect 30270 87390 30322 87442
rect 2158 87278 2210 87330
rect 6638 87278 6690 87330
rect 11230 87278 11282 87330
rect 21870 87278 21922 87330
rect 23214 87278 23266 87330
rect 23886 87278 23938 87330
rect 3390 87166 3442 87218
rect 7870 87166 7922 87218
rect 13582 87166 13634 87218
rect 18846 87166 18898 87218
rect 19966 87166 20018 87218
rect 20750 87166 20802 87218
rect 23550 87166 23602 87218
rect 30606 87166 30658 87218
rect 4466 86998 4518 87050
rect 4570 86998 4622 87050
rect 4674 86998 4726 87050
rect 24466 86998 24518 87050
rect 24570 86998 24622 87050
rect 24674 86998 24726 87050
rect 6414 86830 6466 86882
rect 9886 86830 9938 86882
rect 22878 86830 22930 86882
rect 1598 86718 1650 86770
rect 4174 86718 4226 86770
rect 11454 86718 11506 86770
rect 12462 86718 12514 86770
rect 12910 86718 12962 86770
rect 18846 86718 18898 86770
rect 19854 86718 19906 86770
rect 23438 86718 23490 86770
rect 30606 86718 30658 86770
rect 3726 86606 3778 86658
rect 5966 86606 6018 86658
rect 9438 86606 9490 86658
rect 11006 86606 11058 86658
rect 11790 86606 11842 86658
rect 12350 86606 12402 86658
rect 13470 86606 13522 86658
rect 14590 86606 14642 86658
rect 19294 86606 19346 86658
rect 19630 86606 19682 86658
rect 20526 86606 20578 86658
rect 20862 86606 20914 86658
rect 21870 86606 21922 86658
rect 22766 86606 22818 86658
rect 22990 86606 23042 86658
rect 23550 86606 23602 86658
rect 30270 86606 30322 86658
rect 1262 86494 1314 86546
rect 23998 86494 24050 86546
rect 2830 86382 2882 86434
rect 5294 86382 5346 86434
rect 7534 86382 7586 86434
rect 22542 86382 22594 86434
rect 23438 86382 23490 86434
rect 23886 86382 23938 86434
rect 3806 86214 3858 86266
rect 3910 86214 3962 86266
rect 4014 86214 4066 86266
rect 23806 86214 23858 86266
rect 23910 86214 23962 86266
rect 24014 86214 24066 86266
rect 19966 86046 20018 86098
rect 23326 86046 23378 86098
rect 2718 85934 2770 85986
rect 7086 85934 7138 85986
rect 7982 85934 8034 85986
rect 13022 85934 13074 85986
rect 15150 85934 15202 85986
rect 22318 85934 22370 85986
rect 1262 85822 1314 85874
rect 8430 85822 8482 85874
rect 8878 85822 8930 85874
rect 9438 85822 9490 85874
rect 10222 85822 10274 85874
rect 11006 85822 11058 85874
rect 15486 85822 15538 85874
rect 16046 85822 16098 85874
rect 17166 85822 17218 85874
rect 18174 85822 18226 85874
rect 19630 85822 19682 85874
rect 22878 85822 22930 85874
rect 23102 85822 23154 85874
rect 23550 85822 23602 85874
rect 23774 85822 23826 85874
rect 1038 85710 1090 85762
rect 6750 85710 6802 85762
rect 8990 85710 9042 85762
rect 13470 85710 13522 85762
rect 14590 85710 14642 85762
rect 16158 85710 16210 85762
rect 16606 85710 16658 85762
rect 19070 85710 19122 85762
rect 19406 85710 19458 85762
rect 20750 85710 20802 85762
rect 24110 85710 24162 85762
rect 24446 85710 24498 85762
rect 1822 85598 1874 85650
rect 2158 85598 2210 85650
rect 3166 85598 3218 85650
rect 4286 85598 4338 85650
rect 5518 85598 5570 85650
rect 21870 85598 21922 85650
rect 23886 85598 23938 85650
rect 4466 85430 4518 85482
rect 4570 85430 4622 85482
rect 4674 85430 4726 85482
rect 24466 85430 24518 85482
rect 24570 85430 24622 85482
rect 24674 85430 24726 85482
rect 17390 85262 17442 85314
rect 20414 85262 20466 85314
rect 23102 85262 23154 85314
rect 23550 85262 23602 85314
rect 1038 85150 1090 85202
rect 2830 85150 2882 85202
rect 6750 85150 6802 85202
rect 11230 85150 11282 85202
rect 13918 85150 13970 85202
rect 22990 85150 23042 85202
rect 23886 85150 23938 85202
rect 30270 85150 30322 85202
rect 30606 85150 30658 85202
rect 1374 85038 1426 85090
rect 2270 85038 2322 85090
rect 2606 85038 2658 85090
rect 3502 85038 3554 85090
rect 3838 85038 3890 85090
rect 4846 85038 4898 85090
rect 7198 85038 7250 85090
rect 10894 85038 10946 85090
rect 12462 85038 12514 85090
rect 13246 85038 13298 85090
rect 13806 85038 13858 85090
rect 14590 85038 14642 85090
rect 14926 85038 14978 85090
rect 16046 85038 16098 85090
rect 16830 85038 16882 85090
rect 19742 85038 19794 85090
rect 20190 85038 20242 85090
rect 21086 85038 21138 85090
rect 21422 85038 21474 85090
rect 22542 85038 22594 85090
rect 1822 84926 1874 84978
rect 12910 84926 12962 84978
rect 19406 84926 19458 84978
rect 5518 84814 5570 84866
rect 18510 84814 18562 84866
rect 3806 84646 3858 84698
rect 3910 84646 3962 84698
rect 4014 84646 4066 84698
rect 23806 84646 23858 84698
rect 23910 84646 23962 84698
rect 24014 84646 24066 84698
rect 7422 84366 7474 84418
rect 11342 84366 11394 84418
rect 15038 84366 15090 84418
rect 20638 84366 20690 84418
rect 1486 84254 1538 84306
rect 2046 84254 2098 84306
rect 2830 84254 2882 84306
rect 3166 84254 3218 84306
rect 3390 84254 3442 84306
rect 4174 84254 4226 84306
rect 5294 84254 5346 84306
rect 7870 84254 7922 84306
rect 8206 84254 8258 84306
rect 8878 84254 8930 84306
rect 9662 84254 9714 84306
rect 10558 84254 10610 84306
rect 15374 84254 15426 84306
rect 15934 84254 15986 84306
rect 16494 84254 16546 84306
rect 17054 84254 17106 84306
rect 17278 84254 17330 84306
rect 18062 84254 18114 84306
rect 19070 84254 19122 84306
rect 20974 84254 21026 84306
rect 21422 84254 21474 84306
rect 22094 84254 22146 84306
rect 22654 84254 22706 84306
rect 23662 84254 23714 84306
rect 1150 84142 1202 84194
rect 5854 84142 5906 84194
rect 13022 84142 13074 84194
rect 16046 84142 16098 84194
rect 19294 84142 19346 84194
rect 19630 84142 19682 84194
rect 21646 84142 21698 84194
rect 2158 84030 2210 84082
rect 6974 84030 7026 84082
rect 8430 84030 8482 84082
rect 12798 84030 12850 84082
rect 18734 84030 18786 84082
rect 30270 84030 30322 84082
rect 30606 84030 30658 84082
rect 4466 83862 4518 83914
rect 4570 83862 4622 83914
rect 4674 83862 4726 83914
rect 24466 83862 24518 83914
rect 24570 83862 24622 83914
rect 24674 83862 24726 83914
rect 1374 83694 1426 83746
rect 4286 83694 4338 83746
rect 9886 83694 9938 83746
rect 22094 83694 22146 83746
rect 23662 83694 23714 83746
rect 2382 83582 2434 83634
rect 3950 83582 4002 83634
rect 6078 83582 6130 83634
rect 6526 83582 6578 83634
rect 8878 83582 8930 83634
rect 14926 83582 14978 83634
rect 16718 83582 16770 83634
rect 17726 83582 17778 83634
rect 20862 83582 20914 83634
rect 30606 83582 30658 83634
rect 1038 83470 1090 83522
rect 1822 83470 1874 83522
rect 5406 83470 5458 83522
rect 5854 83470 5906 83522
rect 7310 83470 7362 83522
rect 8094 83470 8146 83522
rect 9214 83470 9266 83522
rect 9662 83470 9714 83522
rect 10334 83470 10386 83522
rect 11118 83470 11170 83522
rect 12014 83470 12066 83522
rect 13918 83470 13970 83522
rect 16046 83470 16098 83522
rect 17054 83470 17106 83522
rect 17502 83470 17554 83522
rect 18398 83470 18450 83522
rect 18734 83470 18786 83522
rect 19742 83470 19794 83522
rect 20414 83470 20466 83522
rect 23326 83470 23378 83522
rect 30270 83470 30322 83522
rect 5070 83358 5122 83410
rect 14478 83358 14530 83410
rect 3502 83246 3554 83298
rect 13358 83246 13410 83298
rect 13470 83246 13522 83298
rect 13694 83246 13746 83298
rect 3806 83078 3858 83130
rect 3910 83078 3962 83130
rect 4014 83078 4066 83130
rect 23806 83078 23858 83130
rect 23910 83078 23962 83130
rect 24014 83078 24066 83130
rect 9886 82910 9938 82962
rect 17726 82910 17778 82962
rect 5854 82798 5906 82850
rect 1598 82686 1650 82738
rect 1934 82686 1986 82738
rect 2830 82686 2882 82738
rect 3166 82686 3218 82738
rect 4174 82686 4226 82738
rect 8318 82686 8370 82738
rect 10558 82686 10610 82738
rect 14478 82686 14530 82738
rect 16046 82686 16098 82738
rect 18286 82686 18338 82738
rect 1150 82574 1202 82626
rect 6190 82574 6242 82626
rect 8766 82574 8818 82626
rect 10894 82574 10946 82626
rect 14142 82574 14194 82626
rect 16494 82574 16546 82626
rect 22878 82574 22930 82626
rect 2158 82462 2210 82514
rect 4958 82462 5010 82514
rect 5294 82462 5346 82514
rect 7422 82462 7474 82514
rect 12126 82462 12178 82514
rect 12910 82462 12962 82514
rect 18510 82462 18562 82514
rect 22542 82462 22594 82514
rect 4466 82294 4518 82346
rect 4570 82294 4622 82346
rect 4674 82294 4726 82346
rect 24466 82294 24518 82346
rect 24570 82294 24622 82346
rect 24674 82294 24726 82346
rect 8318 82126 8370 82178
rect 8990 82126 9042 82178
rect 2158 82014 2210 82066
rect 3726 82014 3778 82066
rect 4734 82014 4786 82066
rect 5182 82014 5234 82066
rect 7310 82014 7362 82066
rect 7982 82014 8034 82066
rect 10222 82014 10274 82066
rect 12014 82014 12066 82066
rect 13022 82014 13074 82066
rect 13470 82014 13522 82066
rect 15710 82014 15762 82066
rect 19966 82014 20018 82066
rect 22766 82014 22818 82066
rect 29822 82014 29874 82066
rect 30270 82014 30322 82066
rect 30606 82014 30658 82066
rect 4062 81902 4114 81954
rect 4510 81902 4562 81954
rect 5742 81902 5794 81954
rect 6750 81902 6802 81954
rect 7534 81902 7586 81954
rect 10670 81902 10722 81954
rect 12350 81902 12402 81954
rect 12798 81902 12850 81954
rect 14254 81902 14306 81954
rect 15038 81902 15090 81954
rect 15486 81902 15538 81954
rect 15822 81902 15874 81954
rect 19406 81902 19458 81954
rect 29486 81902 29538 81954
rect 1710 81790 1762 81842
rect 23214 81790 23266 81842
rect 3278 81678 3330 81730
rect 21086 81678 21138 81730
rect 21646 81678 21698 81730
rect 3806 81510 3858 81562
rect 3910 81510 3962 81562
rect 4014 81510 4066 81562
rect 23806 81510 23858 81562
rect 23910 81510 23962 81562
rect 24014 81510 24066 81562
rect 10894 81230 10946 81282
rect 15710 81230 15762 81282
rect 20862 81230 20914 81282
rect 1710 81118 1762 81170
rect 6190 81118 6242 81170
rect 8542 81118 8594 81170
rect 12910 81118 12962 81170
rect 14590 81118 14642 81170
rect 15038 81118 15090 81170
rect 2046 81006 2098 81058
rect 6638 81006 6690 81058
rect 8878 81006 8930 81058
rect 10558 81006 10610 81058
rect 16046 81006 16098 81058
rect 21198 81006 21250 81058
rect 3278 80894 3330 80946
rect 3950 80894 4002 80946
rect 4286 80894 4338 80946
rect 4958 80894 5010 80946
rect 5294 80894 5346 80946
rect 7870 80894 7922 80946
rect 10110 80894 10162 80946
rect 10782 80894 10834 80946
rect 13470 80894 13522 80946
rect 15150 80894 15202 80946
rect 16158 80894 16210 80946
rect 17278 80894 17330 80946
rect 22430 80894 22482 80946
rect 30270 80894 30322 80946
rect 30606 80894 30658 80946
rect 4466 80726 4518 80778
rect 4570 80726 4622 80778
rect 4674 80726 4726 80778
rect 24466 80726 24518 80778
rect 24570 80726 24622 80778
rect 24674 80726 24726 80778
rect 12910 80558 12962 80610
rect 14030 80558 14082 80610
rect 14926 80558 14978 80610
rect 18846 80558 18898 80610
rect 21422 80558 21474 80610
rect 29822 80558 29874 80610
rect 2494 80446 2546 80498
rect 2942 80446 2994 80498
rect 5070 80446 5122 80498
rect 6078 80446 6130 80498
rect 6526 80446 6578 80498
rect 9886 80446 9938 80498
rect 15038 80446 15090 80498
rect 15262 80446 15314 80498
rect 20414 80446 20466 80498
rect 21870 80446 21922 80498
rect 1934 80334 1986 80386
rect 2382 80334 2434 80386
rect 3614 80334 3666 80386
rect 4510 80334 4562 80386
rect 5518 80334 5570 80386
rect 5854 80334 5906 80386
rect 7086 80334 7138 80386
rect 8094 80334 8146 80386
rect 12350 80334 12402 80386
rect 14478 80334 14530 80386
rect 14814 80334 14866 80386
rect 18398 80334 18450 80386
rect 20862 80334 20914 80386
rect 21198 80334 21250 80386
rect 22654 80334 22706 80386
rect 23550 80334 23602 80386
rect 29486 80334 29538 80386
rect 1486 80222 1538 80274
rect 9550 80222 9602 80274
rect 11118 80110 11170 80162
rect 19966 80110 20018 80162
rect 3806 79942 3858 79994
rect 3910 79942 3962 79994
rect 4014 79942 4066 79994
rect 23806 79942 23858 79994
rect 23910 79942 23962 79994
rect 24014 79942 24066 79994
rect 14366 79774 14418 79826
rect 8430 79662 8482 79714
rect 20638 79662 20690 79714
rect 1262 79550 1314 79602
rect 3390 79550 3442 79602
rect 4286 79550 4338 79602
rect 7198 79550 7250 79602
rect 8766 79550 8818 79602
rect 9214 79550 9266 79602
rect 9998 79550 10050 79602
rect 10670 79550 10722 79602
rect 11454 79550 11506 79602
rect 12238 79550 12290 79602
rect 14366 79550 14418 79602
rect 15598 79550 15650 79602
rect 15934 79550 15986 79602
rect 16382 79550 16434 79602
rect 17278 79550 17330 79602
rect 17838 79550 17890 79602
rect 18622 79550 18674 79602
rect 20974 79550 21026 79602
rect 21422 79550 21474 79602
rect 22318 79550 22370 79602
rect 22654 79550 22706 79602
rect 23774 79550 23826 79602
rect 6750 79438 6802 79490
rect 12126 79438 12178 79490
rect 14030 79438 14082 79490
rect 16606 79438 16658 79490
rect 22094 79438 22146 79490
rect 1710 79326 1762 79378
rect 2830 79326 2882 79378
rect 3614 79326 3666 79378
rect 4062 79326 4114 79378
rect 5630 79326 5682 79378
rect 7758 79326 7810 79378
rect 8094 79326 8146 79378
rect 9438 79326 9490 79378
rect 11902 79326 11954 79378
rect 21646 79326 21698 79378
rect 29486 79326 29538 79378
rect 29822 79326 29874 79378
rect 30270 79326 30322 79378
rect 30606 79326 30658 79378
rect 4466 79158 4518 79210
rect 4570 79158 4622 79210
rect 4674 79158 4726 79210
rect 24466 79158 24518 79210
rect 24570 79158 24622 79210
rect 24674 79158 24726 79210
rect 11454 78990 11506 79042
rect 15934 78990 15986 79042
rect 17726 78990 17778 79042
rect 2382 78878 2434 78930
rect 3950 78878 4002 78930
rect 5518 78878 5570 78930
rect 6862 78878 6914 78930
rect 9550 78878 9602 78930
rect 11678 78878 11730 78930
rect 11902 78878 11954 78930
rect 14814 78878 14866 78930
rect 16718 78878 16770 78930
rect 20302 78878 20354 78930
rect 21310 78878 21362 78930
rect 30606 78878 30658 78930
rect 2718 78766 2770 78818
rect 5854 78766 5906 78818
rect 6414 78766 6466 78818
rect 11118 78766 11170 78818
rect 12686 78766 12738 78818
rect 14254 78766 14306 78818
rect 17054 78766 17106 78818
rect 17502 78766 17554 78818
rect 18174 78766 18226 78818
rect 18734 78766 18786 78818
rect 19742 78766 19794 78818
rect 20750 78766 20802 78818
rect 21086 78766 21138 78818
rect 21982 78766 22034 78818
rect 22318 78766 22370 78818
rect 23326 78766 23378 78818
rect 30270 78766 30322 78818
rect 3502 78654 3554 78706
rect 9102 78654 9154 78706
rect 14366 78654 14418 78706
rect 1150 78542 1202 78594
rect 5070 78542 5122 78594
rect 8094 78542 8146 78594
rect 10670 78542 10722 78594
rect 11454 78542 11506 78594
rect 12238 78542 12290 78594
rect 12350 78542 12402 78594
rect 12574 78542 12626 78594
rect 3806 78374 3858 78426
rect 3910 78374 3962 78426
rect 4014 78374 4066 78426
rect 23806 78374 23858 78426
rect 23910 78374 23962 78426
rect 24014 78374 24066 78426
rect 12126 78206 12178 78258
rect 17614 78206 17666 78258
rect 1262 78094 1314 78146
rect 9438 78094 9490 78146
rect 10110 78094 10162 78146
rect 12238 78094 12290 78146
rect 13022 78094 13074 78146
rect 4174 77982 4226 78034
rect 5630 77982 5682 78034
rect 7870 77982 7922 78034
rect 15486 77982 15538 78034
rect 19182 77982 19234 78034
rect 22430 77982 22482 78034
rect 1710 77870 1762 77922
rect 6078 77870 6130 77922
rect 8318 77870 8370 77922
rect 13358 77870 13410 77922
rect 15934 77870 15986 77922
rect 21870 77870 21922 77922
rect 29486 77870 29538 77922
rect 29822 77870 29874 77922
rect 2830 77758 2882 77810
rect 3278 77758 3330 77810
rect 3614 77758 3666 77810
rect 3950 77758 4002 77810
rect 7198 77758 7250 77810
rect 10558 77758 10610 77810
rect 11678 77758 11730 77810
rect 14590 77758 14642 77810
rect 17054 77758 17106 77810
rect 18734 77758 18786 77810
rect 20750 77758 20802 77810
rect 4466 77590 4518 77642
rect 4570 77590 4622 77642
rect 4674 77590 4726 77642
rect 24466 77590 24518 77642
rect 24570 77590 24622 77642
rect 24674 77590 24726 77642
rect 6638 77422 6690 77474
rect 20190 77422 20242 77474
rect 1038 77310 1090 77362
rect 1710 77310 1762 77362
rect 3390 77310 3442 77362
rect 9214 77310 9266 77362
rect 9886 77310 9938 77362
rect 10894 77310 10946 77362
rect 13470 77310 13522 77362
rect 14814 77310 14866 77362
rect 17390 77310 17442 77362
rect 21198 77310 21250 77362
rect 21646 77310 21698 77362
rect 1374 77198 1426 77250
rect 2046 77198 2098 77250
rect 2382 77198 2434 77250
rect 2718 77198 2770 77250
rect 3166 77198 3218 77250
rect 3838 77198 3890 77250
rect 4398 77198 4450 77250
rect 5406 77198 5458 77250
rect 9550 77198 9602 77250
rect 10334 77198 10386 77250
rect 10782 77198 10834 77250
rect 11566 77198 11618 77250
rect 11902 77198 11954 77250
rect 12910 77198 12962 77250
rect 13806 77198 13858 77250
rect 14366 77198 14418 77250
rect 16046 77198 16098 77250
rect 16830 77198 16882 77250
rect 19966 77198 20018 77250
rect 20638 77198 20690 77250
rect 6190 77086 6242 77138
rect 20974 77086 21026 77138
rect 7758 76974 7810 77026
rect 18510 76974 18562 77026
rect 3806 76806 3858 76858
rect 3910 76806 3962 76858
rect 4014 76806 4066 76858
rect 23806 76806 23858 76858
rect 23910 76806 23962 76858
rect 24014 76806 24066 76858
rect 1934 76526 1986 76578
rect 6638 76526 6690 76578
rect 12910 76526 12962 76578
rect 16494 76526 16546 76578
rect 5070 76414 5122 76466
rect 7086 76414 7138 76466
rect 7422 76414 7474 76466
rect 8094 76414 8146 76466
rect 8878 76414 8930 76466
rect 9774 76414 9826 76466
rect 10446 76414 10498 76466
rect 12126 76414 12178 76466
rect 13246 76414 13298 76466
rect 13694 76414 13746 76466
rect 14590 76414 14642 76466
rect 14926 76414 14978 76466
rect 15934 76414 15986 76466
rect 16942 76414 16994 76466
rect 17278 76414 17330 76466
rect 18174 76414 18226 76466
rect 18622 76414 18674 76466
rect 19518 76414 19570 76466
rect 22318 76414 22370 76466
rect 2382 76302 2434 76354
rect 7646 76302 7698 76354
rect 10894 76302 10946 76354
rect 13918 76302 13970 76354
rect 21870 76302 21922 76354
rect 1038 76190 1090 76242
rect 1374 76190 1426 76242
rect 3502 76190 3554 76242
rect 3950 76190 4002 76242
rect 4286 76190 4338 76242
rect 5294 76190 5346 76242
rect 5630 76190 5682 76242
rect 5966 76190 6018 76242
rect 17502 76190 17554 76242
rect 20750 76190 20802 76242
rect 4466 76022 4518 76074
rect 4570 76022 4622 76074
rect 4674 76022 4726 76074
rect 24466 76022 24518 76074
rect 24570 76022 24622 76074
rect 24674 76022 24726 76074
rect 3166 75854 3218 75906
rect 7086 75854 7138 75906
rect 11678 75854 11730 75906
rect 13022 75854 13074 75906
rect 17502 75854 17554 75906
rect 20078 75854 20130 75906
rect 1038 75742 1090 75794
rect 3614 75742 3666 75794
rect 20414 75742 20466 75794
rect 20750 75742 20802 75794
rect 21758 75742 21810 75794
rect 1374 75630 1426 75682
rect 2158 75630 2210 75682
rect 2606 75630 2658 75682
rect 2942 75630 2994 75682
rect 4174 75630 4226 75682
rect 5182 75630 5234 75682
rect 6638 75630 6690 75682
rect 8206 75630 8258 75682
rect 12014 75630 12066 75682
rect 18622 75630 18674 75682
rect 21086 75630 21138 75682
rect 21534 75630 21586 75682
rect 22430 75630 22482 75682
rect 22990 75630 23042 75682
rect 23774 75630 23826 75682
rect 12574 75518 12626 75570
rect 17054 75518 17106 75570
rect 14142 75406 14194 75458
rect 3806 75238 3858 75290
rect 3910 75238 3962 75290
rect 4014 75238 4066 75290
rect 23806 75238 23858 75290
rect 23910 75238 23962 75290
rect 24014 75238 24066 75290
rect 1822 74958 1874 75010
rect 6078 74958 6130 75010
rect 26910 74958 26962 75010
rect 4398 74846 4450 74898
rect 5406 74846 5458 74898
rect 8318 74846 8370 74898
rect 10558 74846 10610 74898
rect 12126 74846 12178 74898
rect 13134 74846 13186 74898
rect 13582 74846 13634 74898
rect 14254 74846 14306 74898
rect 14926 74846 14978 74898
rect 15822 74846 15874 74898
rect 17054 74846 17106 74898
rect 17614 74846 17666 74898
rect 18398 74846 18450 74898
rect 18846 74846 18898 74898
rect 19742 74846 19794 74898
rect 22878 74846 22930 74898
rect 2270 74734 2322 74786
rect 6526 74734 6578 74786
rect 8094 74734 8146 74786
rect 11006 74734 11058 74786
rect 12798 74734 12850 74786
rect 13806 74734 13858 74786
rect 16718 74734 16770 74786
rect 27694 74734 27746 74786
rect 3390 74622 3442 74674
rect 4062 74622 4114 74674
rect 5182 74622 5234 74674
rect 7646 74622 7698 74674
rect 17726 74622 17778 74674
rect 30270 74622 30322 74674
rect 30606 74622 30658 74674
rect 4466 74454 4518 74506
rect 4570 74454 4622 74506
rect 4674 74454 4726 74506
rect 24466 74454 24518 74506
rect 24570 74454 24622 74506
rect 24674 74454 24726 74506
rect 3950 74286 4002 74338
rect 7534 74286 7586 74338
rect 8206 74286 8258 74338
rect 16046 74286 16098 74338
rect 16718 74286 16770 74338
rect 17054 74286 17106 74338
rect 22990 74286 23042 74338
rect 1038 74174 1090 74226
rect 2158 74174 2210 74226
rect 2942 74174 2994 74226
rect 6526 74174 6578 74226
rect 7198 74174 7250 74226
rect 9438 74174 9490 74226
rect 11790 74174 11842 74226
rect 14814 74174 14866 74226
rect 18622 74174 18674 74226
rect 21758 74174 21810 74226
rect 30606 74174 30658 74226
rect 1374 74062 1426 74114
rect 1934 74062 1986 74114
rect 3278 74062 3330 74114
rect 3838 74062 3890 74114
rect 4622 74062 4674 74114
rect 5070 74062 5122 74114
rect 5966 74062 6018 74114
rect 6862 74062 6914 74114
rect 7982 74062 8034 74114
rect 8318 74062 8370 74114
rect 8990 74062 9042 74114
rect 14478 74062 14530 74114
rect 18062 74062 18114 74114
rect 18398 74062 18450 74114
rect 19294 74062 19346 74114
rect 19742 74062 19794 74114
rect 20638 74062 20690 74114
rect 21422 74062 21474 74114
rect 30270 74062 30322 74114
rect 11454 73950 11506 74002
rect 17614 73950 17666 74002
rect 10670 73838 10722 73890
rect 13022 73838 13074 73890
rect 3806 73670 3858 73722
rect 3910 73670 3962 73722
rect 4014 73670 4066 73722
rect 23806 73670 23858 73722
rect 23910 73670 23962 73722
rect 24014 73670 24066 73722
rect 10558 73502 10610 73554
rect 18398 73502 18450 73554
rect 10222 73390 10274 73442
rect 11342 73390 11394 73442
rect 12798 73390 12850 73442
rect 1822 73278 1874 73330
rect 4174 73278 4226 73330
rect 5854 73278 5906 73330
rect 7198 73278 7250 73330
rect 8094 73278 8146 73330
rect 8542 73278 8594 73330
rect 9326 73278 9378 73330
rect 9774 73278 9826 73330
rect 13134 73278 13186 73330
rect 13694 73278 13746 73330
rect 15038 73278 15090 73330
rect 15822 73278 15874 73330
rect 16830 73278 16882 73330
rect 2270 73166 2322 73218
rect 3838 73166 3890 73218
rect 4958 73166 5010 73218
rect 10782 73166 10834 73218
rect 11230 73166 11282 73218
rect 11902 73166 11954 73218
rect 14254 73166 14306 73218
rect 20638 73166 20690 73218
rect 23326 73166 23378 73218
rect 3390 73054 3442 73106
rect 5294 73054 5346 73106
rect 5630 73054 5682 73106
rect 6302 73054 6354 73106
rect 6638 73054 6690 73106
rect 9214 73054 9266 73106
rect 10670 73054 10722 73106
rect 12238 73054 12290 73106
rect 13806 73054 13858 73106
rect 17278 73054 17330 73106
rect 20974 73054 21026 73106
rect 22990 73054 23042 73106
rect 4466 72886 4518 72938
rect 4570 72886 4622 72938
rect 4674 72886 4726 72938
rect 24466 72886 24518 72938
rect 24570 72886 24622 72938
rect 24674 72886 24726 72938
rect 3054 72718 3106 72770
rect 9438 72718 9490 72770
rect 10334 72718 10386 72770
rect 12798 72718 12850 72770
rect 17390 72718 17442 72770
rect 17726 72718 17778 72770
rect 21534 72718 21586 72770
rect 1038 72606 1090 72658
rect 3502 72606 3554 72658
rect 6302 72606 6354 72658
rect 7870 72606 7922 72658
rect 9886 72606 9938 72658
rect 11678 72606 11730 72658
rect 13918 72606 13970 72658
rect 18846 72606 18898 72658
rect 30606 72606 30658 72658
rect 1374 72494 1426 72546
rect 2382 72494 2434 72546
rect 2942 72494 2994 72546
rect 4286 72494 4338 72546
rect 5070 72494 5122 72546
rect 5854 72494 5906 72546
rect 8206 72494 8258 72546
rect 9550 72494 9602 72546
rect 10110 72494 10162 72546
rect 10334 72494 10386 72546
rect 10670 72494 10722 72546
rect 11230 72494 11282 72546
rect 13470 72494 13522 72546
rect 18398 72494 18450 72546
rect 20078 72494 20130 72546
rect 20862 72494 20914 72546
rect 21310 72494 21362 72546
rect 22206 72494 22258 72546
rect 22654 72494 22706 72546
rect 23662 72494 23714 72546
rect 30270 72494 30322 72546
rect 2046 72382 2098 72434
rect 9326 72382 9378 72434
rect 20526 72382 20578 72434
rect 7422 72270 7474 72322
rect 9102 72270 9154 72322
rect 15038 72270 15090 72322
rect 3806 72102 3858 72154
rect 3910 72102 3962 72154
rect 4014 72102 4066 72154
rect 23806 72102 23858 72154
rect 23910 72102 23962 72154
rect 24014 72102 24066 72154
rect 9774 71934 9826 71986
rect 19966 71934 20018 71986
rect 22654 71934 22706 71986
rect 6078 71822 6130 71874
rect 11342 71822 11394 71874
rect 14590 71822 14642 71874
rect 1262 71710 1314 71762
rect 2718 71710 2770 71762
rect 4286 71710 4338 71762
rect 6414 71710 6466 71762
rect 6974 71710 7026 71762
rect 7646 71710 7698 71762
rect 8094 71710 8146 71762
rect 9214 71710 9266 71762
rect 15038 71710 15090 71762
rect 15486 71710 15538 71762
rect 16718 71710 16770 71762
rect 17614 71710 17666 71762
rect 18286 71710 18338 71762
rect 21086 71710 21138 71762
rect 23214 71710 23266 71762
rect 30382 71710 30434 71762
rect 3166 71598 3218 71650
rect 10894 71598 10946 71650
rect 13918 71598 13970 71650
rect 16046 71598 16098 71650
rect 21422 71598 21474 71650
rect 23438 71598 23490 71650
rect 1038 71486 1090 71538
rect 1710 71486 1762 71538
rect 2046 71486 2098 71538
rect 4958 71486 5010 71538
rect 5294 71486 5346 71538
rect 7086 71486 7138 71538
rect 14254 71486 14306 71538
rect 15598 71486 15650 71538
rect 18846 71486 18898 71538
rect 30606 71486 30658 71538
rect 4466 71318 4518 71370
rect 4570 71318 4622 71370
rect 4674 71318 4726 71370
rect 24466 71318 24518 71370
rect 24570 71318 24622 71370
rect 24674 71318 24726 71370
rect 6078 71150 6130 71202
rect 16046 71150 16098 71202
rect 29822 71150 29874 71202
rect 2494 71038 2546 71090
rect 8878 71038 8930 71090
rect 11006 71038 11058 71090
rect 14814 71038 14866 71090
rect 21534 71038 21586 71090
rect 30606 71038 30658 71090
rect 1822 70926 1874 70978
rect 2270 70926 2322 70978
rect 3166 70926 3218 70978
rect 3502 70926 3554 70978
rect 4510 70926 4562 70978
rect 5518 70926 5570 70978
rect 5854 70926 5906 70978
rect 6638 70926 6690 70978
rect 7310 70926 7362 70978
rect 8094 70926 8146 70978
rect 9102 70926 9154 70978
rect 14366 70926 14418 70978
rect 21086 70926 21138 70978
rect 29486 70926 29538 70978
rect 30270 70926 30322 70978
rect 1486 70814 1538 70866
rect 5070 70814 5122 70866
rect 11342 70814 11394 70866
rect 18958 70814 19010 70866
rect 9774 70702 9826 70754
rect 22766 70702 22818 70754
rect 3806 70534 3858 70586
rect 3910 70534 3962 70586
rect 4014 70534 4066 70586
rect 23806 70534 23858 70586
rect 23910 70534 23962 70586
rect 24014 70534 24066 70586
rect 5630 70366 5682 70418
rect 7198 70254 7250 70306
rect 8990 70254 9042 70306
rect 15374 70254 15426 70306
rect 1262 70142 1314 70194
rect 3502 70142 3554 70194
rect 4062 70142 4114 70194
rect 7310 70142 7362 70194
rect 9326 70142 9378 70194
rect 9886 70142 9938 70194
rect 10446 70142 10498 70194
rect 11230 70142 11282 70194
rect 12014 70142 12066 70194
rect 17726 70142 17778 70194
rect 21198 70142 21250 70194
rect 3278 70030 3330 70082
rect 4286 70030 4338 70082
rect 7758 70030 7810 70082
rect 8094 70030 8146 70082
rect 14478 70030 14530 70082
rect 18174 70030 18226 70082
rect 19742 70030 19794 70082
rect 1710 69918 1762 69970
rect 2830 69918 2882 69970
rect 6750 69918 6802 69970
rect 9998 69918 10050 69970
rect 14814 69918 14866 69970
rect 15822 69918 15874 69970
rect 16942 69918 16994 69970
rect 19294 69918 19346 69970
rect 20078 69918 20130 69970
rect 21758 69918 21810 69970
rect 22878 69918 22930 69970
rect 4466 69750 4518 69802
rect 4570 69750 4622 69802
rect 4674 69750 4726 69802
rect 24466 69750 24518 69802
rect 24570 69750 24622 69802
rect 24674 69750 24726 69802
rect 8318 69582 8370 69634
rect 8990 69582 9042 69634
rect 10110 69582 10162 69634
rect 11902 69582 11954 69634
rect 22430 69582 22482 69634
rect 1038 69470 1090 69522
rect 2942 69470 2994 69522
rect 3390 69470 3442 69522
rect 6078 69470 6130 69522
rect 7982 69470 8034 69522
rect 14590 69470 14642 69522
rect 17278 69470 17330 69522
rect 19518 69470 19570 69522
rect 30606 69470 30658 69522
rect 1374 69358 1426 69410
rect 2382 69358 2434 69410
rect 2830 69358 2882 69410
rect 3950 69358 4002 69410
rect 4958 69358 5010 69410
rect 12238 69358 12290 69410
rect 16942 69358 16994 69410
rect 19182 69358 19234 69410
rect 22878 69358 22930 69410
rect 23774 69358 23826 69410
rect 30270 69358 30322 69410
rect 1934 69246 1986 69298
rect 5742 69246 5794 69298
rect 10558 69246 10610 69298
rect 14142 69246 14194 69298
rect 7310 69134 7362 69186
rect 15710 69134 15762 69186
rect 18510 69134 18562 69186
rect 20750 69134 20802 69186
rect 21310 69134 21362 69186
rect 23438 69134 23490 69186
rect 23774 69134 23826 69186
rect 3806 68966 3858 69018
rect 3910 68966 3962 69018
rect 4014 68966 4066 69018
rect 23806 68966 23858 69018
rect 23910 68966 23962 69018
rect 24014 68966 24066 69018
rect 5182 68686 5234 68738
rect 10558 68686 10610 68738
rect 14478 68686 14530 68738
rect 19966 68686 20018 68738
rect 20638 68686 20690 68738
rect 24334 68686 24386 68738
rect 1934 68574 1986 68626
rect 4174 68574 4226 68626
rect 7310 68574 7362 68626
rect 9774 68574 9826 68626
rect 15262 68574 15314 68626
rect 15710 68574 15762 68626
rect 16158 68574 16210 68626
rect 16830 68574 16882 68626
rect 17278 68574 17330 68626
rect 18398 68574 18450 68626
rect 19294 68574 19346 68626
rect 19630 68574 19682 68626
rect 19742 68574 19794 68626
rect 20078 68574 20130 68626
rect 21086 68574 21138 68626
rect 21422 68574 21474 68626
rect 22318 68574 22370 68626
rect 22878 68574 22930 68626
rect 23662 68574 23714 68626
rect 24222 68574 24274 68626
rect 24670 68574 24722 68626
rect 24782 68574 24834 68626
rect 2270 68462 2322 68514
rect 5630 68462 5682 68514
rect 7758 68462 7810 68514
rect 10894 68462 10946 68514
rect 14142 68462 14194 68514
rect 16270 68462 16322 68514
rect 18958 68462 19010 68514
rect 19070 68462 19122 68514
rect 21646 68462 21698 68514
rect 24446 68462 24498 68514
rect 29822 68462 29874 68514
rect 1038 68350 1090 68402
rect 1374 68350 1426 68402
rect 3502 68350 3554 68402
rect 3950 68350 4002 68402
rect 6750 68350 6802 68402
rect 8990 68350 9042 68402
rect 9438 68350 9490 68402
rect 12126 68350 12178 68402
rect 12910 68350 12962 68402
rect 29486 68350 29538 68402
rect 30270 68350 30322 68402
rect 30606 68350 30658 68402
rect 4466 68182 4518 68234
rect 4570 68182 4622 68234
rect 4674 68182 4726 68234
rect 24466 68182 24518 68234
rect 24570 68182 24622 68234
rect 24674 68182 24726 68234
rect 1822 68014 1874 68066
rect 5966 68014 6018 68066
rect 9998 68014 10050 68066
rect 13134 68014 13186 68066
rect 15822 68014 15874 68066
rect 21422 68014 21474 68066
rect 29822 68014 29874 68066
rect 1038 67902 1090 67954
rect 3390 67902 3442 67954
rect 4958 67902 5010 67954
rect 12126 67902 12178 67954
rect 13582 67902 13634 67954
rect 16158 67902 16210 67954
rect 16830 67902 16882 67954
rect 17838 67902 17890 67954
rect 21870 67902 21922 67954
rect 1374 67790 1426 67842
rect 2158 67790 2210 67842
rect 4510 67790 4562 67842
rect 5294 67790 5346 67842
rect 5854 67790 5906 67842
rect 6638 67790 6690 67842
rect 6974 67790 7026 67842
rect 7198 67790 7250 67842
rect 8094 67790 8146 67842
rect 12462 67790 12514 67842
rect 12910 67790 12962 67842
rect 14142 67790 14194 67842
rect 15262 67790 15314 67842
rect 17278 67790 17330 67842
rect 17614 67790 17666 67842
rect 18398 67790 18450 67842
rect 18846 67790 18898 67842
rect 19966 67790 20018 67842
rect 20750 67790 20802 67842
rect 21198 67790 21250 67842
rect 22430 67790 22482 67842
rect 23438 67790 23490 67842
rect 29598 67790 29650 67842
rect 2942 67678 2994 67730
rect 9550 67678 9602 67730
rect 20414 67678 20466 67730
rect 11118 67566 11170 67618
rect 3806 67398 3858 67450
rect 3910 67398 3962 67450
rect 4014 67398 4066 67450
rect 23806 67398 23858 67450
rect 23910 67398 23962 67450
rect 24014 67398 24066 67450
rect 2718 67118 2770 67170
rect 6974 67118 7026 67170
rect 14142 67118 14194 67170
rect 19406 67118 19458 67170
rect 21086 67118 21138 67170
rect 22654 67118 22706 67170
rect 23102 67118 23154 67170
rect 23214 67118 23266 67170
rect 9662 67006 9714 67058
rect 14590 67006 14642 67058
rect 14926 67006 14978 67058
rect 15822 67006 15874 67058
rect 16158 67006 16210 67058
rect 17166 67006 17218 67058
rect 30382 67006 30434 67058
rect 1486 66894 1538 66946
rect 1822 66894 1874 66946
rect 3054 66894 3106 66946
rect 7310 66894 7362 66946
rect 9998 66894 10050 66946
rect 19070 66894 19122 66946
rect 21422 66894 21474 66946
rect 1150 66782 1202 66834
rect 2158 66782 2210 66834
rect 4286 66782 4338 66834
rect 8542 66782 8594 66834
rect 11230 66782 11282 66834
rect 13470 66782 13522 66834
rect 13806 66782 13858 66834
rect 15150 66782 15202 66834
rect 17838 66782 17890 66834
rect 30606 66782 30658 66834
rect 4466 66614 4518 66666
rect 4570 66614 4622 66666
rect 4674 66614 4726 66666
rect 24466 66614 24518 66666
rect 24570 66614 24622 66666
rect 24674 66614 24726 66666
rect 3278 66446 3330 66498
rect 4286 66446 4338 66498
rect 6078 66446 6130 66498
rect 14702 66446 14754 66498
rect 15822 66446 15874 66498
rect 19182 66446 19234 66498
rect 1598 66334 1650 66386
rect 3614 66334 3666 66386
rect 10334 66334 10386 66386
rect 18174 66334 18226 66386
rect 30606 66334 30658 66386
rect 1262 66222 1314 66274
rect 3950 66222 4002 66274
rect 5406 66222 5458 66274
rect 5854 66222 5906 66274
rect 6638 66222 6690 66274
rect 7310 66222 7362 66274
rect 8094 66222 8146 66274
rect 9662 66222 9714 66274
rect 10110 66222 10162 66274
rect 11006 66222 11058 66274
rect 11342 66222 11394 66274
rect 12350 66222 12402 66274
rect 14254 66222 14306 66274
rect 18510 66222 18562 66274
rect 18958 66222 19010 66274
rect 19854 66222 19906 66274
rect 20190 66222 20242 66274
rect 21198 66222 21250 66274
rect 30270 66222 30322 66274
rect 5070 66110 5122 66162
rect 9326 66110 9378 66162
rect 2830 65998 2882 66050
rect 3806 65830 3858 65882
rect 3910 65830 3962 65882
rect 4014 65830 4066 65882
rect 23806 65830 23858 65882
rect 23910 65830 23962 65882
rect 24014 65830 24066 65882
rect 14590 65662 14642 65714
rect 19854 65662 19906 65714
rect 1934 65550 1986 65602
rect 5854 65550 5906 65602
rect 13022 65550 13074 65602
rect 15822 65550 15874 65602
rect 18286 65550 18338 65602
rect 1262 65438 1314 65490
rect 4398 65438 4450 65490
rect 9326 65438 9378 65490
rect 9886 65438 9938 65490
rect 10670 65438 10722 65490
rect 11006 65438 11058 65490
rect 11230 65438 11282 65490
rect 12126 65438 12178 65490
rect 17390 65438 17442 65490
rect 2382 65326 2434 65378
rect 8990 65326 9042 65378
rect 13358 65326 13410 65378
rect 16270 65326 16322 65378
rect 20974 65326 21026 65378
rect 1038 65214 1090 65266
rect 3502 65214 3554 65266
rect 4062 65214 4114 65266
rect 4958 65214 5010 65266
rect 5294 65214 5346 65266
rect 6302 65214 6354 65266
rect 7422 65214 7474 65266
rect 9998 65214 10050 65266
rect 18734 65214 18786 65266
rect 20638 65214 20690 65266
rect 4466 65046 4518 65098
rect 4570 65046 4622 65098
rect 4674 65046 4726 65098
rect 24466 65046 24518 65098
rect 24570 65046 24622 65098
rect 24674 65046 24726 65098
rect 3054 64878 3106 64930
rect 5966 64878 6018 64930
rect 13582 64878 13634 64930
rect 1710 64766 1762 64818
rect 5630 64766 5682 64818
rect 6974 64766 7026 64818
rect 8990 64766 9042 64818
rect 9998 64766 10050 64818
rect 19070 64766 19122 64818
rect 20078 64766 20130 64818
rect 30606 64766 30658 64818
rect 1374 64654 1426 64706
rect 2382 64654 2434 64706
rect 2830 64654 2882 64706
rect 3614 64654 3666 64706
rect 4286 64654 4338 64706
rect 5070 64654 5122 64706
rect 6526 64654 6578 64706
rect 8206 64654 8258 64706
rect 9326 64654 9378 64706
rect 9886 64654 9938 64706
rect 10446 64654 10498 64706
rect 11006 64654 11058 64706
rect 12126 64654 12178 64706
rect 13134 64654 13186 64706
rect 18846 64654 18898 64706
rect 19630 64654 19682 64706
rect 30270 64654 30322 64706
rect 2046 64542 2098 64594
rect 14702 64430 14754 64482
rect 21310 64430 21362 64482
rect 3806 64262 3858 64314
rect 3910 64262 3962 64314
rect 4014 64262 4066 64314
rect 23806 64262 23858 64314
rect 23910 64262 23962 64314
rect 24014 64262 24066 64314
rect 8206 64094 8258 64146
rect 8878 63982 8930 64034
rect 10782 63982 10834 64034
rect 14254 63982 14306 64034
rect 20974 63982 21026 64034
rect 1262 63870 1314 63922
rect 1822 63870 1874 63922
rect 3502 63870 3554 63922
rect 4174 63870 4226 63922
rect 5182 63870 5234 63922
rect 6526 63870 6578 63922
rect 18174 63870 18226 63922
rect 2382 63758 2434 63810
rect 4958 63758 5010 63810
rect 9326 63758 9378 63810
rect 14702 63758 14754 63810
rect 17390 63758 17442 63810
rect 18734 63758 18786 63810
rect 21310 63758 21362 63810
rect 29822 63758 29874 63810
rect 1038 63646 1090 63698
rect 3950 63646 4002 63698
rect 7086 63646 7138 63698
rect 10446 63646 10498 63698
rect 15822 63646 15874 63698
rect 17726 63646 17778 63698
rect 19854 63646 19906 63698
rect 22542 63646 22594 63698
rect 29486 63646 29538 63698
rect 30270 63646 30322 63698
rect 30606 63646 30658 63698
rect 4466 63478 4518 63530
rect 4570 63478 4622 63530
rect 4674 63478 4726 63530
rect 24466 63478 24518 63530
rect 24570 63478 24622 63530
rect 24674 63478 24726 63530
rect 1262 63310 1314 63362
rect 2942 63310 2994 63362
rect 6302 63310 6354 63362
rect 7982 63310 8034 63362
rect 8318 63310 8370 63362
rect 8878 63310 8930 63362
rect 9214 63310 9266 63362
rect 11902 63310 11954 63362
rect 15150 63310 15202 63362
rect 17502 63310 17554 63362
rect 20078 63310 20130 63362
rect 29822 63310 29874 63362
rect 3390 63198 3442 63250
rect 15934 63198 15986 63250
rect 19070 63198 19122 63250
rect 30606 63198 30658 63250
rect 1486 63086 1538 63138
rect 2382 63086 2434 63138
rect 2718 63086 2770 63138
rect 4174 63086 4226 63138
rect 4958 63086 5010 63138
rect 5742 63086 5794 63138
rect 11230 63086 11282 63138
rect 11678 63086 11730 63138
rect 12350 63086 12402 63138
rect 12910 63086 12962 63138
rect 13918 63086 13970 63138
rect 14926 63086 14978 63138
rect 15262 63086 15314 63138
rect 16942 63086 16994 63138
rect 19518 63086 19570 63138
rect 19966 63086 20018 63138
rect 20750 63086 20802 63138
rect 21086 63086 21138 63138
rect 22094 63086 22146 63138
rect 29486 63086 29538 63138
rect 30270 63086 30322 63138
rect 1934 62974 1986 63026
rect 10894 62974 10946 63026
rect 15710 62974 15762 63026
rect 7422 62862 7474 62914
rect 16046 62862 16098 62914
rect 18622 62862 18674 62914
rect 3806 62694 3858 62746
rect 3910 62694 3962 62746
rect 4014 62694 4066 62746
rect 23806 62694 23858 62746
rect 23910 62694 23962 62746
rect 24014 62694 24066 62746
rect 19630 62526 19682 62578
rect 5630 62414 5682 62466
rect 10894 62414 10946 62466
rect 14254 62414 14306 62466
rect 18062 62414 18114 62466
rect 1150 62302 1202 62354
rect 1486 62302 1538 62354
rect 2046 62302 2098 62354
rect 2830 62302 2882 62354
rect 3390 62302 3442 62354
rect 4286 62302 4338 62354
rect 5966 62302 6018 62354
rect 6414 62302 6466 62354
rect 7310 62302 7362 62354
rect 7646 62302 7698 62354
rect 8654 62302 8706 62354
rect 9550 62302 9602 62354
rect 14590 62302 14642 62354
rect 15038 62302 15090 62354
rect 15822 62302 15874 62354
rect 16270 62302 16322 62354
rect 17278 62302 17330 62354
rect 21086 62302 21138 62354
rect 21534 62302 21586 62354
rect 22318 62302 22370 62354
rect 22654 62302 22706 62354
rect 23774 62302 23826 62354
rect 2158 62190 2210 62242
rect 4958 62190 5010 62242
rect 5294 62190 5346 62242
rect 6638 62190 6690 62242
rect 18398 62190 18450 62242
rect 20638 62190 20690 62242
rect 21646 62190 21698 62242
rect 9214 62078 9266 62130
rect 15262 62078 15314 62130
rect 4466 61910 4518 61962
rect 4570 61910 4622 61962
rect 4674 61910 4726 61962
rect 24466 61910 24518 61962
rect 24570 61910 24622 61962
rect 24674 61910 24726 61962
rect 2158 61742 2210 61794
rect 6078 61742 6130 61794
rect 9998 61742 10050 61794
rect 15710 61742 15762 61794
rect 17614 61742 17666 61794
rect 19182 61742 19234 61794
rect 29822 61742 29874 61794
rect 1038 61630 1090 61682
rect 1374 61630 1426 61682
rect 1822 61630 1874 61682
rect 3502 61630 3554 61682
rect 5070 61630 5122 61682
rect 6526 61630 6578 61682
rect 11566 61630 11618 61682
rect 12574 61630 12626 61682
rect 15374 61630 15426 61682
rect 18174 61630 18226 61682
rect 30606 61630 30658 61682
rect 2942 61518 2994 61570
rect 4622 61518 4674 61570
rect 5406 61518 5458 61570
rect 5966 61518 6018 61570
rect 7310 61518 7362 61570
rect 8206 61518 8258 61570
rect 9438 61518 9490 61570
rect 11118 61518 11170 61570
rect 11902 61518 11954 61570
rect 12462 61518 12514 61570
rect 13022 61518 13074 61570
rect 13582 61518 13634 61570
rect 14590 61518 14642 61570
rect 15598 61518 15650 61570
rect 16046 61518 16098 61570
rect 16830 61518 16882 61570
rect 17054 61518 17106 61570
rect 18622 61518 18674 61570
rect 18958 61518 19010 61570
rect 19742 61518 19794 61570
rect 20414 61518 20466 61570
rect 21198 61518 21250 61570
rect 29598 61518 29650 61570
rect 30270 61518 30322 61570
rect 17726 61406 17778 61458
rect 15934 61294 15986 61346
rect 16718 61294 16770 61346
rect 17166 61294 17218 61346
rect 3806 61126 3858 61178
rect 3910 61126 3962 61178
rect 4014 61126 4066 61178
rect 23806 61126 23858 61178
rect 23910 61126 23962 61178
rect 24014 61126 24066 61178
rect 4286 60958 4338 61010
rect 12126 60958 12178 61010
rect 14814 60958 14866 61010
rect 5630 60846 5682 60898
rect 10558 60846 10610 60898
rect 20638 60846 20690 60898
rect 2606 60734 2658 60786
rect 5966 60734 6018 60786
rect 6414 60734 6466 60786
rect 7310 60734 7362 60786
rect 7646 60734 7698 60786
rect 8654 60734 8706 60786
rect 13134 60734 13186 60786
rect 15374 60734 15426 60786
rect 17614 60734 17666 60786
rect 19294 60734 19346 60786
rect 20974 60734 21026 60786
rect 21422 60734 21474 60786
rect 22654 60734 22706 60786
rect 23662 60734 23714 60786
rect 2158 60622 2210 60674
rect 6638 60622 6690 60674
rect 11006 60622 11058 60674
rect 13694 60622 13746 60674
rect 15934 60622 15986 60674
rect 18174 60622 18226 60674
rect 21646 60622 21698 60674
rect 22094 60622 22146 60674
rect 29822 60622 29874 60674
rect 1038 60510 1090 60562
rect 1374 60510 1426 60562
rect 1822 60510 1874 60562
rect 3166 60510 3218 60562
rect 17054 60510 17106 60562
rect 29486 60510 29538 60562
rect 30270 60510 30322 60562
rect 30606 60510 30658 60562
rect 4466 60342 4518 60394
rect 4570 60342 4622 60394
rect 4674 60342 4726 60394
rect 24466 60342 24518 60394
rect 24570 60342 24622 60394
rect 24674 60342 24726 60394
rect 1150 60174 1202 60226
rect 4062 60174 4114 60226
rect 5182 60174 5234 60226
rect 7422 60174 7474 60226
rect 11118 60174 11170 60226
rect 11902 60174 11954 60226
rect 14814 60174 14866 60226
rect 15934 60174 15986 60226
rect 20638 60174 20690 60226
rect 29822 60174 29874 60226
rect 2382 60062 2434 60114
rect 6302 60062 6354 60114
rect 9886 60062 9938 60114
rect 11566 60062 11618 60114
rect 16942 60062 16994 60114
rect 17950 60062 18002 60114
rect 21870 60062 21922 60114
rect 9550 59950 9602 60002
rect 14254 59950 14306 60002
rect 16606 59950 16658 60002
rect 17278 59950 17330 60002
rect 17838 59950 17890 60002
rect 18510 59950 18562 60002
rect 18958 59950 19010 60002
rect 20078 59950 20130 60002
rect 29486 59950 29538 60002
rect 2718 59838 2770 59890
rect 3614 59838 3666 59890
rect 5854 59838 5906 59890
rect 22206 59838 22258 59890
rect 3806 59558 3858 59610
rect 3910 59558 3962 59610
rect 4014 59558 4066 59610
rect 23806 59558 23858 59610
rect 23910 59558 23962 59610
rect 24014 59558 24066 59610
rect 18510 59390 18562 59442
rect 18958 59278 19010 59330
rect 2158 59166 2210 59218
rect 8318 59166 8370 59218
rect 14702 59166 14754 59218
rect 16830 59166 16882 59218
rect 2494 59054 2546 59106
rect 2830 59054 2882 59106
rect 8766 59054 8818 59106
rect 15038 59054 15090 59106
rect 17390 59054 17442 59106
rect 1038 58942 1090 58994
rect 1374 58942 1426 58994
rect 1822 58942 1874 58994
rect 9886 58942 9938 58994
rect 16270 58942 16322 58994
rect 30270 58942 30322 58994
rect 30606 58942 30658 58994
rect 4466 58774 4518 58826
rect 4570 58774 4622 58826
rect 4674 58774 4726 58826
rect 24466 58774 24518 58826
rect 24570 58774 24622 58826
rect 24674 58774 24726 58826
rect 1374 58606 1426 58658
rect 16718 58606 16770 58658
rect 17054 58606 17106 58658
rect 20638 58606 20690 58658
rect 29822 58606 29874 58658
rect 1038 58494 1090 58546
rect 1710 58494 1762 58546
rect 9998 58494 10050 58546
rect 14030 58494 14082 58546
rect 19406 58494 19458 58546
rect 30606 58494 30658 58546
rect 2046 58382 2098 58434
rect 9662 58382 9714 58434
rect 13694 58382 13746 58434
rect 19070 58382 19122 58434
rect 29486 58382 29538 58434
rect 30270 58382 30322 58434
rect 11230 58158 11282 58210
rect 15262 58158 15314 58210
rect 3806 57990 3858 58042
rect 3910 57990 3962 58042
rect 4014 57990 4066 58042
rect 23806 57990 23858 58042
rect 23910 57990 23962 58042
rect 24014 57990 24066 58042
rect 8094 57710 8146 57762
rect 10334 57710 10386 57762
rect 14590 57710 14642 57762
rect 18958 57710 19010 57762
rect 1374 57598 1426 57650
rect 15038 57598 15090 57650
rect 15374 57598 15426 57650
rect 16270 57598 16322 57650
rect 16718 57598 16770 57650
rect 17726 57598 17778 57650
rect 1038 57486 1090 57538
rect 8542 57486 8594 57538
rect 10782 57486 10834 57538
rect 13582 57486 13634 57538
rect 13918 57486 13970 57538
rect 29822 57486 29874 57538
rect 9662 57374 9714 57426
rect 11902 57374 11954 57426
rect 13246 57374 13298 57426
rect 14254 57374 14306 57426
rect 15598 57374 15650 57426
rect 29486 57374 29538 57426
rect 4466 57206 4518 57258
rect 4570 57206 4622 57258
rect 4674 57206 4726 57258
rect 24466 57206 24518 57258
rect 24570 57206 24622 57258
rect 24674 57206 24726 57258
rect 18958 57038 19010 57090
rect 4846 56926 4898 56978
rect 7086 56926 7138 56978
rect 10110 56926 10162 56978
rect 11118 56926 11170 56978
rect 30606 56926 30658 56978
rect 6638 56814 6690 56866
rect 10446 56814 10498 56866
rect 11006 56814 11058 56866
rect 11678 56814 11730 56866
rect 12350 56814 12402 56866
rect 13134 56814 13186 56866
rect 30382 56814 30434 56866
rect 4398 56702 4450 56754
rect 5966 56590 6018 56642
rect 8206 56590 8258 56642
rect 3806 56422 3858 56474
rect 3910 56422 3962 56474
rect 4014 56422 4066 56474
rect 23806 56422 23858 56474
rect 23910 56422 23962 56474
rect 24014 56422 24066 56474
rect 5854 56142 5906 56194
rect 8990 56142 9042 56194
rect 14478 56142 14530 56194
rect 18958 56142 19010 56194
rect 9438 56030 9490 56082
rect 9886 56030 9938 56082
rect 10670 56030 10722 56082
rect 11230 56030 11282 56082
rect 12126 56030 12178 56082
rect 14030 55918 14082 55970
rect 21310 55918 21362 55970
rect 6302 55806 6354 55858
rect 7422 55806 7474 55858
rect 9998 55806 10050 55858
rect 12910 55806 12962 55858
rect 20974 55806 21026 55858
rect 30270 55806 30322 55858
rect 30606 55806 30658 55858
rect 4466 55638 4518 55690
rect 4570 55638 4622 55690
rect 4674 55638 4726 55690
rect 24466 55638 24518 55690
rect 24570 55638 24622 55690
rect 24674 55638 24726 55690
rect 18958 55470 19010 55522
rect 30494 55470 30546 55522
rect 3502 55358 3554 55410
rect 5070 55358 5122 55410
rect 6078 55358 6130 55410
rect 9774 55358 9826 55410
rect 14142 55358 14194 55410
rect 2942 55246 2994 55298
rect 4622 55246 4674 55298
rect 5406 55246 5458 55298
rect 5854 55246 5906 55298
rect 6526 55246 6578 55298
rect 7310 55246 7362 55298
rect 8094 55246 8146 55298
rect 9326 55246 9378 55298
rect 28366 55246 28418 55298
rect 30158 55246 30210 55298
rect 13694 55134 13746 55186
rect 24782 55134 24834 55186
rect 11006 55022 11058 55074
rect 15262 55022 15314 55074
rect 3806 54854 3858 54906
rect 3910 54854 3962 54906
rect 4014 54854 4066 54906
rect 23806 54854 23858 54906
rect 23910 54854 23962 54906
rect 24014 54854 24066 54906
rect 3726 54686 3778 54738
rect 2158 54574 2210 54626
rect 5742 54574 5794 54626
rect 14142 54574 14194 54626
rect 6078 54462 6130 54514
rect 6526 54462 6578 54514
rect 7422 54462 7474 54514
rect 7758 54462 7810 54514
rect 8766 54462 8818 54514
rect 10446 54462 10498 54514
rect 14590 54462 14642 54514
rect 14926 54462 14978 54514
rect 15822 54462 15874 54514
rect 16158 54462 16210 54514
rect 17166 54462 17218 54514
rect 2494 54350 2546 54402
rect 10894 54350 10946 54402
rect 30606 54350 30658 54402
rect 6750 54238 6802 54290
rect 12126 54238 12178 54290
rect 15150 54238 15202 54290
rect 30270 54238 30322 54290
rect 4466 54070 4518 54122
rect 4570 54070 4622 54122
rect 4674 54070 4726 54122
rect 24466 54070 24518 54122
rect 24570 54070 24622 54122
rect 24674 54070 24726 54122
rect 3502 53790 3554 53842
rect 10558 53790 10610 53842
rect 15598 53790 15650 53842
rect 21758 53790 21810 53842
rect 30606 53790 30658 53842
rect 2942 53678 2994 53730
rect 6750 53678 6802 53730
rect 9550 53678 9602 53730
rect 9886 53678 9938 53730
rect 10334 53678 10386 53730
rect 11118 53678 11170 53730
rect 11678 53678 11730 53730
rect 12574 53678 12626 53730
rect 15262 53678 15314 53730
rect 21422 53678 21474 53730
rect 30382 53678 30434 53730
rect 14030 53566 14082 53618
rect 4622 53454 4674 53506
rect 3806 53286 3858 53338
rect 3910 53286 3962 53338
rect 4014 53286 4066 53338
rect 23806 53286 23858 53338
rect 23910 53286 23962 53338
rect 24014 53286 24066 53338
rect 10894 53118 10946 53170
rect 16046 53118 16098 53170
rect 2606 52894 2658 52946
rect 6974 52894 7026 52946
rect 8094 52894 8146 52946
rect 8430 52894 8482 52946
rect 9214 52894 9266 52946
rect 9662 52894 9714 52946
rect 11230 52894 11282 52946
rect 12014 52894 12066 52946
rect 14478 52894 14530 52946
rect 16494 52894 16546 52946
rect 3054 52782 3106 52834
rect 10110 52782 10162 52834
rect 11790 52782 11842 52834
rect 14926 52782 14978 52834
rect 4286 52670 4338 52722
rect 9102 52670 9154 52722
rect 16830 52670 16882 52722
rect 30270 52670 30322 52722
rect 30606 52670 30658 52722
rect 4466 52502 4518 52554
rect 4570 52502 4622 52554
rect 4674 52502 4726 52554
rect 24466 52502 24518 52554
rect 24570 52502 24622 52554
rect 24674 52502 24726 52554
rect 4510 52334 4562 52386
rect 11118 52334 11170 52386
rect 14926 52334 14978 52386
rect 3278 52222 3330 52274
rect 10110 52222 10162 52274
rect 17054 52222 17106 52274
rect 6862 52110 6914 52162
rect 10446 52110 10498 52162
rect 10894 52110 10946 52162
rect 11566 52110 11618 52162
rect 12126 52110 12178 52162
rect 13134 52110 13186 52162
rect 16830 52110 16882 52162
rect 2942 51998 2994 52050
rect 15374 51998 15426 52050
rect 13806 51886 13858 51938
rect 3806 51718 3858 51770
rect 3910 51718 3962 51770
rect 4014 51718 4066 51770
rect 23806 51718 23858 51770
rect 23910 51718 23962 51770
rect 24014 51718 24066 51770
rect 4958 51438 5010 51490
rect 2718 51326 2770 51378
rect 5294 51326 5346 51378
rect 5854 51326 5906 51378
rect 6414 51326 6466 51378
rect 7086 51326 7138 51378
rect 7982 51326 8034 51378
rect 9326 51326 9378 51378
rect 9886 51326 9938 51378
rect 10670 51326 10722 51378
rect 11230 51326 11282 51378
rect 12014 51326 12066 51378
rect 13134 51326 13186 51378
rect 13694 51326 13746 51378
rect 14254 51326 14306 51378
rect 14814 51326 14866 51378
rect 15822 51326 15874 51378
rect 3054 51214 3106 51266
rect 8990 51214 9042 51266
rect 9998 51214 10050 51266
rect 12798 51214 12850 51266
rect 4286 51102 4338 51154
rect 5966 51102 6018 51154
rect 13806 51102 13858 51154
rect 16942 51102 16994 51154
rect 17278 51102 17330 51154
rect 30270 51102 30322 51154
rect 30606 51102 30658 51154
rect 4466 50934 4518 50986
rect 4570 50934 4622 50986
rect 4674 50934 4726 50986
rect 24466 50934 24518 50986
rect 24570 50934 24622 50986
rect 24674 50934 24726 50986
rect 1150 50766 1202 50818
rect 2494 50766 2546 50818
rect 5070 50766 5122 50818
rect 10782 50766 10834 50818
rect 17950 50766 18002 50818
rect 1486 50654 1538 50706
rect 3614 50654 3666 50706
rect 5518 50654 5570 50706
rect 12798 50654 12850 50706
rect 30606 50654 30658 50706
rect 2046 50542 2098 50594
rect 4398 50542 4450 50594
rect 4958 50542 5010 50594
rect 6078 50542 6130 50594
rect 7086 50542 7138 50594
rect 11230 50542 11282 50594
rect 12126 50542 12178 50594
rect 12574 50542 12626 50594
rect 13246 50542 13298 50594
rect 13806 50542 13858 50594
rect 14030 50542 14082 50594
rect 14814 50542 14866 50594
rect 30382 50542 30434 50594
rect 4062 50430 4114 50482
rect 11790 50430 11842 50482
rect 15262 50430 15314 50482
rect 18398 50430 18450 50482
rect 9662 50318 9714 50370
rect 16830 50318 16882 50370
rect 3806 50150 3858 50202
rect 3910 50150 3962 50202
rect 4014 50150 4066 50202
rect 23806 50150 23858 50202
rect 23910 50150 23962 50202
rect 24014 50150 24066 50202
rect 8542 49982 8594 50034
rect 12126 49982 12178 50034
rect 13246 49982 13298 50034
rect 1486 49758 1538 49810
rect 6974 49758 7026 49810
rect 9886 49758 9938 49810
rect 10558 49758 10610 49810
rect 14814 49758 14866 49810
rect 15822 49758 15874 49810
rect 16158 49758 16210 49810
rect 16830 49758 16882 49810
rect 17390 49758 17442 49810
rect 18398 49758 18450 49810
rect 1934 49646 1986 49698
rect 11006 49646 11058 49698
rect 14478 49646 14530 49698
rect 15374 49646 15426 49698
rect 3166 49534 3218 49586
rect 7422 49534 7474 49586
rect 9998 49534 10050 49586
rect 16382 49534 16434 49586
rect 4466 49366 4518 49418
rect 4570 49366 4622 49418
rect 4674 49366 4726 49418
rect 24466 49366 24518 49418
rect 24570 49366 24622 49418
rect 24674 49366 24726 49418
rect 2270 49198 2322 49250
rect 8206 49198 8258 49250
rect 10446 49198 10498 49250
rect 11566 49198 11618 49250
rect 12686 49198 12738 49250
rect 1374 49086 1426 49138
rect 1598 49086 1650 49138
rect 3726 49086 3778 49138
rect 7086 49086 7138 49138
rect 19742 49086 19794 49138
rect 30606 49086 30658 49138
rect 1934 48974 1986 49026
rect 3054 48974 3106 49026
rect 3614 48974 3666 49026
rect 4174 48974 4226 49026
rect 4846 48974 4898 49026
rect 5854 48974 5906 49026
rect 6638 48974 6690 49026
rect 12126 48974 12178 49026
rect 19406 48974 19458 49026
rect 30270 48974 30322 49026
rect 2718 48862 2770 48914
rect 9998 48862 10050 48914
rect 15262 48862 15314 48914
rect 13806 48750 13858 48802
rect 3806 48582 3858 48634
rect 3910 48582 3962 48634
rect 4014 48582 4066 48634
rect 23806 48582 23858 48634
rect 23910 48582 23962 48634
rect 24014 48582 24066 48634
rect 2158 48414 2210 48466
rect 15934 48414 15986 48466
rect 12238 48302 12290 48354
rect 16606 48302 16658 48354
rect 3726 48190 3778 48242
rect 6638 48190 6690 48242
rect 10782 48190 10834 48242
rect 11902 48190 11954 48242
rect 13358 48190 13410 48242
rect 13470 48190 13522 48242
rect 13582 48190 13634 48242
rect 14366 48190 14418 48242
rect 3390 48078 3442 48130
rect 7086 48078 7138 48130
rect 11342 48078 11394 48130
rect 11454 48078 11506 48130
rect 11678 48078 11730 48130
rect 13022 48078 13074 48130
rect 13246 48078 13298 48130
rect 16942 48078 16994 48130
rect 18958 48078 19010 48130
rect 8318 47966 8370 48018
rect 9102 47966 9154 48018
rect 10222 47966 10274 48018
rect 12126 47966 12178 48018
rect 13806 47966 13858 48018
rect 14814 47966 14866 48018
rect 18174 47966 18226 48018
rect 18622 47966 18674 48018
rect 30270 47966 30322 48018
rect 30606 47966 30658 48018
rect 4466 47798 4518 47850
rect 4570 47798 4622 47850
rect 4674 47798 4726 47850
rect 24466 47798 24518 47850
rect 24570 47798 24622 47850
rect 24674 47798 24726 47850
rect 3278 47630 3330 47682
rect 10222 47630 10274 47682
rect 14814 47630 14866 47682
rect 1934 47518 1986 47570
rect 3726 47518 3778 47570
rect 6526 47518 6578 47570
rect 9214 47518 9266 47570
rect 10670 47518 10722 47570
rect 13470 47518 13522 47570
rect 17726 47518 17778 47570
rect 18174 47518 18226 47570
rect 30606 47518 30658 47570
rect 1710 47406 1762 47458
rect 2718 47406 2770 47458
rect 3054 47406 3106 47458
rect 4286 47406 4338 47458
rect 5406 47406 5458 47458
rect 9550 47406 9602 47458
rect 9998 47406 10050 47458
rect 11230 47406 11282 47458
rect 12238 47406 12290 47458
rect 13022 47406 13074 47458
rect 15934 47406 15986 47458
rect 17054 47406 17106 47458
rect 17502 47406 17554 47458
rect 18734 47406 18786 47458
rect 19742 47406 19794 47458
rect 30270 47406 30322 47458
rect 2270 47294 2322 47346
rect 6078 47294 6130 47346
rect 8206 47294 8258 47346
rect 14366 47294 14418 47346
rect 16718 47294 16770 47346
rect 7646 47182 7698 47234
rect 8094 47182 8146 47234
rect 13134 47182 13186 47234
rect 13358 47182 13410 47234
rect 3806 47014 3858 47066
rect 3910 47014 3962 47066
rect 4014 47014 4066 47066
rect 23806 47014 23858 47066
rect 23910 47014 23962 47066
rect 24014 47014 24066 47066
rect 3166 46846 3218 46898
rect 12910 46846 12962 46898
rect 1486 46622 1538 46674
rect 5182 46622 5234 46674
rect 5854 46622 5906 46674
rect 7198 46622 7250 46674
rect 7534 46622 7586 46674
rect 8318 46622 8370 46674
rect 8990 46622 9042 46674
rect 9886 46622 9938 46674
rect 12014 46622 12066 46674
rect 14478 46622 14530 46674
rect 1934 46510 1986 46562
rect 5070 46510 5122 46562
rect 6750 46510 6802 46562
rect 7758 46510 7810 46562
rect 16382 46510 16434 46562
rect 23550 46510 23602 46562
rect 6190 46398 6242 46450
rect 10446 46398 10498 46450
rect 11566 46398 11618 46450
rect 14030 46398 14082 46450
rect 16046 46398 16098 46450
rect 16606 46398 16658 46450
rect 23214 46398 23266 46450
rect 4466 46230 4518 46282
rect 4570 46230 4622 46282
rect 4674 46230 4726 46282
rect 24466 46230 24518 46282
rect 24570 46230 24622 46282
rect 24674 46230 24726 46282
rect 9662 46062 9714 46114
rect 17838 46062 17890 46114
rect 22654 46062 22706 46114
rect 1598 45950 1650 46002
rect 4846 45950 4898 46002
rect 7086 45950 7138 46002
rect 11342 45950 11394 46002
rect 18846 45950 18898 46002
rect 20078 45950 20130 46002
rect 30606 45950 30658 46002
rect 6526 45838 6578 45890
rect 8206 45838 8258 45890
rect 8878 45838 8930 45890
rect 9102 45838 9154 45890
rect 9662 45838 9714 45890
rect 10670 45838 10722 45890
rect 11118 45838 11170 45890
rect 12014 45838 12066 45890
rect 12350 45838 12402 45890
rect 13358 45838 13410 45890
rect 18958 45838 19010 45890
rect 22318 45838 22370 45890
rect 30270 45838 30322 45890
rect 1262 45726 1314 45778
rect 4398 45726 4450 45778
rect 6638 45726 6690 45778
rect 10334 45726 10386 45778
rect 19742 45726 19794 45778
rect 2830 45614 2882 45666
rect 5966 45614 6018 45666
rect 9438 45614 9490 45666
rect 18174 45614 18226 45666
rect 21310 45614 21362 45666
rect 3806 45446 3858 45498
rect 3910 45446 3962 45498
rect 4014 45446 4066 45498
rect 23806 45446 23858 45498
rect 23910 45446 23962 45498
rect 24014 45446 24066 45498
rect 12126 45278 12178 45330
rect 18958 45278 19010 45330
rect 9774 45166 9826 45218
rect 13470 45166 13522 45218
rect 1262 45054 1314 45106
rect 5854 45054 5906 45106
rect 6526 45054 6578 45106
rect 6862 45054 6914 45106
rect 7534 45054 7586 45106
rect 8206 45054 8258 45106
rect 9214 45054 9266 45106
rect 10446 45054 10498 45106
rect 17390 45054 17442 45106
rect 5518 44942 5570 44994
rect 6078 44942 6130 44994
rect 7086 44942 7138 44994
rect 9662 44942 9714 44994
rect 13806 44942 13858 44994
rect 17838 44942 17890 44994
rect 29822 44942 29874 44994
rect 1710 44830 1762 44882
rect 2830 44830 2882 44882
rect 5630 44830 5682 44882
rect 9886 44830 9938 44882
rect 11006 44830 11058 44882
rect 15038 44830 15090 44882
rect 29486 44830 29538 44882
rect 30270 44830 30322 44882
rect 30606 44830 30658 44882
rect 4466 44662 4518 44714
rect 4570 44662 4622 44714
rect 4674 44662 4726 44714
rect 24466 44662 24518 44714
rect 24570 44662 24622 44714
rect 24674 44662 24726 44714
rect 2942 44494 2994 44546
rect 8206 44494 8258 44546
rect 10894 44494 10946 44546
rect 14814 44494 14866 44546
rect 19854 44494 19906 44546
rect 22654 44494 22706 44546
rect 29822 44494 29874 44546
rect 3390 44382 3442 44434
rect 7086 44382 7138 44434
rect 9438 44382 9490 44434
rect 9886 44382 9938 44434
rect 17278 44382 17330 44434
rect 2382 44270 2434 44322
rect 2830 44270 2882 44322
rect 4174 44270 4226 44322
rect 4958 44270 5010 44322
rect 6638 44270 6690 44322
rect 8990 44270 9042 44322
rect 9102 44270 9154 44322
rect 10222 44270 10274 44322
rect 10782 44270 10834 44322
rect 11566 44270 11618 44322
rect 11902 44270 11954 44322
rect 13022 44270 13074 44322
rect 14366 44270 14418 44322
rect 16830 44270 16882 44322
rect 19294 44270 19346 44322
rect 29598 44270 29650 44322
rect 1934 44158 1986 44210
rect 19406 44158 19458 44210
rect 23102 44158 23154 44210
rect 9326 44046 9378 44098
rect 15934 44046 15986 44098
rect 18510 44046 18562 44098
rect 20974 44046 21026 44098
rect 21534 44046 21586 44098
rect 3806 43878 3858 43930
rect 3910 43878 3962 43930
rect 4014 43878 4066 43930
rect 23806 43878 23858 43930
rect 23910 43878 23962 43930
rect 24014 43878 24066 43930
rect 11566 43710 11618 43762
rect 5294 43598 5346 43650
rect 6862 43598 6914 43650
rect 9326 43598 9378 43650
rect 1598 43486 1650 43538
rect 2046 43486 2098 43538
rect 2606 43486 2658 43538
rect 3166 43486 3218 43538
rect 4174 43486 4226 43538
rect 7758 43486 7810 43538
rect 9998 43486 10050 43538
rect 14478 43486 14530 43538
rect 14814 43486 14866 43538
rect 15710 43486 15762 43538
rect 16046 43486 16098 43538
rect 17166 43486 17218 43538
rect 17726 43486 17778 43538
rect 20974 43486 21026 43538
rect 21422 43486 21474 43538
rect 22094 43486 22146 43538
rect 22654 43486 22706 43538
rect 23662 43486 23714 43538
rect 1150 43374 1202 43426
rect 2158 43374 2210 43426
rect 8206 43374 8258 43426
rect 10334 43374 10386 43426
rect 14030 43374 14082 43426
rect 18286 43374 18338 43426
rect 20638 43374 20690 43426
rect 21646 43374 21698 43426
rect 5742 43262 5794 43314
rect 15038 43262 15090 43314
rect 19406 43262 19458 43314
rect 29486 43262 29538 43314
rect 29822 43262 29874 43314
rect 30270 43262 30322 43314
rect 30606 43262 30658 43314
rect 4466 43094 4518 43146
rect 4570 43094 4622 43146
rect 4674 43094 4726 43146
rect 24466 43094 24518 43146
rect 24570 43094 24622 43146
rect 24674 43094 24726 43146
rect 6190 42926 6242 42978
rect 15150 42926 15202 42978
rect 18846 42926 18898 42978
rect 2942 42814 2994 42866
rect 9326 42814 9378 42866
rect 10334 42814 10386 42866
rect 22766 42814 22818 42866
rect 30606 42814 30658 42866
rect 2382 42702 2434 42754
rect 2830 42702 2882 42754
rect 3390 42702 3442 42754
rect 4062 42702 4114 42754
rect 4958 42702 5010 42754
rect 5742 42702 5794 42754
rect 9662 42702 9714 42754
rect 10110 42702 10162 42754
rect 10782 42702 10834 42754
rect 11454 42702 11506 42754
rect 12350 42702 12402 42754
rect 13134 42702 13186 42754
rect 13918 42702 13970 42754
rect 14478 42702 14530 42754
rect 15262 42702 15314 42754
rect 15710 42702 15762 42754
rect 18286 42702 18338 42754
rect 18622 42702 18674 42754
rect 19406 42702 19458 42754
rect 19854 42702 19906 42754
rect 20862 42702 20914 42754
rect 23214 42702 23266 42754
rect 30270 42702 30322 42754
rect 1934 42590 1986 42642
rect 16158 42590 16210 42642
rect 17838 42590 17890 42642
rect 7310 42478 7362 42530
rect 21534 42478 21586 42530
rect 3806 42310 3858 42362
rect 3910 42310 3962 42362
rect 4014 42310 4066 42362
rect 23806 42310 23858 42362
rect 23910 42310 23962 42362
rect 24014 42310 24066 42362
rect 10334 42142 10386 42194
rect 13806 42142 13858 42194
rect 8990 42030 9042 42082
rect 11902 42030 11954 42082
rect 15374 42030 15426 42082
rect 16494 42030 16546 42082
rect 1598 41918 1650 41970
rect 1934 41918 1986 41970
rect 2718 41918 2770 41970
rect 3166 41918 3218 41970
rect 4174 41918 4226 41970
rect 4958 41918 5010 41970
rect 5294 41918 5346 41970
rect 5742 41918 5794 41970
rect 6526 41918 6578 41970
rect 7198 41918 7250 41970
rect 7982 41918 8034 41970
rect 8654 41918 8706 41970
rect 19630 41918 19682 41970
rect 20638 41918 20690 41970
rect 20974 41918 21026 41970
rect 21422 41918 21474 41970
rect 22654 41918 22706 41970
rect 23662 41918 23714 41970
rect 1150 41806 1202 41858
rect 9214 41806 9266 41858
rect 9550 41806 9602 41858
rect 11454 41806 11506 41858
rect 15038 41806 15090 41858
rect 16942 41806 16994 41858
rect 18958 41806 19010 41858
rect 19294 41806 19346 41858
rect 21646 41806 21698 41858
rect 22094 41806 22146 41858
rect 29822 41806 29874 41858
rect 2158 41694 2210 41746
rect 5966 41694 6018 41746
rect 18062 41694 18114 41746
rect 19966 41694 20018 41746
rect 29486 41694 29538 41746
rect 4466 41526 4518 41578
rect 4570 41526 4622 41578
rect 4674 41526 4726 41578
rect 24466 41526 24518 41578
rect 24570 41526 24622 41578
rect 24674 41526 24726 41578
rect 3278 41358 3330 41410
rect 4398 41358 4450 41410
rect 5854 41358 5906 41410
rect 11006 41358 11058 41410
rect 19070 41358 19122 41410
rect 21758 41358 21810 41410
rect 22878 41358 22930 41410
rect 14814 41246 14866 41298
rect 19518 41246 19570 41298
rect 29822 41246 29874 41298
rect 30270 41246 30322 41298
rect 30606 41246 30658 41298
rect 4846 41134 4898 41186
rect 5294 41134 5346 41186
rect 5630 41134 5682 41186
rect 6526 41134 6578 41186
rect 7086 41134 7138 41186
rect 7870 41134 7922 41186
rect 10334 41134 10386 41186
rect 10782 41134 10834 41186
rect 11454 41134 11506 41186
rect 12014 41134 12066 41186
rect 12238 41134 12290 41186
rect 13022 41134 13074 41186
rect 14478 41134 14530 41186
rect 18510 41134 18562 41186
rect 18846 41134 18898 41186
rect 20190 41134 20242 41186
rect 21086 41134 21138 41186
rect 23326 41134 23378 41186
rect 29486 41134 29538 41186
rect 2830 41022 2882 41074
rect 9998 41022 10050 41074
rect 18062 41022 18114 41074
rect 16046 40910 16098 40962
rect 3806 40742 3858 40794
rect 3910 40742 3962 40794
rect 4014 40742 4066 40794
rect 23806 40742 23858 40794
rect 23910 40742 23962 40794
rect 24014 40742 24066 40794
rect 5854 40574 5906 40626
rect 8430 40574 8482 40626
rect 8990 40574 9042 40626
rect 14590 40574 14642 40626
rect 1710 40462 1762 40514
rect 6862 40462 6914 40514
rect 10558 40462 10610 40514
rect 13022 40462 13074 40514
rect 20638 40462 20690 40514
rect 3278 40350 3330 40402
rect 5182 40350 5234 40402
rect 16494 40350 16546 40402
rect 16942 40350 16994 40402
rect 17838 40350 17890 40402
rect 18174 40350 18226 40402
rect 19182 40350 19234 40402
rect 20974 40350 21026 40402
rect 21534 40350 21586 40402
rect 22206 40350 22258 40402
rect 22766 40350 22818 40402
rect 23662 40350 23714 40402
rect 30270 40350 30322 40402
rect 2046 40238 2098 40290
rect 5070 40238 5122 40290
rect 10110 40238 10162 40290
rect 13470 40238 13522 40290
rect 16158 40238 16210 40290
rect 17166 40238 17218 40290
rect 21646 40238 21698 40290
rect 29822 40238 29874 40290
rect 6190 40126 6242 40178
rect 7310 40126 7362 40178
rect 29486 40126 29538 40178
rect 30606 40126 30658 40178
rect 4466 39958 4518 40010
rect 4570 39958 4622 40010
rect 4674 39958 4726 40010
rect 24466 39958 24518 40010
rect 24570 39958 24622 40010
rect 24674 39958 24726 40010
rect 2830 39790 2882 39842
rect 6526 39790 6578 39842
rect 1598 39678 1650 39730
rect 5406 39678 5458 39730
rect 7086 39678 7138 39730
rect 7646 39678 7698 39730
rect 10894 39678 10946 39730
rect 11902 39678 11954 39730
rect 4958 39566 5010 39618
rect 11230 39566 11282 39618
rect 11678 39566 11730 39618
rect 12350 39566 12402 39618
rect 12910 39566 12962 39618
rect 13918 39566 13970 39618
rect 1262 39454 1314 39506
rect 7870 39342 7922 39394
rect 8206 39342 8258 39394
rect 3806 39174 3858 39226
rect 3910 39174 3962 39226
rect 4014 39174 4066 39226
rect 23806 39174 23858 39226
rect 23910 39174 23962 39226
rect 24014 39174 24066 39226
rect 2830 39006 2882 39058
rect 9886 39006 9938 39058
rect 12126 39006 12178 39058
rect 1262 38894 1314 38946
rect 8318 38894 8370 38946
rect 10558 38894 10610 38946
rect 5518 38782 5570 38834
rect 14030 38782 14082 38834
rect 14478 38782 14530 38834
rect 15374 38782 15426 38834
rect 15710 38782 15762 38834
rect 16718 38782 16770 38834
rect 20862 38782 20914 38834
rect 1598 38670 1650 38722
rect 6078 38670 6130 38722
rect 8766 38670 8818 38722
rect 10894 38670 10946 38722
rect 13694 38670 13746 38722
rect 14702 38670 14754 38722
rect 21422 38670 21474 38722
rect 7198 38558 7250 38610
rect 22542 38558 22594 38610
rect 4466 38390 4518 38442
rect 4570 38390 4622 38442
rect 4674 38390 4726 38442
rect 24466 38390 24518 38442
rect 24570 38390 24622 38442
rect 24674 38390 24726 38442
rect 6078 38222 6130 38274
rect 9886 38222 9938 38274
rect 11006 38222 11058 38274
rect 12126 38222 12178 38274
rect 13246 38222 13298 38274
rect 15486 38222 15538 38274
rect 18622 38222 18674 38274
rect 1934 38110 1986 38162
rect 14254 38110 14306 38162
rect 20078 38110 20130 38162
rect 21310 38110 21362 38162
rect 1374 37998 1426 38050
rect 18734 37998 18786 38050
rect 19518 37998 19570 38050
rect 19854 37998 19906 38050
rect 1486 37886 1538 37938
rect 5630 37886 5682 37938
rect 9438 37886 9490 37938
rect 11678 37886 11730 37938
rect 13918 37886 13970 37938
rect 19182 37886 19234 37938
rect 20078 37886 20130 37938
rect 20862 37886 20914 37938
rect 3054 37774 3106 37826
rect 7198 37774 7250 37826
rect 18622 37774 18674 37826
rect 19070 37774 19122 37826
rect 22430 37774 22482 37826
rect 3806 37606 3858 37658
rect 3910 37606 3962 37658
rect 4014 37606 4066 37658
rect 23806 37606 23858 37658
rect 23910 37606 23962 37658
rect 24014 37606 24066 37658
rect 2718 37326 2770 37378
rect 1934 37214 1986 37266
rect 6862 37214 6914 37266
rect 7198 37214 7250 37266
rect 8654 37214 8706 37266
rect 9438 37214 9490 37266
rect 10110 37214 10162 37266
rect 14702 37214 14754 37266
rect 15038 37214 15090 37266
rect 15934 37214 15986 37266
rect 16270 37214 16322 37266
rect 17278 37214 17330 37266
rect 18062 37214 18114 37266
rect 20862 37214 20914 37266
rect 6414 37102 6466 37154
rect 7422 37102 7474 37154
rect 7870 37102 7922 37154
rect 14254 37102 14306 37154
rect 18398 37102 18450 37154
rect 2158 36990 2210 37042
rect 3166 36990 3218 37042
rect 4286 36990 4338 37042
rect 10670 36990 10722 37042
rect 11790 36990 11842 37042
rect 15262 36990 15314 37042
rect 19630 36990 19682 37042
rect 21422 36990 21474 37042
rect 22542 36990 22594 37042
rect 4466 36822 4518 36874
rect 4570 36822 4622 36874
rect 4674 36822 4726 36874
rect 24466 36822 24518 36874
rect 24570 36822 24622 36874
rect 24674 36822 24726 36874
rect 2494 36654 2546 36706
rect 16046 36654 16098 36706
rect 17950 36654 18002 36706
rect 23662 36654 23714 36706
rect 7310 36542 7362 36594
rect 11342 36542 11394 36594
rect 11790 36542 11842 36594
rect 14814 36542 14866 36594
rect 19630 36542 19682 36594
rect 19966 36542 20018 36594
rect 21310 36542 21362 36594
rect 23998 36542 24050 36594
rect 1486 36430 1538 36482
rect 1822 36430 1874 36482
rect 2270 36430 2322 36482
rect 2942 36430 2994 36482
rect 3502 36430 3554 36482
rect 3726 36430 3778 36482
rect 4510 36430 4562 36482
rect 5182 36430 5234 36482
rect 6078 36430 6130 36482
rect 6750 36430 6802 36482
rect 7534 36430 7586 36482
rect 7870 36430 7922 36482
rect 8318 36430 8370 36482
rect 10334 36430 10386 36482
rect 10670 36430 10722 36482
rect 11118 36430 11170 36482
rect 12350 36430 12402 36482
rect 13358 36430 13410 36482
rect 14366 36430 14418 36482
rect 20862 36430 20914 36482
rect 18398 36318 18450 36370
rect 16830 36206 16882 36258
rect 19070 36206 19122 36258
rect 19406 36206 19458 36258
rect 22542 36206 22594 36258
rect 3806 36038 3858 36090
rect 3910 36038 3962 36090
rect 4014 36038 4066 36090
rect 23806 36038 23858 36090
rect 23910 36038 23962 36090
rect 24014 36038 24066 36090
rect 15038 35870 15090 35922
rect 16942 35870 16994 35922
rect 19294 35870 19346 35922
rect 1150 35758 1202 35810
rect 12238 35758 12290 35810
rect 20974 35758 21026 35810
rect 1486 35646 1538 35698
rect 2046 35646 2098 35698
rect 2718 35646 2770 35698
rect 3278 35646 3330 35698
rect 4174 35646 4226 35698
rect 5742 35646 5794 35698
rect 6190 35646 6242 35698
rect 6862 35646 6914 35698
rect 7422 35646 7474 35698
rect 8430 35646 8482 35698
rect 9214 35646 9266 35698
rect 10222 35646 10274 35698
rect 10558 35646 10610 35698
rect 11342 35646 11394 35698
rect 11790 35646 11842 35698
rect 13470 35646 13522 35698
rect 16382 35646 16434 35698
rect 17166 35646 17218 35698
rect 17726 35646 17778 35698
rect 21422 35646 21474 35698
rect 21758 35646 21810 35698
rect 22542 35646 22594 35698
rect 22990 35646 23042 35698
rect 24110 35646 24162 35698
rect 30270 35646 30322 35698
rect 5406 35534 5458 35586
rect 6414 35534 6466 35586
rect 16046 35534 16098 35586
rect 16606 35534 16658 35586
rect 18062 35534 18114 35586
rect 19742 35534 19794 35586
rect 2158 35422 2210 35474
rect 11230 35422 11282 35474
rect 13918 35422 13970 35474
rect 15710 35422 15762 35474
rect 15934 35422 15986 35474
rect 17166 35422 17218 35474
rect 19854 35422 19906 35474
rect 19966 35422 20018 35474
rect 21982 35422 22034 35474
rect 30606 35422 30658 35474
rect 4466 35254 4518 35306
rect 4570 35254 4622 35306
rect 4674 35254 4726 35306
rect 24466 35254 24518 35306
rect 24570 35254 24622 35306
rect 24674 35254 24726 35306
rect 3726 35086 3778 35138
rect 13918 35086 13970 35138
rect 20302 35086 20354 35138
rect 21758 35086 21810 35138
rect 30270 35086 30322 35138
rect 6078 34974 6130 35026
rect 6526 34974 6578 35026
rect 9102 34974 9154 35026
rect 11342 34974 11394 35026
rect 12462 34974 12514 35026
rect 17502 34974 17554 35026
rect 17838 34974 17890 35026
rect 19182 34974 19234 35026
rect 20750 34974 20802 35026
rect 24782 34974 24834 35026
rect 30606 34974 30658 35026
rect 1710 34862 1762 34914
rect 2718 34862 2770 34914
rect 3278 34862 3330 34914
rect 3838 34850 3890 34902
rect 4286 34862 4338 34914
rect 4734 34862 4786 34914
rect 5518 34862 5570 34914
rect 5854 34862 5906 34914
rect 7086 34862 7138 34914
rect 7310 34862 7362 34914
rect 8094 34862 8146 34914
rect 9214 34862 9266 34914
rect 9774 34862 9826 34914
rect 13246 34862 13298 34914
rect 13806 34862 13858 34914
rect 14366 34862 14418 34914
rect 14926 34862 14978 34914
rect 15934 34862 15986 34914
rect 17166 34862 17218 34914
rect 17278 34862 17330 34914
rect 18062 34862 18114 34914
rect 21198 34862 21250 34914
rect 21534 34862 21586 34914
rect 22430 34862 22482 34914
rect 22766 34862 22818 34914
rect 23774 34862 23826 34914
rect 24670 34862 24722 34914
rect 25454 34862 25506 34914
rect 5070 34750 5122 34802
rect 10894 34750 10946 34802
rect 12910 34750 12962 34802
rect 16718 34750 16770 34802
rect 18174 34750 18226 34802
rect 18734 34750 18786 34802
rect 10110 34638 10162 34690
rect 16830 34638 16882 34690
rect 25790 34638 25842 34690
rect 3806 34470 3858 34522
rect 3910 34470 3962 34522
rect 4014 34470 4066 34522
rect 23806 34470 23858 34522
rect 23910 34470 23962 34522
rect 24014 34470 24066 34522
rect 7870 34302 7922 34354
rect 2382 34190 2434 34242
rect 6302 34190 6354 34242
rect 16830 34190 16882 34242
rect 20974 34190 21026 34242
rect 3950 34078 4002 34130
rect 9102 34078 9154 34130
rect 9662 34078 9714 34130
rect 10446 34078 10498 34130
rect 10782 34078 10834 34130
rect 11902 34078 11954 34130
rect 14702 34078 14754 34130
rect 17278 34078 17330 34130
rect 17614 34078 17666 34130
rect 18846 34078 18898 34130
rect 19854 34078 19906 34130
rect 21422 34078 21474 34130
rect 21758 34078 21810 34130
rect 22654 34078 22706 34130
rect 22990 34078 23042 34130
rect 23998 34078 24050 34130
rect 24894 34078 24946 34130
rect 25454 34078 25506 34130
rect 30270 34078 30322 34130
rect 3502 33966 3554 34018
rect 6638 33966 6690 34018
rect 8766 33966 8818 34018
rect 9774 33966 9826 34018
rect 17838 33966 17890 34018
rect 18286 33966 18338 34018
rect 21982 33966 22034 34018
rect 24670 33966 24722 34018
rect 12798 33854 12850 33906
rect 15262 33854 15314 33906
rect 16382 33854 16434 33906
rect 25790 33854 25842 33906
rect 30606 33854 30658 33906
rect 4466 33686 4518 33738
rect 4570 33686 4622 33738
rect 4674 33686 4726 33738
rect 24466 33686 24518 33738
rect 24570 33686 24622 33738
rect 24674 33686 24726 33738
rect 6302 33518 6354 33570
rect 17726 33518 17778 33570
rect 19070 33518 19122 33570
rect 21758 33518 21810 33570
rect 1822 33406 1874 33458
rect 2158 33406 2210 33458
rect 2606 33406 2658 33458
rect 3614 33406 3666 33458
rect 7422 33406 7474 33458
rect 11678 33406 11730 33458
rect 14702 33406 14754 33458
rect 18286 33406 18338 33458
rect 19294 33406 19346 33458
rect 19630 33406 19682 33458
rect 20750 33406 20802 33458
rect 30606 33406 30658 33458
rect 2942 33294 2994 33346
rect 3390 33294 3442 33346
rect 4286 33294 4338 33346
rect 4622 33294 4674 33346
rect 4846 33294 4898 33346
rect 5630 33294 5682 33346
rect 14142 33294 14194 33346
rect 17054 33294 17106 33346
rect 17502 33294 17554 33346
rect 18062 33294 18114 33346
rect 18510 33294 18562 33346
rect 18958 33294 19010 33346
rect 19518 33294 19570 33346
rect 21086 33294 21138 33346
rect 21534 33294 21586 33346
rect 22318 33294 22370 33346
rect 22766 33294 22818 33346
rect 23774 33294 23826 33346
rect 30382 33294 30434 33346
rect 7870 33182 7922 33234
rect 11230 33182 11282 33234
rect 16718 33182 16770 33234
rect 16830 33182 16882 33234
rect 17614 33182 17666 33234
rect 18734 33182 18786 33234
rect 19854 33182 19906 33234
rect 29598 33182 29650 33234
rect 12798 33070 12850 33122
rect 15822 33070 15874 33122
rect 20078 33070 20130 33122
rect 29710 33070 29762 33122
rect 3806 32902 3858 32954
rect 3910 32902 3962 32954
rect 4014 32902 4066 32954
rect 23806 32902 23858 32954
rect 23910 32902 23962 32954
rect 24014 32902 24066 32954
rect 1150 32734 1202 32786
rect 7982 32734 8034 32786
rect 9886 32734 9938 32786
rect 13694 32734 13746 32786
rect 19294 32734 19346 32786
rect 23438 32734 23490 32786
rect 6414 32622 6466 32674
rect 15150 32622 15202 32674
rect 21086 32622 21138 32674
rect 2830 32510 2882 32562
rect 11454 32510 11506 32562
rect 13022 32510 13074 32562
rect 15598 32510 15650 32562
rect 15934 32510 15986 32562
rect 16606 32510 16658 32562
rect 17278 32510 17330 32562
rect 18174 32510 18226 32562
rect 18734 32510 18786 32562
rect 18958 32510 19010 32562
rect 19406 32510 19458 32562
rect 20526 32510 20578 32562
rect 20974 32510 21026 32562
rect 21198 32510 21250 32562
rect 21870 32510 21922 32562
rect 2382 32398 2434 32450
rect 11006 32398 11058 32450
rect 12910 32398 12962 32450
rect 16158 32398 16210 32450
rect 6862 32286 6914 32338
rect 14030 32286 14082 32338
rect 19518 32286 19570 32338
rect 22318 32286 22370 32338
rect 4466 32118 4518 32170
rect 4570 32118 4622 32170
rect 4674 32118 4726 32170
rect 24466 32118 24518 32170
rect 24570 32118 24622 32170
rect 24674 32118 24726 32170
rect 13806 31950 13858 32002
rect 18062 31950 18114 32002
rect 18286 31950 18338 32002
rect 22094 31950 22146 32002
rect 30270 31950 30322 32002
rect 2942 31838 2994 31890
rect 5630 31838 5682 31890
rect 6750 31838 6802 31890
rect 9550 31838 9602 31890
rect 10670 31838 10722 31890
rect 11902 31838 11954 31890
rect 14926 31838 14978 31890
rect 16046 31838 16098 31890
rect 17390 31838 17442 31890
rect 19070 31838 19122 31890
rect 23214 31838 23266 31890
rect 30606 31838 30658 31890
rect 2382 31726 2434 31778
rect 2718 31726 2770 31778
rect 3614 31726 3666 31778
rect 4174 31726 4226 31778
rect 4958 31726 5010 31778
rect 16158 31726 16210 31778
rect 17054 31726 17106 31778
rect 17614 31726 17666 31778
rect 19294 31726 19346 31778
rect 19518 31726 19570 31778
rect 21534 31726 21586 31778
rect 1934 31614 1986 31666
rect 7198 31614 7250 31666
rect 9102 31614 9154 31666
rect 11566 31614 11618 31666
rect 15374 31614 15426 31666
rect 18174 31614 18226 31666
rect 19630 31614 19682 31666
rect 13134 31502 13186 31554
rect 17054 31502 17106 31554
rect 18622 31502 18674 31554
rect 18734 31502 18786 31554
rect 3806 31334 3858 31386
rect 3910 31334 3962 31386
rect 4014 31334 4066 31386
rect 23806 31334 23858 31386
rect 23910 31334 23962 31386
rect 24014 31334 24066 31386
rect 3166 31166 3218 31218
rect 5070 31166 5122 31218
rect 8990 31166 9042 31218
rect 15150 31166 15202 31218
rect 18510 31166 18562 31218
rect 7422 31054 7474 31106
rect 17166 31054 17218 31106
rect 1598 30942 1650 30994
rect 6750 30942 6802 30994
rect 10446 30942 10498 30994
rect 13022 30942 13074 30994
rect 15486 30942 15538 30994
rect 16606 30942 16658 30994
rect 17054 30942 17106 30994
rect 17278 30942 17330 30994
rect 18062 30942 18114 30994
rect 19742 30942 19794 30994
rect 20078 30942 20130 30994
rect 30382 30942 30434 30994
rect 2046 30830 2098 30882
rect 6190 30830 6242 30882
rect 11006 30830 11058 30882
rect 13358 30830 13410 30882
rect 15710 30830 15762 30882
rect 16046 30830 16098 30882
rect 17726 30830 17778 30882
rect 19294 30830 19346 30882
rect 19518 30830 19570 30882
rect 7870 30718 7922 30770
rect 12126 30718 12178 30770
rect 14590 30718 14642 30770
rect 18846 30718 18898 30770
rect 20078 30718 20130 30770
rect 30606 30718 30658 30770
rect 4466 30550 4518 30602
rect 4570 30550 4622 30602
rect 4674 30550 4726 30602
rect 24466 30550 24518 30602
rect 24570 30550 24622 30602
rect 24674 30550 24726 30602
rect 7086 30382 7138 30434
rect 10222 30382 10274 30434
rect 12798 30382 12850 30434
rect 16270 30382 16322 30434
rect 17838 30382 17890 30434
rect 18846 30382 18898 30434
rect 20750 30382 20802 30434
rect 2718 30270 2770 30322
rect 3726 30270 3778 30322
rect 15934 30270 15986 30322
rect 16046 30270 16098 30322
rect 17054 30270 17106 30322
rect 21310 30270 21362 30322
rect 21422 30270 21474 30322
rect 30606 30270 30658 30322
rect 3054 30158 3106 30210
rect 3502 30158 3554 30210
rect 4286 30158 4338 30210
rect 4846 30158 4898 30210
rect 5742 30158 5794 30210
rect 6638 30158 6690 30210
rect 9774 30158 9826 30210
rect 11790 30158 11842 30210
rect 12238 30158 12290 30210
rect 12574 30158 12626 30210
rect 13470 30158 13522 30210
rect 13806 30158 13858 30210
rect 14814 30158 14866 30210
rect 17278 30158 17330 30210
rect 17838 30158 17890 30210
rect 20302 30158 20354 30210
rect 20862 30158 20914 30210
rect 20974 30158 21026 30210
rect 21646 30158 21698 30210
rect 30270 30158 30322 30210
rect 18398 30046 18450 30098
rect 8206 29934 8258 29986
rect 11342 29934 11394 29986
rect 17614 29934 17666 29986
rect 19966 29934 20018 29986
rect 3806 29766 3858 29818
rect 3910 29766 3962 29818
rect 4014 29766 4066 29818
rect 23806 29766 23858 29818
rect 23910 29766 23962 29818
rect 24014 29766 24066 29818
rect 1150 29598 1202 29650
rect 5070 29598 5122 29650
rect 20750 29598 20802 29650
rect 2718 29486 2770 29538
rect 6638 29486 6690 29538
rect 7534 29486 7586 29538
rect 16830 29486 16882 29538
rect 10558 29374 10610 29426
rect 14366 29374 14418 29426
rect 17166 29374 17218 29426
rect 17614 29374 17666 29426
rect 18286 29374 18338 29426
rect 18846 29374 18898 29426
rect 19854 29374 19906 29426
rect 20638 29374 20690 29426
rect 21310 29374 21362 29426
rect 21870 29374 21922 29426
rect 22206 29374 22258 29426
rect 30270 29374 30322 29426
rect 2270 29262 2322 29314
rect 6190 29262 6242 29314
rect 7982 29262 8034 29314
rect 11006 29262 11058 29314
rect 14814 29262 14866 29314
rect 17838 29262 17890 29314
rect 20974 29262 21026 29314
rect 21534 29262 21586 29314
rect 22542 29262 22594 29314
rect 9102 29150 9154 29202
rect 12126 29150 12178 29202
rect 15934 29150 15986 29202
rect 21422 29150 21474 29202
rect 22094 29150 22146 29202
rect 30606 29150 30658 29202
rect 4466 28982 4518 29034
rect 4570 28982 4622 29034
rect 4674 28982 4726 29034
rect 24466 28982 24518 29034
rect 24570 28982 24622 29034
rect 24674 28982 24726 29034
rect 2158 28814 2210 28866
rect 3278 28814 3330 28866
rect 7310 28814 7362 28866
rect 17502 28814 17554 28866
rect 18622 28814 18674 28866
rect 21310 28814 21362 28866
rect 8318 28702 8370 28754
rect 9886 28702 9938 28754
rect 13918 28702 13970 28754
rect 19630 28702 19682 28754
rect 30270 28702 30322 28754
rect 30606 28702 30658 28754
rect 1710 28590 1762 28642
rect 5182 28590 5234 28642
rect 6078 28590 6130 28642
rect 6862 28590 6914 28642
rect 7534 28590 7586 28642
rect 7982 28590 8034 28642
rect 9214 28590 9266 28642
rect 9774 28590 9826 28642
rect 10446 28590 10498 28642
rect 10894 28590 10946 28642
rect 11118 28590 11170 28642
rect 11790 28595 11842 28647
rect 13246 28590 13298 28642
rect 13806 28590 13858 28642
rect 14590 28590 14642 28642
rect 15038 28590 15090 28642
rect 15934 28590 15986 28642
rect 19966 28590 20018 28642
rect 8878 28478 8930 28530
rect 12910 28478 12962 28530
rect 19070 28478 19122 28530
rect 19742 28478 19794 28530
rect 20862 28478 20914 28530
rect 20078 28366 20130 28418
rect 22430 28366 22482 28418
rect 3806 28198 3858 28250
rect 3910 28198 3962 28250
rect 4014 28198 4066 28250
rect 23806 28198 23858 28250
rect 23910 28198 23962 28250
rect 24014 28198 24066 28250
rect 19966 28030 20018 28082
rect 21870 28030 21922 28082
rect 1150 27918 1202 27970
rect 6302 27918 6354 27970
rect 8318 27918 8370 27970
rect 20862 27918 20914 27970
rect 21982 27918 22034 27970
rect 1598 27806 1650 27858
rect 2046 27806 2098 27858
rect 2718 27806 2770 27858
rect 3278 27806 3330 27858
rect 4174 27806 4226 27858
rect 8654 27806 8706 27858
rect 9102 27806 9154 27858
rect 10558 27806 10610 27858
rect 11454 27806 11506 27858
rect 14478 27806 14530 27858
rect 14926 27806 14978 27858
rect 15822 27806 15874 27858
rect 16158 27806 16210 27858
rect 17166 27806 17218 27858
rect 18398 27806 18450 27858
rect 20638 27806 20690 27858
rect 21086 27806 21138 27858
rect 21310 27806 21362 27858
rect 21646 27806 21698 27858
rect 29598 27806 29650 27858
rect 30270 27806 30322 27858
rect 6638 27694 6690 27746
rect 9774 27694 9826 27746
rect 14142 27694 14194 27746
rect 18734 27694 18786 27746
rect 29710 27694 29762 27746
rect 2158 27582 2210 27634
rect 7870 27582 7922 27634
rect 9326 27582 9378 27634
rect 15150 27582 15202 27634
rect 20750 27582 20802 27634
rect 30606 27582 30658 27634
rect 4466 27414 4518 27466
rect 4570 27414 4622 27466
rect 4674 27414 4726 27466
rect 24466 27414 24518 27466
rect 24570 27414 24622 27466
rect 24674 27414 24726 27466
rect 18622 27246 18674 27298
rect 19182 27246 19234 27298
rect 21086 27246 21138 27298
rect 30270 27246 30322 27298
rect 1486 27134 1538 27186
rect 2494 27134 2546 27186
rect 7310 27134 7362 27186
rect 8318 27134 8370 27186
rect 9886 27134 9938 27186
rect 10334 27134 10386 27186
rect 14702 27134 14754 27186
rect 15150 27134 15202 27186
rect 16158 27134 16210 27186
rect 16942 27134 16994 27186
rect 18510 27134 18562 27186
rect 19294 27134 19346 27186
rect 19630 27134 19682 27186
rect 19742 27134 19794 27186
rect 30606 27134 30658 27186
rect 1822 27022 1874 27074
rect 2382 27022 2434 27074
rect 3166 27022 3218 27074
rect 3726 27022 3778 27074
rect 4510 27022 4562 27074
rect 5182 27022 5234 27074
rect 6078 27022 6130 27074
rect 6750 27022 6802 27074
rect 7534 27022 7586 27074
rect 7870 27022 7922 27074
rect 9214 27022 9266 27074
rect 9774 27022 9826 27074
rect 10894 27022 10946 27074
rect 11902 27022 11954 27074
rect 13022 27022 13074 27074
rect 13918 27022 13970 27074
rect 15262 27022 15314 27074
rect 15710 27022 15762 27074
rect 16830 27022 16882 27074
rect 17614 27022 17666 27074
rect 8878 26910 8930 26962
rect 21198 26910 21250 26962
rect 21310 26910 21362 26962
rect 21646 26910 21698 26962
rect 21758 26910 21810 26962
rect 17950 26798 18002 26850
rect 18622 26798 18674 26850
rect 19182 26798 19234 26850
rect 3806 26630 3858 26682
rect 3910 26630 3962 26682
rect 4014 26630 4066 26682
rect 23806 26630 23858 26682
rect 23910 26630 23962 26682
rect 24014 26630 24066 26682
rect 2830 26462 2882 26514
rect 16158 26462 16210 26514
rect 20750 26462 20802 26514
rect 1262 26350 1314 26402
rect 8766 26350 8818 26402
rect 13918 26350 13970 26402
rect 6638 26238 6690 26290
rect 8318 26238 8370 26290
rect 9102 26238 9154 26290
rect 9550 26238 9602 26290
rect 10334 26238 10386 26290
rect 10894 26238 10946 26290
rect 11902 26238 11954 26290
rect 14478 26238 14530 26290
rect 17166 26238 17218 26290
rect 22318 26238 22370 26290
rect 1598 26126 1650 26178
rect 7198 26014 7250 26066
rect 9774 26014 9826 26066
rect 14030 26014 14082 26066
rect 15038 26014 15090 26066
rect 16606 26014 16658 26066
rect 16718 26014 16770 26066
rect 16830 26014 16882 26066
rect 21870 26014 21922 26066
rect 4466 25846 4518 25898
rect 4570 25846 4622 25898
rect 4674 25846 4726 25898
rect 24466 25846 24518 25898
rect 24570 25846 24622 25898
rect 24674 25846 24726 25898
rect 4174 25678 4226 25730
rect 6190 25678 6242 25730
rect 7310 25678 7362 25730
rect 15598 25678 15650 25730
rect 17278 25678 17330 25730
rect 17726 25678 17778 25730
rect 17950 25678 18002 25730
rect 20750 25678 20802 25730
rect 22318 25678 22370 25730
rect 30270 25678 30322 25730
rect 3726 25566 3778 25618
rect 5182 25566 5234 25618
rect 9550 25566 9602 25618
rect 12910 25566 12962 25618
rect 16046 25566 16098 25618
rect 18062 25566 18114 25618
rect 30606 25566 30658 25618
rect 2158 25454 2210 25506
rect 2942 25454 2994 25506
rect 3166 25454 3218 25506
rect 4286 25454 4338 25506
rect 4846 25454 4898 25506
rect 5742 25454 5794 25506
rect 9102 25454 9154 25506
rect 12238 25454 12290 25506
rect 12798 25454 12850 25506
rect 13470 25454 13522 25506
rect 13918 25454 13970 25506
rect 14926 25454 14978 25506
rect 15710 25454 15762 25506
rect 15822 25454 15874 25506
rect 16270 25454 16322 25506
rect 16718 25454 16770 25506
rect 16942 25454 16994 25506
rect 17166 25454 17218 25506
rect 17390 25454 17442 25506
rect 21870 25454 21922 25506
rect 22542 25454 22594 25506
rect 22766 25454 22818 25506
rect 11902 25342 11954 25394
rect 20302 25342 20354 25394
rect 10670 25230 10722 25282
rect 22206 25230 22258 25282
rect 3806 25062 3858 25114
rect 3910 25062 3962 25114
rect 4014 25062 4066 25114
rect 23806 25062 23858 25114
rect 23910 25062 23962 25114
rect 24014 25062 24066 25114
rect 2830 24894 2882 24946
rect 6750 24894 6802 24946
rect 8094 24894 8146 24946
rect 14590 24894 14642 24946
rect 15598 24894 15650 24946
rect 21422 24894 21474 24946
rect 22206 24894 22258 24946
rect 5182 24782 5234 24834
rect 10558 24782 10610 24834
rect 13022 24782 13074 24834
rect 20862 24782 20914 24834
rect 21646 24782 21698 24834
rect 1262 24670 1314 24722
rect 7310 24670 7362 24722
rect 17278 24670 17330 24722
rect 20638 24670 20690 24722
rect 22094 24670 22146 24722
rect 30270 24670 30322 24722
rect 1598 24558 1650 24610
rect 5518 24558 5570 24610
rect 7534 24558 7586 24610
rect 8990 24558 9042 24610
rect 13358 24558 13410 24610
rect 16718 24558 16770 24610
rect 20974 24558 21026 24610
rect 21870 24558 21922 24610
rect 8430 24446 8482 24498
rect 10110 24446 10162 24498
rect 30606 24446 30658 24498
rect 4466 24278 4518 24330
rect 4570 24278 4622 24330
rect 4674 24278 4726 24330
rect 24466 24278 24518 24330
rect 24570 24278 24622 24330
rect 24674 24278 24726 24330
rect 1374 24110 1426 24162
rect 7422 24110 7474 24162
rect 1038 23998 1090 24050
rect 2942 23998 2994 24050
rect 3390 23998 3442 24050
rect 6190 23998 6242 24050
rect 10782 23998 10834 24050
rect 14814 23998 14866 24050
rect 19854 23998 19906 24050
rect 20302 23998 20354 24050
rect 21646 23998 21698 24050
rect 30270 23998 30322 24050
rect 30606 23998 30658 24050
rect 2382 23886 2434 23938
rect 2718 23886 2770 23938
rect 4062 23886 4114 23938
rect 4958 23886 5010 23938
rect 14478 23886 14530 23938
rect 19406 23886 19458 23938
rect 19630 23886 19682 23938
rect 23550 23886 23602 23938
rect 1934 23774 1986 23826
rect 5854 23774 5906 23826
rect 10446 23774 10498 23826
rect 20414 23774 20466 23826
rect 21198 23774 21250 23826
rect 23326 23774 23378 23826
rect 12014 23662 12066 23714
rect 16046 23662 16098 23714
rect 19518 23662 19570 23714
rect 20526 23662 20578 23714
rect 22766 23662 22818 23714
rect 23214 23662 23266 23714
rect 3806 23494 3858 23546
rect 3910 23494 3962 23546
rect 4014 23494 4066 23546
rect 23806 23494 23858 23546
rect 23910 23494 23962 23546
rect 24014 23494 24066 23546
rect 4286 23326 4338 23378
rect 6750 23326 6802 23378
rect 11678 23326 11730 23378
rect 16046 23326 16098 23378
rect 5182 23214 5234 23266
rect 14030 23214 14082 23266
rect 1262 23102 1314 23154
rect 2718 23102 2770 23154
rect 7646 23102 7698 23154
rect 8094 23102 8146 23154
rect 9438 23102 9490 23154
rect 10222 23102 10274 23154
rect 11006 23102 11058 23154
rect 14590 23102 14642 23154
rect 15262 23102 15314 23154
rect 15486 23102 15538 23154
rect 16830 23102 16882 23154
rect 17278 23102 17330 23154
rect 17502 23102 17554 23154
rect 18398 23102 18450 23154
rect 22430 23102 22482 23154
rect 23102 23102 23154 23154
rect 23214 23102 23266 23154
rect 23326 23102 23378 23154
rect 23662 23102 23714 23154
rect 23886 23102 23938 23154
rect 30270 23102 30322 23154
rect 7198 22990 7250 23042
rect 8654 22990 8706 23042
rect 10894 22990 10946 23042
rect 12014 22990 12066 23042
rect 13134 22990 13186 23042
rect 13246 22990 13298 23042
rect 13694 22990 13746 23042
rect 14366 22990 14418 23042
rect 14926 22990 14978 23042
rect 15598 22990 15650 23042
rect 16718 22990 16770 23042
rect 18846 22990 18898 23042
rect 21870 22990 21922 23042
rect 24222 22990 24274 23042
rect 1038 22878 1090 22930
rect 1710 22878 1762 22930
rect 2046 22878 2098 22930
rect 3166 22878 3218 22930
rect 5630 22878 5682 22930
rect 8206 22878 8258 22930
rect 13470 22878 13522 22930
rect 13918 22878 13970 22930
rect 14814 22878 14866 22930
rect 17614 22878 17666 22930
rect 19966 22878 20018 22930
rect 20750 22878 20802 22930
rect 23214 22878 23266 22930
rect 24110 22878 24162 22930
rect 30606 22878 30658 22930
rect 4466 22710 4518 22762
rect 4570 22710 4622 22762
rect 4674 22710 4726 22762
rect 24466 22710 24518 22762
rect 24570 22710 24622 22762
rect 24674 22710 24726 22762
rect 3726 22542 3778 22594
rect 4286 22542 4338 22594
rect 14926 22542 14978 22594
rect 16942 22542 16994 22594
rect 18062 22542 18114 22594
rect 23438 22542 23490 22594
rect 30270 22542 30322 22594
rect 2606 22430 2658 22482
rect 5406 22430 5458 22482
rect 7086 22430 7138 22482
rect 10446 22430 10498 22482
rect 12798 22430 12850 22482
rect 16158 22430 16210 22482
rect 20750 22430 20802 22482
rect 21198 22430 21250 22482
rect 30606 22430 30658 22482
rect 14366 22318 14418 22370
rect 14814 22318 14866 22370
rect 15038 22318 15090 22370
rect 15598 22318 15650 22370
rect 15934 22318 15986 22370
rect 20078 22318 20130 22370
rect 20526 22318 20578 22370
rect 21982 22318 22034 22370
rect 22766 22318 22818 22370
rect 23326 22318 23378 22370
rect 23550 22318 23602 22370
rect 2158 22206 2210 22258
rect 5854 22206 5906 22258
rect 6638 22206 6690 22258
rect 10110 22206 10162 22258
rect 12350 22206 12402 22258
rect 16158 22206 16210 22258
rect 17054 22206 17106 22258
rect 17614 22206 17666 22258
rect 19742 22206 19794 22258
rect 23774 22206 23826 22258
rect 8206 22094 8258 22146
rect 11678 22094 11730 22146
rect 13918 22094 13970 22146
rect 16718 22094 16770 22146
rect 19182 22094 19234 22146
rect 3806 21926 3858 21978
rect 3910 21926 3962 21978
rect 4014 21926 4066 21978
rect 23806 21926 23858 21978
rect 23910 21926 23962 21978
rect 24014 21926 24066 21978
rect 2942 21758 2994 21810
rect 5742 21758 5794 21810
rect 22542 21758 22594 21810
rect 23102 21758 23154 21810
rect 1374 21646 1426 21698
rect 16830 21646 16882 21698
rect 20974 21646 21026 21698
rect 7310 21534 7362 21586
rect 8094 21534 8146 21586
rect 13134 21534 13186 21586
rect 13582 21534 13634 21586
rect 14254 21534 14306 21586
rect 14814 21534 14866 21586
rect 15822 21534 15874 21586
rect 17166 21534 17218 21586
rect 17726 21534 17778 21586
rect 18398 21534 18450 21586
rect 19070 21534 19122 21586
rect 19854 21534 19906 21586
rect 20862 21534 20914 21586
rect 22990 21534 23042 21586
rect 1822 21422 1874 21474
rect 6862 21422 6914 21474
rect 7870 21422 7922 21474
rect 12798 21422 12850 21474
rect 16494 21422 16546 21474
rect 21422 21422 21474 21474
rect 3726 21310 3778 21362
rect 4062 21310 4114 21362
rect 8542 21310 8594 21362
rect 13806 21310 13858 21362
rect 16382 21310 16434 21362
rect 17838 21310 17890 21362
rect 30270 21310 30322 21362
rect 30606 21310 30658 21362
rect 4466 21142 4518 21194
rect 4570 21142 4622 21194
rect 4674 21142 4726 21194
rect 24466 21142 24518 21194
rect 24570 21142 24622 21194
rect 24674 21142 24726 21194
rect 16830 20974 16882 21026
rect 20750 20974 20802 21026
rect 3726 20862 3778 20914
rect 6078 20862 6130 20914
rect 9998 20862 10050 20914
rect 11678 20862 11730 20914
rect 12686 20862 12738 20914
rect 16158 20862 16210 20914
rect 18062 20862 18114 20914
rect 19518 20862 19570 20914
rect 21198 20862 21250 20914
rect 30606 20862 30658 20914
rect 1710 20750 1762 20802
rect 2606 20750 2658 20802
rect 3054 20750 3106 20802
rect 3838 20750 3890 20802
rect 4286 20750 4338 20802
rect 5518 20750 5570 20802
rect 5966 20750 6018 20802
rect 6526 20750 6578 20802
rect 7310 20750 7362 20802
rect 8094 20750 8146 20802
rect 11230 20750 11282 20802
rect 12126 20750 12178 20802
rect 12462 20750 12514 20802
rect 13134 20750 13186 20802
rect 13918 20750 13970 20802
rect 14702 20750 14754 20802
rect 15934 20750 15986 20802
rect 18398 20750 18450 20802
rect 21310 20750 21362 20802
rect 21534 20750 21586 20802
rect 21758 20750 21810 20802
rect 30270 20750 30322 20802
rect 4734 20638 4786 20690
rect 5070 20638 5122 20690
rect 9662 20638 9714 20690
rect 19182 20638 19234 20690
rect 15374 20526 15426 20578
rect 15598 20526 15650 20578
rect 16046 20526 16098 20578
rect 21982 20526 22034 20578
rect 3806 20358 3858 20410
rect 3910 20358 3962 20410
rect 4014 20358 4066 20410
rect 23806 20358 23858 20410
rect 23910 20358 23962 20410
rect 24014 20358 24066 20410
rect 14814 20190 14866 20242
rect 20638 20190 20690 20242
rect 1150 20078 1202 20130
rect 17166 20078 17218 20130
rect 17614 20078 17666 20130
rect 20750 20078 20802 20130
rect 1486 19966 1538 20018
rect 2046 19966 2098 20018
rect 3166 19966 3218 20018
rect 3390 19966 3442 20018
rect 4174 19966 4226 20018
rect 5406 19966 5458 20018
rect 5854 19966 5906 20018
rect 6750 19966 6802 20018
rect 7310 19966 7362 20018
rect 8094 19966 8146 20018
rect 8990 19966 9042 20018
rect 9438 19966 9490 20018
rect 10110 19966 10162 20018
rect 10670 19966 10722 20018
rect 11678 19966 11730 20018
rect 13134 19966 13186 20018
rect 15598 19966 15650 20018
rect 18398 19966 18450 20018
rect 2606 19854 2658 19906
rect 5070 19854 5122 19906
rect 8654 19854 8706 19906
rect 13694 19854 13746 19906
rect 16046 19854 16098 19906
rect 17726 19854 17778 19906
rect 19966 19854 20018 19906
rect 2158 19742 2210 19794
rect 6078 19742 6130 19794
rect 9662 19742 9714 19794
rect 18846 19742 18898 19794
rect 4466 19574 4518 19626
rect 4570 19574 4622 19626
rect 4674 19574 4726 19626
rect 24466 19574 24518 19626
rect 24570 19574 24622 19626
rect 24674 19574 24726 19626
rect 8206 19406 8258 19458
rect 15150 19406 15202 19458
rect 16270 19406 16322 19458
rect 17390 19406 17442 19458
rect 18510 19406 18562 19458
rect 19854 19406 19906 19458
rect 19966 19406 20018 19458
rect 30270 19406 30322 19458
rect 1262 19294 1314 19346
rect 1598 19294 1650 19346
rect 1934 19294 1986 19346
rect 2942 19294 2994 19346
rect 5518 19294 5570 19346
rect 7086 19294 7138 19346
rect 9998 19294 10050 19346
rect 11566 19294 11618 19346
rect 12574 19294 12626 19346
rect 15710 19294 15762 19346
rect 15934 19294 15986 19346
rect 16158 19294 16210 19346
rect 20078 19294 20130 19346
rect 30606 19294 30658 19346
rect 2382 19182 2434 19234
rect 2718 19182 2770 19234
rect 3502 19182 3554 19234
rect 3950 19182 4002 19234
rect 4958 19182 5010 19234
rect 5742 19182 5794 19234
rect 9550 19182 9602 19234
rect 11118 19182 11170 19234
rect 11902 19182 11954 19234
rect 12350 19182 12402 19234
rect 13134 19182 13186 19234
rect 13582 19182 13634 19234
rect 14590 19182 14642 19234
rect 16942 19182 16994 19234
rect 6638 19070 6690 19122
rect 15262 19070 15314 19122
rect 3806 18790 3858 18842
rect 3910 18790 3962 18842
rect 4014 18790 4066 18842
rect 23806 18790 23858 18842
rect 23910 18790 23962 18842
rect 24014 18790 24066 18842
rect 16830 18622 16882 18674
rect 17278 18622 17330 18674
rect 18286 18622 18338 18674
rect 6638 18510 6690 18562
rect 8654 18510 8706 18562
rect 13022 18510 13074 18562
rect 15262 18510 15314 18562
rect 17502 18510 17554 18562
rect 18062 18510 18114 18562
rect 1710 18398 1762 18450
rect 3278 18398 3330 18450
rect 4174 18398 4226 18450
rect 8206 18398 8258 18450
rect 8990 18398 9042 18450
rect 9438 18398 9490 18450
rect 9886 18398 9938 18450
rect 10670 18398 10722 18450
rect 11006 18398 11058 18450
rect 12014 18398 12066 18450
rect 14590 18398 14642 18450
rect 17950 18398 18002 18450
rect 30270 18398 30322 18450
rect 2158 18286 2210 18338
rect 3950 18286 4002 18338
rect 6974 18286 7026 18338
rect 13470 18286 13522 18338
rect 15598 18286 15650 18338
rect 17502 18286 17554 18338
rect 4958 18174 5010 18226
rect 5294 18174 5346 18226
rect 5630 18174 5682 18226
rect 5966 18174 6018 18226
rect 9998 18174 10050 18226
rect 30606 18174 30658 18226
rect 4466 18006 4518 18058
rect 4570 18006 4622 18058
rect 4674 18006 4726 18058
rect 24466 18006 24518 18058
rect 24570 18006 24622 18058
rect 24674 18006 24726 18058
rect 1150 17838 1202 17890
rect 2270 17838 2322 17890
rect 5518 17838 5570 17890
rect 7758 17838 7810 17890
rect 9550 17838 9602 17890
rect 10670 17838 10722 17890
rect 11902 17838 11954 17890
rect 13022 17838 13074 17890
rect 13806 17838 13858 17890
rect 16046 17838 16098 17890
rect 16942 17838 16994 17890
rect 30270 17838 30322 17890
rect 4286 17726 4338 17778
rect 6638 17726 6690 17778
rect 13694 17726 13746 17778
rect 13918 17726 13970 17778
rect 14926 17726 14978 17778
rect 17054 17726 17106 17778
rect 18286 17726 18338 17778
rect 18622 17726 18674 17778
rect 18958 17726 19010 17778
rect 19966 17726 20018 17778
rect 30606 17726 30658 17778
rect 2718 17614 2770 17666
rect 6190 17614 6242 17666
rect 9102 17614 9154 17666
rect 11342 17614 11394 17666
rect 14478 17614 14530 17666
rect 16718 17614 16770 17666
rect 19406 17614 19458 17666
rect 19742 17614 19794 17666
rect 20638 17614 20690 17666
rect 21198 17614 21250 17666
rect 21982 17614 22034 17666
rect 3950 17502 4002 17554
rect 3806 17222 3858 17274
rect 3910 17222 3962 17274
rect 4014 17222 4066 17274
rect 23806 17222 23858 17274
rect 23910 17222 23962 17274
rect 24014 17222 24066 17274
rect 1150 17054 1202 17106
rect 6974 17054 7026 17106
rect 9438 17054 9490 17106
rect 12910 17054 12962 17106
rect 19742 17054 19794 17106
rect 2718 16942 2770 16994
rect 5406 16942 5458 16994
rect 7870 16942 7922 16994
rect 11566 16942 11618 16994
rect 4286 16830 4338 16882
rect 9998 16830 10050 16882
rect 14590 16830 14642 16882
rect 18062 16830 18114 16882
rect 2270 16718 2322 16770
rect 3278 16718 3330 16770
rect 3950 16718 4002 16770
rect 5742 16718 5794 16770
rect 8206 16718 8258 16770
rect 14142 16718 14194 16770
rect 18510 16718 18562 16770
rect 3614 16606 3666 16658
rect 11118 16606 11170 16658
rect 30270 16606 30322 16658
rect 30606 16606 30658 16658
rect 4466 16438 4518 16490
rect 4570 16438 4622 16490
rect 4674 16438 4726 16490
rect 24466 16438 24518 16490
rect 24570 16438 24622 16490
rect 24674 16438 24726 16490
rect 2158 16270 2210 16322
rect 3278 16270 3330 16322
rect 4622 16270 4674 16322
rect 4958 16270 5010 16322
rect 5966 16270 6018 16322
rect 7086 16270 7138 16322
rect 7982 16270 8034 16322
rect 9550 16270 9602 16322
rect 16718 16270 16770 16322
rect 19854 16270 19906 16322
rect 20974 16270 21026 16322
rect 30270 16270 30322 16322
rect 3950 16158 4002 16210
rect 11230 16158 11282 16210
rect 11566 16158 11618 16210
rect 12910 16158 12962 16210
rect 17390 16158 17442 16210
rect 22654 16158 22706 16210
rect 30606 16158 30658 16210
rect 1710 16046 1762 16098
rect 4286 16046 4338 16098
rect 5518 16046 5570 16098
rect 8318 16046 8370 16098
rect 8990 16046 9042 16098
rect 12238 16046 12290 16098
rect 12798 16046 12850 16098
rect 13470 16046 13522 16098
rect 14030 16046 14082 16098
rect 14926 16046 14978 16098
rect 17054 16046 17106 16098
rect 17726 16046 17778 16098
rect 23102 16046 23154 16098
rect 11902 15934 11954 15986
rect 19406 15934 19458 15986
rect 10670 15822 10722 15874
rect 21534 15822 21586 15874
rect 3806 15654 3858 15706
rect 3910 15654 3962 15706
rect 4014 15654 4066 15706
rect 23806 15654 23858 15706
rect 23910 15654 23962 15706
rect 24014 15654 24066 15706
rect 2830 15486 2882 15538
rect 5070 15486 5122 15538
rect 1262 15374 1314 15426
rect 6638 15374 6690 15426
rect 14478 15374 14530 15426
rect 21198 15374 21250 15426
rect 3614 15262 3666 15314
rect 8766 15262 8818 15314
rect 9326 15262 9378 15314
rect 10110 15262 10162 15314
rect 10670 15262 10722 15314
rect 11566 15262 11618 15314
rect 15934 15262 15986 15314
rect 18062 15262 18114 15314
rect 30382 15262 30434 15314
rect 1598 15150 1650 15202
rect 3278 15150 3330 15202
rect 4062 15150 4114 15202
rect 4398 15150 4450 15202
rect 8430 15150 8482 15202
rect 9438 15150 9490 15202
rect 12910 15150 12962 15202
rect 14030 15150 14082 15202
rect 15038 15150 15090 15202
rect 16270 15150 16322 15202
rect 18622 15150 18674 15202
rect 21646 15150 21698 15202
rect 6190 15038 6242 15090
rect 7758 15038 7810 15090
rect 8094 15038 8146 15090
rect 15374 15038 15426 15090
rect 17502 15038 17554 15090
rect 19742 15038 19794 15090
rect 22766 15038 22818 15090
rect 30606 15038 30658 15090
rect 4466 14870 4518 14922
rect 4570 14870 4622 14922
rect 4674 14870 4726 14922
rect 24466 14870 24518 14922
rect 24570 14870 24622 14922
rect 24674 14870 24726 14922
rect 6078 14702 6130 14754
rect 12462 14702 12514 14754
rect 13918 14702 13970 14754
rect 17726 14702 17778 14754
rect 30270 14702 30322 14754
rect 3726 14590 3778 14642
rect 5070 14590 5122 14642
rect 8878 14590 8930 14642
rect 9550 14590 9602 14642
rect 11342 14590 11394 14642
rect 21758 14590 21810 14642
rect 30606 14590 30658 14642
rect 1710 14478 1762 14530
rect 2718 14478 2770 14530
rect 3278 14478 3330 14530
rect 3838 14478 3890 14530
rect 4398 14478 4450 14530
rect 5518 14478 5570 14530
rect 5854 14478 5906 14530
rect 6638 14478 6690 14530
rect 7310 14478 7362 14530
rect 8094 14478 8146 14530
rect 9102 14478 9154 14530
rect 9886 14478 9938 14530
rect 13358 14478 13410 14530
rect 13694 14478 13746 14530
rect 14590 14478 14642 14530
rect 15038 14478 15090 14530
rect 15934 14478 15986 14530
rect 17166 14478 17218 14530
rect 17502 14478 17554 14530
rect 18174 14478 18226 14530
rect 18734 14478 18786 14530
rect 19742 14478 19794 14530
rect 21086 14478 21138 14530
rect 21534 14478 21586 14530
rect 22430 14478 22482 14530
rect 22766 14478 22818 14530
rect 23774 14478 23826 14530
rect 4734 14366 4786 14418
rect 10894 14366 10946 14418
rect 12910 14366 12962 14418
rect 16718 14366 16770 14418
rect 20750 14366 20802 14418
rect 3806 14086 3858 14138
rect 3910 14086 3962 14138
rect 4014 14086 4066 14138
rect 23806 14086 23858 14138
rect 23910 14086 23962 14138
rect 24014 14086 24066 14138
rect 7870 13918 7922 13970
rect 15038 13918 15090 13970
rect 18174 13918 18226 13970
rect 8318 13806 8370 13858
rect 30158 13806 30210 13858
rect 1262 13694 1314 13746
rect 2270 13694 2322 13746
rect 3502 13694 3554 13746
rect 4062 13694 4114 13746
rect 5294 13694 5346 13746
rect 6302 13694 6354 13746
rect 8654 13694 8706 13746
rect 9102 13694 9154 13746
rect 9998 13694 10050 13746
rect 10334 13694 10386 13746
rect 11342 13694 11394 13746
rect 13470 13694 13522 13746
rect 16606 13694 16658 13746
rect 21198 13694 21250 13746
rect 21534 13694 21586 13746
rect 22206 13694 22258 13746
rect 22766 13694 22818 13746
rect 23774 13694 23826 13746
rect 2942 13582 2994 13634
rect 4398 13582 4450 13634
rect 4958 13582 5010 13634
rect 6750 13582 6802 13634
rect 9326 13582 9378 13634
rect 11902 13582 11954 13634
rect 12238 13582 12290 13634
rect 13918 13582 13970 13634
rect 16942 13582 16994 13634
rect 20750 13582 20802 13634
rect 21758 13582 21810 13634
rect 3390 13470 3442 13522
rect 4466 13302 4518 13354
rect 4570 13302 4622 13354
rect 4674 13302 4726 13354
rect 24466 13302 24518 13354
rect 24570 13302 24622 13354
rect 24674 13302 24726 13354
rect 8878 13134 8930 13186
rect 11902 13134 11954 13186
rect 13022 13134 13074 13186
rect 14142 13134 14194 13186
rect 18734 13134 18786 13186
rect 21422 13134 21474 13186
rect 30270 13134 30322 13186
rect 3726 13022 3778 13074
rect 5070 13022 5122 13074
rect 6078 13022 6130 13074
rect 9214 13022 9266 13074
rect 10782 13022 10834 13074
rect 17054 13022 17106 13074
rect 17726 13022 17778 13074
rect 22542 13022 22594 13074
rect 30606 13022 30658 13074
rect 1710 12910 1762 12962
rect 2494 12910 2546 12962
rect 3054 12910 3106 12962
rect 3950 12910 4002 12962
rect 4398 12910 4450 12962
rect 5406 12910 5458 12962
rect 5854 12910 5906 12962
rect 6750 12910 6802 12962
rect 7086 12910 7138 12962
rect 8094 12910 8146 12962
rect 17390 12910 17442 12962
rect 18174 12910 18226 12962
rect 18622 12910 18674 12962
rect 19406 12910 19458 12962
rect 19966 12910 20018 12962
rect 20750 12910 20802 12962
rect 4734 12798 4786 12850
rect 10334 12798 10386 12850
rect 12574 12798 12626 12850
rect 22990 12798 23042 12850
rect 3806 12518 3858 12570
rect 3910 12518 3962 12570
rect 4014 12518 4066 12570
rect 23806 12518 23858 12570
rect 23910 12518 23962 12570
rect 24014 12518 24066 12570
rect 3390 12350 3442 12402
rect 7870 12350 7922 12402
rect 10110 12350 10162 12402
rect 18286 12350 18338 12402
rect 20750 12350 20802 12402
rect 14478 12238 14530 12290
rect 1822 12126 1874 12178
rect 6302 12126 6354 12178
rect 8430 12126 8482 12178
rect 11230 12126 11282 12178
rect 12126 12126 12178 12178
rect 16718 12126 16770 12178
rect 22430 12126 22482 12178
rect 30382 12126 30434 12178
rect 2270 12014 2322 12066
rect 4958 12014 5010 12066
rect 10894 12014 10946 12066
rect 14030 12014 14082 12066
rect 3838 11902 3890 11954
rect 4174 11902 4226 11954
rect 5294 11902 5346 11954
rect 6750 11902 6802 11954
rect 8990 11902 9042 11954
rect 10558 11902 10610 11954
rect 11566 11902 11618 11954
rect 11902 11902 11954 11954
rect 12910 11902 12962 11954
rect 17166 11902 17218 11954
rect 21870 11902 21922 11954
rect 30606 11902 30658 11954
rect 4466 11734 4518 11786
rect 4570 11734 4622 11786
rect 4674 11734 4726 11786
rect 24466 11734 24518 11786
rect 24570 11734 24622 11786
rect 24674 11734 24726 11786
rect 2830 11566 2882 11618
rect 3390 11566 3442 11618
rect 7310 11566 7362 11618
rect 11454 11566 11506 11618
rect 19182 11566 19234 11618
rect 30270 11566 30322 11618
rect 1598 11454 1650 11506
rect 4622 11454 4674 11506
rect 6078 11454 6130 11506
rect 7758 11454 7810 11506
rect 8878 11454 8930 11506
rect 10110 11454 10162 11506
rect 13918 11454 13970 11506
rect 18174 11454 18226 11506
rect 30606 11454 30658 11506
rect 4958 11342 5010 11394
rect 8094 11342 8146 11394
rect 9102 11342 9154 11394
rect 10446 11342 10498 11394
rect 11006 11342 11058 11394
rect 13470 11342 13522 11394
rect 18510 11342 18562 11394
rect 18958 11342 19010 11394
rect 19742 11342 19794 11394
rect 20414 11342 20466 11394
rect 21198 11342 21250 11394
rect 1262 11230 1314 11282
rect 5742 11230 5794 11282
rect 12574 11118 12626 11170
rect 15038 11118 15090 11170
rect 3806 10950 3858 11002
rect 3910 10950 3962 11002
rect 4014 10950 4066 11002
rect 23806 10950 23858 11002
rect 23910 10950 23962 11002
rect 24014 10950 24066 11002
rect 2830 10782 2882 10834
rect 7198 10782 7250 10834
rect 18510 10782 18562 10834
rect 1262 10670 1314 10722
rect 3502 10558 3554 10610
rect 4174 10558 4226 10610
rect 5630 10558 5682 10610
rect 8766 10558 8818 10610
rect 9662 10558 9714 10610
rect 11006 10558 11058 10610
rect 11566 10558 11618 10610
rect 13022 10558 13074 10610
rect 13694 10558 13746 10610
rect 16942 10558 16994 10610
rect 22318 10558 22370 10610
rect 1598 10446 1650 10498
rect 3950 10446 4002 10498
rect 5966 10446 6018 10498
rect 7646 10446 7698 10498
rect 10446 10446 10498 10498
rect 10894 10446 10946 10498
rect 11902 10446 11954 10498
rect 12798 10446 12850 10498
rect 14142 10446 14194 10498
rect 15710 10446 15762 10498
rect 17278 10446 17330 10498
rect 20750 10446 20802 10498
rect 21870 10446 21922 10498
rect 3278 10334 3330 10386
rect 7982 10334 8034 10386
rect 15262 10334 15314 10386
rect 16046 10334 16098 10386
rect 17390 10334 17442 10386
rect 4466 10166 4518 10218
rect 4570 10166 4622 10218
rect 4674 10166 4726 10218
rect 24466 10166 24518 10218
rect 24570 10166 24622 10218
rect 24674 10166 24726 10218
rect 1150 9998 1202 10050
rect 2270 9998 2322 10050
rect 5966 9998 6018 10050
rect 10334 9998 10386 10050
rect 12014 9998 12066 10050
rect 14926 9998 14978 10050
rect 16718 9998 16770 10050
rect 19742 9998 19794 10050
rect 21198 9998 21250 10050
rect 4734 9886 4786 9938
rect 7086 9886 7138 9938
rect 8878 9886 8930 9938
rect 9550 9886 9602 9938
rect 14590 9886 14642 9938
rect 15262 9886 15314 9938
rect 18510 9886 18562 9938
rect 6526 9774 6578 9826
rect 9102 9774 9154 9826
rect 9774 9774 9826 9826
rect 10670 9774 10722 9826
rect 11342 9774 11394 9826
rect 11790 9774 11842 9826
rect 12574 9774 12626 9826
rect 13022 9774 13074 9826
rect 14030 9774 14082 9826
rect 15486 9774 15538 9826
rect 17054 9774 17106 9826
rect 18062 9774 18114 9826
rect 20638 9774 20690 9826
rect 21086 9762 21138 9814
rect 21870 9774 21922 9826
rect 22206 9774 22258 9826
rect 22430 9774 22482 9826
rect 23326 9774 23378 9826
rect 2718 9662 2770 9714
rect 4398 9662 4450 9714
rect 11006 9662 11058 9714
rect 20190 9662 20242 9714
rect 8206 9550 8258 9602
rect 3806 9382 3858 9434
rect 3910 9382 3962 9434
rect 4014 9382 4066 9434
rect 23806 9382 23858 9434
rect 23910 9382 23962 9434
rect 24014 9382 24066 9434
rect 4286 9214 4338 9266
rect 22430 9214 22482 9266
rect 13582 9102 13634 9154
rect 17278 9102 17330 9154
rect 18846 9102 18898 9154
rect 24558 9102 24610 9154
rect 1374 8990 1426 9042
rect 2046 8990 2098 9042
rect 2718 8990 2770 9042
rect 5294 8990 5346 9042
rect 5966 8990 6018 9042
rect 6862 8990 6914 9042
rect 7310 8990 7362 9042
rect 8430 8990 8482 9042
rect 9438 8990 9490 9042
rect 10558 8990 10610 9042
rect 12126 8990 12178 9042
rect 13918 8990 13970 9042
rect 14366 8990 14418 9042
rect 15150 8990 15202 9042
rect 15598 8990 15650 9042
rect 16606 8990 16658 9042
rect 20862 8990 20914 9042
rect 1038 8878 1090 8930
rect 1710 8878 1762 8930
rect 3166 8878 3218 8930
rect 6414 8878 6466 8930
rect 7870 8878 7922 8930
rect 14590 8878 14642 8930
rect 18510 8878 18562 8930
rect 21198 8878 21250 8930
rect 24110 8878 24162 8930
rect 4958 8766 5010 8818
rect 5630 8766 5682 8818
rect 7422 8766 7474 8818
rect 11006 8766 11058 8818
rect 12798 8766 12850 8818
rect 13134 8766 13186 8818
rect 19742 8766 19794 8818
rect 20078 8766 20130 8818
rect 22990 8766 23042 8818
rect 4466 8598 4518 8650
rect 4570 8598 4622 8650
rect 4674 8598 4726 8650
rect 24466 8598 24518 8650
rect 24570 8598 24622 8650
rect 24674 8598 24726 8650
rect 11118 8430 11170 8482
rect 20750 8430 20802 8482
rect 1038 8318 1090 8370
rect 1822 8318 1874 8370
rect 4062 8318 4114 8370
rect 6638 8318 6690 8370
rect 7310 8318 7362 8370
rect 7646 8318 7698 8370
rect 7982 8318 8034 8370
rect 9998 8318 10050 8370
rect 12574 8318 12626 8370
rect 13022 8318 13074 8370
rect 15150 8318 15202 8370
rect 15486 8318 15538 8370
rect 15822 8318 15874 8370
rect 17950 8318 18002 8370
rect 19518 8318 19570 8370
rect 21758 8318 21810 8370
rect 1374 8206 1426 8258
rect 2158 8206 2210 8258
rect 3502 8206 3554 8258
rect 3950 8206 4002 8258
rect 4734 8206 4786 8258
rect 5070 8206 5122 8258
rect 6078 8206 6130 8258
rect 6974 8206 7026 8258
rect 8206 8206 8258 8258
rect 11902 8206 11954 8258
rect 12350 8206 12402 8258
rect 13582 8206 13634 8258
rect 14590 8206 14642 8258
rect 16158 8206 16210 8258
rect 18398 8206 18450 8258
rect 19182 8206 19234 8258
rect 3054 8094 3106 8146
rect 9550 8094 9602 8146
rect 11566 8094 11618 8146
rect 21422 8094 21474 8146
rect 16830 7982 16882 8034
rect 22990 7982 23042 8034
rect 3806 7814 3858 7866
rect 3910 7814 3962 7866
rect 4014 7814 4066 7866
rect 23806 7814 23858 7866
rect 23910 7814 23962 7866
rect 24014 7814 24066 7866
rect 3390 7646 3442 7698
rect 12126 7646 12178 7698
rect 6750 7534 6802 7586
rect 10558 7534 10610 7586
rect 14590 7534 14642 7586
rect 18398 7534 18450 7586
rect 19966 7534 20018 7586
rect 20638 7534 20690 7586
rect 1822 7422 1874 7474
rect 5294 7422 5346 7474
rect 5742 7422 5794 7474
rect 7198 7422 7250 7474
rect 7646 7425 7698 7477
rect 8766 7422 8818 7474
rect 9774 7422 9826 7474
rect 15038 7422 15090 7474
rect 15374 7422 15426 7474
rect 16270 7422 16322 7474
rect 16718 7422 16770 7474
rect 17614 7422 17666 7474
rect 20974 7422 21026 7474
rect 21422 7422 21474 7474
rect 22318 7422 22370 7474
rect 22878 7422 22930 7474
rect 23662 7422 23714 7474
rect 2270 7310 2322 7362
rect 4958 7310 5010 7362
rect 5966 7310 6018 7362
rect 8206 7310 8258 7362
rect 13246 7310 13298 7362
rect 15598 7310 15650 7362
rect 18846 7310 18898 7362
rect 21646 7310 21698 7362
rect 7758 7198 7810 7250
rect 11006 7198 11058 7250
rect 13582 7198 13634 7250
rect 13918 7198 13970 7250
rect 14254 7198 14306 7250
rect 4466 7030 4518 7082
rect 4570 7030 4622 7082
rect 4674 7030 4726 7082
rect 24466 7030 24518 7082
rect 24570 7030 24622 7082
rect 24674 7030 24726 7082
rect 6638 6862 6690 6914
rect 8318 6862 8370 6914
rect 11342 6862 11394 6914
rect 13918 6862 13970 6914
rect 1710 6750 1762 6802
rect 2382 6750 2434 6802
rect 3054 6750 3106 6802
rect 4062 6750 4114 6802
rect 7310 6750 7362 6802
rect 8878 6750 8930 6802
rect 10334 6750 10386 6802
rect 19070 6750 19122 6802
rect 20078 6750 20130 6802
rect 21422 6750 21474 6802
rect 1374 6638 1426 6690
rect 2158 6638 2210 6690
rect 3390 6638 3442 6690
rect 3950 6638 4002 6690
rect 4734 6638 4786 6690
rect 5070 6638 5122 6690
rect 6078 6638 6130 6690
rect 6974 6638 7026 6690
rect 7646 6638 7698 6690
rect 7982 6638 8034 6690
rect 9102 6638 9154 6690
rect 10110 6638 10162 6690
rect 12462 6638 12514 6690
rect 13358 6638 13410 6690
rect 13694 6638 13746 6690
rect 14366 6638 14418 6690
rect 14926 6638 14978 6690
rect 15934 6638 15986 6690
rect 16942 6638 16994 6690
rect 18062 6638 18114 6690
rect 18622 6638 18674 6690
rect 19182 6638 19234 6690
rect 19742 6638 19794 6690
rect 20750 6638 20802 6690
rect 21310 6638 21362 6690
rect 22094 6638 22146 6690
rect 22430 6638 22482 6690
rect 23438 6638 23490 6690
rect 10894 6526 10946 6578
rect 12910 6526 12962 6578
rect 20414 6526 20466 6578
rect 3806 6246 3858 6298
rect 3910 6246 3962 6298
rect 4014 6246 4066 6298
rect 23806 6246 23858 6298
rect 23910 6246 23962 6298
rect 24014 6246 24066 6298
rect 20750 6078 20802 6130
rect 22990 6078 23042 6130
rect 10110 5966 10162 6018
rect 14814 5966 14866 6018
rect 1262 5854 1314 5906
rect 2270 5854 2322 5906
rect 3838 5854 3890 5906
rect 5070 5854 5122 5906
rect 6974 5854 7026 5906
rect 7870 5854 7922 5906
rect 8430 5854 8482 5906
rect 9214 5854 9266 5906
rect 9662 5854 9714 5906
rect 12014 5854 12066 5906
rect 13470 5854 13522 5906
rect 14142 5854 14194 5906
rect 15262 5854 15314 5906
rect 15598 5854 15650 5906
rect 16830 5854 16882 5906
rect 17838 5854 17890 5906
rect 18622 5854 18674 5906
rect 19630 5854 19682 5906
rect 22318 5854 22370 5906
rect 24558 5854 24610 5906
rect 25342 5854 25394 5906
rect 1038 5742 1090 5794
rect 5966 5742 6018 5794
rect 9102 5742 9154 5794
rect 12238 5742 12290 5794
rect 15822 5742 15874 5794
rect 16270 5742 16322 5794
rect 19406 5742 19458 5794
rect 21870 5742 21922 5794
rect 24110 5742 24162 5794
rect 25790 5742 25842 5794
rect 26910 5742 26962 5794
rect 2718 5630 2770 5682
rect 5294 5630 5346 5682
rect 5630 5630 5682 5682
rect 10558 5630 10610 5682
rect 10894 5630 10946 5682
rect 11230 5630 11282 5682
rect 11566 5630 11618 5682
rect 13246 5630 13298 5682
rect 13918 5630 13970 5682
rect 18398 5630 18450 5682
rect 4466 5462 4518 5514
rect 4570 5462 4622 5514
rect 4674 5462 4726 5514
rect 24466 5462 24518 5514
rect 24570 5462 24622 5514
rect 24674 5462 24726 5514
rect 1038 5294 1090 5346
rect 1374 5294 1426 5346
rect 2046 5294 2098 5346
rect 2382 5294 2434 5346
rect 2718 5294 2770 5346
rect 5406 5294 5458 5346
rect 7086 5294 7138 5346
rect 7982 5294 8034 5346
rect 10670 5294 10722 5346
rect 15374 5294 15426 5346
rect 18734 5294 18786 5346
rect 23326 5294 23378 5346
rect 23998 5294 24050 5346
rect 24446 5294 24498 5346
rect 26350 5294 26402 5346
rect 1710 5182 1762 5234
rect 4958 5182 5010 5234
rect 6414 5182 6466 5234
rect 6750 5182 6802 5234
rect 8318 5182 8370 5234
rect 9550 5182 9602 5234
rect 12238 5182 12290 5234
rect 15038 5182 15090 5234
rect 16158 5182 16210 5234
rect 17502 5182 17554 5234
rect 19406 5182 19458 5234
rect 20414 5182 20466 5234
rect 22990 5182 23042 5234
rect 23662 5182 23714 5234
rect 25118 5182 25170 5234
rect 3390 5070 3442 5122
rect 4174 5070 4226 5122
rect 5630 5070 5682 5122
rect 6078 5070 6130 5122
rect 11230 5070 11282 5122
rect 11566 5070 11618 5122
rect 12126 5070 12178 5122
rect 12686 5070 12738 5122
rect 13246 5070 13298 5122
rect 14254 5070 14306 5122
rect 15822 5070 15874 5122
rect 19742 5070 19794 5122
rect 20302 5070 20354 5122
rect 21086 5070 21138 5122
rect 21534 5070 21586 5122
rect 22430 5070 22482 5122
rect 9102 4958 9154 5010
rect 17166 4958 17218 5010
rect 3806 4678 3858 4730
rect 3910 4678 3962 4730
rect 4014 4678 4066 4730
rect 23806 4678 23858 4730
rect 23910 4678 23962 4730
rect 24014 4678 24066 4730
rect 4286 4510 4338 4562
rect 15598 4510 15650 4562
rect 17838 4510 17890 4562
rect 22430 4510 22482 4562
rect 22990 4510 23042 4562
rect 10110 4398 10162 4450
rect 1374 4286 1426 4338
rect 2046 4286 2098 4338
rect 2718 4286 2770 4338
rect 5182 4286 5234 4338
rect 6974 4286 7026 4338
rect 7870 4286 7922 4338
rect 9214 4286 9266 4338
rect 9774 4286 9826 4338
rect 10558 4286 10610 4338
rect 11566 4286 11618 4338
rect 12238 4286 12290 4338
rect 13358 4286 13410 4338
rect 14030 4286 14082 4338
rect 16270 4286 16322 4338
rect 18286 4286 18338 4338
rect 19294 4286 19346 4338
rect 19630 4286 19682 4338
rect 20862 4286 20914 4338
rect 24670 4286 24722 4338
rect 1038 4174 1090 4226
rect 1710 4174 1762 4226
rect 3166 4174 3218 4226
rect 5406 4174 5458 4226
rect 6078 4174 6130 4226
rect 8654 4174 8706 4226
rect 9102 4174 9154 4226
rect 10894 4174 10946 4226
rect 11902 4174 11954 4226
rect 16606 4174 16658 4226
rect 18958 4174 19010 4226
rect 19966 4174 20018 4226
rect 21198 4174 21250 4226
rect 24110 4174 24162 4226
rect 25118 4174 25170 4226
rect 26350 4174 26402 4226
rect 5742 4062 5794 4114
rect 11230 4062 11282 4114
rect 13134 4062 13186 4114
rect 14478 4062 14530 4114
rect 18622 4062 18674 4114
rect 25454 4062 25506 4114
rect 4466 3894 4518 3946
rect 4570 3894 4622 3946
rect 4674 3894 4726 3946
rect 24466 3894 24518 3946
rect 24570 3894 24622 3946
rect 24674 3894 24726 3946
rect 1038 3726 1090 3778
rect 1374 3726 1426 3778
rect 1710 3726 1762 3778
rect 2046 3726 2098 3778
rect 2718 3726 2770 3778
rect 5406 3726 5458 3778
rect 7310 3726 7362 3778
rect 7646 3726 7698 3778
rect 9774 3726 9826 3778
rect 10894 3726 10946 3778
rect 13582 3726 13634 3778
rect 15822 3726 15874 3778
rect 17054 3726 17106 3778
rect 18734 3726 18786 3778
rect 21422 3726 21474 3778
rect 22542 3726 22594 3778
rect 23550 3726 23602 3778
rect 24558 3726 24610 3778
rect 24894 3726 24946 3778
rect 25566 3726 25618 3778
rect 2382 3614 2434 3666
rect 4958 3614 5010 3666
rect 25230 3670 25282 3722
rect 26238 3726 26290 3778
rect 26574 3726 26626 3778
rect 6414 3614 6466 3666
rect 8318 3614 8370 3666
rect 15486 3614 15538 3666
rect 17726 3614 17778 3666
rect 23886 3614 23938 3666
rect 25902 3614 25954 3666
rect 3390 3502 3442 3554
rect 4174 3502 4226 3554
rect 5630 3502 5682 3554
rect 6078 3502 6130 3554
rect 8094 3502 8146 3554
rect 11454 3507 11506 3559
rect 12350 3502 12402 3554
rect 12910 3502 12962 3554
rect 13694 3502 13746 3554
rect 14254 3502 14306 3554
rect 14590 3502 14642 3554
rect 15150 3502 15202 3554
rect 16046 3502 16098 3554
rect 16830 3502 16882 3554
rect 18174 3502 18226 3554
rect 18510 3502 18562 3554
rect 19182 3502 19234 3554
rect 19966 3502 20018 3554
rect 20750 3502 20802 3554
rect 26798 3502 26850 3554
rect 9326 3390 9378 3442
rect 22990 3390 23042 3442
rect 3806 3110 3858 3162
rect 3910 3110 3962 3162
rect 4014 3110 4066 3162
rect 23806 3110 23858 3162
rect 23910 3110 23962 3162
rect 24014 3110 24066 3162
rect 3390 2942 3442 2994
rect 6862 2942 6914 2994
rect 15262 2942 15314 2994
rect 18174 2942 18226 2994
rect 20750 2942 20802 2994
rect 22990 2942 23042 2994
rect 10894 2830 10946 2882
rect 11230 2830 11282 2882
rect 13694 2830 13746 2882
rect 16606 2830 16658 2882
rect 24558 2830 24610 2882
rect 1710 2718 1762 2770
rect 3838 2718 3890 2770
rect 5294 2718 5346 2770
rect 7758 2718 7810 2770
rect 8654 2718 8706 2770
rect 9438 2718 9490 2770
rect 10110 2718 10162 2770
rect 10558 2718 10610 2770
rect 12014 2718 12066 2770
rect 13022 2718 13074 2770
rect 15710 2718 15762 2770
rect 18622 2718 18674 2770
rect 19630 2718 19682 2770
rect 22318 2718 22370 2770
rect 25454 2718 25506 2770
rect 26126 2718 26178 2770
rect 26686 2718 26738 2770
rect 27358 2718 27410 2770
rect 2158 2606 2210 2658
rect 4174 2606 4226 2658
rect 5742 2606 5794 2658
rect 9886 2606 9938 2658
rect 12798 2606 12850 2658
rect 14030 2606 14082 2658
rect 16046 2606 16098 2658
rect 17054 2606 17106 2658
rect 18958 2606 19010 2658
rect 11566 2494 11618 2546
rect 12238 2494 12290 2546
rect 19294 2494 19346 2546
rect 21870 2494 21922 2546
rect 24110 2494 24162 2546
rect 25118 2494 25170 2546
rect 25790 2494 25842 2546
rect 26462 2494 26514 2546
rect 27134 2494 27186 2546
rect 4466 2326 4518 2378
rect 4570 2326 4622 2378
rect 4674 2326 4726 2378
rect 24466 2326 24518 2378
rect 24570 2326 24622 2378
rect 24674 2326 24726 2378
rect 1150 2158 1202 2210
rect 1486 2158 1538 2210
rect 1822 2158 1874 2210
rect 2494 2158 2546 2210
rect 4958 2158 5010 2210
rect 6078 2158 6130 2210
rect 7198 2158 7250 2210
rect 7982 2158 8034 2210
rect 8318 2158 8370 2210
rect 9214 2158 9266 2210
rect 11678 2158 11730 2210
rect 13918 2158 13970 2210
rect 15038 2158 15090 2210
rect 15374 2158 15426 2210
rect 15710 2158 15762 2210
rect 18174 2158 18226 2210
rect 19294 2158 19346 2210
rect 20414 2158 20466 2210
rect 21534 2158 21586 2210
rect 22094 2158 22146 2210
rect 24670 2158 24722 2210
rect 27806 2158 27858 2210
rect 28478 2158 28530 2210
rect 2158 2046 2210 2098
rect 3838 2046 3890 2098
rect 7646 2046 7698 2098
rect 9550 2046 9602 2098
rect 10446 2046 10498 2098
rect 12798 2046 12850 2098
rect 14702 2046 14754 2098
rect 16046 2046 16098 2098
rect 16830 2046 16882 2098
rect 17166 2046 17218 2098
rect 23214 2046 23266 2098
rect 25902 2046 25954 2098
rect 26798 2046 26850 2098
rect 27470 2046 27522 2098
rect 28142 2046 28194 2098
rect 2718 1934 2770 1986
rect 3390 1934 3442 1986
rect 5630 1934 5682 1986
rect 12350 1934 12402 1986
rect 14366 1934 14418 1986
rect 17614 1934 17666 1986
rect 19854 1934 19906 1986
rect 23662 1934 23714 1986
rect 27022 1934 27074 1986
rect 10110 1822 10162 1874
rect 26238 1822 26290 1874
rect 3806 1542 3858 1594
rect 3910 1542 3962 1594
rect 4014 1542 4066 1594
rect 23806 1542 23858 1594
rect 23910 1542 23962 1594
rect 24014 1542 24066 1594
rect 3390 1374 3442 1426
rect 7982 1374 8034 1426
rect 11790 1374 11842 1426
rect 14254 1374 14306 1426
rect 19406 1374 19458 1426
rect 20190 1374 20242 1426
rect 23998 1374 24050 1426
rect 1822 1262 1874 1314
rect 6414 1262 6466 1314
rect 17838 1262 17890 1314
rect 25566 1262 25618 1314
rect 3838 1150 3890 1202
rect 5630 1150 5682 1202
rect 9326 1150 9378 1202
rect 10222 1150 10274 1202
rect 12686 1150 12738 1202
rect 14814 1150 14866 1202
rect 15486 1150 15538 1202
rect 21758 1150 21810 1202
rect 22542 1150 22594 1202
rect 23326 1150 23378 1202
rect 26350 1150 26402 1202
rect 28030 1150 28082 1202
rect 28590 1150 28642 1202
rect 29262 1150 29314 1202
rect 2270 1038 2322 1090
rect 4174 1038 4226 1090
rect 4846 1038 4898 1090
rect 6862 1038 6914 1090
rect 10670 1038 10722 1090
rect 18174 1038 18226 1090
rect 21422 1038 21474 1090
rect 25230 1038 25282 1090
rect 26126 1038 26178 1090
rect 27694 1038 27746 1090
rect 28366 1038 28418 1090
rect 5182 926 5234 978
rect 5854 926 5906 978
rect 9550 926 9602 978
rect 13134 926 13186 978
rect 15038 926 15090 978
rect 15710 926 15762 978
rect 16606 926 16658 978
rect 16942 926 16994 978
rect 22318 926 22370 978
rect 22990 926 23042 978
rect 26798 926 26850 978
rect 27134 926 27186 978
rect 29038 926 29090 978
rect 4466 758 4518 810
rect 4570 758 4622 810
rect 4674 758 4726 810
rect 24466 758 24518 810
rect 24570 758 24622 810
rect 24674 758 24726 810
<< metal2 >>
rect 5376 114800 5488 114912
rect 5600 114800 5712 114912
rect 5824 114800 5936 114912
rect 6048 114800 6160 114912
rect 6272 114800 6384 114912
rect 6496 114800 6608 114912
rect 6720 114800 6832 114912
rect 6944 114800 7056 114912
rect 7168 114800 7280 114912
rect 7392 114800 7504 114912
rect 7616 114800 7728 114912
rect 7840 114800 7952 114912
rect 8064 114800 8176 114912
rect 8288 114800 8400 114912
rect 8512 114800 8624 114912
rect 8736 114800 8848 114912
rect 8960 114800 9072 114912
rect 9184 114800 9296 114912
rect 9408 114800 9520 114912
rect 9632 114800 9744 114912
rect 9856 114800 9968 114912
rect 10080 114800 10192 114912
rect 10304 114800 10416 114912
rect 10528 114800 10640 114912
rect 10752 114800 10864 114912
rect 10976 114800 11088 114912
rect 11200 114800 11312 114912
rect 11424 114800 11536 114912
rect 11648 114800 11760 114912
rect 11872 114800 11984 114912
rect 12096 114800 12208 114912
rect 12320 114800 12432 114912
rect 12544 114800 12656 114912
rect 12768 114800 12880 114912
rect 12992 114800 13104 114912
rect 13216 114800 13328 114912
rect 13440 114800 13552 114912
rect 13664 114800 13776 114912
rect 13888 114800 14000 114912
rect 14112 114800 14224 114912
rect 14336 114800 14448 114912
rect 14560 114800 14672 114912
rect 14784 114800 14896 114912
rect 15008 114800 15120 114912
rect 15232 114800 15344 114912
rect 15456 114800 15568 114912
rect 15680 114800 15792 114912
rect 15904 114800 16016 114912
rect 16128 114800 16240 114912
rect 16352 114800 16464 114912
rect 16576 114800 16688 114912
rect 16800 114800 16912 114912
rect 17024 114800 17136 114912
rect 17248 114800 17360 114912
rect 17472 114800 17584 114912
rect 17696 114800 17808 114912
rect 17920 114800 18032 114912
rect 18144 114800 18256 114912
rect 18368 114800 18480 114912
rect 18592 114800 18704 114912
rect 18816 114800 18928 114912
rect 19040 114800 19152 114912
rect 19264 114800 19376 114912
rect 19488 114800 19600 114912
rect 19712 114800 19824 114912
rect 19936 114800 20048 114912
rect 20160 114800 20272 114912
rect 20384 114800 20496 114912
rect 20608 114800 20720 114912
rect 20832 114800 20944 114912
rect 21056 114800 21168 114912
rect 21280 114800 21392 114912
rect 21504 114800 21616 114912
rect 21728 114800 21840 114912
rect 21952 114800 22064 114912
rect 22176 114800 22288 114912
rect 22400 114800 22512 114912
rect 22624 114800 22736 114912
rect 22848 114800 22960 114912
rect 23072 114800 23184 114912
rect 23296 114800 23408 114912
rect 23520 114800 23632 114912
rect 23744 114800 23856 114912
rect 23968 114800 24080 114912
rect 24192 114800 24304 114912
rect 24416 114800 24528 114912
rect 24640 114800 24752 114912
rect 24864 114800 24976 114912
rect 25088 114800 25200 114912
rect 25312 114800 25424 114912
rect 25536 114800 25648 114912
rect 25760 114800 25872 114912
rect 25984 114800 26096 114912
rect 140 114212 196 114222
rect 140 96516 196 114156
rect 4844 114212 4900 114222
rect 1932 113988 1988 113998
rect 812 113764 868 113774
rect 588 111972 644 111982
rect 588 110964 644 111916
rect 588 109228 644 110908
rect 812 111860 868 113708
rect 1484 113540 1540 113550
rect 1484 113446 1540 113484
rect 1260 113316 1316 113326
rect 1260 113222 1316 113260
rect 1484 113204 1540 113214
rect 1484 112418 1540 113148
rect 1484 112366 1486 112418
rect 1538 112366 1540 112418
rect 1484 112354 1540 112366
rect 588 109172 756 109228
rect 476 108388 532 108398
rect 364 106260 420 106270
rect 140 96450 196 96460
rect 252 99988 308 99998
rect 140 85764 196 85774
rect 140 76580 196 85708
rect 252 83748 308 99932
rect 252 83682 308 83692
rect 364 83300 420 106204
rect 476 97860 532 108332
rect 476 92820 532 97804
rect 476 92754 532 92764
rect 588 100548 644 100558
rect 588 90692 644 100492
rect 700 98532 756 109172
rect 812 102228 868 111804
rect 1148 112306 1204 112318
rect 1148 112254 1150 112306
rect 1202 112254 1204 112306
rect 1148 109508 1204 112254
rect 1820 112308 1876 112318
rect 1820 112214 1876 112252
rect 1708 112196 1764 112206
rect 1596 111860 1652 111870
rect 1596 111766 1652 111804
rect 1260 111636 1316 111646
rect 1260 111542 1316 111580
rect 1484 111524 1540 111534
rect 1148 109442 1204 109452
rect 1260 110962 1316 110974
rect 1260 110910 1262 110962
rect 1314 110910 1316 110962
rect 1260 109506 1316 110910
rect 1484 110852 1540 111468
rect 1260 109454 1262 109506
rect 1314 109454 1316 109506
rect 1260 109228 1316 109454
rect 924 109172 1316 109228
rect 1372 110178 1428 110190
rect 1372 110126 1374 110178
rect 1426 110126 1428 110178
rect 924 104916 980 109172
rect 1260 108610 1316 108622
rect 1260 108558 1262 108610
rect 1314 108558 1316 108610
rect 1260 108052 1316 108558
rect 1260 107986 1316 107996
rect 1260 107826 1316 107838
rect 1260 107774 1262 107826
rect 1314 107774 1316 107826
rect 1260 107492 1316 107774
rect 924 104850 980 104860
rect 1036 107436 1316 107492
rect 1036 103236 1092 107436
rect 1148 107268 1204 107278
rect 1372 107268 1428 110126
rect 1484 109620 1540 110796
rect 1596 110964 1652 110974
rect 1596 110850 1652 110908
rect 1596 110798 1598 110850
rect 1650 110798 1652 110850
rect 1596 110786 1652 110798
rect 1708 110628 1764 112140
rect 1596 110572 1764 110628
rect 1596 110180 1652 110572
rect 1932 110516 1988 113932
rect 4464 113708 4728 113718
rect 4520 113652 4568 113708
rect 4624 113652 4672 113708
rect 4464 113642 4728 113652
rect 4844 113538 4900 114156
rect 5404 113876 5460 114800
rect 5404 113810 5460 113820
rect 4844 113486 4846 113538
rect 4898 113486 4900 113538
rect 4844 113474 4900 113486
rect 5180 113652 5236 113662
rect 5180 113538 5236 113596
rect 5180 113486 5182 113538
rect 5234 113486 5236 113538
rect 5180 113474 5236 113486
rect 2940 113426 2996 113438
rect 2940 113374 2942 113426
rect 2994 113374 2996 113426
rect 2604 113204 2660 113214
rect 2604 113202 2772 113204
rect 2604 113150 2606 113202
rect 2658 113150 2772 113202
rect 2604 113148 2772 113150
rect 2604 113138 2660 113148
rect 2716 112530 2772 113148
rect 2716 112478 2718 112530
rect 2770 112478 2772 112530
rect 2156 112308 2212 112318
rect 2156 112306 2436 112308
rect 2156 112254 2158 112306
rect 2210 112254 2436 112306
rect 2156 112252 2436 112254
rect 2156 112242 2212 112252
rect 1708 110460 1988 110516
rect 1708 110402 1764 110460
rect 1708 110350 1710 110402
rect 1762 110350 1764 110402
rect 1708 110338 1764 110350
rect 1596 110124 1764 110180
rect 1484 109564 1652 109620
rect 1596 109282 1652 109564
rect 1596 109230 1598 109282
rect 1650 109230 1652 109282
rect 1596 109218 1652 109230
rect 1148 107266 1428 107268
rect 1148 107214 1150 107266
rect 1202 107214 1428 107266
rect 1148 107212 1428 107214
rect 1596 107380 1652 107390
rect 1148 107202 1204 107212
rect 1484 107042 1540 107054
rect 1484 106990 1486 107042
rect 1538 106990 1540 107042
rect 1372 106596 1428 106606
rect 1260 106260 1316 106270
rect 1260 106166 1316 106204
rect 1260 105476 1316 105486
rect 1036 103170 1092 103180
rect 1148 105474 1316 105476
rect 1148 105422 1262 105474
rect 1314 105422 1316 105474
rect 1148 105420 1316 105422
rect 812 102162 868 102172
rect 1036 102900 1092 102910
rect 700 98466 756 98476
rect 1036 101220 1092 102844
rect 1148 102340 1204 105420
rect 1260 105410 1316 105420
rect 1148 102274 1204 102284
rect 1260 104916 1316 104926
rect 1260 104802 1316 104860
rect 1260 104750 1262 104802
rect 1314 104750 1316 104802
rect 1260 103234 1316 104750
rect 1372 104580 1428 106540
rect 1372 104514 1428 104524
rect 1372 103908 1428 103918
rect 1372 103814 1428 103852
rect 1260 103182 1262 103234
rect 1314 103182 1316 103234
rect 1260 102338 1316 103182
rect 1260 102286 1262 102338
rect 1314 102286 1316 102338
rect 1036 97468 1092 101164
rect 1260 100772 1316 102286
rect 1260 100706 1316 100716
rect 1372 101554 1428 101566
rect 1372 101502 1374 101554
rect 1426 101502 1428 101554
rect 1260 100548 1316 100558
rect 1260 100454 1316 100492
rect 1260 99988 1316 99998
rect 1372 99988 1428 101502
rect 1316 99932 1428 99988
rect 1260 99894 1316 99932
rect 1372 98868 1428 98878
rect 588 90626 644 90636
rect 700 97412 1092 97468
rect 1148 97634 1204 97646
rect 1148 97582 1150 97634
rect 1202 97582 1204 97634
rect 364 83234 420 83244
rect 588 90356 644 90366
rect 588 80052 644 90300
rect 700 86772 756 97412
rect 1036 95170 1092 95182
rect 1036 95118 1038 95170
rect 1090 95118 1092 95170
rect 1036 93042 1092 95118
rect 1036 92990 1038 93042
rect 1090 92990 1092 93042
rect 1036 92708 1092 92990
rect 1036 92642 1092 92652
rect 1148 92148 1204 97582
rect 1260 96292 1316 96302
rect 1260 94612 1316 96236
rect 1260 93714 1316 94556
rect 1260 93662 1262 93714
rect 1314 93662 1316 93714
rect 1260 93650 1316 93662
rect 1372 95954 1428 98812
rect 1372 95902 1374 95954
rect 1426 95902 1428 95954
rect 1036 92092 1204 92148
rect 812 91252 868 91262
rect 812 86996 868 91196
rect 1036 89012 1092 92092
rect 1372 92036 1428 95902
rect 1484 95844 1540 106990
rect 1596 106596 1652 107324
rect 1596 106530 1652 106540
rect 1708 106036 1764 110124
rect 2268 110066 2324 110078
rect 2268 110014 2270 110066
rect 2322 110014 2324 110066
rect 1820 109732 1876 109742
rect 1820 109228 1876 109676
rect 1820 109172 2100 109228
rect 1932 107044 1988 107054
rect 1820 107042 1988 107044
rect 1820 106990 1934 107042
rect 1986 106990 1988 107042
rect 1820 106988 1988 106990
rect 1820 106260 1876 106988
rect 1932 106978 1988 106988
rect 1820 106194 1876 106204
rect 1932 106372 1988 106382
rect 1932 106036 1988 106316
rect 1708 105980 1988 106036
rect 1596 105586 1652 105598
rect 1596 105534 1598 105586
rect 1650 105534 1652 105586
rect 1596 104692 1652 105534
rect 1596 104626 1652 104636
rect 1708 104580 1764 104590
rect 1708 104486 1764 104524
rect 1596 104020 1652 104030
rect 1596 103926 1652 103964
rect 1596 103010 1652 103022
rect 1596 102958 1598 103010
rect 1650 102958 1652 103010
rect 1596 102788 1652 102958
rect 1596 102722 1652 102732
rect 1708 102452 1764 102462
rect 1820 102452 1876 105980
rect 2044 105476 2100 109172
rect 2268 109060 2324 110014
rect 2268 108994 2324 109004
rect 2380 108836 2436 112252
rect 2716 111636 2772 112478
rect 2716 111570 2772 111580
rect 2828 111522 2884 111534
rect 2828 111470 2830 111522
rect 2882 111470 2884 111522
rect 2828 110964 2884 111470
rect 2828 110898 2884 110908
rect 2828 110740 2884 110750
rect 2156 108780 2436 108836
rect 2492 110738 2884 110740
rect 2492 110686 2830 110738
rect 2882 110686 2884 110738
rect 2492 110684 2884 110686
rect 2156 106484 2212 108780
rect 2268 108610 2324 108622
rect 2268 108558 2270 108610
rect 2322 108558 2324 108610
rect 2268 107716 2324 108558
rect 2268 107650 2324 107660
rect 2380 107826 2436 107838
rect 2380 107774 2382 107826
rect 2434 107774 2436 107826
rect 2380 106932 2436 107774
rect 2380 106866 2436 106876
rect 2156 106418 2212 106428
rect 2380 106484 2436 106494
rect 2156 106260 2212 106270
rect 2156 106166 2212 106204
rect 2156 105924 2212 105934
rect 2156 105812 2324 105868
rect 2044 105410 2100 105420
rect 2156 105362 2212 105374
rect 2156 105310 2158 105362
rect 2210 105310 2212 105362
rect 2156 104132 2212 105310
rect 2044 104076 2156 104132
rect 1764 102396 1876 102452
rect 1932 103460 1988 103470
rect 1708 102358 1764 102396
rect 1932 99314 1988 103404
rect 1932 99262 1934 99314
rect 1986 99262 1988 99314
rect 1932 99250 1988 99262
rect 1596 99090 1652 99102
rect 1596 99038 1598 99090
rect 1650 99038 1652 99090
rect 1596 96852 1652 99038
rect 1820 98532 1876 98542
rect 2044 98532 2100 104076
rect 2156 104066 2212 104076
rect 2156 103796 2212 103806
rect 2268 103796 2324 105812
rect 2156 103794 2324 103796
rect 2156 103742 2158 103794
rect 2210 103742 2324 103794
rect 2156 103740 2324 103742
rect 2156 103730 2212 103740
rect 2156 101554 2212 101566
rect 2156 101502 2158 101554
rect 2210 101502 2212 101554
rect 2156 99986 2212 101502
rect 2156 99934 2158 99986
rect 2210 99934 2212 99986
rect 2156 99652 2212 99934
rect 2156 99586 2212 99596
rect 2268 98868 2324 103740
rect 2380 102900 2436 106428
rect 2380 102834 2436 102844
rect 2380 100996 2436 101006
rect 2380 100902 2436 100940
rect 2268 98802 2324 98812
rect 2380 100772 2436 100782
rect 2380 98644 2436 100716
rect 2380 98578 2436 98588
rect 1820 98530 2100 98532
rect 1820 98478 1822 98530
rect 1874 98478 2100 98530
rect 1820 98476 2100 98478
rect 1820 98466 1876 98476
rect 2380 98308 2436 98318
rect 2268 98196 2324 98206
rect 2156 98140 2268 98196
rect 1708 97860 1764 97870
rect 1708 97766 1764 97804
rect 2156 96964 2212 98140
rect 2268 98102 2324 98140
rect 2380 97636 2436 98252
rect 2156 96898 2212 96908
rect 2268 97580 2436 97636
rect 1596 96786 1652 96796
rect 2156 96404 2212 96414
rect 1708 96180 1764 96190
rect 1708 96086 1764 96124
rect 1484 95778 1540 95788
rect 1708 95956 1764 95966
rect 1484 95284 1540 95294
rect 1484 95190 1540 95228
rect 1484 94388 1540 94398
rect 1484 92930 1540 94332
rect 1484 92878 1486 92930
rect 1538 92878 1540 92930
rect 1484 92866 1540 92878
rect 1596 93044 1652 93054
rect 1372 91980 1540 92036
rect 1148 91924 1204 91934
rect 1148 91922 1428 91924
rect 1148 91870 1150 91922
rect 1202 91870 1428 91922
rect 1148 91868 1428 91870
rect 1148 91858 1204 91868
rect 1260 91252 1316 91262
rect 1260 91158 1316 91196
rect 1148 90356 1204 90394
rect 1148 90290 1204 90300
rect 1036 88946 1092 88956
rect 1148 90132 1204 90142
rect 1148 87220 1204 90076
rect 1148 87154 1204 87164
rect 1260 88114 1316 88126
rect 1260 88062 1262 88114
rect 1314 88062 1316 88114
rect 1260 86996 1316 88062
rect 812 86940 1316 86996
rect 700 86706 756 86716
rect 1036 85764 1092 85802
rect 1036 85698 1092 85708
rect 588 79986 644 79996
rect 700 85652 756 85662
rect 588 79828 644 79838
rect 588 77028 644 79772
rect 700 78932 756 85596
rect 1148 85428 1204 86940
rect 1260 86546 1316 86558
rect 1260 86494 1262 86546
rect 1314 86494 1316 86546
rect 1260 86324 1316 86494
rect 1372 86548 1428 91868
rect 1484 91252 1540 91980
rect 1484 91186 1540 91196
rect 1484 90692 1540 90702
rect 1484 89794 1540 90636
rect 1596 89906 1652 92988
rect 1708 91700 1764 95900
rect 1932 95732 1988 95742
rect 1932 95282 1988 95676
rect 1932 95230 1934 95282
rect 1986 95230 1988 95282
rect 1820 94724 1876 94734
rect 1820 94610 1876 94668
rect 1820 94558 1822 94610
rect 1874 94558 1876 94610
rect 1820 94546 1876 94558
rect 1932 94500 1988 95230
rect 1932 92930 1988 94444
rect 2044 95058 2100 95070
rect 2044 95006 2046 95058
rect 2098 95006 2100 95058
rect 2044 94276 2100 95006
rect 2156 94388 2212 96348
rect 2156 94322 2212 94332
rect 2268 94498 2324 97580
rect 2268 94446 2270 94498
rect 2322 94446 2324 94498
rect 2044 94210 2100 94220
rect 2156 94164 2212 94174
rect 2156 93714 2212 94108
rect 2156 93662 2158 93714
rect 2210 93662 2212 93714
rect 2044 93044 2100 93054
rect 2044 92950 2100 92988
rect 1932 92878 1934 92930
rect 1986 92878 1988 92930
rect 1932 92866 1988 92878
rect 2156 92036 2212 93662
rect 2268 93492 2324 94446
rect 2492 95282 2548 110684
rect 2828 110674 2884 110684
rect 2716 110290 2772 110302
rect 2716 110238 2718 110290
rect 2770 110238 2772 110290
rect 2604 109060 2660 109070
rect 2604 105924 2660 109004
rect 2716 106484 2772 110238
rect 2940 109732 2996 113374
rect 3164 113428 3220 113438
rect 3164 112306 3220 113372
rect 5516 113428 5572 113438
rect 5516 113334 5572 113372
rect 3164 112254 3166 112306
rect 3218 112254 3220 112306
rect 3164 111524 3220 112254
rect 3164 111458 3220 111468
rect 3388 113316 3444 113326
rect 3388 111412 3444 113260
rect 4172 113090 4228 113102
rect 4172 113038 4174 113090
rect 4226 113038 4228 113090
rect 3804 112924 4068 112934
rect 3860 112868 3908 112924
rect 3964 112868 4012 112924
rect 3804 112858 4068 112868
rect 3836 111860 3892 111870
rect 3612 111858 3892 111860
rect 3612 111806 3838 111858
rect 3890 111806 3892 111858
rect 3612 111804 3892 111806
rect 3500 111636 3556 111646
rect 3500 111542 3556 111580
rect 3388 111356 3556 111412
rect 3388 110738 3444 110750
rect 3388 110686 3390 110738
rect 3442 110686 3444 110738
rect 3388 110404 3444 110686
rect 3388 110338 3444 110348
rect 3500 110180 3556 111356
rect 3388 110124 3556 110180
rect 2940 109666 2996 109676
rect 3276 109956 3332 109966
rect 2828 109172 2884 109182
rect 2828 109170 3108 109172
rect 2828 109118 2830 109170
rect 2882 109118 3108 109170
rect 2828 109116 3108 109118
rect 2828 109106 2884 109116
rect 2940 108610 2996 108622
rect 2940 108558 2942 108610
rect 2994 108558 2996 108610
rect 2940 108052 2996 108558
rect 2940 107826 2996 107996
rect 2940 107774 2942 107826
rect 2994 107774 2996 107826
rect 2940 107762 2996 107774
rect 2716 106418 2772 106428
rect 2828 107042 2884 107054
rect 2828 106990 2830 107042
rect 2882 106990 2884 107042
rect 2828 106260 2884 106990
rect 2828 106194 2884 106204
rect 2940 106484 2996 106494
rect 2940 106258 2996 106428
rect 2940 106206 2942 106258
rect 2994 106206 2996 106258
rect 2940 106194 2996 106206
rect 2604 105858 2660 105868
rect 2716 106148 2772 106158
rect 2604 105586 2660 105598
rect 2604 105534 2606 105586
rect 2658 105534 2660 105586
rect 2604 104244 2660 105534
rect 2716 105252 2772 106092
rect 2716 105186 2772 105196
rect 2604 104178 2660 104188
rect 2828 104466 2884 104478
rect 2828 104414 2830 104466
rect 2882 104414 2884 104466
rect 2604 104020 2660 104030
rect 2604 103926 2660 103964
rect 2828 103124 2884 104414
rect 2604 103068 2884 103124
rect 2604 98308 2660 103068
rect 2828 102900 2884 102910
rect 2716 102898 2884 102900
rect 2716 102846 2830 102898
rect 2882 102846 2884 102898
rect 2716 102844 2884 102846
rect 2716 99764 2772 102844
rect 2828 102834 2884 102844
rect 2940 102116 2996 102126
rect 2940 102022 2996 102060
rect 2940 101780 2996 101790
rect 2940 101554 2996 101724
rect 2940 101502 2942 101554
rect 2994 101502 2996 101554
rect 2940 101490 2996 101502
rect 2828 100772 2884 100782
rect 2828 100678 2884 100716
rect 2940 100212 2996 100222
rect 2940 99986 2996 100156
rect 2940 99934 2942 99986
rect 2994 99934 2996 99986
rect 2940 99922 2996 99934
rect 2716 99708 2996 99764
rect 2604 98242 2660 98252
rect 2828 99540 2884 99550
rect 2828 98196 2884 99484
rect 2828 98130 2884 98140
rect 2828 97412 2884 97422
rect 2492 95230 2494 95282
rect 2546 95230 2548 95282
rect 2492 94108 2548 95230
rect 2380 94052 2548 94108
rect 2604 97410 2884 97412
rect 2604 97358 2830 97410
rect 2882 97358 2884 97410
rect 2604 97356 2884 97358
rect 2380 93716 2436 94052
rect 2380 93650 2436 93660
rect 2268 93436 2548 93492
rect 2492 93042 2548 93436
rect 2492 92990 2494 93042
rect 2546 92990 2548 93042
rect 2492 92978 2548 92990
rect 2604 92820 2660 97356
rect 2828 97346 2884 97356
rect 2716 96852 2772 96862
rect 2716 95956 2772 96796
rect 2940 96404 2996 99708
rect 2940 96338 2996 96348
rect 3052 96068 3108 109116
rect 3276 108836 3332 109900
rect 3388 109282 3444 110124
rect 3612 110068 3668 111804
rect 3836 111794 3892 111804
rect 3804 111356 4068 111366
rect 3860 111300 3908 111356
rect 3964 111300 4012 111356
rect 3804 111290 4068 111300
rect 3724 111076 3780 111086
rect 3724 110850 3780 111020
rect 3724 110798 3726 110850
rect 3778 110798 3780 110850
rect 3724 110786 3780 110798
rect 4060 110740 4116 110750
rect 4060 110646 4116 110684
rect 3948 110516 4004 110526
rect 3948 110180 4004 110460
rect 3948 110114 4004 110124
rect 3500 110012 3668 110068
rect 3500 109396 3556 110012
rect 3836 109956 3892 109966
rect 3500 109330 3556 109340
rect 3612 109954 3892 109956
rect 3612 109902 3838 109954
rect 3890 109902 3892 109954
rect 3612 109900 3892 109902
rect 3388 109230 3390 109282
rect 3442 109230 3444 109282
rect 3388 109218 3444 109230
rect 3388 108836 3444 108846
rect 3276 108834 3444 108836
rect 3276 108782 3390 108834
rect 3442 108782 3444 108834
rect 3276 108780 3444 108782
rect 3388 108770 3444 108780
rect 3612 108724 3668 109900
rect 3836 109890 3892 109900
rect 3804 109788 4068 109798
rect 3860 109732 3908 109788
rect 3964 109732 4012 109788
rect 3804 109722 4068 109732
rect 4172 109620 4228 113038
rect 4956 112644 5012 112654
rect 4844 112420 4900 112430
rect 4284 112306 4340 112318
rect 4284 112254 4286 112306
rect 4338 112254 4340 112306
rect 4284 111188 4340 112254
rect 4464 112140 4728 112150
rect 4520 112084 4568 112140
rect 4624 112084 4672 112140
rect 4464 112074 4728 112084
rect 4284 111122 4340 111132
rect 4396 111972 4452 111982
rect 4396 110850 4452 111916
rect 4844 111076 4900 112364
rect 4844 111010 4900 111020
rect 4396 110798 4398 110850
rect 4450 110798 4452 110850
rect 4396 110786 4452 110798
rect 4844 110740 4900 110750
rect 4464 110572 4728 110582
rect 4284 110516 4340 110526
rect 4520 110516 4568 110572
rect 4624 110516 4672 110572
rect 4464 110506 4728 110516
rect 4284 109844 4340 110460
rect 4284 109778 4340 109788
rect 4396 110292 4452 110302
rect 4060 109564 4228 109620
rect 3836 109396 3892 109406
rect 3724 109284 3780 109322
rect 3724 109218 3780 109228
rect 3612 108658 3668 108668
rect 3276 108612 3332 108622
rect 3500 108612 3556 108622
rect 3276 107716 3332 108556
rect 3388 108610 3556 108612
rect 3388 108558 3502 108610
rect 3554 108558 3556 108610
rect 3388 108556 3556 108558
rect 3388 108388 3444 108556
rect 3500 108546 3556 108556
rect 3836 108500 3892 109340
rect 3948 108948 4004 108958
rect 3948 108612 4004 108892
rect 4060 108836 4116 109564
rect 4172 109394 4228 109406
rect 4172 109342 4174 109394
rect 4226 109342 4228 109394
rect 4172 109060 4228 109342
rect 4396 109282 4452 110236
rect 4620 110290 4676 110302
rect 4620 110238 4622 110290
rect 4674 110238 4676 110290
rect 4620 109620 4676 110238
rect 4620 109554 4676 109564
rect 4396 109230 4398 109282
rect 4450 109230 4452 109282
rect 4396 109218 4452 109230
rect 4172 108994 4228 109004
rect 4464 109004 4728 109014
rect 4520 108948 4568 109004
rect 4624 108948 4672 109004
rect 4464 108938 4728 108948
rect 4844 108948 4900 110684
rect 4956 110290 5012 112588
rect 5516 112532 5572 112542
rect 5068 112308 5124 112318
rect 5068 112214 5124 112252
rect 5404 112306 5460 112318
rect 5404 112254 5406 112306
rect 5458 112254 5460 112306
rect 5068 111860 5124 111870
rect 5068 111766 5124 111804
rect 5404 111412 5460 112254
rect 5516 111748 5572 112476
rect 5628 112084 5684 114800
rect 5852 113876 5908 114800
rect 5852 113810 5908 113820
rect 5852 113428 5908 113438
rect 5852 113334 5908 113372
rect 6076 113316 6132 114800
rect 6300 113988 6356 114800
rect 6300 113922 6356 113932
rect 6076 113250 6132 113260
rect 6300 113314 6356 113326
rect 6300 113262 6302 113314
rect 6354 113262 6356 113314
rect 6076 112868 6132 112878
rect 6076 112418 6132 112812
rect 6300 112532 6356 113262
rect 6300 112466 6356 112476
rect 6076 112366 6078 112418
rect 6130 112366 6132 112418
rect 6076 112354 6132 112366
rect 5740 112308 5796 112318
rect 5740 112214 5796 112252
rect 6524 112084 6580 114800
rect 6748 113764 6804 114800
rect 6972 114100 7028 114800
rect 6972 114044 7140 114100
rect 6748 113708 7028 113764
rect 6860 113426 6916 113438
rect 6860 113374 6862 113426
rect 6914 113374 6916 113426
rect 5628 112028 5908 112084
rect 5628 111748 5684 111758
rect 5516 111746 5684 111748
rect 5516 111694 5630 111746
rect 5682 111694 5684 111746
rect 5516 111692 5684 111694
rect 5628 111682 5684 111692
rect 5404 111346 5460 111356
rect 5516 110964 5572 110974
rect 5516 110870 5572 110908
rect 5740 110738 5796 110750
rect 5740 110686 5742 110738
rect 5794 110686 5796 110738
rect 4956 110238 4958 110290
rect 5010 110238 5012 110290
rect 4956 110226 5012 110238
rect 5404 110628 5460 110638
rect 5292 109956 5348 109966
rect 5292 109862 5348 109900
rect 5404 109844 5460 110572
rect 5628 110068 5684 110078
rect 5628 109974 5684 110012
rect 5740 109956 5796 110686
rect 5740 109890 5796 109900
rect 5404 109778 5460 109788
rect 5404 109508 5460 109518
rect 4844 108882 4900 108892
rect 4956 109396 5012 109406
rect 4060 108770 4116 108780
rect 4844 108724 4900 108734
rect 3948 108610 4228 108612
rect 3948 108558 3950 108610
rect 4002 108558 4228 108610
rect 3948 108556 4228 108558
rect 3948 108546 4004 108556
rect 3388 108322 3444 108332
rect 3612 108444 3892 108500
rect 3500 108052 3556 108062
rect 3500 107828 3556 107996
rect 3500 107762 3556 107772
rect 3612 107826 3668 108444
rect 3804 108220 4068 108230
rect 3860 108164 3908 108220
rect 3964 108164 4012 108220
rect 3804 108154 4068 108164
rect 3612 107774 3614 107826
rect 3666 107774 3668 107826
rect 3612 107762 3668 107774
rect 4060 107828 4116 107838
rect 4172 107828 4228 108556
rect 4396 108500 4452 108510
rect 4620 108500 4676 108510
rect 4396 108498 4620 108500
rect 4396 108446 4398 108498
rect 4450 108446 4620 108498
rect 4396 108444 4620 108446
rect 4396 108434 4452 108444
rect 4620 108434 4676 108444
rect 4732 108498 4788 108510
rect 4732 108446 4734 108498
rect 4786 108446 4788 108498
rect 4732 108276 4788 108446
rect 4732 108210 4788 108220
rect 4060 107826 4228 107828
rect 4060 107774 4062 107826
rect 4114 107774 4228 107826
rect 4060 107772 4228 107774
rect 4060 107762 4116 107772
rect 3388 107716 3444 107726
rect 3276 107714 3444 107716
rect 3276 107662 3390 107714
rect 3442 107662 3444 107714
rect 3276 107660 3444 107662
rect 3388 107650 3444 107660
rect 4396 107714 4452 107726
rect 4396 107662 4398 107714
rect 4450 107662 4452 107714
rect 4396 107604 4452 107662
rect 4396 107538 4452 107548
rect 4464 107436 4728 107446
rect 4520 107380 4568 107436
rect 4624 107380 4672 107436
rect 3612 107324 4228 107380
rect 4464 107370 4728 107380
rect 3500 107156 3556 107166
rect 3388 107042 3444 107054
rect 3388 106990 3390 107042
rect 3442 106990 3444 107042
rect 3388 106820 3444 106990
rect 3388 106754 3444 106764
rect 3276 106036 3332 106046
rect 3388 106036 3444 106046
rect 3332 106034 3444 106036
rect 3332 105982 3390 106034
rect 3442 105982 3444 106034
rect 3332 105980 3444 105982
rect 3276 105970 3332 105980
rect 3388 105970 3444 105980
rect 3164 105252 3220 105262
rect 3164 99540 3220 105196
rect 3276 104636 3444 104692
rect 3276 104244 3332 104636
rect 3388 104468 3444 104636
rect 3500 104690 3556 107100
rect 3612 107044 3668 107324
rect 3612 106260 3668 106988
rect 4060 107154 4116 107166
rect 4060 107102 4062 107154
rect 4114 107102 4116 107154
rect 4060 106820 4116 107102
rect 4172 107042 4228 107324
rect 4172 106990 4174 107042
rect 4226 106990 4228 107042
rect 4172 106978 4228 106990
rect 4732 107044 4788 107054
rect 4732 106950 4788 106988
rect 4620 106932 4676 106942
rect 4060 106764 4228 106820
rect 3804 106652 4068 106662
rect 3860 106596 3908 106652
rect 3964 106596 4012 106652
rect 3804 106586 4068 106596
rect 4172 106484 4228 106764
rect 3612 106166 3668 106204
rect 3724 106428 4228 106484
rect 3724 105476 3780 106428
rect 4508 106372 4564 106382
rect 4060 106316 4508 106372
rect 4060 106258 4116 106316
rect 4508 106306 4564 106316
rect 4060 106206 4062 106258
rect 4114 106206 4116 106258
rect 4060 106194 4116 106206
rect 4396 106148 4452 106158
rect 4620 106148 4676 106876
rect 4396 106146 4676 106148
rect 4396 106094 4398 106146
rect 4450 106094 4676 106146
rect 4396 106092 4676 106094
rect 4172 106036 4228 106046
rect 4060 105812 4116 105822
rect 3500 104638 3502 104690
rect 3554 104638 3556 104690
rect 3500 104626 3556 104638
rect 3612 105420 3780 105476
rect 3836 105476 3892 105486
rect 3612 104468 3668 105420
rect 3724 105252 3780 105262
rect 3836 105252 3892 105420
rect 4060 105476 4116 105756
rect 4060 105410 4116 105420
rect 3724 105250 3892 105252
rect 3724 105198 3726 105250
rect 3778 105198 3892 105250
rect 3724 105196 3892 105198
rect 3724 105186 3780 105196
rect 4172 105140 4228 105980
rect 4396 106036 4452 106092
rect 4396 105970 4452 105980
rect 4284 105924 4340 105934
rect 4284 105588 4340 105868
rect 4464 105868 4728 105878
rect 4520 105812 4568 105868
rect 4624 105812 4672 105868
rect 4464 105802 4728 105812
rect 4732 105588 4788 105598
rect 4284 105532 4676 105588
rect 4396 105364 4452 105374
rect 4396 105362 4564 105364
rect 4396 105310 4398 105362
rect 4450 105310 4564 105362
rect 4396 105308 4564 105310
rect 4396 105298 4452 105308
rect 4508 105252 4564 105308
rect 4508 105186 4564 105196
rect 3804 105084 4068 105094
rect 4172 105084 4452 105140
rect 3860 105028 3908 105084
rect 3964 105028 4012 105084
rect 3804 105018 4068 105028
rect 4060 104804 4116 104814
rect 3724 104580 3780 104590
rect 3724 104486 3780 104524
rect 4060 104578 4116 104748
rect 4284 104692 4340 104702
rect 4060 104526 4062 104578
rect 4114 104526 4116 104578
rect 4060 104514 4116 104526
rect 4172 104690 4340 104692
rect 4172 104638 4286 104690
rect 4338 104638 4340 104690
rect 4172 104636 4340 104638
rect 3388 104412 3668 104468
rect 4172 104468 4228 104636
rect 4284 104626 4340 104636
rect 4396 104468 4452 105084
rect 4620 104804 4676 105532
rect 4732 105494 4788 105532
rect 4620 104738 4676 104748
rect 4172 104402 4228 104412
rect 4284 104412 4452 104468
rect 3276 104188 3444 104244
rect 3388 103122 3444 104188
rect 4172 104132 4228 104142
rect 3724 103684 3780 103694
rect 3388 103070 3390 103122
rect 3442 103070 3444 103122
rect 3388 103058 3444 103070
rect 3612 103682 3780 103684
rect 3612 103630 3726 103682
rect 3778 103630 3780 103682
rect 3612 103628 3780 103630
rect 3276 102452 3332 102462
rect 3276 101444 3332 102396
rect 3500 101554 3556 101566
rect 3500 101502 3502 101554
rect 3554 101502 3556 101554
rect 3388 101444 3444 101454
rect 3276 101442 3444 101444
rect 3276 101390 3390 101442
rect 3442 101390 3444 101442
rect 3276 101388 3444 101390
rect 3388 101378 3444 101388
rect 3500 99988 3556 101502
rect 3612 100548 3668 103628
rect 3724 103618 3780 103628
rect 3804 103516 4068 103526
rect 3860 103460 3908 103516
rect 3964 103460 4012 103516
rect 3804 103450 4068 103460
rect 3724 103348 3780 103358
rect 3724 103010 3780 103292
rect 3948 103236 4004 103246
rect 3724 102958 3726 103010
rect 3778 102958 3780 103010
rect 3724 102946 3780 102958
rect 3836 103124 3892 103134
rect 3836 102788 3892 103068
rect 3836 102722 3892 102732
rect 3948 102338 4004 103180
rect 4060 102898 4116 102910
rect 4060 102846 4062 102898
rect 4114 102846 4116 102898
rect 4060 102788 4116 102846
rect 4060 102722 4116 102732
rect 3948 102286 3950 102338
rect 4002 102286 4004 102338
rect 3948 102274 4004 102286
rect 3804 101948 4068 101958
rect 3860 101892 3908 101948
rect 3964 101892 4012 101948
rect 3804 101882 4068 101892
rect 4060 101554 4116 101566
rect 4060 101502 4062 101554
rect 4114 101502 4116 101554
rect 4060 100996 4116 101502
rect 4060 100930 4116 100940
rect 3836 100772 3892 100782
rect 3836 100678 3892 100716
rect 3612 100482 3668 100492
rect 3804 100380 4068 100390
rect 3860 100324 3908 100380
rect 3964 100324 4012 100380
rect 3804 100314 4068 100324
rect 4060 100100 4116 100110
rect 3612 99988 3668 99998
rect 3500 99986 3668 99988
rect 3500 99934 3614 99986
rect 3666 99934 3668 99986
rect 3500 99932 3668 99934
rect 3388 99764 3444 99774
rect 3164 99474 3220 99484
rect 3276 99762 3444 99764
rect 3276 99710 3390 99762
rect 3442 99710 3444 99762
rect 3276 99708 3444 99710
rect 3276 99316 3332 99708
rect 3388 99698 3444 99708
rect 3276 99250 3332 99260
rect 3164 99204 3220 99214
rect 3164 99110 3220 99148
rect 3500 99092 3556 99932
rect 3612 99652 3668 99932
rect 4060 99986 4116 100044
rect 4060 99934 4062 99986
rect 4114 99934 4116 99986
rect 4060 99922 4116 99934
rect 3612 99586 3668 99596
rect 3276 99036 3556 99092
rect 3836 99202 3892 99214
rect 3836 99150 3838 99202
rect 3890 99150 3892 99202
rect 3164 96626 3220 96638
rect 3164 96574 3166 96626
rect 3218 96574 3220 96626
rect 3164 96292 3220 96574
rect 3164 96226 3220 96236
rect 2716 95890 2772 95900
rect 2828 96012 3108 96068
rect 2828 95284 2884 96012
rect 2940 95844 2996 95854
rect 2940 95842 3220 95844
rect 2940 95790 2942 95842
rect 2994 95790 3220 95842
rect 2940 95788 3220 95790
rect 2940 95778 2996 95788
rect 2884 95228 2996 95284
rect 2828 95218 2884 95228
rect 2716 95172 2772 95182
rect 2716 94498 2772 95116
rect 2716 94446 2718 94498
rect 2770 94446 2772 94498
rect 2716 94434 2772 94446
rect 2828 94610 2884 94622
rect 2828 94558 2830 94610
rect 2882 94558 2884 94610
rect 2380 92764 2660 92820
rect 1932 91980 2212 92036
rect 2268 92148 2324 92158
rect 2380 92148 2436 92764
rect 2380 92092 2548 92148
rect 2268 92034 2324 92092
rect 2268 91982 2270 92034
rect 2322 91982 2324 92034
rect 1708 91644 1876 91700
rect 1708 91474 1764 91486
rect 1708 91422 1710 91474
rect 1762 91422 1764 91474
rect 1708 90132 1764 91422
rect 1708 90066 1764 90076
rect 1596 89854 1598 89906
rect 1650 89854 1652 89906
rect 1596 89842 1652 89854
rect 1484 89742 1486 89794
rect 1538 89742 1540 89794
rect 1484 89730 1540 89742
rect 1708 88452 1764 88462
rect 1820 88452 1876 91644
rect 1932 88676 1988 91980
rect 2268 91970 2324 91982
rect 2380 91476 2436 91486
rect 2268 90356 2324 90366
rect 2156 90354 2324 90356
rect 2156 90302 2270 90354
rect 2322 90302 2324 90354
rect 2156 90300 2324 90302
rect 1932 88620 2100 88676
rect 1708 88450 1876 88452
rect 1708 88398 1710 88450
rect 1762 88398 1876 88450
rect 1708 88396 1876 88398
rect 1708 87108 1764 88396
rect 1820 87556 1876 87566
rect 1820 87462 1876 87500
rect 1708 87042 1764 87052
rect 1372 86482 1428 86492
rect 1484 86772 1540 86782
rect 1260 86258 1316 86268
rect 924 85372 1204 85428
rect 1260 85874 1316 85886
rect 1260 85822 1262 85874
rect 1314 85822 1316 85874
rect 700 78866 756 78876
rect 812 80948 868 80958
rect 588 76962 644 76972
rect 140 76514 196 76524
rect 252 76804 308 76814
rect 252 75684 308 76748
rect 140 75628 308 75684
rect 28 75460 84 75470
rect 28 68068 84 75404
rect 140 69412 196 75628
rect 812 75236 868 80892
rect 924 80836 980 85372
rect 1036 85202 1092 85214
rect 1036 85150 1038 85202
rect 1090 85150 1092 85202
rect 1036 83748 1092 85150
rect 1148 84980 1204 84990
rect 1148 84194 1204 84924
rect 1148 84142 1150 84194
rect 1202 84142 1204 84194
rect 1148 84084 1204 84142
rect 1148 84018 1204 84028
rect 1260 83748 1316 85822
rect 1484 85652 1540 86716
rect 1596 86772 1652 86810
rect 1596 86706 1652 86716
rect 1484 85586 1540 85596
rect 1596 86548 1652 86558
rect 1484 85428 1540 85438
rect 1372 85090 1428 85102
rect 1372 85038 1374 85090
rect 1426 85038 1428 85090
rect 1372 84756 1428 85038
rect 1372 84690 1428 84700
rect 1484 84306 1540 85372
rect 1484 84254 1486 84306
rect 1538 84254 1540 84306
rect 1484 84242 1540 84254
rect 1484 84084 1540 84094
rect 1372 83748 1428 83758
rect 1036 83692 1204 83748
rect 1260 83746 1428 83748
rect 1260 83694 1374 83746
rect 1426 83694 1428 83746
rect 1260 83692 1428 83694
rect 924 80770 980 80780
rect 1036 83522 1092 83534
rect 1036 83470 1038 83522
rect 1090 83470 1092 83522
rect 1036 80276 1092 83470
rect 1148 82852 1204 83692
rect 1372 83682 1428 83692
rect 1148 82796 1428 82852
rect 1148 82626 1204 82638
rect 1148 82574 1150 82626
rect 1202 82574 1204 82626
rect 1148 82068 1204 82574
rect 1148 82002 1204 82012
rect 1036 80210 1092 80220
rect 1260 79602 1316 79614
rect 1260 79550 1262 79602
rect 1314 79550 1316 79602
rect 1260 79492 1316 79550
rect 1260 79426 1316 79436
rect 924 79156 980 79166
rect 924 76692 980 79100
rect 1148 78594 1204 78606
rect 1148 78542 1150 78594
rect 1202 78542 1204 78594
rect 1036 77362 1092 77374
rect 1036 77310 1038 77362
rect 1090 77310 1092 77362
rect 1036 76804 1092 77310
rect 1036 76738 1092 76748
rect 924 76626 980 76636
rect 1036 76244 1092 76254
rect 924 76242 1092 76244
rect 924 76190 1038 76242
rect 1090 76190 1092 76242
rect 924 76188 1092 76190
rect 924 75460 980 76188
rect 1036 76178 1092 76188
rect 924 75394 980 75404
rect 1036 75794 1092 75806
rect 1036 75742 1038 75794
rect 1090 75742 1092 75794
rect 812 75170 868 75180
rect 1036 74900 1092 75742
rect 588 74844 1092 74900
rect 140 69346 196 69356
rect 252 74228 308 74238
rect 140 68068 196 68078
rect 28 68012 140 68068
rect 140 68002 196 68012
rect 140 67844 196 67854
rect 140 63140 196 67788
rect 252 66724 308 74172
rect 252 66658 308 66668
rect 364 68404 420 68414
rect 140 63074 196 63084
rect 252 66052 308 66062
rect 252 55468 308 65996
rect 364 62692 420 68348
rect 364 62626 420 62636
rect 476 67956 532 67966
rect 476 62244 532 67900
rect 588 67172 644 74844
rect 1036 74228 1092 74238
rect 1036 74134 1092 74172
rect 1036 72658 1092 72670
rect 1036 72606 1038 72658
rect 1090 72606 1092 72658
rect 1036 71764 1092 72606
rect 1148 72436 1204 78542
rect 1260 78148 1316 78158
rect 1260 78054 1316 78092
rect 1372 77476 1428 82796
rect 1484 82068 1540 84028
rect 1596 82738 1652 86492
rect 1932 86324 1988 86334
rect 1820 85652 1876 85662
rect 1596 82686 1598 82738
rect 1650 82686 1652 82738
rect 1596 82674 1652 82686
rect 1708 85650 1876 85652
rect 1708 85598 1822 85650
rect 1874 85598 1876 85650
rect 1708 85596 1876 85598
rect 1708 82740 1764 85596
rect 1820 85586 1876 85596
rect 1820 84980 1876 84990
rect 1820 84886 1876 84924
rect 1932 84756 1988 86268
rect 2044 85428 2100 88620
rect 2156 87332 2212 90300
rect 2268 90290 2324 90300
rect 2268 89796 2324 89806
rect 2380 89796 2436 91420
rect 2268 89794 2436 89796
rect 2268 89742 2270 89794
rect 2322 89742 2436 89794
rect 2268 89740 2436 89742
rect 2268 89730 2324 89740
rect 2156 87238 2212 87276
rect 2268 89236 2324 89246
rect 2044 85362 2100 85372
rect 2156 85650 2212 85662
rect 2156 85598 2158 85650
rect 2210 85598 2212 85650
rect 1820 84700 1988 84756
rect 2044 85092 2100 85102
rect 1820 83748 1876 84700
rect 1820 83522 1876 83692
rect 1820 83470 1822 83522
rect 1874 83470 1876 83522
rect 1820 83458 1876 83470
rect 2044 84306 2100 85036
rect 2044 84254 2046 84306
rect 2098 84254 2100 84306
rect 1932 83412 1988 83422
rect 1932 82740 1988 83356
rect 1708 82674 1764 82684
rect 1820 82738 1988 82740
rect 1820 82686 1934 82738
rect 1986 82686 1988 82738
rect 1820 82684 1988 82686
rect 1484 80274 1540 82012
rect 1484 80222 1486 80274
rect 1538 80222 1540 80274
rect 1484 79044 1540 80222
rect 1484 78978 1540 78988
rect 1596 82292 1652 82302
rect 1260 77420 1428 77476
rect 1260 75684 1316 77420
rect 1372 77252 1428 77262
rect 1372 77250 1540 77252
rect 1372 77198 1374 77250
rect 1426 77198 1540 77250
rect 1372 77196 1540 77198
rect 1372 77186 1428 77196
rect 1372 76244 1428 76254
rect 1372 76150 1428 76188
rect 1484 75908 1540 77196
rect 1484 75842 1540 75852
rect 1260 75618 1316 75628
rect 1372 75684 1428 75694
rect 1372 75682 1540 75684
rect 1372 75630 1374 75682
rect 1426 75630 1540 75682
rect 1372 75628 1540 75630
rect 1372 75618 1428 75628
rect 1260 75460 1316 75470
rect 1260 74004 1316 75404
rect 1372 74116 1428 74126
rect 1372 74022 1428 74060
rect 1260 73938 1316 73948
rect 1148 72370 1204 72380
rect 1372 72546 1428 72558
rect 1372 72494 1374 72546
rect 1426 72494 1428 72546
rect 1260 71764 1316 71774
rect 588 67106 644 67116
rect 700 71708 1092 71764
rect 1148 71762 1316 71764
rect 1148 71710 1262 71762
rect 1314 71710 1316 71762
rect 1148 71708 1316 71710
rect 476 62178 532 62188
rect 588 66836 644 66846
rect 588 62020 644 66780
rect 700 65828 756 71708
rect 1036 71538 1092 71550
rect 1036 71486 1038 71538
rect 1090 71486 1092 71538
rect 1036 70756 1092 71486
rect 700 65762 756 65772
rect 812 70700 1092 70756
rect 812 64036 868 70700
rect 924 70532 980 70542
rect 924 66948 980 70476
rect 1036 69522 1092 69534
rect 1036 69470 1038 69522
rect 1090 69470 1092 69522
rect 1036 68628 1092 69470
rect 1036 68562 1092 68572
rect 1036 68404 1092 68414
rect 1036 68310 1092 68348
rect 1036 67956 1092 67966
rect 1036 67862 1092 67900
rect 1148 67284 1204 71708
rect 1260 71698 1316 71708
rect 1260 71540 1316 71550
rect 1260 70644 1316 71484
rect 1372 70756 1428 72494
rect 1484 71092 1540 75628
rect 1484 71026 1540 71036
rect 1372 70690 1428 70700
rect 1484 70866 1540 70878
rect 1484 70814 1486 70866
rect 1538 70814 1540 70866
rect 1260 70578 1316 70588
rect 1484 70644 1540 70814
rect 1484 70578 1540 70588
rect 1260 70420 1316 70430
rect 1260 70194 1316 70364
rect 1260 70142 1262 70194
rect 1314 70142 1316 70194
rect 1260 69300 1316 70142
rect 1372 69412 1428 69422
rect 1372 69318 1428 69356
rect 1260 69234 1316 69244
rect 1596 68628 1652 82236
rect 1708 81842 1764 81854
rect 1708 81790 1710 81842
rect 1762 81790 1764 81842
rect 1708 81170 1764 81790
rect 1708 81118 1710 81170
rect 1762 81118 1764 81170
rect 1708 79604 1764 81118
rect 1820 79716 1876 82684
rect 1932 82674 1988 82684
rect 2044 82404 2100 84254
rect 2156 84308 2212 85598
rect 2268 85316 2324 89180
rect 2268 85250 2324 85260
rect 2380 85428 2436 85438
rect 2268 85090 2324 85102
rect 2268 85038 2270 85090
rect 2322 85038 2324 85090
rect 2268 84980 2324 85038
rect 2268 84914 2324 84924
rect 2156 84252 2324 84308
rect 2156 84084 2212 84094
rect 2156 83990 2212 84028
rect 1932 82348 2100 82404
rect 2156 82514 2212 82526
rect 2156 82462 2158 82514
rect 2210 82462 2212 82514
rect 1932 80836 1988 82348
rect 2156 82292 2212 82462
rect 2268 82516 2324 84252
rect 2380 83860 2436 85372
rect 2492 84980 2548 92092
rect 2716 92146 2772 92158
rect 2716 92094 2718 92146
rect 2770 92094 2772 92146
rect 2716 91140 2772 92094
rect 2828 91476 2884 94558
rect 2940 93714 2996 95228
rect 2940 93662 2942 93714
rect 2994 93662 2996 93714
rect 2940 93650 2996 93662
rect 3052 95282 3108 95294
rect 3052 95230 3054 95282
rect 3106 95230 3108 95282
rect 2828 91410 2884 91420
rect 3052 92930 3108 95230
rect 3052 92878 3054 92930
rect 3106 92878 3108 92930
rect 2716 90690 2772 91084
rect 2828 91140 2884 91150
rect 3052 91140 3108 92878
rect 2828 91138 2996 91140
rect 2828 91086 2830 91138
rect 2882 91086 2996 91138
rect 2828 91084 2996 91086
rect 2828 91074 2884 91084
rect 2716 90638 2718 90690
rect 2770 90638 2772 90690
rect 2716 90626 2772 90638
rect 2716 90132 2772 90142
rect 2604 89572 2660 89582
rect 2604 89478 2660 89516
rect 2716 89236 2772 90076
rect 2716 89170 2772 89180
rect 2604 89012 2660 89022
rect 2604 88918 2660 88956
rect 2940 88452 2996 91084
rect 3052 91074 3108 91084
rect 3164 90804 3220 95788
rect 3276 93828 3332 99036
rect 3836 98980 3892 99150
rect 3836 98914 3892 98924
rect 3804 98812 4068 98822
rect 3860 98756 3908 98812
rect 3964 98756 4012 98812
rect 3804 98746 4068 98756
rect 4172 98532 4228 104076
rect 4284 100772 4340 104412
rect 4464 104300 4728 104310
rect 4520 104244 4568 104300
rect 4624 104244 4672 104300
rect 4464 104234 4728 104244
rect 4844 104244 4900 108668
rect 4844 104178 4900 104188
rect 4732 104018 4788 104030
rect 4732 103966 4734 104018
rect 4786 103966 4788 104018
rect 4396 103796 4452 103806
rect 4396 103702 4452 103740
rect 4396 103012 4452 103022
rect 4396 102918 4452 102956
rect 4732 102900 4788 103966
rect 4732 102834 4788 102844
rect 4464 102732 4728 102742
rect 4520 102676 4568 102732
rect 4624 102676 4672 102732
rect 4464 102666 4728 102676
rect 4844 102338 4900 102350
rect 4844 102286 4846 102338
rect 4898 102286 4900 102338
rect 4396 101444 4452 101454
rect 4396 101350 4452 101388
rect 4844 101444 4900 102286
rect 4464 101164 4728 101174
rect 4520 101108 4568 101164
rect 4624 101108 4672 101164
rect 4464 101098 4728 101108
rect 4732 100772 4788 100782
rect 4284 100770 4788 100772
rect 4284 100718 4734 100770
rect 4786 100718 4788 100770
rect 4284 100716 4788 100718
rect 4396 99876 4452 99886
rect 4284 99874 4452 99876
rect 4284 99822 4398 99874
rect 4450 99822 4452 99874
rect 4284 99820 4452 99822
rect 4284 99428 4340 99820
rect 4396 99810 4452 99820
rect 4732 99876 4788 100716
rect 4732 99810 4788 99820
rect 4464 99596 4728 99606
rect 4520 99540 4568 99596
rect 4624 99540 4672 99596
rect 4464 99530 4728 99540
rect 4284 99362 4340 99372
rect 4396 99316 4452 99326
rect 4396 99222 4452 99260
rect 4060 98476 4228 98532
rect 4284 98980 4340 98990
rect 3388 98194 3444 98206
rect 3388 98142 3390 98194
rect 3442 98142 3444 98194
rect 3388 94724 3444 98142
rect 4060 98084 4116 98476
rect 4172 98308 4228 98318
rect 4172 98214 4228 98252
rect 4284 98306 4340 98924
rect 4284 98254 4286 98306
rect 4338 98254 4340 98306
rect 4284 98242 4340 98254
rect 4396 98756 4452 98766
rect 4396 98308 4452 98700
rect 4732 98420 4788 98430
rect 4844 98420 4900 101388
rect 4788 98364 4900 98420
rect 4732 98354 4788 98364
rect 4396 98242 4452 98252
rect 4956 98308 5012 109340
rect 5404 109282 5460 109452
rect 5404 109230 5406 109282
rect 5458 109230 5460 109282
rect 5404 109218 5460 109230
rect 5740 109284 5796 109322
rect 5740 109218 5796 109228
rect 5292 109172 5348 109182
rect 5068 108836 5124 108846
rect 5068 108610 5124 108780
rect 5068 108558 5070 108610
rect 5122 108558 5124 108610
rect 5068 108546 5124 108558
rect 5180 107828 5236 107838
rect 5180 107734 5236 107772
rect 5292 107716 5348 109116
rect 5740 108722 5796 108734
rect 5740 108670 5742 108722
rect 5794 108670 5796 108722
rect 5628 108612 5684 108622
rect 5628 108518 5684 108556
rect 5516 107940 5572 107950
rect 5404 107716 5460 107726
rect 5292 107714 5460 107716
rect 5292 107662 5406 107714
rect 5458 107662 5460 107714
rect 5292 107660 5460 107662
rect 5404 107650 5460 107660
rect 5404 107156 5460 107166
rect 5404 107062 5460 107100
rect 5068 106932 5124 106942
rect 5516 106932 5572 107884
rect 5740 107940 5796 108670
rect 5740 107874 5796 107884
rect 5852 107268 5908 112028
rect 5068 106930 5236 106932
rect 5068 106878 5070 106930
rect 5122 106878 5236 106930
rect 5068 106876 5236 106878
rect 5068 106866 5124 106876
rect 5068 104690 5124 104702
rect 5068 104638 5070 104690
rect 5122 104638 5124 104690
rect 5068 103348 5124 104638
rect 5068 103282 5124 103292
rect 5068 103122 5124 103134
rect 5068 103070 5070 103122
rect 5122 103070 5124 103122
rect 5068 102452 5124 103070
rect 5068 102386 5124 102396
rect 5180 102116 5236 106876
rect 5292 106876 5572 106932
rect 5628 107212 5908 107268
rect 5964 112028 6580 112084
rect 6636 113092 6692 113102
rect 5292 105252 5348 106876
rect 5516 106708 5572 106718
rect 5292 105186 5348 105196
rect 5404 106596 5460 106606
rect 5404 106370 5460 106540
rect 5404 106318 5406 106370
rect 5458 106318 5460 106370
rect 5292 105028 5348 105038
rect 5292 104578 5348 104972
rect 5292 104526 5294 104578
rect 5346 104526 5348 104578
rect 5292 104514 5348 104526
rect 5292 102900 5348 102910
rect 5292 102806 5348 102844
rect 5404 102564 5460 106318
rect 5516 106148 5572 106652
rect 5516 106082 5572 106092
rect 5404 102498 5460 102508
rect 5516 105252 5572 105262
rect 5404 102340 5460 102350
rect 5068 102060 5236 102116
rect 5292 102338 5460 102340
rect 5292 102286 5406 102338
rect 5458 102286 5460 102338
rect 5292 102284 5460 102286
rect 5068 98868 5124 102060
rect 5292 102004 5348 102284
rect 5404 102274 5460 102284
rect 5292 101938 5348 101948
rect 5180 101892 5236 101902
rect 5180 101554 5236 101836
rect 5180 101502 5182 101554
rect 5234 101502 5236 101554
rect 5180 101490 5236 101502
rect 5404 101444 5460 101454
rect 5404 101350 5460 101388
rect 5292 101332 5348 101342
rect 5292 100770 5348 101276
rect 5516 101220 5572 105196
rect 5628 103124 5684 107212
rect 5740 107042 5796 107054
rect 5740 106990 5742 107042
rect 5794 106990 5796 107042
rect 5740 105924 5796 106990
rect 5740 105858 5796 105868
rect 5852 106034 5908 106046
rect 5852 105982 5854 106034
rect 5906 105982 5908 106034
rect 5852 105588 5908 105982
rect 5740 105532 5908 105588
rect 5740 103572 5796 105532
rect 5964 105476 6020 112028
rect 6188 111858 6244 111870
rect 6188 111806 6190 111858
rect 6242 111806 6244 111858
rect 5740 103348 5796 103516
rect 5740 103282 5796 103292
rect 5852 105420 6020 105476
rect 6076 110850 6132 110862
rect 6076 110798 6078 110850
rect 6130 110798 6132 110850
rect 6076 109506 6132 110798
rect 6188 110516 6244 111806
rect 6636 111412 6692 113036
rect 6860 112532 6916 113374
rect 6860 112466 6916 112476
rect 6860 112308 6916 112318
rect 6188 110450 6244 110460
rect 6300 111356 6692 111412
rect 6748 112306 6916 112308
rect 6748 112254 6862 112306
rect 6914 112254 6916 112306
rect 6748 112252 6916 112254
rect 6300 110292 6356 111356
rect 6412 111188 6468 111198
rect 6412 110962 6468 111132
rect 6412 110910 6414 110962
rect 6466 110910 6468 110962
rect 6412 110898 6468 110910
rect 6748 110852 6804 112252
rect 6860 112242 6916 112252
rect 6524 110796 6804 110852
rect 6860 110964 6916 110974
rect 6076 109454 6078 109506
rect 6130 109454 6132 109506
rect 6076 108276 6132 109454
rect 6188 110236 6356 110292
rect 6412 110516 6468 110526
rect 6188 108722 6244 110236
rect 6412 110180 6468 110460
rect 6188 108670 6190 108722
rect 6242 108670 6244 108722
rect 6188 108658 6244 108670
rect 6300 110066 6356 110078
rect 6300 110014 6302 110066
rect 6354 110014 6356 110066
rect 6076 107492 6132 108220
rect 6300 108164 6356 110014
rect 6412 109228 6468 110124
rect 6524 109394 6580 110796
rect 6636 110516 6692 110526
rect 6636 110290 6692 110460
rect 6636 110238 6638 110290
rect 6690 110238 6692 110290
rect 6636 110226 6692 110238
rect 6524 109342 6526 109394
rect 6578 109342 6580 109394
rect 6524 109330 6580 109342
rect 6636 109956 6692 109966
rect 6412 109172 6580 109228
rect 6300 108098 6356 108108
rect 5628 103068 5796 103124
rect 5628 102900 5684 102910
rect 5628 102806 5684 102844
rect 5740 101444 5796 103068
rect 5852 103012 5908 105420
rect 5964 105250 6020 105262
rect 5964 105198 5966 105250
rect 6018 105198 6020 105250
rect 5964 104020 6020 105198
rect 6076 104802 6132 107436
rect 6300 107940 6356 107950
rect 6076 104750 6078 104802
rect 6130 104750 6132 104802
rect 6076 104244 6132 104750
rect 6076 104178 6132 104188
rect 6188 106818 6244 106830
rect 6188 106766 6190 106818
rect 6242 106766 6244 106818
rect 5964 103954 6020 103964
rect 5964 103684 6020 103694
rect 5964 103682 6132 103684
rect 5964 103630 5966 103682
rect 6018 103630 6132 103682
rect 5964 103628 6132 103630
rect 5964 103618 6020 103628
rect 5964 103012 6020 103022
rect 5852 103010 6020 103012
rect 5852 102958 5966 103010
rect 6018 102958 6020 103010
rect 5852 102956 6020 102958
rect 5964 102946 6020 102956
rect 6076 102676 6132 103628
rect 6188 103124 6244 106766
rect 6300 106596 6356 107884
rect 6300 106530 6356 106540
rect 6412 107604 6468 107614
rect 6412 104690 6468 107548
rect 6412 104638 6414 104690
rect 6466 104638 6468 104690
rect 6412 104626 6468 104638
rect 6412 104020 6468 104030
rect 6300 103348 6356 103358
rect 6300 103234 6356 103292
rect 6300 103182 6302 103234
rect 6354 103182 6356 103234
rect 6300 103170 6356 103182
rect 6188 103058 6244 103068
rect 5964 102620 6132 102676
rect 6412 102676 6468 103964
rect 5740 101378 5796 101388
rect 5852 102452 5908 102462
rect 5852 102228 5908 102396
rect 5852 101554 5908 102172
rect 5964 101780 6020 102620
rect 6412 102610 6468 102620
rect 6524 102508 6580 109172
rect 6636 105924 6692 109900
rect 6860 109394 6916 110908
rect 6860 109342 6862 109394
rect 6914 109342 6916 109394
rect 6748 108724 6804 108734
rect 6748 108610 6804 108668
rect 6748 108558 6750 108610
rect 6802 108558 6804 108610
rect 6748 108546 6804 108558
rect 6860 108612 6916 109342
rect 6748 107602 6804 107614
rect 6748 107550 6750 107602
rect 6802 107550 6804 107602
rect 6748 106708 6804 107550
rect 6748 106642 6804 106652
rect 6860 106372 6916 108556
rect 6636 105858 6692 105868
rect 6748 106316 6916 106372
rect 6636 105362 6692 105374
rect 6636 105310 6638 105362
rect 6690 105310 6692 105362
rect 6636 104020 6692 105310
rect 6748 104692 6804 106316
rect 6972 106260 7028 113708
rect 7084 113204 7140 114044
rect 7084 113138 7140 113148
rect 7196 112644 7252 114800
rect 7420 112980 7476 114800
rect 7420 112914 7476 112924
rect 7196 112578 7252 112588
rect 7644 112532 7700 114800
rect 7420 112476 7700 112532
rect 7308 111522 7364 111534
rect 7308 111470 7310 111522
rect 7362 111470 7364 111522
rect 7084 110740 7140 110750
rect 7084 110738 7252 110740
rect 7084 110686 7086 110738
rect 7138 110686 7252 110738
rect 7084 110684 7252 110686
rect 7084 110674 7140 110684
rect 7084 109396 7140 109406
rect 7084 109282 7140 109340
rect 7084 109230 7086 109282
rect 7138 109230 7140 109282
rect 7084 109218 7140 109230
rect 7084 108836 7140 108846
rect 7084 107940 7140 108780
rect 7196 108500 7252 110684
rect 7196 108434 7252 108444
rect 7084 107884 7252 107940
rect 6860 106204 7028 106260
rect 7084 107716 7140 107726
rect 6860 105028 6916 106204
rect 6972 106036 7028 106046
rect 6972 105942 7028 105980
rect 6972 105812 7028 105822
rect 6972 105588 7028 105756
rect 6972 105494 7028 105532
rect 6860 104962 6916 104972
rect 6972 104692 7028 104702
rect 6748 104690 7028 104692
rect 6748 104638 6974 104690
rect 7026 104638 7028 104690
rect 6748 104636 7028 104638
rect 6972 104580 7028 104636
rect 6972 104514 7028 104524
rect 7084 104578 7140 107660
rect 7196 107268 7252 107884
rect 7308 107604 7364 111470
rect 7308 107538 7364 107548
rect 7308 107268 7364 107278
rect 7196 107266 7364 107268
rect 7196 107214 7310 107266
rect 7362 107214 7364 107266
rect 7196 107212 7364 107214
rect 7196 106148 7252 107212
rect 7308 107156 7364 107212
rect 7308 107090 7364 107100
rect 7196 106082 7252 106092
rect 7308 106932 7364 106942
rect 7084 104526 7086 104578
rect 7138 104526 7140 104578
rect 7084 104244 7140 104526
rect 6972 104188 7140 104244
rect 7308 104356 7364 106876
rect 7420 104468 7476 112476
rect 7644 111860 7700 111870
rect 7532 111076 7588 111086
rect 7532 110962 7588 111020
rect 7532 110910 7534 110962
rect 7586 110910 7588 110962
rect 7532 110898 7588 110910
rect 7644 109394 7700 111804
rect 7756 111748 7812 111758
rect 7756 111654 7812 111692
rect 7868 111524 7924 114800
rect 8092 113540 8148 114800
rect 8092 113474 8148 113484
rect 7980 113092 8036 113102
rect 7980 112998 8036 113036
rect 8092 112756 8148 112766
rect 7980 112308 8036 112318
rect 7980 112214 8036 112252
rect 8092 111970 8148 112700
rect 8092 111918 8094 111970
rect 8146 111918 8148 111970
rect 8092 111906 8148 111918
rect 7644 109342 7646 109394
rect 7698 109342 7700 109394
rect 7644 109330 7700 109342
rect 7756 111468 7924 111524
rect 7980 111524 8036 111534
rect 7756 109228 7812 111468
rect 7980 110964 8036 111468
rect 7980 110898 8036 110908
rect 8092 110962 8148 110974
rect 8092 110910 8094 110962
rect 8146 110910 8148 110962
rect 7644 109172 7812 109228
rect 7868 109954 7924 109966
rect 7868 109902 7870 109954
rect 7922 109902 7924 109954
rect 7868 109228 7924 109902
rect 8092 109396 8148 110910
rect 8092 109302 8148 109340
rect 7868 109172 8036 109228
rect 7644 106596 7700 109172
rect 7868 108610 7924 108622
rect 7868 108558 7870 108610
rect 7922 108558 7924 108610
rect 7868 108500 7924 108558
rect 7868 108434 7924 108444
rect 7756 108164 7812 108174
rect 7756 106932 7812 108108
rect 7868 107716 7924 107726
rect 7868 107622 7924 107660
rect 7756 106838 7812 106876
rect 7644 106540 7924 106596
rect 7644 106260 7700 106270
rect 7644 106166 7700 106204
rect 7532 106036 7588 106046
rect 7532 104690 7588 105980
rect 7532 104638 7534 104690
rect 7586 104638 7588 104690
rect 7532 104626 7588 104638
rect 7420 104402 7476 104412
rect 6636 103964 6804 104020
rect 6636 103794 6692 103806
rect 6636 103742 6638 103794
rect 6690 103742 6692 103794
rect 6636 103684 6692 103742
rect 6748 103796 6804 103964
rect 6748 103730 6804 103740
rect 6636 103618 6692 103628
rect 6748 103124 6804 103134
rect 6748 103030 6804 103068
rect 6076 102450 6132 102462
rect 6076 102398 6078 102450
rect 6130 102398 6132 102450
rect 6076 102340 6132 102398
rect 6300 102452 6580 102508
rect 6972 102452 7028 104188
rect 7308 104132 7364 104300
rect 7308 104076 7476 104132
rect 7084 104020 7140 104030
rect 7084 103926 7140 103964
rect 7308 103908 7364 103918
rect 7196 103122 7252 103134
rect 7196 103070 7198 103122
rect 7250 103070 7252 103122
rect 7084 102452 7140 102462
rect 6076 102274 6132 102284
rect 6188 102338 6244 102350
rect 6188 102286 6190 102338
rect 6242 102286 6244 102338
rect 5964 101724 6132 101780
rect 5852 101502 5854 101554
rect 5906 101502 5908 101554
rect 5516 101154 5572 101164
rect 5292 100718 5294 100770
rect 5346 100718 5348 100770
rect 5292 100706 5348 100718
rect 5516 100548 5572 100558
rect 5180 100324 5236 100334
rect 5180 100098 5236 100268
rect 5180 100046 5182 100098
rect 5234 100046 5236 100098
rect 5180 100034 5236 100046
rect 5516 99204 5572 100492
rect 5628 100436 5684 100446
rect 5628 99874 5684 100380
rect 5628 99822 5630 99874
rect 5682 99822 5684 99874
rect 5628 99810 5684 99822
rect 5852 99652 5908 101502
rect 6076 101444 6132 101724
rect 6076 101378 6132 101388
rect 6076 101220 6132 101230
rect 5852 99586 5908 99596
rect 5964 100882 6020 100894
rect 5964 100830 5966 100882
rect 6018 100830 6020 100882
rect 5964 99204 6020 100830
rect 5516 99148 5684 99204
rect 5068 98802 5124 98812
rect 5180 98980 5236 98990
rect 5516 98980 5572 98990
rect 4956 98242 5012 98252
rect 4508 98196 4564 98206
rect 4508 98194 4900 98196
rect 4508 98142 4510 98194
rect 4562 98142 4900 98194
rect 4508 98140 4900 98142
rect 4508 98130 4564 98140
rect 4060 98028 4228 98084
rect 4060 97748 4116 97758
rect 4060 97654 4116 97692
rect 4172 97636 4228 98028
rect 4464 98028 4728 98038
rect 4520 97972 4568 98028
rect 4624 97972 4672 98028
rect 4464 97962 4728 97972
rect 4508 97860 4564 97870
rect 4844 97860 4900 98140
rect 4844 97804 5012 97860
rect 4396 97636 4452 97646
rect 4172 97634 4452 97636
rect 4172 97582 4398 97634
rect 4450 97582 4452 97634
rect 4172 97580 4452 97582
rect 3804 97244 4068 97254
rect 3860 97188 3908 97244
rect 3964 97188 4012 97244
rect 3804 97178 4068 97188
rect 3500 96964 3556 96974
rect 3500 95956 3556 96908
rect 4172 96066 4228 97580
rect 4396 97570 4452 97580
rect 4508 97524 4564 97804
rect 4508 97458 4564 97468
rect 4844 97634 4900 97646
rect 4844 97582 4846 97634
rect 4898 97582 4900 97634
rect 4844 97524 4900 97582
rect 4844 97458 4900 97468
rect 4172 96014 4174 96066
rect 4226 96014 4228 96066
rect 4172 96002 4228 96014
rect 4284 96626 4340 96638
rect 4284 96574 4286 96626
rect 4338 96574 4340 96626
rect 3724 95956 3780 95966
rect 3500 95890 3556 95900
rect 3612 95954 3780 95956
rect 3612 95902 3726 95954
rect 3778 95902 3780 95954
rect 3612 95900 3780 95902
rect 3612 95732 3668 95900
rect 3724 95890 3780 95900
rect 3612 95666 3668 95676
rect 3804 95676 4068 95686
rect 3860 95620 3908 95676
rect 3964 95620 4012 95676
rect 3804 95610 4068 95620
rect 4172 95284 4228 95294
rect 4060 95172 4116 95182
rect 3388 94668 3668 94724
rect 3388 94498 3444 94510
rect 3388 94446 3390 94498
rect 3442 94446 3444 94498
rect 3388 94388 3444 94446
rect 3388 94322 3444 94332
rect 3612 94052 3668 94668
rect 4060 94500 4116 95116
rect 4060 94406 4116 94444
rect 3804 94108 4068 94118
rect 3860 94052 3908 94108
rect 3964 94052 4012 94108
rect 3804 94042 4068 94052
rect 3612 93986 3668 93996
rect 3276 93762 3332 93772
rect 3500 93828 3556 93838
rect 3500 93714 3556 93772
rect 3500 93662 3502 93714
rect 3554 93662 3556 93714
rect 3500 93650 3556 93662
rect 3948 93716 4004 93726
rect 3948 93622 4004 93660
rect 3388 93490 3444 93502
rect 3388 93438 3390 93490
rect 3442 93438 3444 93490
rect 3388 93380 3444 93438
rect 3276 93324 3444 93380
rect 3276 91028 3332 93324
rect 4172 92930 4228 95228
rect 4172 92878 4174 92930
rect 4226 92878 4228 92930
rect 3804 92540 4068 92550
rect 3860 92484 3908 92540
rect 3964 92484 4012 92540
rect 3804 92474 4068 92484
rect 3276 90962 3332 90972
rect 3388 91138 3444 91150
rect 3388 91086 3390 91138
rect 3442 91086 3444 91138
rect 3164 90748 3332 90804
rect 3164 90580 3220 90590
rect 3052 89682 3108 89694
rect 3052 89630 3054 89682
rect 3106 89630 3108 89682
rect 3052 89572 3108 89630
rect 3164 89684 3220 90524
rect 3164 89618 3220 89628
rect 3052 89506 3108 89516
rect 3164 89012 3220 89022
rect 3164 88898 3220 88956
rect 3164 88846 3166 88898
rect 3218 88846 3220 88898
rect 3164 88834 3220 88846
rect 2940 88396 3108 88452
rect 2828 88004 2884 88014
rect 2828 88002 2996 88004
rect 2828 87950 2830 88002
rect 2882 87950 2996 88002
rect 2828 87948 2996 87950
rect 2828 87938 2884 87948
rect 2716 87556 2772 87566
rect 2604 87220 2660 87230
rect 2604 86884 2660 87164
rect 2604 85652 2660 86828
rect 2716 86772 2772 87500
rect 2716 86212 2772 86716
rect 2716 85986 2772 86156
rect 2716 85934 2718 85986
rect 2770 85934 2772 85986
rect 2716 85922 2772 85934
rect 2828 86434 2884 86446
rect 2828 86382 2830 86434
rect 2882 86382 2884 86434
rect 2828 85708 2884 86382
rect 2604 85586 2660 85596
rect 2716 85652 2884 85708
rect 2604 85092 2660 85130
rect 2604 85026 2660 85036
rect 2492 84914 2548 84924
rect 2380 83804 2548 83860
rect 2380 83636 2436 83646
rect 2380 83542 2436 83580
rect 2268 82450 2324 82460
rect 2156 82226 2212 82236
rect 2044 82180 2100 82190
rect 2044 81058 2100 82124
rect 2156 82066 2212 82078
rect 2156 82014 2158 82066
rect 2210 82014 2212 82066
rect 2156 81844 2212 82014
rect 2156 81778 2212 81788
rect 2044 81006 2046 81058
rect 2098 81006 2100 81058
rect 2044 80994 2100 81006
rect 1932 80780 2100 80836
rect 1932 80386 1988 80398
rect 1932 80334 1934 80386
rect 1986 80334 1988 80386
rect 1932 80052 1988 80334
rect 2044 80388 2100 80780
rect 2492 80724 2548 83804
rect 2716 82628 2772 85652
rect 2828 85204 2884 85214
rect 2828 85110 2884 85148
rect 2828 84308 2884 84318
rect 2828 84214 2884 84252
rect 2828 82740 2884 82750
rect 2828 82646 2884 82684
rect 2044 80322 2100 80332
rect 2156 80668 2548 80724
rect 2604 82572 2772 82628
rect 1932 79986 1988 79996
rect 1820 79660 2100 79716
rect 1708 79548 1876 79604
rect 1820 79492 1876 79548
rect 1932 79492 1988 79502
rect 1820 79436 1932 79492
rect 1708 79378 1764 79390
rect 1708 79326 1710 79378
rect 1762 79326 1764 79378
rect 1708 78932 1764 79326
rect 1708 78596 1764 78876
rect 1708 77922 1764 78540
rect 1932 78260 1988 79436
rect 1708 77870 1710 77922
rect 1762 77870 1764 77922
rect 1708 77858 1764 77870
rect 1820 78148 1876 78158
rect 1708 77362 1764 77374
rect 1708 77310 1710 77362
rect 1762 77310 1764 77362
rect 1708 72660 1764 77310
rect 1820 75010 1876 78092
rect 1932 76578 1988 78204
rect 2044 77588 2100 79660
rect 2044 77522 2100 77532
rect 1932 76526 1934 76578
rect 1986 76526 1988 76578
rect 1932 76514 1988 76526
rect 2044 77250 2100 77262
rect 2044 77198 2046 77250
rect 2098 77198 2100 77250
rect 1820 74958 1822 75010
rect 1874 74958 1876 75010
rect 1820 73330 1876 74958
rect 1932 75796 1988 75806
rect 1932 74114 1988 75740
rect 1932 74062 1934 74114
rect 1986 74062 1988 74114
rect 1932 74050 1988 74062
rect 1820 73278 1822 73330
rect 1874 73278 1876 73330
rect 1820 72884 1876 73278
rect 2044 73220 2100 77198
rect 2156 77252 2212 80668
rect 2492 80500 2548 80510
rect 2492 80406 2548 80444
rect 2380 80388 2436 80398
rect 2380 80294 2436 80332
rect 2156 77186 2212 77196
rect 2268 80164 2324 80174
rect 2156 76580 2212 76590
rect 2156 75682 2212 76524
rect 2156 75630 2158 75682
rect 2210 75630 2212 75682
rect 2156 75572 2212 75630
rect 2268 75684 2324 80108
rect 2492 79380 2548 79390
rect 2380 78930 2436 78942
rect 2380 78878 2382 78930
rect 2434 78878 2436 78930
rect 2380 78708 2436 78878
rect 2380 78642 2436 78652
rect 2380 77252 2436 77262
rect 2380 77158 2436 77196
rect 2380 76356 2436 76366
rect 2380 76262 2436 76300
rect 2492 76020 2548 79324
rect 2604 77252 2660 82572
rect 2716 82292 2772 82302
rect 2716 78818 2772 82236
rect 2940 80498 2996 87948
rect 3052 82740 3108 88396
rect 3276 88340 3332 90748
rect 3164 88284 3332 88340
rect 3164 86884 3220 88284
rect 3276 88116 3332 88126
rect 3276 88022 3332 88060
rect 3388 87668 3444 91086
rect 3804 90972 4068 90982
rect 3860 90916 3908 90972
rect 3964 90916 4012 90972
rect 3804 90906 4068 90916
rect 4060 90356 4116 90366
rect 4060 90018 4116 90300
rect 4060 89966 4062 90018
rect 4114 89966 4116 90018
rect 4060 89954 4116 89966
rect 3500 89796 3556 89806
rect 3724 89796 3780 89806
rect 3500 89794 3724 89796
rect 3500 89742 3502 89794
rect 3554 89742 3724 89794
rect 3500 89740 3724 89742
rect 3500 89730 3556 89740
rect 3724 89730 3780 89740
rect 3836 89794 3892 89806
rect 3836 89742 3838 89794
rect 3890 89742 3892 89794
rect 3836 89572 3892 89742
rect 3612 89516 3892 89572
rect 3612 89236 3668 89516
rect 3804 89404 4068 89414
rect 3860 89348 3908 89404
rect 3964 89348 4012 89404
rect 3804 89338 4068 89348
rect 3612 89180 3780 89236
rect 3612 88228 3668 88238
rect 3612 88134 3668 88172
rect 3724 88116 3780 89180
rect 4172 89124 4228 92878
rect 4284 90020 4340 96574
rect 4464 96460 4728 96470
rect 4520 96404 4568 96460
rect 4624 96404 4672 96460
rect 4464 96394 4728 96404
rect 4956 96404 5012 97804
rect 4956 96338 5012 96348
rect 5068 97746 5124 97758
rect 5068 97694 5070 97746
rect 5122 97694 5124 97746
rect 4732 96180 4788 96190
rect 4732 96178 5012 96180
rect 4732 96126 4734 96178
rect 4786 96126 5012 96178
rect 4732 96124 5012 96126
rect 4732 96114 4788 96124
rect 4620 96066 4676 96078
rect 4620 96014 4622 96066
rect 4674 96014 4676 96066
rect 4620 95956 4676 96014
rect 4620 95172 4676 95900
rect 4620 95106 4676 95116
rect 4464 94892 4728 94902
rect 4520 94836 4568 94892
rect 4624 94836 4672 94892
rect 4464 94826 4728 94836
rect 4396 94724 4452 94734
rect 4396 93826 4452 94668
rect 4844 94612 4900 94622
rect 4844 94498 4900 94556
rect 4844 94446 4846 94498
rect 4898 94446 4900 94498
rect 4844 94164 4900 94446
rect 4844 94098 4900 94108
rect 4396 93774 4398 93826
rect 4450 93774 4452 93826
rect 4396 93762 4452 93774
rect 4464 93324 4728 93334
rect 4520 93268 4568 93324
rect 4624 93268 4672 93324
rect 4464 93258 4728 93268
rect 4956 93042 5012 96124
rect 4956 92990 4958 93042
rect 5010 92990 5012 93042
rect 4956 92978 5012 92990
rect 5068 92932 5124 97694
rect 5068 92866 5124 92876
rect 4956 92708 5012 92718
rect 4844 92484 4900 92494
rect 4464 91756 4728 91766
rect 4520 91700 4568 91756
rect 4624 91700 4672 91756
rect 4464 91690 4728 91700
rect 4620 91476 4676 91486
rect 4620 91382 4676 91420
rect 4464 90188 4728 90198
rect 4520 90132 4568 90188
rect 4624 90132 4672 90188
rect 4464 90122 4728 90132
rect 4284 89964 4564 90020
rect 4508 89906 4564 89964
rect 4508 89854 4510 89906
rect 4562 89854 4564 89906
rect 4508 89842 4564 89854
rect 4172 89058 4228 89068
rect 4284 88788 4340 88798
rect 4172 88786 4340 88788
rect 4172 88734 4286 88786
rect 4338 88734 4340 88786
rect 4172 88732 4340 88734
rect 3724 88050 3780 88060
rect 4060 88226 4116 88238
rect 4060 88174 4062 88226
rect 4114 88174 4116 88226
rect 4060 88116 4116 88174
rect 4060 88050 4116 88060
rect 3804 87836 4068 87846
rect 3860 87780 3908 87836
rect 3964 87780 4012 87836
rect 3804 87770 4068 87780
rect 3388 87602 3444 87612
rect 3388 87218 3444 87230
rect 3388 87166 3390 87218
rect 3442 87166 3444 87218
rect 3388 87108 3444 87166
rect 3388 87052 3668 87108
rect 3164 86828 3332 86884
rect 3164 85652 3220 85662
rect 3164 85558 3220 85596
rect 3164 84532 3220 84542
rect 3164 84306 3220 84476
rect 3164 84254 3166 84306
rect 3218 84254 3220 84306
rect 3164 84242 3220 84254
rect 3276 84308 3332 86828
rect 3500 85092 3556 85102
rect 3500 84998 3556 85036
rect 3276 84242 3332 84252
rect 3388 84306 3444 84318
rect 3388 84254 3390 84306
rect 3442 84254 3444 84306
rect 3052 82674 3108 82684
rect 3164 84084 3220 84094
rect 3164 82738 3220 84028
rect 3164 82686 3166 82738
rect 3218 82686 3220 82738
rect 2940 80446 2942 80498
rect 2994 80446 2996 80498
rect 2940 80434 2996 80446
rect 3052 81732 3108 81742
rect 2828 79380 2884 79390
rect 2828 79286 2884 79324
rect 2716 78766 2718 78818
rect 2770 78766 2772 78818
rect 2716 78148 2772 78766
rect 2716 78082 2772 78092
rect 2940 78708 2996 78718
rect 2828 77810 2884 77822
rect 2828 77758 2830 77810
rect 2882 77758 2884 77810
rect 2716 77252 2772 77262
rect 2604 77250 2772 77252
rect 2604 77198 2718 77250
rect 2770 77198 2772 77250
rect 2604 77196 2772 77198
rect 2716 77186 2772 77196
rect 2716 76916 2772 76926
rect 2268 75618 2324 75628
rect 2380 75964 2548 76020
rect 2604 76692 2660 76702
rect 2156 75506 2212 75516
rect 2268 74900 2324 74910
rect 2268 74786 2324 74844
rect 2268 74734 2270 74786
rect 2322 74734 2324 74786
rect 2268 74722 2324 74734
rect 2044 73154 2100 73164
rect 2156 74226 2212 74238
rect 2156 74174 2158 74226
rect 2210 74174 2212 74226
rect 1820 72818 1876 72828
rect 2044 72772 2100 72782
rect 1708 72604 1988 72660
rect 1820 72436 1876 72446
rect 1708 71538 1764 71550
rect 1708 71486 1710 71538
rect 1762 71486 1764 71538
rect 1708 70196 1764 71486
rect 1820 70978 1876 72380
rect 1820 70926 1822 70978
rect 1874 70926 1876 70978
rect 1820 70914 1876 70926
rect 1932 70868 1988 72604
rect 2044 72434 2100 72716
rect 2044 72382 2046 72434
rect 2098 72382 2100 72434
rect 2044 71876 2100 72382
rect 2156 72436 2212 74174
rect 2268 73556 2324 73566
rect 2268 73218 2324 73500
rect 2268 73166 2270 73218
rect 2322 73166 2324 73218
rect 2268 73154 2324 73166
rect 2156 72370 2212 72380
rect 2268 72660 2324 72670
rect 2044 71764 2100 71820
rect 2044 71708 2212 71764
rect 1932 70802 1988 70812
rect 2044 71538 2100 71550
rect 2044 71486 2046 71538
rect 2098 71486 2100 71538
rect 1708 70130 1764 70140
rect 1820 70644 1876 70654
rect 1708 69970 1764 69982
rect 1708 69918 1710 69970
rect 1762 69918 1764 69970
rect 1708 69636 1764 69918
rect 1708 69570 1764 69580
rect 1148 67218 1204 67228
rect 1260 68572 1652 68628
rect 1820 69300 1876 70588
rect 2044 70532 2100 71486
rect 2156 71540 2212 71708
rect 2156 71474 2212 71484
rect 2268 71316 2324 72604
rect 2380 72546 2436 75964
rect 2604 75682 2660 76636
rect 2604 75630 2606 75682
rect 2658 75630 2660 75682
rect 2604 75618 2660 75630
rect 2492 75572 2548 75582
rect 2492 72772 2548 75516
rect 2716 73948 2772 76860
rect 2492 72706 2548 72716
rect 2604 73892 2772 73948
rect 2380 72494 2382 72546
rect 2434 72494 2436 72546
rect 2380 72482 2436 72494
rect 2604 72548 2660 73892
rect 2828 72772 2884 77758
rect 2940 77140 2996 78652
rect 3052 77924 3108 81676
rect 3164 80164 3220 82686
rect 3276 81732 3332 81742
rect 3276 81638 3332 81676
rect 3388 81620 3444 84254
rect 3388 81554 3444 81564
rect 3500 83298 3556 83310
rect 3500 83246 3502 83298
rect 3554 83246 3556 83298
rect 3164 80098 3220 80108
rect 3276 80946 3332 80958
rect 3276 80894 3278 80946
rect 3330 80894 3332 80946
rect 3276 78036 3332 80894
rect 3388 79602 3444 79614
rect 3388 79550 3390 79602
rect 3442 79550 3444 79602
rect 3388 79380 3444 79550
rect 3388 79314 3444 79324
rect 3500 79044 3556 83246
rect 3612 82964 3668 87052
rect 4172 86996 4228 88732
rect 4284 88722 4340 88732
rect 4464 88620 4728 88630
rect 4520 88564 4568 88620
rect 4624 88564 4672 88620
rect 4464 88554 4728 88564
rect 4284 88338 4340 88350
rect 4284 88286 4286 88338
rect 4338 88286 4340 88338
rect 4284 87444 4340 88286
rect 4844 88226 4900 92428
rect 4956 91476 5012 92652
rect 5068 92372 5124 92382
rect 5180 92372 5236 98924
rect 5404 98978 5572 98980
rect 5404 98926 5518 98978
rect 5570 98926 5572 98978
rect 5404 98924 5572 98926
rect 5292 98644 5348 98654
rect 5292 98530 5348 98588
rect 5292 98478 5294 98530
rect 5346 98478 5348 98530
rect 5292 98420 5348 98478
rect 5292 98354 5348 98364
rect 5292 98196 5348 98206
rect 5292 96516 5348 98140
rect 5292 96450 5348 96460
rect 5404 96292 5460 98924
rect 5516 98914 5572 98924
rect 5628 97634 5684 99148
rect 5964 99138 6020 99148
rect 5740 98308 5796 98318
rect 5740 98214 5796 98252
rect 5628 97582 5630 97634
rect 5682 97582 5684 97634
rect 5516 96964 5572 96974
rect 5516 96870 5572 96908
rect 5628 96292 5684 97582
rect 6076 97524 6132 101164
rect 6188 100770 6244 102286
rect 6188 100718 6190 100770
rect 6242 100718 6244 100770
rect 6188 100548 6244 100718
rect 6188 100482 6244 100492
rect 6188 99652 6244 99662
rect 6188 99090 6244 99596
rect 6188 99038 6190 99090
rect 6242 99038 6244 99090
rect 6188 99026 6244 99038
rect 6188 97748 6244 97758
rect 6188 97634 6244 97692
rect 6188 97582 6190 97634
rect 6242 97582 6244 97634
rect 6188 97570 6244 97582
rect 5964 96626 6020 96638
rect 5964 96574 5966 96626
rect 6018 96574 6020 96626
rect 5292 96236 5460 96292
rect 5516 96236 5684 96292
rect 5740 96516 5796 96526
rect 5292 93042 5348 96236
rect 5404 96068 5460 96078
rect 5516 96068 5572 96236
rect 5404 96066 5572 96068
rect 5404 96014 5406 96066
rect 5458 96014 5572 96066
rect 5404 96012 5572 96014
rect 5740 96066 5796 96460
rect 5740 96014 5742 96066
rect 5794 96014 5796 96066
rect 5404 96002 5460 96012
rect 5516 95060 5572 95070
rect 5292 92990 5294 93042
rect 5346 92990 5348 93042
rect 5292 92978 5348 92990
rect 5404 95058 5572 95060
rect 5404 95006 5518 95058
rect 5570 95006 5572 95058
rect 5404 95004 5572 95006
rect 5068 92370 5236 92372
rect 5068 92318 5070 92370
rect 5122 92318 5236 92370
rect 5068 92316 5236 92318
rect 5292 92708 5348 92718
rect 5068 92306 5124 92316
rect 5292 92260 5348 92652
rect 5404 92484 5460 95004
rect 5516 94994 5572 95004
rect 5740 94724 5796 96014
rect 5740 94658 5796 94668
rect 5964 94724 6020 96574
rect 6076 95396 6132 97468
rect 6076 95330 6132 95340
rect 6300 94724 6356 102452
rect 6972 102450 7140 102452
rect 6972 102398 7086 102450
rect 7138 102398 7140 102450
rect 6972 102396 7140 102398
rect 6636 102338 6692 102350
rect 6636 102286 6638 102338
rect 6690 102286 6692 102338
rect 6412 101556 6468 101566
rect 6412 101332 6468 101500
rect 6412 101330 6580 101332
rect 6412 101278 6414 101330
rect 6466 101278 6580 101330
rect 6412 101276 6580 101278
rect 6412 101266 6468 101276
rect 6412 98868 6468 98878
rect 6412 97636 6468 98812
rect 6524 98084 6580 101276
rect 6636 101220 6692 102286
rect 6636 101154 6692 101164
rect 6972 100882 7028 102396
rect 7084 102386 7140 102396
rect 7196 102340 7252 103070
rect 7308 103010 7364 103852
rect 7308 102958 7310 103010
rect 7362 102958 7364 103010
rect 7308 102946 7364 102958
rect 7196 102274 7252 102284
rect 7420 101444 7476 104076
rect 7868 102452 7924 106540
rect 7980 103122 8036 109172
rect 8316 109172 8372 114800
rect 8540 113764 8596 114800
rect 8540 113698 8596 113708
rect 8316 109106 8372 109116
rect 8428 112530 8484 112542
rect 8428 112478 8430 112530
rect 8482 112478 8484 112530
rect 8428 111636 8484 112478
rect 8316 108498 8372 108510
rect 8316 108446 8318 108498
rect 8370 108446 8372 108498
rect 8316 107602 8372 108446
rect 8316 107550 8318 107602
rect 8370 107550 8372 107602
rect 8316 106932 8372 107550
rect 8316 106838 8372 106876
rect 8428 106260 8484 111580
rect 8540 112308 8596 112318
rect 8540 106820 8596 112252
rect 8764 111636 8820 114800
rect 8988 114324 9044 114800
rect 8988 114258 9044 114268
rect 9100 114436 9156 114446
rect 9100 112980 9156 114380
rect 9212 114100 9268 114800
rect 9212 114034 9268 114044
rect 9212 113204 9268 113214
rect 9212 113202 9380 113204
rect 9212 113150 9214 113202
rect 9266 113150 9380 113202
rect 9212 113148 9380 113150
rect 9212 113138 9268 113148
rect 9324 112980 9380 113148
rect 9100 112924 9268 112980
rect 9100 112308 9156 112318
rect 9100 112214 9156 112252
rect 8764 111570 8820 111580
rect 8876 112084 8932 112094
rect 8876 110516 8932 112028
rect 9212 111970 9268 112924
rect 9324 112914 9380 112924
rect 9436 112084 9492 114800
rect 9660 113988 9716 114800
rect 9884 114772 9940 114800
rect 9884 114706 9940 114716
rect 9660 113922 9716 113932
rect 9212 111918 9214 111970
rect 9266 111918 9268 111970
rect 9212 111906 9268 111918
rect 9324 112028 9492 112084
rect 9660 113426 9716 113438
rect 9660 113374 9662 113426
rect 9714 113374 9716 113426
rect 9660 112084 9716 113374
rect 10108 112644 10164 114800
rect 10220 114212 10276 114222
rect 10220 113092 10276 114156
rect 10332 113652 10388 114800
rect 10556 114436 10612 114800
rect 10556 114370 10612 114380
rect 10332 113586 10388 113596
rect 10780 113428 10836 114800
rect 10220 113026 10276 113036
rect 10332 113372 10836 113428
rect 10108 112578 10164 112588
rect 10220 112532 10276 112542
rect 10220 112418 10276 112476
rect 10220 112366 10222 112418
rect 10274 112366 10276 112418
rect 10220 112354 10276 112366
rect 8876 110450 8932 110460
rect 8988 111746 9044 111758
rect 8988 111694 8990 111746
rect 9042 111694 9044 111746
rect 8876 110178 8932 110190
rect 8876 110126 8878 110178
rect 8930 110126 8932 110178
rect 8652 109284 8708 109294
rect 8876 109228 8932 110126
rect 8652 107714 8708 109228
rect 8652 107662 8654 107714
rect 8706 107662 8708 107714
rect 8652 107650 8708 107662
rect 8764 109172 8932 109228
rect 8540 106754 8596 106764
rect 8428 106194 8484 106204
rect 8092 106034 8148 106046
rect 8092 105982 8094 106034
rect 8146 105982 8148 106034
rect 8092 105588 8148 105982
rect 8092 105028 8148 105532
rect 8316 105924 8372 105934
rect 8092 104962 8148 104972
rect 8204 105250 8260 105262
rect 8204 105198 8206 105250
rect 8258 105198 8260 105250
rect 8092 104690 8148 104702
rect 8092 104638 8094 104690
rect 8146 104638 8148 104690
rect 8092 104468 8148 104638
rect 8092 104402 8148 104412
rect 8204 103908 8260 105198
rect 7980 103070 7982 103122
rect 8034 103070 8036 103122
rect 7980 103058 8036 103070
rect 8092 103852 8260 103908
rect 7980 102452 8036 102462
rect 7868 102450 8036 102452
rect 7868 102398 7982 102450
rect 8034 102398 8036 102450
rect 7868 102396 8036 102398
rect 7980 102386 8036 102396
rect 6972 100830 6974 100882
rect 7026 100830 7028 100882
rect 6636 100770 6692 100782
rect 6636 100718 6638 100770
rect 6690 100718 6692 100770
rect 6636 100660 6692 100718
rect 6636 100594 6692 100604
rect 6748 99762 6804 99774
rect 6748 99710 6750 99762
rect 6802 99710 6804 99762
rect 6524 98018 6580 98028
rect 6636 99314 6692 99326
rect 6636 99262 6638 99314
rect 6690 99262 6692 99314
rect 6412 97300 6468 97580
rect 6412 97234 6468 97244
rect 6524 97860 6580 97870
rect 5964 94668 6356 94724
rect 6412 96516 6468 96526
rect 6412 96180 6468 96460
rect 6412 94836 6468 96124
rect 6524 95844 6580 97804
rect 6636 96964 6692 99262
rect 6748 97468 6804 99710
rect 6972 98756 7028 100830
rect 6972 98690 7028 98700
rect 7196 101388 7476 101444
rect 6860 98196 6916 98206
rect 6860 98102 6916 98140
rect 7084 97634 7140 97646
rect 7084 97582 7086 97634
rect 7138 97582 7140 97634
rect 7084 97524 7140 97582
rect 6748 97412 6916 97468
rect 7084 97458 7140 97468
rect 6636 96898 6692 96908
rect 6748 96068 6804 96078
rect 6748 95974 6804 96012
rect 6524 95788 6804 95844
rect 6636 95172 6692 95182
rect 6636 95078 6692 95116
rect 6412 94780 6692 94836
rect 5516 94276 5572 94286
rect 5516 94274 5908 94276
rect 5516 94222 5518 94274
rect 5570 94222 5908 94274
rect 5516 94220 5908 94222
rect 5516 94210 5572 94220
rect 5404 92418 5460 92428
rect 5516 94052 5572 94062
rect 4956 91410 5012 91420
rect 5180 92204 5348 92260
rect 5404 92260 5460 92270
rect 4956 91252 5012 91262
rect 4956 91158 5012 91196
rect 4844 88174 4846 88226
rect 4898 88174 4900 88226
rect 4844 88162 4900 88174
rect 5068 89012 5124 89022
rect 5180 89012 5236 92204
rect 5404 92166 5460 92204
rect 5292 91922 5348 91934
rect 5292 91870 5294 91922
rect 5346 91870 5348 91922
rect 5292 91812 5348 91870
rect 5516 91812 5572 93996
rect 5740 93716 5796 93754
rect 5740 93650 5796 93660
rect 5740 93492 5796 93502
rect 5628 92932 5684 92942
rect 5628 92838 5684 92876
rect 5740 92484 5796 93436
rect 5740 92418 5796 92428
rect 5740 92036 5796 92046
rect 5292 91756 5684 91812
rect 5404 90244 5460 90254
rect 5124 88956 5236 89012
rect 5292 89794 5348 89806
rect 5292 89742 5294 89794
rect 5346 89742 5348 89794
rect 4284 87378 4340 87388
rect 4060 86940 4228 86996
rect 4464 87052 4728 87062
rect 4520 86996 4568 87052
rect 4624 86996 4672 87052
rect 4464 86986 4728 86996
rect 3948 86884 4004 86894
rect 3724 86660 3780 86670
rect 3724 86566 3780 86604
rect 3948 86548 4004 86828
rect 4060 86548 4116 86940
rect 4172 86772 4228 86782
rect 4172 86770 4900 86772
rect 4172 86718 4174 86770
rect 4226 86718 4900 86770
rect 4172 86716 4900 86718
rect 4172 86706 4228 86716
rect 4060 86492 4228 86548
rect 3948 86482 4004 86492
rect 3804 86268 4068 86278
rect 3860 86212 3908 86268
rect 3964 86212 4012 86268
rect 3804 86202 4068 86212
rect 3948 86100 4004 86110
rect 3836 85090 3892 85102
rect 3836 85038 3838 85090
rect 3890 85038 3892 85090
rect 3836 84868 3892 85038
rect 3948 84868 4004 86044
rect 4172 84980 4228 86492
rect 4844 85708 4900 86716
rect 4284 85652 4340 85662
rect 4844 85652 5012 85708
rect 4284 85558 4340 85596
rect 4464 85484 4728 85494
rect 4520 85428 4568 85484
rect 4624 85428 4672 85484
rect 4464 85418 4728 85428
rect 4844 85090 4900 85102
rect 4844 85038 4846 85090
rect 4898 85038 4900 85090
rect 4172 84924 4452 84980
rect 3948 84812 4340 84868
rect 3836 84802 3892 84812
rect 3804 84700 4068 84710
rect 3860 84644 3908 84700
rect 3964 84644 4012 84700
rect 3804 84634 4068 84644
rect 4172 84308 4228 84318
rect 3948 83634 4004 83646
rect 3948 83582 3950 83634
rect 4002 83582 4004 83634
rect 3948 83524 4004 83582
rect 3948 83458 4004 83468
rect 3804 83132 4068 83142
rect 3860 83076 3908 83132
rect 3964 83076 4012 83132
rect 3804 83066 4068 83076
rect 3612 82908 4116 82964
rect 3724 82068 3780 82078
rect 3724 81974 3780 82012
rect 4060 81954 4116 82908
rect 4060 81902 4062 81954
rect 4114 81902 4116 81954
rect 4060 81890 4116 81902
rect 4172 82738 4228 84252
rect 4284 83746 4340 84812
rect 4396 84084 4452 84924
rect 4844 84308 4900 85038
rect 4844 84242 4900 84252
rect 4396 84018 4452 84028
rect 4464 83916 4728 83926
rect 4520 83860 4568 83916
rect 4624 83860 4672 83916
rect 4464 83850 4728 83860
rect 4284 83694 4286 83746
rect 4338 83694 4340 83746
rect 4284 83682 4340 83694
rect 4956 82740 5012 85652
rect 5068 83636 5124 88956
rect 5292 88226 5348 89742
rect 5292 88174 5294 88226
rect 5346 88174 5348 88226
rect 5292 88004 5348 88174
rect 5292 87938 5348 87948
rect 5404 86660 5460 90188
rect 5628 89124 5684 91756
rect 5740 90916 5796 91980
rect 5740 90850 5796 90860
rect 5852 89348 5908 94220
rect 5964 93380 6020 94668
rect 6188 94500 6244 94510
rect 6188 93716 6244 94444
rect 5964 93314 6020 93324
rect 6076 93602 6132 93614
rect 6076 93550 6078 93602
rect 6130 93550 6132 93602
rect 5964 92820 6020 92830
rect 5964 92726 6020 92764
rect 6076 92596 6132 93550
rect 6076 92530 6132 92540
rect 5964 92484 6020 92494
rect 5964 90692 6020 92428
rect 6188 92146 6244 93660
rect 6188 92094 6190 92146
rect 6242 92094 6244 92146
rect 6188 91476 6244 92094
rect 6076 90692 6132 90702
rect 5964 90690 6132 90692
rect 5964 90638 6078 90690
rect 6130 90638 6132 90690
rect 5964 90636 6132 90638
rect 6076 90626 6132 90636
rect 6188 90244 6244 91420
rect 6188 90178 6244 90188
rect 6300 94164 6356 94174
rect 6300 90020 6356 94108
rect 6412 91700 6468 94780
rect 6636 94722 6692 94780
rect 6636 94670 6638 94722
rect 6690 94670 6692 94722
rect 6636 94658 6692 94670
rect 6636 92932 6692 92942
rect 6636 92838 6692 92876
rect 6748 92596 6804 95788
rect 6748 92530 6804 92540
rect 6860 92372 6916 97412
rect 7084 96626 7140 96638
rect 7084 96574 7086 96626
rect 7138 96574 7140 96626
rect 7084 95620 7140 96574
rect 7084 95554 7140 95564
rect 7084 95396 7140 95406
rect 7084 95302 7140 95340
rect 7084 94500 7140 94510
rect 7084 94406 7140 94444
rect 6636 92316 6916 92372
rect 6972 94276 7028 94286
rect 6636 92260 6692 92316
rect 6972 92260 7028 94220
rect 7084 93268 7140 93278
rect 7084 93154 7140 93212
rect 7084 93102 7086 93154
rect 7138 93102 7140 93154
rect 7084 93090 7140 93102
rect 6524 92204 6692 92260
rect 6748 92204 7028 92260
rect 7084 92596 7140 92606
rect 6524 91924 6580 92204
rect 6636 92036 6692 92046
rect 6636 91942 6692 91980
rect 6524 91858 6580 91868
rect 6412 91644 6692 91700
rect 6524 91476 6580 91486
rect 6524 91362 6580 91420
rect 6524 91310 6526 91362
rect 6578 91310 6580 91362
rect 6524 91298 6580 91310
rect 6524 91140 6580 91150
rect 6524 90578 6580 91084
rect 6524 90526 6526 90578
rect 6578 90526 6580 90578
rect 6524 90514 6580 90526
rect 5852 89282 5908 89292
rect 5964 89964 6356 90020
rect 5852 89124 5908 89134
rect 5628 89122 5908 89124
rect 5628 89070 5854 89122
rect 5906 89070 5908 89122
rect 5628 89068 5908 89070
rect 5852 89058 5908 89068
rect 5964 88900 6020 89964
rect 6188 89796 6244 89806
rect 6188 89794 6356 89796
rect 6188 89742 6190 89794
rect 6242 89742 6356 89794
rect 6188 89740 6356 89742
rect 6188 89730 6244 89740
rect 6188 89348 6244 89358
rect 6188 89010 6244 89292
rect 6188 88958 6190 89010
rect 6242 88958 6244 89010
rect 6188 88946 6244 88958
rect 5740 88844 6020 88900
rect 5460 86604 5684 86660
rect 5404 86594 5460 86604
rect 5292 86434 5348 86446
rect 5292 86382 5294 86434
rect 5346 86382 5348 86434
rect 5292 85988 5348 86382
rect 5292 85922 5348 85932
rect 5516 85652 5572 85662
rect 5068 83570 5124 83580
rect 5180 85650 5572 85652
rect 5180 85598 5518 85650
rect 5570 85598 5572 85650
rect 5180 85596 5572 85598
rect 4172 82686 4174 82738
rect 4226 82686 4228 82738
rect 3612 81732 3668 81742
rect 3612 80388 3668 81676
rect 3804 81564 4068 81574
rect 3860 81508 3908 81564
rect 3964 81508 4012 81564
rect 3804 81498 4068 81508
rect 4172 81284 4228 82686
rect 4844 82684 5012 82740
rect 5068 83410 5124 83422
rect 5068 83358 5070 83410
rect 5122 83358 5124 83410
rect 4464 82348 4728 82358
rect 4520 82292 4568 82348
rect 4624 82292 4672 82348
rect 4464 82282 4728 82292
rect 4732 82066 4788 82078
rect 4732 82014 4734 82066
rect 4786 82014 4788 82066
rect 4508 81954 4564 81966
rect 4508 81902 4510 81954
rect 4562 81902 4564 81954
rect 4508 81732 4564 81902
rect 4508 81666 4564 81676
rect 3948 80948 4004 80958
rect 3948 80854 4004 80892
rect 3612 80294 3668 80332
rect 4172 80276 4228 81228
rect 4284 80948 4340 80958
rect 4508 80948 4564 80958
rect 4284 80946 4508 80948
rect 4284 80894 4286 80946
rect 4338 80894 4508 80946
rect 4284 80892 4508 80894
rect 4732 80948 4788 82014
rect 4844 81508 4900 82684
rect 4956 82514 5012 82526
rect 4956 82462 4958 82514
rect 5010 82462 5012 82514
rect 4956 81844 5012 82462
rect 5068 82068 5124 83358
rect 5068 82002 5124 82012
rect 5180 82066 5236 85596
rect 5516 85586 5572 85596
rect 5628 85092 5684 86604
rect 5404 85036 5684 85092
rect 5292 84308 5348 84318
rect 5404 84308 5460 85036
rect 5292 84306 5460 84308
rect 5292 84254 5294 84306
rect 5346 84254 5460 84306
rect 5292 84252 5460 84254
rect 5516 84866 5572 84878
rect 5516 84814 5518 84866
rect 5570 84814 5572 84866
rect 5292 82740 5348 84252
rect 5404 83972 5460 83982
rect 5404 83522 5460 83916
rect 5404 83470 5406 83522
rect 5458 83470 5460 83522
rect 5404 83458 5460 83470
rect 5292 82674 5348 82684
rect 5292 82514 5348 82526
rect 5292 82462 5294 82514
rect 5346 82462 5348 82514
rect 5292 82404 5348 82462
rect 5292 82338 5348 82348
rect 5180 82014 5182 82066
rect 5234 82014 5236 82066
rect 5180 82002 5236 82014
rect 4956 81788 5236 81844
rect 4844 81442 4900 81452
rect 4732 80892 4900 80948
rect 4284 80882 4340 80892
rect 4508 80882 4564 80892
rect 4464 80780 4728 80790
rect 4520 80724 4568 80780
rect 4624 80724 4672 80780
rect 4464 80714 4728 80724
rect 4508 80386 4564 80398
rect 4508 80334 4510 80386
rect 4562 80334 4564 80386
rect 4508 80276 4564 80334
rect 4172 80220 4564 80276
rect 3804 79996 4068 80006
rect 3860 79940 3908 79996
rect 3964 79940 4012 79996
rect 3804 79930 4068 79940
rect 3388 78988 3556 79044
rect 3612 79378 3668 79390
rect 3612 79326 3614 79378
rect 3666 79326 3668 79378
rect 3388 78148 3444 78988
rect 3500 78706 3556 78718
rect 3500 78654 3502 78706
rect 3554 78654 3556 78706
rect 3500 78372 3556 78654
rect 3500 78306 3556 78316
rect 3612 78148 3668 79326
rect 4060 79378 4116 79390
rect 4060 79326 4062 79378
rect 4114 79326 4116 79378
rect 4060 79156 4116 79326
rect 4060 79090 4116 79100
rect 3948 78930 4004 78942
rect 3948 78878 3950 78930
rect 4002 78878 4004 78930
rect 3948 78820 4004 78878
rect 3948 78754 4004 78764
rect 3804 78428 4068 78438
rect 3860 78372 3908 78428
rect 3964 78372 4012 78428
rect 3804 78362 4068 78372
rect 4172 78372 4228 80220
rect 4172 78306 4228 78316
rect 4284 79602 4340 79614
rect 4284 79550 4286 79602
rect 4338 79550 4340 79602
rect 3388 78092 3556 78148
rect 3612 78092 4228 78148
rect 3052 77858 3108 77868
rect 3164 77980 3332 78036
rect 3500 78036 3556 78092
rect 3500 77980 3892 78036
rect 3052 77588 3108 77598
rect 3052 77252 3108 77532
rect 3164 77476 3220 77980
rect 3388 77924 3444 77934
rect 3444 77868 3556 77924
rect 3388 77858 3444 77868
rect 3276 77812 3332 77822
rect 3276 77718 3332 77756
rect 3164 77420 3332 77476
rect 3164 77252 3220 77262
rect 3052 77250 3220 77252
rect 3052 77198 3166 77250
rect 3218 77198 3220 77250
rect 3052 77196 3220 77198
rect 2940 77084 3108 77140
rect 2940 75684 2996 75694
rect 2940 75590 2996 75628
rect 2940 74788 2996 74798
rect 2940 74226 2996 74732
rect 2940 74174 2942 74226
rect 2994 74174 2996 74226
rect 2940 74162 2996 74174
rect 3052 73948 3108 77084
rect 3164 76916 3220 77196
rect 3164 76850 3220 76860
rect 3164 76468 3220 76478
rect 3164 75906 3220 76412
rect 3164 75854 3166 75906
rect 3218 75854 3220 75906
rect 3164 75842 3220 75854
rect 3276 74114 3332 77420
rect 3388 77362 3444 77374
rect 3388 77310 3390 77362
rect 3442 77310 3444 77362
rect 3388 77252 3444 77310
rect 3388 77186 3444 77196
rect 3500 76916 3556 77868
rect 3612 77812 3668 77850
rect 3612 77746 3668 77756
rect 3836 77250 3892 77980
rect 4172 78034 4228 78092
rect 4172 77982 4174 78034
rect 4226 77982 4228 78034
rect 4172 77970 4228 77982
rect 3948 77810 4004 77822
rect 3948 77758 3950 77810
rect 4002 77758 4004 77810
rect 3948 77364 4004 77758
rect 4172 77812 4228 77822
rect 4284 77812 4340 79550
rect 4464 79212 4728 79222
rect 4520 79156 4568 79212
rect 4624 79156 4672 79212
rect 4464 79146 4728 79156
rect 4228 77756 4340 77812
rect 4172 77746 4228 77756
rect 4844 77700 4900 80892
rect 4956 80946 5012 80958
rect 4956 80894 4958 80946
rect 5010 80894 5012 80946
rect 4956 79828 5012 80894
rect 5068 80724 5124 80734
rect 5068 80498 5124 80668
rect 5068 80446 5070 80498
rect 5122 80446 5124 80498
rect 5068 80434 5124 80446
rect 4956 79762 5012 79772
rect 5068 78594 5124 78606
rect 5068 78542 5070 78594
rect 5122 78542 5124 78594
rect 4464 77644 4728 77654
rect 4844 77644 5012 77700
rect 4520 77588 4568 77644
rect 4624 77588 4672 77644
rect 4464 77578 4728 77588
rect 3948 77298 4004 77308
rect 4844 77364 4900 77374
rect 3836 77198 3838 77250
rect 3890 77198 3892 77250
rect 3836 77186 3892 77198
rect 4396 77250 4452 77262
rect 4396 77198 4398 77250
rect 4450 77198 4452 77250
rect 4396 77140 4452 77198
rect 4396 77074 4452 77084
rect 3388 76860 3556 76916
rect 4172 77028 4228 77038
rect 3804 76860 4068 76870
rect 3388 76692 3444 76860
rect 3860 76804 3908 76860
rect 3964 76804 4012 76860
rect 3804 76794 4068 76804
rect 3388 76636 3668 76692
rect 3500 76242 3556 76254
rect 3500 76190 3502 76242
rect 3554 76190 3556 76242
rect 3276 74062 3278 74114
rect 3330 74062 3332 74114
rect 3276 74050 3332 74062
rect 3388 74674 3444 74686
rect 3388 74622 3390 74674
rect 3442 74622 3444 74674
rect 3052 73892 3220 73948
rect 3388 73892 3444 74622
rect 2604 72482 2660 72492
rect 2716 72716 2884 72772
rect 2940 73332 2996 73342
rect 2716 72212 2772 72716
rect 2156 71260 2324 71316
rect 2380 72156 2772 72212
rect 2828 72548 2884 72558
rect 2156 70532 2212 71260
rect 2268 70980 2324 70990
rect 2268 70886 2324 70924
rect 2156 70476 2324 70532
rect 2044 70466 2100 70476
rect 2044 70196 2100 70206
rect 1932 69300 1988 69310
rect 1820 69298 1988 69300
rect 1820 69246 1934 69298
rect 1986 69246 1988 69298
rect 1820 69244 1988 69246
rect 924 66882 980 66892
rect 1148 66836 1204 66846
rect 1148 66742 1204 66780
rect 1260 66612 1316 68572
rect 1372 68402 1428 68414
rect 1372 68350 1374 68402
rect 1426 68350 1428 68402
rect 1372 68068 1428 68350
rect 1820 68404 1876 69244
rect 1932 69234 1988 69244
rect 1932 68628 1988 68638
rect 1932 68534 1988 68572
rect 1820 68348 1988 68404
rect 1372 68002 1428 68012
rect 1820 68068 1876 68078
rect 1820 67974 1876 68012
rect 1372 67842 1428 67854
rect 1372 67790 1374 67842
rect 1426 67790 1428 67842
rect 1372 66724 1428 67790
rect 1820 67284 1876 67294
rect 1484 66948 1540 66958
rect 1484 66854 1540 66892
rect 1820 66946 1876 67228
rect 1820 66894 1822 66946
rect 1874 66894 1876 66946
rect 1820 66882 1876 66894
rect 1372 66668 1764 66724
rect 1260 66556 1540 66612
rect 1260 66388 1316 66398
rect 1260 66274 1316 66332
rect 1260 66222 1262 66274
rect 1314 66222 1316 66274
rect 1260 66210 1316 66222
rect 1260 65490 1316 65502
rect 1260 65438 1262 65490
rect 1314 65438 1316 65490
rect 1036 65268 1092 65278
rect 812 63970 868 63980
rect 924 65266 1092 65268
rect 924 65214 1038 65266
rect 1090 65214 1092 65266
rect 924 65212 1092 65214
rect 924 63700 980 65212
rect 1036 65202 1092 65212
rect 1260 64148 1316 65438
rect 1260 64082 1316 64092
rect 1372 64706 1428 64718
rect 1372 64654 1374 64706
rect 1426 64654 1428 64706
rect 1260 63922 1316 63934
rect 1260 63870 1262 63922
rect 1314 63870 1316 63922
rect 588 61954 644 61964
rect 700 63644 980 63700
rect 1036 63698 1092 63710
rect 1036 63646 1038 63698
rect 1090 63646 1092 63698
rect 700 61348 756 63644
rect 1036 62188 1092 63646
rect 1260 63362 1316 63870
rect 1260 63310 1262 63362
rect 1314 63310 1316 63362
rect 1260 63298 1316 63310
rect 1372 63364 1428 64654
rect 1372 63298 1428 63308
rect 1484 63138 1540 66556
rect 1596 66500 1652 66510
rect 1596 66386 1652 66444
rect 1596 66334 1598 66386
rect 1650 66334 1652 66386
rect 1596 66322 1652 66334
rect 1708 66164 1764 66668
rect 1596 66108 1764 66164
rect 1820 66388 1876 66398
rect 1596 64596 1652 66108
rect 1820 65604 1876 66332
rect 1932 66052 1988 68348
rect 2044 66724 2100 70140
rect 2268 68514 2324 70476
rect 2380 69410 2436 72156
rect 2716 71762 2772 71774
rect 2716 71710 2718 71762
rect 2770 71710 2772 71762
rect 2492 71090 2548 71102
rect 2492 71038 2494 71090
rect 2546 71038 2548 71090
rect 2492 70644 2548 71038
rect 2492 70578 2548 70588
rect 2604 70868 2660 70878
rect 2380 69358 2382 69410
rect 2434 69358 2436 69410
rect 2380 69346 2436 69358
rect 2492 69972 2548 69982
rect 2268 68462 2270 68514
rect 2322 68462 2324 68514
rect 2268 68450 2324 68462
rect 2156 67842 2212 67854
rect 2156 67790 2158 67842
rect 2210 67790 2212 67842
rect 2156 67620 2212 67790
rect 2156 67554 2212 67564
rect 2492 67284 2548 69916
rect 2268 67228 2548 67284
rect 2044 66658 2100 66668
rect 2156 66834 2212 66846
rect 2156 66782 2158 66834
rect 2210 66782 2212 66834
rect 2156 66612 2212 66782
rect 2156 66546 2212 66556
rect 2156 66276 2212 66286
rect 1932 65996 2100 66052
rect 1932 65604 1988 65614
rect 1820 65548 1932 65604
rect 1932 65510 1988 65548
rect 1596 64530 1652 64540
rect 1708 64818 1764 64830
rect 1708 64766 1710 64818
rect 1762 64766 1764 64818
rect 1708 64036 1764 64766
rect 2044 64596 2100 65996
rect 1708 63970 1764 63980
rect 1932 64594 2100 64596
rect 1932 64542 2046 64594
rect 2098 64542 2100 64594
rect 1932 64540 2100 64542
rect 1484 63086 1486 63138
rect 1538 63086 1540 63138
rect 1484 63074 1540 63086
rect 1820 63922 1876 63934
rect 1820 63870 1822 63922
rect 1874 63870 1876 63922
rect 1820 63140 1876 63870
rect 1820 63074 1876 63084
rect 1932 63026 1988 64540
rect 2044 64530 2100 64540
rect 1932 62974 1934 63026
rect 1986 62974 1988 63026
rect 700 61282 756 61292
rect 812 62132 1092 62188
rect 1148 62354 1204 62366
rect 1148 62302 1150 62354
rect 1202 62302 1204 62354
rect 1148 62132 1204 62302
rect 1484 62354 1540 62366
rect 1484 62302 1486 62354
rect 1538 62302 1540 62354
rect 1484 62188 1540 62302
rect 700 60900 756 60910
rect 700 57876 756 60844
rect 812 60452 868 62132
rect 1148 62066 1204 62076
rect 1260 62132 1540 62188
rect 1932 62244 1988 62974
rect 2044 62356 2100 62366
rect 2044 62262 2100 62300
rect 1932 62178 1988 62188
rect 2156 62242 2212 66220
rect 2268 64708 2324 67228
rect 2380 67060 2436 67070
rect 2380 65378 2436 67004
rect 2380 65326 2382 65378
rect 2434 65326 2436 65378
rect 2380 65314 2436 65326
rect 2492 66948 2548 66958
rect 2492 65268 2548 66892
rect 2604 66164 2660 70812
rect 2716 67170 2772 71710
rect 2828 70868 2884 72492
rect 2828 70802 2884 70812
rect 2940 72546 2996 73276
rect 3052 72772 3108 72782
rect 3052 72678 3108 72716
rect 2940 72494 2942 72546
rect 2994 72494 2996 72546
rect 2940 70980 2996 72494
rect 3164 71650 3220 73892
rect 3164 71598 3166 71650
rect 3218 71598 3220 71650
rect 3164 71586 3220 71598
rect 3276 73836 3444 73892
rect 2828 69972 2884 69982
rect 2828 69878 2884 69916
rect 2940 69748 2996 70924
rect 3164 70980 3220 70990
rect 3276 70980 3332 73836
rect 3164 70978 3332 70980
rect 3164 70926 3166 70978
rect 3218 70926 3332 70978
rect 3164 70924 3332 70926
rect 3388 73106 3444 73118
rect 3388 73054 3390 73106
rect 3442 73054 3444 73106
rect 3164 70914 3220 70924
rect 3276 70756 3332 70766
rect 3276 70082 3332 70700
rect 3276 70030 3278 70082
rect 3330 70030 3332 70082
rect 3276 70018 3332 70030
rect 2828 69692 2996 69748
rect 2828 69410 2884 69692
rect 2940 69524 2996 69534
rect 2940 69522 3332 69524
rect 2940 69470 2942 69522
rect 2994 69470 3332 69522
rect 2940 69468 3332 69470
rect 2940 69458 2996 69468
rect 2828 69358 2830 69410
rect 2882 69358 2884 69410
rect 2828 69346 2884 69358
rect 2940 69300 2996 69310
rect 2940 68628 2996 69244
rect 2940 67730 2996 68572
rect 2940 67678 2942 67730
rect 2994 67678 2996 67730
rect 2940 67620 2996 67678
rect 2940 67564 3220 67620
rect 2716 67118 2718 67170
rect 2770 67118 2772 67170
rect 2716 66388 2772 67118
rect 3052 66948 3108 66958
rect 3052 66854 3108 66892
rect 2716 66322 2772 66332
rect 3052 66612 3108 66622
rect 2604 66108 2772 66164
rect 2492 65212 2660 65268
rect 2492 65044 2548 65054
rect 2380 64708 2436 64718
rect 2268 64706 2436 64708
rect 2268 64654 2382 64706
rect 2434 64654 2436 64706
rect 2268 64652 2436 64654
rect 2380 64642 2436 64652
rect 2380 63812 2436 63822
rect 2380 63718 2436 63756
rect 2380 63140 2436 63150
rect 2492 63140 2548 64988
rect 2380 63138 2548 63140
rect 2380 63086 2382 63138
rect 2434 63086 2548 63138
rect 2380 63084 2548 63086
rect 2380 63074 2436 63084
rect 2156 62190 2158 62242
rect 2210 62190 2212 62242
rect 2156 62178 2212 62190
rect 1036 61684 1092 61694
rect 812 60386 868 60396
rect 924 61682 1092 61684
rect 924 61630 1038 61682
rect 1090 61630 1092 61682
rect 924 61628 1092 61630
rect 924 60004 980 61628
rect 1036 61618 1092 61628
rect 924 59938 980 59948
rect 1036 60562 1092 60574
rect 1036 60510 1038 60562
rect 1090 60510 1092 60562
rect 1036 59556 1092 60510
rect 1148 60228 1204 60238
rect 1260 60228 1316 62132
rect 2156 61796 2212 61806
rect 2156 61702 2212 61740
rect 1372 61684 1428 61694
rect 1372 61590 1428 61628
rect 1820 61684 1876 61694
rect 1820 61590 1876 61628
rect 1484 61460 1540 61470
rect 1372 60564 1428 60574
rect 1372 60470 1428 60508
rect 1148 60226 1316 60228
rect 1148 60174 1150 60226
rect 1202 60174 1316 60226
rect 1148 60172 1316 60174
rect 1148 60162 1204 60172
rect 1036 59490 1092 59500
rect 1484 59444 1540 61404
rect 1260 59388 1540 59444
rect 1596 61348 1652 61358
rect 1036 58996 1092 59006
rect 924 58994 1092 58996
rect 924 58942 1038 58994
rect 1090 58942 1092 58994
rect 924 58940 1092 58942
rect 924 58660 980 58940
rect 1036 58930 1092 58940
rect 924 58594 980 58604
rect 1036 58546 1092 58558
rect 1036 58494 1038 58546
rect 1090 58494 1092 58546
rect 1036 58212 1092 58494
rect 1260 58436 1316 59388
rect 1372 58996 1428 59006
rect 1596 58996 1652 61292
rect 2604 61012 2660 65212
rect 2716 64708 2772 66108
rect 2828 66050 2884 66062
rect 2828 65998 2830 66050
rect 2882 65998 2884 66050
rect 2828 65044 2884 65998
rect 2828 64978 2884 64988
rect 3052 64930 3108 66556
rect 3052 64878 3054 64930
rect 3106 64878 3108 64930
rect 3052 64866 3108 64878
rect 2828 64708 2884 64718
rect 2716 64706 2884 64708
rect 2716 64654 2830 64706
rect 2882 64654 2884 64706
rect 2716 64652 2884 64654
rect 2828 64372 2884 64652
rect 2716 64316 2884 64372
rect 2716 63138 2772 64316
rect 2716 63086 2718 63138
rect 2770 63086 2772 63138
rect 2716 62356 2772 63086
rect 2716 62290 2772 62300
rect 2828 63924 2884 63934
rect 2828 62354 2884 63868
rect 2940 63364 2996 63374
rect 2940 63270 2996 63308
rect 2828 62302 2830 62354
rect 2882 62302 2884 62354
rect 2828 62290 2884 62302
rect 2940 63140 2996 63150
rect 2268 60956 2660 61012
rect 2940 61570 2996 63084
rect 3164 63140 3220 67564
rect 3276 66498 3332 69468
rect 3388 69522 3444 73054
rect 3500 72658 3556 76190
rect 3612 75794 3668 76636
rect 3612 75742 3614 75794
rect 3666 75742 3668 75794
rect 3612 75730 3668 75742
rect 3948 76242 4004 76254
rect 3948 76190 3950 76242
rect 4002 76190 4004 76242
rect 3948 75684 4004 76190
rect 3948 75618 4004 75628
rect 4172 75682 4228 76972
rect 4172 75630 4174 75682
rect 4226 75630 4228 75682
rect 4172 75618 4228 75630
rect 4284 76242 4340 76254
rect 4284 76190 4286 76242
rect 4338 76190 4340 76242
rect 4172 75460 4228 75470
rect 3804 75292 4068 75302
rect 3860 75236 3908 75292
rect 3964 75236 4012 75292
rect 3804 75226 4068 75236
rect 3836 74900 3892 74910
rect 3836 74676 3892 74844
rect 3836 74610 3892 74620
rect 4060 74674 4116 74686
rect 4060 74622 4062 74674
rect 4114 74622 4116 74674
rect 4060 74564 4116 74622
rect 4060 74498 4116 74508
rect 3948 74452 4004 74462
rect 3948 74338 4004 74396
rect 3948 74286 3950 74338
rect 4002 74286 4004 74338
rect 3948 74274 4004 74286
rect 3836 74228 3892 74238
rect 3836 74114 3892 74172
rect 3836 74062 3838 74114
rect 3890 74062 3892 74114
rect 3836 74050 3892 74062
rect 3612 74004 3668 74014
rect 3612 73220 3668 73948
rect 3804 73724 4068 73734
rect 3860 73668 3908 73724
rect 3964 73668 4012 73724
rect 3804 73658 4068 73668
rect 4172 73330 4228 75404
rect 4284 75124 4340 76190
rect 4464 76076 4728 76086
rect 4520 76020 4568 76076
rect 4624 76020 4672 76076
rect 4464 76010 4728 76020
rect 4284 75058 4340 75068
rect 4396 75012 4452 75022
rect 4172 73278 4174 73330
rect 4226 73278 4228 73330
rect 4172 73266 4228 73278
rect 4284 74900 4340 74910
rect 4284 74116 4340 74844
rect 4396 74898 4452 74956
rect 4396 74846 4398 74898
rect 4450 74846 4452 74898
rect 4396 74834 4452 74846
rect 4464 74508 4728 74518
rect 4520 74452 4568 74508
rect 4624 74452 4672 74508
rect 4464 74442 4728 74452
rect 3836 73220 3892 73230
rect 3612 73218 3892 73220
rect 3612 73166 3838 73218
rect 3890 73166 3892 73218
rect 3612 73164 3892 73166
rect 3836 73154 3892 73164
rect 3500 72606 3502 72658
rect 3554 72606 3556 72658
rect 3500 72594 3556 72606
rect 4284 72546 4340 74060
rect 4620 74116 4676 74126
rect 4844 74116 4900 77308
rect 4956 75460 5012 77644
rect 5068 77364 5124 78542
rect 5068 77298 5124 77308
rect 5180 77252 5236 81788
rect 5404 81732 5460 81742
rect 5292 80946 5348 80958
rect 5292 80894 5294 80946
rect 5346 80894 5348 80946
rect 5292 77364 5348 80894
rect 5404 79380 5460 81676
rect 5516 80386 5572 84814
rect 5516 80334 5518 80386
rect 5570 80334 5572 80386
rect 5516 80322 5572 80334
rect 5628 84084 5684 84094
rect 5628 82852 5684 84028
rect 5628 79604 5684 82796
rect 5740 81954 5796 88844
rect 6300 88228 6356 89740
rect 6636 89236 6692 91644
rect 6748 89906 6804 92204
rect 7084 92148 7140 92540
rect 6860 92092 7140 92148
rect 6860 90578 6916 92092
rect 7084 91588 7140 91598
rect 6860 90526 6862 90578
rect 6914 90526 6916 90578
rect 6860 90356 6916 90526
rect 6860 90290 6916 90300
rect 6972 91532 7084 91588
rect 6748 89854 6750 89906
rect 6802 89854 6804 89906
rect 6748 89842 6804 89854
rect 6636 89180 6804 89236
rect 6636 89012 6692 89022
rect 6636 88918 6692 88956
rect 6748 88788 6804 89180
rect 6860 88900 6916 88910
rect 6860 88806 6916 88844
rect 6636 88732 6804 88788
rect 6412 88228 6468 88238
rect 6300 88226 6468 88228
rect 6300 88174 6414 88226
rect 6466 88174 6468 88226
rect 6300 88172 6468 88174
rect 6300 87556 6356 87566
rect 5964 87500 6300 87556
rect 5964 86658 6020 87500
rect 6300 87462 6356 87500
rect 5964 86606 5966 86658
rect 6018 86606 6020 86658
rect 5852 84308 5908 84318
rect 5852 84194 5908 84252
rect 5852 84142 5854 84194
rect 5906 84142 5908 84194
rect 5852 84130 5908 84142
rect 5964 84084 6020 86606
rect 5964 84018 6020 84028
rect 6188 87332 6244 87342
rect 6188 85876 6244 87276
rect 6412 87220 6468 88172
rect 6636 87330 6692 88732
rect 6636 87278 6638 87330
rect 6690 87278 6692 87330
rect 6636 87266 6692 87278
rect 6076 83636 6132 83646
rect 5964 83634 6132 83636
rect 5964 83582 6078 83634
rect 6130 83582 6132 83634
rect 5964 83580 6132 83582
rect 5852 83522 5908 83534
rect 5852 83470 5854 83522
rect 5906 83470 5908 83522
rect 5852 83300 5908 83470
rect 5852 83234 5908 83244
rect 5852 82852 5908 82862
rect 5852 82758 5908 82796
rect 5740 81902 5742 81954
rect 5794 81902 5796 81954
rect 5740 80724 5796 81902
rect 5740 80658 5796 80668
rect 5852 80386 5908 80398
rect 5852 80334 5854 80386
rect 5906 80334 5908 80386
rect 5852 80164 5908 80334
rect 5852 80098 5908 80108
rect 5628 79548 5908 79604
rect 5404 79314 5460 79324
rect 5628 79380 5684 79390
rect 5852 79380 5908 79548
rect 5628 79378 5796 79380
rect 5628 79326 5630 79378
rect 5682 79326 5796 79378
rect 5628 79324 5796 79326
rect 5628 79314 5684 79324
rect 5516 78930 5572 78942
rect 5516 78878 5518 78930
rect 5570 78878 5572 78930
rect 5292 77298 5348 77308
rect 5404 78372 5460 78382
rect 5404 78148 5460 78316
rect 5180 77186 5236 77196
rect 5404 77250 5460 78092
rect 5404 77198 5406 77250
rect 5458 77198 5460 77250
rect 5068 76466 5124 76478
rect 5404 76468 5460 77198
rect 5068 76414 5070 76466
rect 5122 76414 5124 76466
rect 5068 76356 5124 76414
rect 5068 76290 5124 76300
rect 5180 76412 5460 76468
rect 5180 75684 5236 76412
rect 4956 75394 5012 75404
rect 5068 75682 5236 75684
rect 5068 75630 5182 75682
rect 5234 75630 5236 75682
rect 5068 75628 5236 75630
rect 5068 74340 5124 75628
rect 5180 75618 5236 75628
rect 5292 76242 5348 76254
rect 5292 76190 5294 76242
rect 5346 76190 5348 76242
rect 5292 74900 5348 76190
rect 5404 74900 5460 74910
rect 5292 74898 5460 74900
rect 5292 74846 5406 74898
rect 5458 74846 5460 74898
rect 5292 74844 5460 74846
rect 5404 74834 5460 74844
rect 4620 74114 4900 74116
rect 4620 74062 4622 74114
rect 4674 74062 4900 74114
rect 4620 74060 4900 74062
rect 4956 74284 5124 74340
rect 5180 74674 5236 74686
rect 5180 74622 5182 74674
rect 5234 74622 5236 74674
rect 4620 74050 4676 74060
rect 4956 73444 5012 74284
rect 5068 74116 5124 74126
rect 5068 74022 5124 74060
rect 4956 73388 5124 73444
rect 4956 73220 5012 73230
rect 4956 73126 5012 73164
rect 4464 72940 4728 72950
rect 4520 72884 4568 72940
rect 4624 72884 4672 72940
rect 4464 72874 4728 72884
rect 4284 72494 4286 72546
rect 4338 72494 4340 72546
rect 4284 72482 4340 72494
rect 4396 72548 4452 72558
rect 3804 72156 4068 72166
rect 3860 72100 3908 72156
rect 3964 72100 4012 72156
rect 3804 72090 4068 72100
rect 4284 71764 4340 71774
rect 4284 71670 4340 71708
rect 4396 71540 4452 72492
rect 5068 72548 5124 73388
rect 5180 73108 5236 74622
rect 5180 73042 5236 73052
rect 5292 73106 5348 73118
rect 5292 73054 5294 73106
rect 5346 73054 5348 73106
rect 5292 72772 5348 73054
rect 5292 72706 5348 72716
rect 5068 72454 5124 72492
rect 5180 71876 5236 71886
rect 4956 71540 5012 71550
rect 4284 71484 4452 71540
rect 4844 71538 5012 71540
rect 4844 71486 4958 71538
rect 5010 71486 5012 71538
rect 4844 71484 5012 71486
rect 4284 71204 4340 71484
rect 4464 71372 4728 71382
rect 4520 71316 4568 71372
rect 4624 71316 4672 71372
rect 4464 71306 4728 71316
rect 4284 71148 4564 71204
rect 3500 70980 3556 70990
rect 4508 70980 4564 71148
rect 3556 70924 3668 70980
rect 3500 70886 3556 70924
rect 3500 70644 3556 70654
rect 3500 70194 3556 70588
rect 3500 70142 3502 70194
rect 3554 70142 3556 70194
rect 3500 70130 3556 70142
rect 3388 69470 3390 69522
rect 3442 69470 3444 69522
rect 3388 69458 3444 69470
rect 3612 69412 3668 70924
rect 4508 70886 4564 70924
rect 3804 70588 4068 70598
rect 3860 70532 3908 70588
rect 3964 70532 4012 70588
rect 3804 70522 4068 70532
rect 4284 70532 4340 70542
rect 4060 70196 4116 70206
rect 4060 70194 4228 70196
rect 4060 70142 4062 70194
rect 4114 70142 4228 70194
rect 4060 70140 4228 70142
rect 4060 70130 4116 70140
rect 3948 69412 4004 69422
rect 3612 69410 4004 69412
rect 3612 69358 3950 69410
rect 4002 69358 4004 69410
rect 3612 69356 4004 69358
rect 3948 69346 4004 69356
rect 3388 69300 3444 69310
rect 3388 69188 3444 69244
rect 3836 69188 3892 69198
rect 3388 69132 3836 69188
rect 3836 69122 3892 69132
rect 3804 69020 4068 69030
rect 3860 68964 3908 69020
rect 3964 68964 4012 69020
rect 3804 68954 4068 68964
rect 4172 68852 4228 70140
rect 4284 70082 4340 70476
rect 4284 70030 4286 70082
rect 4338 70030 4340 70082
rect 4284 70018 4340 70030
rect 4464 69804 4728 69814
rect 4520 69748 4568 69804
rect 4624 69748 4672 69804
rect 4464 69738 4728 69748
rect 4172 68786 4228 68796
rect 4172 68626 4228 68638
rect 4172 68574 4174 68626
rect 4226 68574 4228 68626
rect 3500 68402 3556 68414
rect 3500 68350 3502 68402
rect 3554 68350 3556 68402
rect 3388 67954 3444 67966
rect 3388 67902 3390 67954
rect 3442 67902 3444 67954
rect 3388 67284 3444 67902
rect 3388 67218 3444 67228
rect 3500 66724 3556 68350
rect 3948 68402 4004 68414
rect 3948 68350 3950 68402
rect 4002 68350 4004 68402
rect 3948 67732 4004 68350
rect 3948 67666 4004 67676
rect 3804 67452 4068 67462
rect 3860 67396 3908 67452
rect 3964 67396 4012 67452
rect 3804 67386 4068 67396
rect 3276 66446 3278 66498
rect 3330 66446 3332 66498
rect 3276 66434 3332 66446
rect 3388 66668 3556 66724
rect 3388 65940 3444 66668
rect 4172 66500 4228 68574
rect 4844 68516 4900 71484
rect 4956 71474 5012 71484
rect 4844 68450 4900 68460
rect 4956 70980 5012 70990
rect 4956 69410 5012 70924
rect 5068 70868 5124 70878
rect 5180 70868 5236 71820
rect 5292 71538 5348 71550
rect 5292 71486 5294 71538
rect 5346 71486 5348 71538
rect 5292 71316 5348 71486
rect 5292 71250 5348 71260
rect 5516 71204 5572 78878
rect 5628 78260 5684 78270
rect 5628 78034 5684 78204
rect 5628 77982 5630 78034
rect 5682 77982 5684 78034
rect 5628 77924 5684 77982
rect 5628 77858 5684 77868
rect 5740 76468 5796 79324
rect 5852 79314 5908 79324
rect 5852 78818 5908 78830
rect 5852 78766 5854 78818
rect 5906 78766 5908 78818
rect 5852 76916 5908 78766
rect 5852 76850 5908 76860
rect 5964 76468 6020 83580
rect 6076 83570 6132 83580
rect 6188 82626 6244 85820
rect 6300 87164 6468 87220
rect 6300 84196 6356 87164
rect 6412 86996 6468 87006
rect 6412 86882 6468 86940
rect 6412 86830 6414 86882
rect 6466 86830 6468 86882
rect 6412 85204 6468 86830
rect 6748 86884 6804 86894
rect 6748 86212 6804 86828
rect 6748 85762 6804 86156
rect 6748 85710 6750 85762
rect 6802 85710 6804 85762
rect 6412 85138 6468 85148
rect 6524 85652 6580 85662
rect 6300 84130 6356 84140
rect 6524 83634 6580 85596
rect 6748 85202 6804 85710
rect 6748 85150 6750 85202
rect 6802 85150 6804 85202
rect 6748 85138 6804 85150
rect 6972 84420 7028 91532
rect 7084 91494 7140 91532
rect 7084 90804 7140 90814
rect 7084 90466 7140 90748
rect 7084 90414 7086 90466
rect 7138 90414 7140 90466
rect 7084 90402 7140 90414
rect 7196 90132 7252 101388
rect 7532 101330 7588 101342
rect 7532 101278 7534 101330
rect 7586 101278 7588 101330
rect 7308 100882 7364 100894
rect 7308 100830 7310 100882
rect 7362 100830 7364 100882
rect 7308 100772 7364 100830
rect 7308 100706 7364 100716
rect 7420 100548 7476 100558
rect 7308 98756 7364 98766
rect 7308 97748 7364 98700
rect 7420 98644 7476 100492
rect 7532 98868 7588 101278
rect 7644 100770 7700 100782
rect 7644 100718 7646 100770
rect 7698 100718 7700 100770
rect 7644 100324 7700 100718
rect 7644 100258 7700 100268
rect 8092 99988 8148 103852
rect 8204 103682 8260 103694
rect 8204 103630 8206 103682
rect 8258 103630 8260 103682
rect 8204 100772 8260 103630
rect 8316 103348 8372 105868
rect 8540 104580 8596 104590
rect 8316 103292 8484 103348
rect 8428 102900 8484 103292
rect 8540 103122 8596 104524
rect 8764 104468 8820 109172
rect 8988 108948 9044 111694
rect 8988 108882 9044 108892
rect 9100 110962 9156 110974
rect 9100 110910 9102 110962
rect 9154 110910 9156 110962
rect 9100 109394 9156 110910
rect 9212 110292 9268 110302
rect 9212 110198 9268 110236
rect 9100 109342 9102 109394
rect 9154 109342 9156 109394
rect 8876 108612 8932 108622
rect 8876 108518 8932 108556
rect 9100 108500 9156 109342
rect 9212 108836 9268 108846
rect 9212 108742 9268 108780
rect 8988 107716 9044 107726
rect 8876 107714 9044 107716
rect 8876 107662 8990 107714
rect 9042 107662 9044 107714
rect 8876 107660 9044 107662
rect 8876 106932 8932 107660
rect 8988 107650 9044 107660
rect 8876 106838 8932 106876
rect 9100 106708 9156 108444
rect 9324 108164 9380 112028
rect 9660 112018 9716 112028
rect 9324 108098 9380 108108
rect 9436 111860 9492 111870
rect 9324 107828 9380 107838
rect 9324 107734 9380 107772
rect 8876 106652 9156 106708
rect 8876 104692 8932 106652
rect 9212 106036 9268 106046
rect 9100 106034 9268 106036
rect 9100 105982 9214 106034
rect 9266 105982 9268 106034
rect 9100 105980 9268 105982
rect 9100 105812 9156 105980
rect 9212 105970 9268 105980
rect 9100 105746 9156 105756
rect 9212 105700 9268 105710
rect 9436 105700 9492 111804
rect 10332 111860 10388 113372
rect 11004 113316 11060 114800
rect 11228 113428 11284 114800
rect 10668 113260 11060 113316
rect 11116 113372 11284 113428
rect 10668 113204 10724 113260
rect 10332 111794 10388 111804
rect 10444 113148 10724 113204
rect 10220 111748 10276 111758
rect 9660 111634 9716 111646
rect 9660 111582 9662 111634
rect 9714 111582 9716 111634
rect 9660 111076 9716 111582
rect 9996 111634 10052 111646
rect 9996 111582 9998 111634
rect 10050 111582 10052 111634
rect 9660 111074 9940 111076
rect 9660 111022 9662 111074
rect 9714 111022 9940 111074
rect 9660 111020 9940 111022
rect 9660 111010 9716 111020
rect 9548 110066 9604 110078
rect 9548 110014 9550 110066
rect 9602 110014 9604 110066
rect 9548 109172 9604 110014
rect 9884 109396 9940 111020
rect 9996 110964 10052 111582
rect 9996 110962 10164 110964
rect 9996 110910 9998 110962
rect 10050 110910 10164 110962
rect 9996 110908 10164 110910
rect 9996 110898 10052 110908
rect 9996 110404 10052 110414
rect 9996 110310 10052 110348
rect 10108 110180 10164 110908
rect 10220 110850 10276 111692
rect 10220 110798 10222 110850
rect 10274 110798 10276 110850
rect 10220 110786 10276 110798
rect 10332 110180 10388 110190
rect 10108 110124 10332 110180
rect 10332 110086 10388 110124
rect 9884 109330 9940 109340
rect 10220 109956 10276 109966
rect 9548 109106 9604 109116
rect 9660 109170 9716 109182
rect 9660 109118 9662 109170
rect 9714 109118 9716 109170
rect 9548 108948 9604 108958
rect 9548 108834 9604 108892
rect 9548 108782 9550 108834
rect 9602 108782 9604 108834
rect 9548 108770 9604 108782
rect 9548 106932 9604 106942
rect 9548 106838 9604 106876
rect 9660 106260 9716 109118
rect 10220 108834 10276 109900
rect 10444 109228 10500 113148
rect 10780 113092 10836 113102
rect 10780 113090 11060 113092
rect 10780 113038 10782 113090
rect 10834 113038 11060 113090
rect 10780 113036 11060 113038
rect 10780 113026 10836 113036
rect 10668 112532 10724 112542
rect 10556 111748 10612 111758
rect 10556 111654 10612 111692
rect 10668 111300 10724 112476
rect 10780 112530 10836 112542
rect 10780 112478 10782 112530
rect 10834 112478 10836 112530
rect 10780 112196 10836 112478
rect 10780 112130 10836 112140
rect 10892 111972 10948 111982
rect 10892 111878 10948 111916
rect 10892 111412 10948 111422
rect 10668 111244 10836 111300
rect 10668 111076 10724 111086
rect 10556 110964 10612 110974
rect 10556 110870 10612 110908
rect 10220 108782 10222 108834
rect 10274 108782 10276 108834
rect 10220 108770 10276 108782
rect 10332 109172 10500 109228
rect 9996 108724 10052 108734
rect 9884 108612 9940 108622
rect 9884 108518 9940 108556
rect 9884 107940 9940 107950
rect 9772 107828 9828 107838
rect 9772 107734 9828 107772
rect 9884 107042 9940 107884
rect 9996 107828 10052 108668
rect 10332 108164 10388 109172
rect 10556 108948 10612 108958
rect 10556 108834 10612 108892
rect 10556 108782 10558 108834
rect 10610 108782 10612 108834
rect 10556 108770 10612 108782
rect 10668 108388 10724 111020
rect 10780 109956 10836 111244
rect 10892 110962 10948 111356
rect 10892 110910 10894 110962
rect 10946 110910 10948 110962
rect 10892 110898 10948 110910
rect 10892 110740 10948 110750
rect 10892 110178 10948 110684
rect 10892 110126 10894 110178
rect 10946 110126 10948 110178
rect 10892 110114 10948 110126
rect 10780 109900 10948 109956
rect 10780 109172 10836 109182
rect 10780 109078 10836 109116
rect 10892 108724 10948 109900
rect 11004 109228 11060 113036
rect 11116 112532 11172 113372
rect 11228 113204 11284 113214
rect 11228 113202 11396 113204
rect 11228 113150 11230 113202
rect 11282 113150 11396 113202
rect 11228 113148 11396 113150
rect 11228 113138 11284 113148
rect 11116 112466 11172 112476
rect 11340 112420 11396 113148
rect 11340 112354 11396 112364
rect 11228 112308 11284 112318
rect 11116 112306 11284 112308
rect 11116 112254 11230 112306
rect 11282 112254 11284 112306
rect 11116 112252 11284 112254
rect 11116 109394 11172 112252
rect 11228 112242 11284 112252
rect 11228 111636 11284 111646
rect 11228 111542 11284 111580
rect 11228 110738 11284 110750
rect 11228 110686 11230 110738
rect 11282 110686 11284 110738
rect 11228 109956 11284 110686
rect 11228 109890 11284 109900
rect 11340 110290 11396 110302
rect 11340 110238 11342 110290
rect 11394 110238 11396 110290
rect 11116 109342 11118 109394
rect 11170 109342 11172 109394
rect 11116 109330 11172 109342
rect 11004 109172 11284 109228
rect 10892 108668 11172 108724
rect 10892 108500 10948 108510
rect 10668 108322 10724 108332
rect 10780 108498 10948 108500
rect 10780 108446 10894 108498
rect 10946 108446 10948 108498
rect 10780 108444 10948 108446
rect 9996 107762 10052 107772
rect 10108 108108 10388 108164
rect 9884 106990 9886 107042
rect 9938 106990 9940 107042
rect 9884 106978 9940 106990
rect 9996 107602 10052 107614
rect 9996 107550 9998 107602
rect 10050 107550 10052 107602
rect 9996 107044 10052 107550
rect 10108 107266 10164 108108
rect 10444 107716 10500 107726
rect 10444 107622 10500 107660
rect 10108 107214 10110 107266
rect 10162 107214 10164 107266
rect 10108 107202 10164 107214
rect 9996 106988 10164 107044
rect 9212 105698 9492 105700
rect 9212 105646 9214 105698
rect 9266 105646 9492 105698
rect 9212 105644 9492 105646
rect 9548 106204 9716 106260
rect 9212 105634 9268 105644
rect 9548 105588 9604 106204
rect 9996 106148 10052 106158
rect 9996 106054 10052 106092
rect 9324 105532 9604 105588
rect 9660 106034 9716 106046
rect 9660 105982 9662 106034
rect 9714 105982 9716 106034
rect 8988 105476 9044 105486
rect 9324 105476 9380 105532
rect 8988 105474 9380 105476
rect 8988 105422 8990 105474
rect 9042 105422 9380 105474
rect 8988 105420 9380 105422
rect 8988 105410 9044 105420
rect 9660 105362 9716 105982
rect 10108 105868 10164 106988
rect 10780 106932 10836 108444
rect 10892 108434 10948 108444
rect 11004 107828 11060 107838
rect 11004 107734 11060 107772
rect 10780 106838 10836 106876
rect 11116 106260 11172 108668
rect 11228 108610 11284 109172
rect 11228 108558 11230 108610
rect 11282 108558 11284 108610
rect 11228 108546 11284 108558
rect 11340 107156 11396 110238
rect 11452 109282 11508 114800
rect 11564 113428 11620 113438
rect 11564 113334 11620 113372
rect 11676 112756 11732 114800
rect 11900 114436 11956 114800
rect 11900 114370 11956 114380
rect 12124 114212 12180 114800
rect 12124 114146 12180 114156
rect 12348 113876 12404 114800
rect 12348 113810 12404 113820
rect 12460 114548 12516 114558
rect 11900 113764 11956 113774
rect 11676 112690 11732 112700
rect 11788 113314 11844 113326
rect 11788 113262 11790 113314
rect 11842 113262 11844 113314
rect 11564 112420 11620 112430
rect 11564 112326 11620 112364
rect 11788 111972 11844 113262
rect 11900 112532 11956 113708
rect 12460 113428 12516 114492
rect 12572 113652 12628 114800
rect 12572 113586 12628 113596
rect 12572 113428 12628 113438
rect 12460 113426 12628 113428
rect 12460 113374 12574 113426
rect 12626 113374 12628 113426
rect 12460 113372 12628 113374
rect 12572 113362 12628 113372
rect 12236 113092 12292 113102
rect 11900 112466 11956 112476
rect 12012 112980 12068 112990
rect 11900 112306 11956 112318
rect 11900 112254 11902 112306
rect 11954 112254 11956 112306
rect 11900 112084 11956 112254
rect 11900 112018 11956 112028
rect 11564 111916 11844 111972
rect 11564 111634 11620 111916
rect 11732 111804 11844 111916
rect 12012 111746 12068 112924
rect 12012 111694 12014 111746
rect 12066 111694 12068 111746
rect 12012 111682 12068 111694
rect 12124 112644 12180 112654
rect 11564 111582 11566 111634
rect 11618 111582 11620 111634
rect 11564 111074 11620 111582
rect 12124 111188 12180 112588
rect 12236 112418 12292 113036
rect 12796 112980 12852 114800
rect 13020 113540 13076 114800
rect 13020 113474 13076 113484
rect 13244 113092 13300 114800
rect 13244 113026 13300 113036
rect 12796 112914 12852 112924
rect 12236 112366 12238 112418
rect 12290 112366 12292 112418
rect 12236 112354 12292 112366
rect 12908 112306 12964 112318
rect 12908 112254 12910 112306
rect 12962 112254 12964 112306
rect 11564 111022 11566 111074
rect 11618 111022 11620 111074
rect 11564 110964 11620 111022
rect 11564 110898 11620 110908
rect 11788 111132 12180 111188
rect 12236 112084 12292 112094
rect 12236 111188 12292 112028
rect 11452 109230 11454 109282
rect 11506 109230 11508 109282
rect 11452 109218 11508 109230
rect 11564 110516 11620 110526
rect 11564 108836 11620 110460
rect 11788 109282 11844 111132
rect 12236 111122 12292 111132
rect 12460 112084 12516 112094
rect 12460 111858 12516 112028
rect 12460 111806 12462 111858
rect 12514 111806 12516 111858
rect 12012 110964 12068 110974
rect 12012 110962 12404 110964
rect 12012 110910 12014 110962
rect 12066 110910 12404 110962
rect 12012 110908 12404 110910
rect 12012 110898 12068 110908
rect 12236 110738 12292 110750
rect 12236 110686 12238 110738
rect 12290 110686 12292 110738
rect 12236 110404 12292 110686
rect 12236 110338 12292 110348
rect 11788 109230 11790 109282
rect 11842 109230 11844 109282
rect 11788 109218 11844 109230
rect 12124 109284 12180 109322
rect 12124 109218 12180 109228
rect 11340 107090 11396 107100
rect 11452 108780 11620 108836
rect 11676 109172 11732 109182
rect 11004 106204 11172 106260
rect 10332 106036 10388 106046
rect 10332 106034 10500 106036
rect 10332 105982 10334 106034
rect 10386 105982 10500 106034
rect 10332 105980 10500 105982
rect 10332 105970 10388 105980
rect 9660 105310 9662 105362
rect 9714 105310 9716 105362
rect 9212 104692 9268 104702
rect 8876 104690 9268 104692
rect 8876 104638 9214 104690
rect 9266 104638 9268 104690
rect 8876 104636 9268 104638
rect 8764 104412 9156 104468
rect 8540 103070 8542 103122
rect 8594 103070 8596 103122
rect 8540 103058 8596 103070
rect 8876 103348 8932 103358
rect 8316 102844 8484 102900
rect 8316 102450 8372 102844
rect 8316 102398 8318 102450
rect 8370 102398 8372 102450
rect 8316 102386 8372 102398
rect 8204 100706 8260 100716
rect 8652 102340 8708 102350
rect 8652 101442 8708 102284
rect 8652 101390 8654 101442
rect 8706 101390 8708 101442
rect 8652 100548 8708 101390
rect 8652 100482 8708 100492
rect 8876 100100 8932 103292
rect 8988 102452 9044 102462
rect 8988 101554 9044 102396
rect 9100 102450 9156 104412
rect 9100 102398 9102 102450
rect 9154 102398 9156 102450
rect 9100 102386 9156 102398
rect 8988 101502 8990 101554
rect 9042 101502 9044 101554
rect 8988 101490 9044 101502
rect 8988 100100 9044 100110
rect 8092 99922 8148 99932
rect 8540 100098 9044 100100
rect 8540 100046 8990 100098
rect 9042 100046 9044 100098
rect 8540 100044 9044 100046
rect 8316 99204 8372 99214
rect 8092 99202 8372 99204
rect 8092 99150 8318 99202
rect 8370 99150 8372 99202
rect 8092 99148 8372 99150
rect 7756 99092 7812 99102
rect 8092 99092 8148 99148
rect 8316 99138 8372 99148
rect 7756 99090 8148 99092
rect 7756 99038 7758 99090
rect 7810 99038 8148 99090
rect 7756 99036 8148 99038
rect 7756 99026 7812 99036
rect 7532 98802 7588 98812
rect 7980 98756 8036 99036
rect 8204 98980 8260 98990
rect 8204 98886 8260 98924
rect 7756 98700 8036 98756
rect 8092 98868 8148 98878
rect 7420 98588 7700 98644
rect 7308 97468 7364 97692
rect 7420 98420 7476 98430
rect 7420 97636 7476 98364
rect 7420 97570 7476 97580
rect 7644 97524 7700 98588
rect 7756 97634 7812 98700
rect 7980 98308 8036 98318
rect 7980 98214 8036 98252
rect 8092 98084 8148 98812
rect 7980 98028 8148 98084
rect 7980 97636 8036 98028
rect 8092 97860 8148 97870
rect 8092 97858 8372 97860
rect 8092 97806 8094 97858
rect 8146 97806 8372 97858
rect 8092 97804 8372 97806
rect 8092 97794 8148 97804
rect 7756 97582 7758 97634
rect 7810 97582 7812 97634
rect 7756 97570 7812 97582
rect 7868 97634 8036 97636
rect 7868 97582 7982 97634
rect 8034 97582 8036 97634
rect 7868 97580 8036 97582
rect 7308 97412 7588 97468
rect 7644 97458 7700 97468
rect 7420 97188 7476 97198
rect 7308 96404 7364 96414
rect 7308 96178 7364 96348
rect 7308 96126 7310 96178
rect 7362 96126 7364 96178
rect 7308 96114 7364 96126
rect 7308 95620 7364 95630
rect 7308 93716 7364 95564
rect 7420 93828 7476 97132
rect 7532 93940 7588 97412
rect 7756 97412 7812 97422
rect 7756 96962 7812 97356
rect 7756 96910 7758 96962
rect 7810 96910 7812 96962
rect 7756 96898 7812 96910
rect 7868 96740 7924 97580
rect 7980 97570 8036 97580
rect 8204 97636 8260 97646
rect 8204 97542 8260 97580
rect 7644 96684 7924 96740
rect 8092 97524 8148 97534
rect 7644 96066 7700 96684
rect 7644 96014 7646 96066
rect 7698 96014 7700 96066
rect 7644 96002 7700 96014
rect 7756 96236 8036 96292
rect 7756 96066 7812 96236
rect 7756 96014 7758 96066
rect 7810 96014 7812 96066
rect 7756 96002 7812 96014
rect 7868 96066 7924 96078
rect 7868 96014 7870 96066
rect 7922 96014 7924 96066
rect 7868 95956 7924 96014
rect 7980 96068 8036 96236
rect 8092 96290 8148 97468
rect 8204 96852 8260 96862
rect 8204 96738 8260 96796
rect 8204 96686 8206 96738
rect 8258 96686 8260 96738
rect 8204 96674 8260 96686
rect 8316 96516 8372 97804
rect 8092 96238 8094 96290
rect 8146 96238 8148 96290
rect 8092 96226 8148 96238
rect 8204 96460 8372 96516
rect 8428 97300 8484 97310
rect 8204 96068 8260 96460
rect 7980 96012 8260 96068
rect 7868 95900 8036 95956
rect 7532 93884 7924 93940
rect 7420 93772 7700 93828
rect 7308 93660 7588 93716
rect 7084 90076 7252 90132
rect 7308 93490 7364 93502
rect 7308 93438 7310 93490
rect 7362 93438 7364 93490
rect 7084 87556 7140 90076
rect 7196 89908 7252 89918
rect 7196 89814 7252 89852
rect 7308 89010 7364 93438
rect 7308 88958 7310 89010
rect 7362 88958 7364 89010
rect 7308 88946 7364 88958
rect 7420 90692 7476 90702
rect 7308 88114 7364 88126
rect 7308 88062 7310 88114
rect 7362 88062 7364 88114
rect 7140 87500 7252 87556
rect 7084 87490 7140 87500
rect 6524 83582 6526 83634
rect 6578 83582 6580 83634
rect 6524 83570 6580 83582
rect 6748 84364 7028 84420
rect 7084 86772 7140 86782
rect 7084 85986 7140 86716
rect 7084 85934 7086 85986
rect 7138 85934 7140 85986
rect 6188 82574 6190 82626
rect 6242 82574 6244 82626
rect 6188 82562 6244 82574
rect 6748 82180 6804 84364
rect 6748 82114 6804 82124
rect 6860 84196 6916 84206
rect 6748 81954 6804 81966
rect 6748 81902 6750 81954
rect 6802 81902 6804 81954
rect 6412 81620 6468 81630
rect 6188 81170 6244 81182
rect 6188 81118 6190 81170
rect 6242 81118 6244 81170
rect 6188 80836 6244 81118
rect 6188 80770 6244 80780
rect 6412 81060 6468 81564
rect 6748 81284 6804 81902
rect 6748 81218 6804 81228
rect 6412 80724 6468 81004
rect 6636 81060 6692 81070
rect 6636 80966 6692 81004
rect 6300 80668 6468 80724
rect 6636 80836 6692 80846
rect 6076 80498 6132 80510
rect 6076 80446 6078 80498
rect 6130 80446 6132 80498
rect 6076 80276 6132 80446
rect 6076 80210 6132 80220
rect 6188 80164 6244 80174
rect 6076 78708 6132 78718
rect 6076 78372 6132 78652
rect 6076 77922 6132 78316
rect 6076 77870 6078 77922
rect 6130 77870 6132 77922
rect 6076 77858 6132 77870
rect 6188 77364 6244 80108
rect 5740 76402 5796 76412
rect 5852 76412 6020 76468
rect 6076 77308 6244 77364
rect 5628 76242 5684 76254
rect 5628 76190 5630 76242
rect 5682 76190 5684 76242
rect 5628 74340 5684 76190
rect 5852 75796 5908 76412
rect 5964 76244 6020 76254
rect 5964 76150 6020 76188
rect 5852 75730 5908 75740
rect 6076 75572 6132 77308
rect 6188 77138 6244 77150
rect 6188 77086 6190 77138
rect 6242 77086 6244 77138
rect 6188 75908 6244 77086
rect 6188 75842 6244 75852
rect 5628 74274 5684 74284
rect 5740 75516 6132 75572
rect 6188 75684 6244 75694
rect 5068 70866 5236 70868
rect 5068 70814 5070 70866
rect 5122 70814 5236 70866
rect 5068 70812 5236 70814
rect 5404 71148 5572 71204
rect 5628 73106 5684 73118
rect 5628 73054 5630 73106
rect 5682 73054 5684 73106
rect 5628 71204 5684 73054
rect 5068 70756 5124 70812
rect 5068 70690 5124 70700
rect 4956 69358 4958 69410
rect 5010 69358 5012 69410
rect 4956 68292 5012 69358
rect 5292 70644 5348 70654
rect 5180 68964 5236 68974
rect 5180 68738 5236 68908
rect 5180 68686 5182 68738
rect 5234 68686 5236 68738
rect 5180 68674 5236 68686
rect 4464 68236 4728 68246
rect 4520 68180 4568 68236
rect 4624 68180 4672 68236
rect 4464 68170 4728 68180
rect 4844 68236 5012 68292
rect 4508 67844 4564 67854
rect 4508 67750 4564 67788
rect 4284 66836 4340 66846
rect 4284 66742 4340 66780
rect 4464 66668 4728 66678
rect 4520 66612 4568 66668
rect 4624 66612 4672 66668
rect 4464 66602 4728 66612
rect 4284 66500 4340 66510
rect 4172 66498 4340 66500
rect 4172 66446 4286 66498
rect 4338 66446 4340 66498
rect 4172 66444 4340 66446
rect 4284 66434 4340 66444
rect 3612 66388 3668 66398
rect 3612 66294 3668 66332
rect 3948 66276 4004 66286
rect 3948 66182 4004 66220
rect 3388 65884 3668 65940
rect 3500 65268 3556 65278
rect 3388 65266 3556 65268
rect 3388 65214 3502 65266
rect 3554 65214 3556 65266
rect 3388 65212 3556 65214
rect 3388 63250 3444 65212
rect 3500 65202 3556 65212
rect 3612 64706 3668 65884
rect 3804 65884 4068 65894
rect 3860 65828 3908 65884
rect 3964 65828 4012 65884
rect 3804 65818 4068 65828
rect 4396 65492 4452 65502
rect 4844 65492 4900 68236
rect 5292 68068 5348 70588
rect 5404 70308 5460 71148
rect 5628 71138 5684 71148
rect 5516 70978 5572 70990
rect 5516 70926 5518 70978
rect 5570 70926 5572 70978
rect 5516 70420 5572 70926
rect 5628 70420 5684 70430
rect 5516 70418 5684 70420
rect 5516 70366 5630 70418
rect 5682 70366 5684 70418
rect 5516 70364 5684 70366
rect 5628 70354 5684 70364
rect 5404 70242 5460 70252
rect 5740 69524 5796 75516
rect 6188 75236 6244 75628
rect 5964 75180 6244 75236
rect 5852 75124 5908 75134
rect 5852 73330 5908 75068
rect 5964 74788 6020 75180
rect 6076 75012 6132 75022
rect 6300 75012 6356 80668
rect 6524 80500 6580 80510
rect 6524 80406 6580 80444
rect 6412 79380 6468 79390
rect 6412 78818 6468 79324
rect 6636 79156 6692 80780
rect 6748 79492 6804 79502
rect 6748 79398 6804 79436
rect 6412 78766 6414 78818
rect 6466 78766 6468 78818
rect 6412 77924 6468 78766
rect 6412 77858 6468 77868
rect 6524 79100 6692 79156
rect 6524 75908 6580 79100
rect 6860 78932 6916 84140
rect 6972 84082 7028 84094
rect 6972 84030 6974 84082
rect 7026 84030 7028 84082
rect 6972 83524 7028 84030
rect 6972 83458 7028 83468
rect 7084 82404 7140 85934
rect 7196 85090 7252 87500
rect 7308 86884 7364 88062
rect 7308 86818 7364 86828
rect 7420 85708 7476 90636
rect 7532 90578 7588 93660
rect 7532 90526 7534 90578
rect 7586 90526 7588 90578
rect 7532 90514 7588 90526
rect 7644 89908 7700 93772
rect 7756 91924 7812 91934
rect 7756 91830 7812 91868
rect 7868 91364 7924 93884
rect 7980 92260 8036 95900
rect 8092 95170 8148 95182
rect 8092 95118 8094 95170
rect 8146 95118 8148 95170
rect 8092 92372 8148 95118
rect 8428 94612 8484 97244
rect 8540 95620 8596 100044
rect 8988 100034 9044 100044
rect 9100 98194 9156 98206
rect 9100 98142 9102 98194
rect 9154 98142 9156 98194
rect 8540 95554 8596 95564
rect 8652 97636 8708 97646
rect 8540 95282 8596 95294
rect 8540 95230 8542 95282
rect 8594 95230 8596 95282
rect 8540 94836 8596 95230
rect 8540 94770 8596 94780
rect 8428 94556 8596 94612
rect 8204 94500 8260 94510
rect 8204 93154 8260 94444
rect 8428 93940 8484 93950
rect 8204 93102 8206 93154
rect 8258 93102 8260 93154
rect 8204 93090 8260 93102
rect 8316 93268 8372 93278
rect 8316 92932 8372 93212
rect 8316 92866 8372 92876
rect 8204 92372 8260 92382
rect 8092 92316 8204 92372
rect 7980 92194 8036 92204
rect 8204 92258 8260 92316
rect 8204 92206 8206 92258
rect 8258 92206 8260 92258
rect 8204 92194 8260 92206
rect 8428 92148 8484 93884
rect 8540 93826 8596 94556
rect 8540 93774 8542 93826
rect 8594 93774 8596 93826
rect 8540 93044 8596 93774
rect 8540 92978 8596 92988
rect 8540 92148 8596 92158
rect 8428 92146 8596 92148
rect 8428 92094 8542 92146
rect 8594 92094 8596 92146
rect 8428 92092 8596 92094
rect 8540 92082 8596 92092
rect 8316 91924 8372 91934
rect 8204 91588 8260 91598
rect 8204 91494 8260 91532
rect 7868 91308 8260 91364
rect 8092 90578 8148 90590
rect 8092 90526 8094 90578
rect 8146 90526 8148 90578
rect 7644 89852 8036 89908
rect 7532 89684 7588 89694
rect 7532 89590 7588 89628
rect 7868 89572 7924 89582
rect 7868 89478 7924 89516
rect 7868 87218 7924 87230
rect 7868 87166 7870 87218
rect 7922 87166 7924 87218
rect 7196 85038 7198 85090
rect 7250 85038 7252 85090
rect 7196 85026 7252 85038
rect 7308 85652 7476 85708
rect 7532 86434 7588 86446
rect 7532 86382 7534 86434
rect 7586 86382 7588 86434
rect 7308 83522 7364 85652
rect 7420 84644 7476 84654
rect 7420 84418 7476 84588
rect 7420 84366 7422 84418
rect 7474 84366 7476 84418
rect 7420 84354 7476 84366
rect 7532 84308 7588 86382
rect 7532 84242 7588 84252
rect 7868 84306 7924 87166
rect 7980 85986 8036 89852
rect 8092 89348 8148 90526
rect 8092 89282 8148 89292
rect 7980 85934 7982 85986
rect 8034 85934 8036 85986
rect 7980 85922 8036 85934
rect 8092 89010 8148 89022
rect 8092 88958 8094 89010
rect 8146 88958 8148 89010
rect 7868 84254 7870 84306
rect 7922 84254 7924 84306
rect 7868 84242 7924 84254
rect 8092 85316 8148 88958
rect 8092 84084 8148 85260
rect 8204 84868 8260 91308
rect 8316 85876 8372 91868
rect 8540 91924 8596 91934
rect 8428 85876 8484 85886
rect 8316 85874 8484 85876
rect 8316 85822 8430 85874
rect 8482 85822 8484 85874
rect 8316 85820 8484 85822
rect 8428 85810 8484 85820
rect 8204 84306 8260 84812
rect 8204 84254 8206 84306
rect 8258 84254 8260 84306
rect 8204 84242 8260 84254
rect 8428 84084 8484 84094
rect 8092 84018 8148 84028
rect 8204 84082 8484 84084
rect 8204 84030 8430 84082
rect 8482 84030 8484 84082
rect 8204 84028 8484 84030
rect 7308 83470 7310 83522
rect 7362 83470 7364 83522
rect 7308 83458 7364 83470
rect 7868 83972 7924 83982
rect 7420 82516 7476 82526
rect 7084 82338 7140 82348
rect 7196 82514 7476 82516
rect 7196 82462 7422 82514
rect 7474 82462 7476 82514
rect 7196 82460 7476 82462
rect 7084 82180 7140 82190
rect 7084 80388 7140 82124
rect 7196 80500 7252 82460
rect 7420 82450 7476 82460
rect 7196 80434 7252 80444
rect 7308 82066 7364 82078
rect 7308 82014 7310 82066
rect 7362 82014 7364 82066
rect 6748 78930 6916 78932
rect 6748 78878 6862 78930
rect 6914 78878 6916 78930
rect 6748 78876 6916 78878
rect 6636 77476 6692 77486
rect 6636 77382 6692 77420
rect 6636 76804 6692 76814
rect 6636 76580 6692 76748
rect 6636 76486 6692 76524
rect 6524 75842 6580 75852
rect 6636 75796 6692 75806
rect 6636 75682 6692 75740
rect 6636 75630 6638 75682
rect 6690 75630 6692 75682
rect 6636 75618 6692 75630
rect 6076 75010 6356 75012
rect 6076 74958 6078 75010
rect 6130 74958 6356 75010
rect 6076 74956 6356 74958
rect 6076 74946 6132 74956
rect 5964 74732 6244 74788
rect 5852 73278 5854 73330
rect 5906 73278 5908 73330
rect 5852 73266 5908 73278
rect 5964 74114 6020 74126
rect 5964 74062 5966 74114
rect 6018 74062 6020 74114
rect 5852 72996 5908 73006
rect 5852 72546 5908 72940
rect 5852 72494 5854 72546
rect 5906 72494 5908 72546
rect 5852 72482 5908 72494
rect 5852 71876 5908 71886
rect 5964 71876 6020 74062
rect 5908 71820 6020 71876
rect 6076 71876 6132 71886
rect 5852 71810 5908 71820
rect 6076 71782 6132 71820
rect 6076 71204 6132 71214
rect 6188 71204 6244 74732
rect 6300 73948 6356 74956
rect 6524 74788 6580 74798
rect 6748 74788 6804 78876
rect 6860 78866 6916 78876
rect 6972 80386 7140 80388
rect 6972 80334 7086 80386
rect 7138 80334 7140 80386
rect 6972 80332 7140 80334
rect 6524 74786 6804 74788
rect 6524 74734 6526 74786
rect 6578 74734 6804 74786
rect 6524 74732 6804 74734
rect 6860 78148 6916 78158
rect 6524 74676 6580 74732
rect 6860 74676 6916 78092
rect 6524 74610 6580 74620
rect 6748 74620 6916 74676
rect 6972 76580 7028 80332
rect 7084 80322 7140 80332
rect 7196 79602 7252 79614
rect 7196 79550 7198 79602
rect 7250 79550 7252 79602
rect 7196 79380 7252 79550
rect 7196 79314 7252 79324
rect 7308 78932 7364 82014
rect 7868 82068 7924 83916
rect 8092 83522 8148 83534
rect 8092 83470 8094 83522
rect 8146 83470 8148 83522
rect 7868 82002 7924 82012
rect 7980 82066 8036 82078
rect 7980 82014 7982 82066
rect 8034 82014 8036 82066
rect 7532 81954 7588 81966
rect 7532 81902 7534 81954
rect 7586 81902 7588 81954
rect 7308 78866 7364 78876
rect 7420 81396 7476 81406
rect 7084 78484 7140 78494
rect 7084 78036 7140 78428
rect 7084 77970 7140 77980
rect 6524 74226 6580 74238
rect 6524 74174 6526 74226
rect 6578 74174 6580 74226
rect 6300 73892 6468 73948
rect 6412 73220 6468 73892
rect 6524 73444 6580 74174
rect 6524 73378 6580 73388
rect 6412 73164 6580 73220
rect 6300 73108 6356 73118
rect 6300 73106 6468 73108
rect 6300 73054 6302 73106
rect 6354 73054 6468 73106
rect 6300 73052 6468 73054
rect 6300 73042 6356 73052
rect 6300 72660 6356 72670
rect 6300 72566 6356 72604
rect 6412 71988 6468 73052
rect 6300 71932 6468 71988
rect 6300 71652 6356 71932
rect 6412 71764 6468 71774
rect 6412 71670 6468 71708
rect 6300 71586 6356 71596
rect 6076 71202 6244 71204
rect 6076 71150 6078 71202
rect 6130 71150 6244 71202
rect 6076 71148 6244 71150
rect 6300 71428 6356 71438
rect 6076 71138 6132 71148
rect 5852 70978 5908 70990
rect 5852 70926 5854 70978
rect 5906 70926 5908 70978
rect 5852 70868 5908 70926
rect 5852 70802 5908 70812
rect 5740 69468 5908 69524
rect 5740 69298 5796 69310
rect 5740 69246 5742 69298
rect 5794 69246 5796 69298
rect 5740 69188 5796 69246
rect 5740 69122 5796 69132
rect 5628 68740 5684 68750
rect 5628 68514 5684 68684
rect 5628 68462 5630 68514
rect 5682 68462 5684 68514
rect 5628 68450 5684 68462
rect 5292 68012 5572 68068
rect 4956 67956 5012 67966
rect 4956 67862 5012 67900
rect 5292 67844 5348 67854
rect 5292 67750 5348 67788
rect 5404 66836 5460 66846
rect 5180 66276 5236 66286
rect 5068 66220 5180 66276
rect 5068 66162 5124 66220
rect 5180 66210 5236 66220
rect 5404 66274 5460 66780
rect 5404 66222 5406 66274
rect 5458 66222 5460 66274
rect 5404 66210 5460 66222
rect 5068 66110 5070 66162
rect 5122 66110 5124 66162
rect 5068 66098 5124 66110
rect 4844 65436 5124 65492
rect 4396 65398 4452 65436
rect 4060 65268 4116 65278
rect 3612 64654 3614 64706
rect 3666 64654 3668 64706
rect 3612 64642 3668 64654
rect 3948 65266 4116 65268
rect 3948 65214 4062 65266
rect 4114 65214 4116 65266
rect 3948 65212 4116 65214
rect 3948 64484 4004 65212
rect 4060 65202 4116 65212
rect 4956 65266 5012 65278
rect 4956 65214 4958 65266
rect 5010 65214 5012 65266
rect 4464 65100 4728 65110
rect 4520 65044 4568 65100
rect 4624 65044 4672 65100
rect 4464 65034 4728 65044
rect 4956 64932 5012 65214
rect 4956 64866 5012 64876
rect 3948 64418 4004 64428
rect 4284 64708 4340 64718
rect 3804 64316 4068 64326
rect 3860 64260 3908 64316
rect 3964 64260 4012 64316
rect 3804 64250 4068 64260
rect 4172 64036 4228 64046
rect 3500 63924 3556 63934
rect 3500 63830 3556 63868
rect 4172 63922 4228 63980
rect 4172 63870 4174 63922
rect 4226 63870 4228 63922
rect 4172 63858 4228 63870
rect 3948 63700 4004 63710
rect 3388 63198 3390 63250
rect 3442 63198 3444 63250
rect 3388 63186 3444 63198
rect 3612 63698 4004 63700
rect 3612 63646 3950 63698
rect 4002 63646 4004 63698
rect 3612 63644 4004 63646
rect 3164 63074 3220 63084
rect 3388 62916 3444 62926
rect 3388 62354 3444 62860
rect 3388 62302 3390 62354
rect 3442 62302 3444 62354
rect 3388 62290 3444 62302
rect 3612 61908 3668 63644
rect 3948 63634 4004 63644
rect 4172 63140 4228 63150
rect 4284 63140 4340 64652
rect 5068 64706 5124 65436
rect 5292 65266 5348 65278
rect 5292 65214 5294 65266
rect 5346 65214 5348 65266
rect 5068 64654 5070 64706
rect 5122 64654 5124 64706
rect 4956 64596 5012 64606
rect 4956 63810 5012 64540
rect 4956 63758 4958 63810
rect 5010 63758 5012 63810
rect 4956 63746 5012 63758
rect 5068 64372 5124 64654
rect 5068 63588 5124 64316
rect 5180 64820 5236 64830
rect 5180 63922 5236 64764
rect 5180 63870 5182 63922
rect 5234 63870 5236 63922
rect 5180 63858 5236 63870
rect 4464 63532 4728 63542
rect 4520 63476 4568 63532
rect 4624 63476 4672 63532
rect 4464 63466 4728 63476
rect 4956 63532 5124 63588
rect 4956 63140 5012 63532
rect 5292 63364 5348 65214
rect 5292 63298 5348 63308
rect 4172 63138 4340 63140
rect 4172 63086 4174 63138
rect 4226 63086 4340 63138
rect 4172 63084 4340 63086
rect 4844 63138 5012 63140
rect 4844 63086 4958 63138
rect 5010 63086 5012 63138
rect 4844 63084 5012 63086
rect 4172 62916 4228 63084
rect 4172 62850 4228 62860
rect 3804 62748 4068 62758
rect 3860 62692 3908 62748
rect 3964 62692 4012 62748
rect 3804 62682 4068 62692
rect 4172 62692 4228 62702
rect 3612 61842 3668 61852
rect 3500 61684 3556 61694
rect 3500 61590 3556 61628
rect 2940 61518 2942 61570
rect 2994 61518 2996 61570
rect 2156 60676 2212 60686
rect 2156 60582 2212 60620
rect 1820 60564 1876 60574
rect 1820 60470 1876 60508
rect 2156 59220 2212 59230
rect 2268 59220 2324 60956
rect 2604 60786 2660 60798
rect 2604 60734 2606 60786
rect 2658 60734 2660 60786
rect 2380 60114 2436 60126
rect 2380 60062 2382 60114
rect 2434 60062 2436 60114
rect 2380 60004 2436 60062
rect 2380 59938 2436 59948
rect 2604 59892 2660 60734
rect 2604 59826 2660 59836
rect 2716 59892 2772 59902
rect 2940 59892 2996 61518
rect 3804 61180 4068 61190
rect 3860 61124 3908 61180
rect 3964 61124 4012 61180
rect 3804 61114 4068 61124
rect 3164 60564 3220 60574
rect 3164 60470 3220 60508
rect 4060 60228 4116 60238
rect 4172 60228 4228 62636
rect 4284 62356 4340 62366
rect 4844 62356 4900 63084
rect 4956 63074 5012 63084
rect 4284 62354 4900 62356
rect 4284 62302 4286 62354
rect 4338 62302 4900 62354
rect 4284 62300 4900 62302
rect 4956 62468 5012 62478
rect 4284 62290 4340 62300
rect 4956 62242 5012 62412
rect 4956 62190 4958 62242
rect 5010 62190 5012 62242
rect 4956 62178 5012 62190
rect 5292 62244 5348 62282
rect 5292 62178 5348 62188
rect 4284 62132 4340 62142
rect 4284 61010 4340 62076
rect 5068 62020 5124 62030
rect 4464 61964 4728 61974
rect 4520 61908 4568 61964
rect 4624 61908 4672 61964
rect 4464 61898 4728 61908
rect 5068 61682 5124 61964
rect 5068 61630 5070 61682
rect 5122 61630 5124 61682
rect 5068 61618 5124 61630
rect 4620 61572 4676 61582
rect 4620 61478 4676 61516
rect 5404 61572 5460 61582
rect 5404 61478 5460 61516
rect 4284 60958 4286 61010
rect 4338 60958 4340 61010
rect 4284 60946 4340 60958
rect 4464 60396 4728 60406
rect 4520 60340 4568 60396
rect 4624 60340 4672 60396
rect 4464 60330 4728 60340
rect 4060 60226 4228 60228
rect 4060 60174 4062 60226
rect 4114 60174 4228 60226
rect 4060 60172 4228 60174
rect 5180 60228 5236 60238
rect 4060 60162 4116 60172
rect 5180 60134 5236 60172
rect 2716 59890 2996 59892
rect 2716 59838 2718 59890
rect 2770 59838 2996 59890
rect 2716 59836 2996 59838
rect 3612 59892 3668 59902
rect 2716 59668 2772 59836
rect 3612 59798 3668 59836
rect 2156 59218 2324 59220
rect 2156 59166 2158 59218
rect 2210 59166 2324 59218
rect 2156 59164 2324 59166
rect 2380 59612 2772 59668
rect 3804 59612 4068 59622
rect 2156 59154 2212 59164
rect 1372 58902 1428 58940
rect 1484 58940 1652 58996
rect 1820 58996 1876 59006
rect 1372 58660 1428 58670
rect 1372 58566 1428 58604
rect 1260 58380 1428 58436
rect 1036 58146 1092 58156
rect 700 57820 1092 57876
rect 1036 57538 1092 57820
rect 1372 57650 1428 58380
rect 1372 57598 1374 57650
rect 1426 57598 1428 57650
rect 1372 57586 1428 57598
rect 1036 57486 1038 57538
rect 1090 57486 1092 57538
rect 1036 57474 1092 57486
rect 1260 56756 1316 56766
rect 252 55412 644 55468
rect 252 41412 308 41422
rect 252 31668 308 41356
rect 588 38668 644 55412
rect 1148 50820 1204 50830
rect 1148 50726 1204 50764
rect 812 50708 868 50718
rect 700 45892 756 45902
rect 700 40964 756 45836
rect 700 40898 756 40908
rect 588 38612 756 38668
rect 252 31602 308 31612
rect 364 29652 420 29662
rect 364 26292 420 29596
rect 364 26226 420 26236
rect 700 25620 756 38612
rect 364 25564 756 25620
rect 364 19908 420 25564
rect 812 25284 868 50652
rect 1036 50036 1092 50046
rect 1036 48356 1092 49980
rect 1260 49924 1316 56700
rect 1484 55468 1540 58940
rect 1820 58902 1876 58940
rect 1260 49858 1316 49868
rect 1372 55412 1540 55468
rect 1596 58772 1652 58782
rect 1036 48290 1092 48300
rect 1148 49588 1204 49598
rect 1148 45444 1204 49532
rect 1372 49364 1428 55412
rect 1484 53956 1540 53966
rect 1484 52724 1540 53900
rect 1596 52836 1652 58716
rect 1708 58546 1764 58558
rect 1708 58494 1710 58546
rect 1762 58494 1764 58546
rect 1708 57764 1764 58494
rect 2044 58436 2100 58446
rect 2044 58342 2100 58380
rect 1708 57698 1764 57708
rect 1932 58100 1988 58110
rect 1932 55412 1988 58044
rect 1596 52770 1652 52780
rect 1820 54964 1876 54974
rect 1484 52658 1540 52668
rect 1484 50708 1540 50718
rect 1484 50614 1540 50652
rect 1260 49308 1428 49364
rect 1484 49810 1540 49822
rect 1484 49758 1486 49810
rect 1538 49758 1540 49810
rect 1260 45780 1316 49308
rect 1372 49138 1428 49150
rect 1372 49086 1374 49138
rect 1426 49086 1428 49138
rect 1372 48580 1428 49086
rect 1372 48514 1428 48524
rect 1484 46788 1540 49758
rect 1596 49138 1652 49150
rect 1596 49086 1598 49138
rect 1650 49086 1652 49138
rect 1596 48468 1652 49086
rect 1596 48402 1652 48412
rect 1708 48356 1764 48366
rect 1708 48244 1764 48300
rect 1484 46674 1540 46732
rect 1484 46622 1486 46674
rect 1538 46622 1540 46674
rect 1484 46610 1540 46622
rect 1596 48188 1764 48244
rect 1596 46002 1652 48188
rect 1708 47458 1764 47470
rect 1708 47406 1710 47458
rect 1762 47406 1764 47458
rect 1708 46564 1764 47406
rect 1708 46498 1764 46508
rect 1820 46564 1876 54908
rect 1932 49698 1988 55356
rect 2156 54628 2212 54638
rect 2156 54534 2212 54572
rect 2044 50596 2100 50606
rect 2044 50502 2100 50540
rect 1932 49646 1934 49698
rect 1986 49646 1988 49698
rect 1932 49634 1988 49646
rect 2268 49252 2324 49262
rect 2268 49158 2324 49196
rect 1932 49028 1988 49038
rect 1932 48934 1988 48972
rect 2156 48468 2212 48478
rect 2156 48374 2212 48412
rect 2268 48132 2324 48142
rect 2044 48020 2100 48030
rect 1932 47572 1988 47582
rect 1932 47478 1988 47516
rect 1932 46564 1988 46574
rect 1820 46562 1988 46564
rect 1820 46510 1934 46562
rect 1986 46510 1988 46562
rect 1820 46508 1988 46510
rect 1820 46116 1876 46508
rect 1932 46498 1988 46508
rect 2044 46116 2100 47964
rect 2268 47796 2324 48076
rect 2268 47730 2324 47740
rect 1820 46050 1876 46060
rect 1932 46060 2100 46116
rect 2268 47572 2324 47582
rect 2268 47346 2324 47516
rect 2268 47294 2270 47346
rect 2322 47294 2324 47346
rect 1596 45950 1598 46002
rect 1650 45950 1652 46002
rect 1596 45892 1652 45950
rect 1596 45826 1652 45836
rect 1260 45778 1428 45780
rect 1260 45726 1262 45778
rect 1314 45726 1428 45778
rect 1260 45724 1428 45726
rect 1260 45714 1316 45724
rect 1148 45378 1204 45388
rect 1260 45108 1316 45118
rect 1372 45108 1428 45724
rect 1260 45106 1428 45108
rect 1260 45054 1262 45106
rect 1314 45054 1428 45106
rect 1260 45052 1428 45054
rect 1260 45042 1316 45052
rect 1260 44212 1316 44222
rect 1260 43652 1316 44156
rect 1148 43426 1204 43438
rect 1148 43374 1150 43426
rect 1202 43374 1204 43426
rect 1148 41860 1204 43374
rect 1036 41858 1204 41860
rect 1036 41806 1150 41858
rect 1202 41806 1204 41858
rect 1036 41804 1204 41806
rect 364 19842 420 19852
rect 700 25228 868 25284
rect 924 40852 980 40862
rect 588 19796 644 19806
rect 476 12852 532 12862
rect 364 11956 420 11966
rect 252 9940 308 9950
rect 252 5684 308 9884
rect 252 5618 308 5628
rect 364 4228 420 11900
rect 476 5348 532 12796
rect 476 5282 532 5292
rect 364 4162 420 4172
rect 588 2212 644 19740
rect 700 17444 756 25228
rect 924 25172 980 40796
rect 1036 35252 1092 41804
rect 1148 41794 1204 41804
rect 1260 39732 1316 43596
rect 1148 39676 1316 39732
rect 1148 39396 1204 39676
rect 1148 39330 1204 39340
rect 1260 39508 1316 39518
rect 1260 38946 1316 39452
rect 1260 38894 1262 38946
rect 1314 38894 1316 38946
rect 1260 38882 1316 38894
rect 1372 38050 1428 45052
rect 1708 45444 1764 45454
rect 1596 44884 1652 44894
rect 1484 44660 1540 44670
rect 1484 44100 1540 44604
rect 1484 39732 1540 44044
rect 1596 43538 1652 44828
rect 1708 44882 1764 45388
rect 1708 44830 1710 44882
rect 1762 44830 1764 44882
rect 1708 44772 1764 44830
rect 1708 44706 1764 44716
rect 1932 44548 1988 46060
rect 2268 45892 2324 47294
rect 1596 43486 1598 43538
rect 1650 43486 1652 43538
rect 1596 43474 1652 43486
rect 1708 44492 1988 44548
rect 2044 45836 2324 45892
rect 1596 41970 1652 41982
rect 1596 41918 1598 41970
rect 1650 41918 1652 41970
rect 1596 41636 1652 41918
rect 1596 41570 1652 41580
rect 1708 40514 1764 44492
rect 1932 44212 1988 44222
rect 2044 44212 2100 45836
rect 2380 45780 2436 59612
rect 3860 59556 3908 59612
rect 3964 59556 4012 59612
rect 3804 59546 4068 59556
rect 2492 59108 2548 59118
rect 2492 59014 2548 59052
rect 2828 59108 2884 59118
rect 2828 59014 2884 59052
rect 4464 58828 4728 58838
rect 4520 58772 4568 58828
rect 4624 58772 4672 58828
rect 4464 58762 4728 58772
rect 3804 58044 4068 58054
rect 3860 57988 3908 58044
rect 3964 57988 4012 58044
rect 3804 57978 4068 57988
rect 4464 57260 4728 57270
rect 4520 57204 4568 57260
rect 4624 57204 4672 57260
rect 4464 57194 4728 57204
rect 4844 56978 4900 56990
rect 4844 56926 4846 56978
rect 4898 56926 4900 56978
rect 2940 56756 2996 56766
rect 2492 55860 2548 55870
rect 2492 54402 2548 55804
rect 2492 54350 2494 54402
rect 2546 54350 2548 54402
rect 2492 54338 2548 54350
rect 2940 55298 2996 56700
rect 4396 56756 4452 56766
rect 3804 56476 4068 56486
rect 3860 56420 3908 56476
rect 3964 56420 4012 56476
rect 3804 56410 4068 56420
rect 3500 56308 3556 56318
rect 2940 55246 2942 55298
rect 2994 55246 2996 55298
rect 2940 54628 2996 55246
rect 2940 53730 2996 54572
rect 2940 53678 2942 53730
rect 2994 53678 2996 53730
rect 2492 53508 2548 53518
rect 2492 50818 2548 53452
rect 2492 50766 2494 50818
rect 2546 50766 2548 50818
rect 2492 50708 2548 50766
rect 2492 50642 2548 50652
rect 2604 52948 2660 52958
rect 2940 52948 2996 53678
rect 2604 52946 2996 52948
rect 2604 52894 2606 52946
rect 2658 52894 2996 52946
rect 2604 52892 2996 52894
rect 3276 55860 3332 55870
rect 2604 50484 2660 52892
rect 3052 52834 3108 52846
rect 3052 52782 3054 52834
rect 3106 52782 3108 52834
rect 3052 52164 3108 52782
rect 3276 52500 3332 55804
rect 3500 55410 3556 56252
rect 4396 56196 4452 56700
rect 4396 56130 4452 56140
rect 4844 56644 4900 56926
rect 4464 55692 4728 55702
rect 4520 55636 4568 55692
rect 4624 55636 4672 55692
rect 4464 55626 4728 55636
rect 3500 55358 3502 55410
rect 3554 55358 3556 55410
rect 3500 55346 3556 55358
rect 4620 55300 4676 55310
rect 4620 55206 4676 55244
rect 3804 54908 4068 54918
rect 3860 54852 3908 54908
rect 3964 54852 4012 54908
rect 3804 54842 4068 54852
rect 3724 54740 3780 54750
rect 3724 54646 3780 54684
rect 4464 54124 4728 54134
rect 4520 54068 4568 54124
rect 4624 54068 4672 54124
rect 4464 54058 4728 54068
rect 3500 53842 3556 53854
rect 3500 53790 3502 53842
rect 3554 53790 3556 53842
rect 3500 53508 3556 53790
rect 3500 53442 3556 53452
rect 4620 53508 4676 53518
rect 4620 53414 4676 53452
rect 3804 53340 4068 53350
rect 3860 53284 3908 53340
rect 3964 53284 4012 53340
rect 3804 53274 4068 53284
rect 4284 52724 4340 52734
rect 4284 52630 4340 52668
rect 4464 52556 4728 52566
rect 4520 52500 4568 52556
rect 4624 52500 4672 52556
rect 3276 52444 3444 52500
rect 4464 52490 4728 52500
rect 2940 52050 2996 52062
rect 2940 51998 2942 52050
rect 2994 51998 2996 52050
rect 2716 51380 2772 51390
rect 2716 51378 2884 51380
rect 2716 51326 2718 51378
rect 2770 51326 2884 51378
rect 2716 51324 2884 51326
rect 2716 51314 2772 51324
rect 2492 50428 2660 50484
rect 2828 50596 2884 51324
rect 2492 48020 2548 50428
rect 2604 50036 2660 50046
rect 2604 48132 2660 49980
rect 2716 48916 2772 48926
rect 2716 48822 2772 48860
rect 2604 48066 2660 48076
rect 2716 48692 2772 48702
rect 2492 47954 2548 47964
rect 2716 47684 2772 48636
rect 2828 48356 2884 50540
rect 2940 49588 2996 51998
rect 3052 51266 3108 52108
rect 3052 51214 3054 51266
rect 3106 51214 3108 51266
rect 3052 50428 3108 51214
rect 3276 52274 3332 52286
rect 3276 52222 3278 52274
rect 3330 52222 3332 52274
rect 3052 50372 3220 50428
rect 3164 49812 3220 50372
rect 3276 50036 3332 52222
rect 3276 49970 3332 49980
rect 3388 51268 3444 52444
rect 4508 52388 4564 52398
rect 4508 52294 4564 52332
rect 4844 52276 4900 56588
rect 4844 52210 4900 52220
rect 5068 55412 5124 55422
rect 3804 51772 4068 51782
rect 3860 51716 3908 51772
rect 3964 51716 4012 51772
rect 3804 51706 4068 51716
rect 4956 51492 5012 51502
rect 5068 51492 5124 55356
rect 5404 55298 5460 55310
rect 5404 55246 5406 55298
rect 5458 55246 5460 55298
rect 5404 54740 5460 55246
rect 5404 54674 5460 54684
rect 5292 53508 5348 53518
rect 4956 51490 5236 51492
rect 4956 51438 4958 51490
rect 5010 51438 5236 51490
rect 4956 51436 5236 51438
rect 4956 51426 5012 51436
rect 3164 49756 3332 49812
rect 3164 49588 3220 49598
rect 2940 49522 2996 49532
rect 3052 49586 3220 49588
rect 3052 49534 3166 49586
rect 3218 49534 3220 49586
rect 3052 49532 3220 49534
rect 3052 49028 3108 49532
rect 3164 49522 3220 49532
rect 3276 49140 3332 49756
rect 3276 49074 3332 49084
rect 2828 48290 2884 48300
rect 2940 49026 3108 49028
rect 2940 48974 3054 49026
rect 3106 48974 3108 49026
rect 2940 48972 3108 48974
rect 2716 47628 2884 47684
rect 2716 47460 2772 47470
rect 2716 47236 2772 47404
rect 2716 47170 2772 47180
rect 2828 46900 2884 47628
rect 2940 47572 2996 48972
rect 3052 48962 3108 48972
rect 3276 48580 3332 48590
rect 2940 47506 2996 47516
rect 3052 48020 3108 48030
rect 3052 47458 3108 47964
rect 3276 47682 3332 48524
rect 3388 48130 3444 51212
rect 4284 51156 4340 51166
rect 4284 51062 4340 51100
rect 4464 50988 4728 50998
rect 4520 50932 4568 50988
rect 4624 50932 4672 50988
rect 4464 50922 4728 50932
rect 5068 50820 5124 50830
rect 5068 50726 5124 50764
rect 3612 50708 3668 50718
rect 3612 50706 4228 50708
rect 3612 50654 3614 50706
rect 3666 50654 4228 50706
rect 3612 50652 4228 50654
rect 3612 50642 3668 50652
rect 4172 50596 4228 50652
rect 4396 50596 4452 50606
rect 4172 50594 4452 50596
rect 4172 50542 4398 50594
rect 4450 50542 4452 50594
rect 4172 50540 4452 50542
rect 4396 50530 4452 50540
rect 4956 50596 5012 50606
rect 4060 50484 4116 50522
rect 4956 50502 5012 50540
rect 4060 50418 4116 50428
rect 5180 50428 5236 51436
rect 5292 51378 5348 53452
rect 5516 53284 5572 68012
rect 5852 67844 5908 69468
rect 6076 69522 6132 69534
rect 6076 69470 6078 69522
rect 6130 69470 6132 69522
rect 5964 68852 6020 68862
rect 5964 68066 6020 68796
rect 5964 68014 5966 68066
rect 6018 68014 6020 68066
rect 5964 68002 6020 68014
rect 6076 67844 6132 69470
rect 5740 67842 5908 67844
rect 5740 67790 5854 67842
rect 5906 67790 5908 67842
rect 5740 67788 5908 67790
rect 5628 64818 5684 64830
rect 5628 64766 5630 64818
rect 5682 64766 5684 64818
rect 5628 63700 5684 64766
rect 5740 64708 5796 67788
rect 5852 67778 5908 67788
rect 5964 67788 6132 67844
rect 6188 68180 6244 68190
rect 5964 66612 6020 67788
rect 5964 66546 6020 66556
rect 6076 67620 6132 67630
rect 6076 66498 6132 67564
rect 6076 66446 6078 66498
rect 6130 66446 6132 66498
rect 6076 66434 6132 66446
rect 5964 66388 6020 66398
rect 5852 66276 5908 66286
rect 5852 66182 5908 66220
rect 5852 65604 5908 65614
rect 5852 65510 5908 65548
rect 5964 64930 6020 66332
rect 5964 64878 5966 64930
rect 6018 64878 6020 64930
rect 5964 64866 6020 64878
rect 6076 65940 6132 65950
rect 5740 64642 5796 64652
rect 5628 63634 5684 63644
rect 5628 63252 5684 63262
rect 5628 62466 5684 63196
rect 5740 63140 5796 63150
rect 5740 63046 5796 63084
rect 6076 62916 6132 65884
rect 5628 62414 5630 62466
rect 5682 62414 5684 62466
rect 5628 62020 5684 62414
rect 5628 60898 5684 61964
rect 5628 60846 5630 60898
rect 5682 60846 5684 60898
rect 5628 60834 5684 60846
rect 5740 62860 6132 62916
rect 5740 60900 5796 62860
rect 6076 62468 6132 62478
rect 5964 62356 6020 62366
rect 5964 62262 6020 62300
rect 6076 62188 6132 62412
rect 5964 62132 6132 62188
rect 5964 61570 6020 62132
rect 6076 61796 6132 61806
rect 6076 61702 6132 61740
rect 5964 61518 5966 61570
rect 6018 61518 6020 61570
rect 5964 61506 6020 61518
rect 5740 60844 5908 60900
rect 5852 60116 5908 60844
rect 5964 60786 6020 60798
rect 5964 60734 5966 60786
rect 6018 60734 6020 60786
rect 5964 60228 6020 60734
rect 5964 60162 6020 60172
rect 5628 60060 5908 60116
rect 5628 54740 5684 60060
rect 5852 59892 5908 59902
rect 5852 59798 5908 59836
rect 6188 56868 6244 68124
rect 6300 65940 6356 71372
rect 6524 68852 6580 73164
rect 6636 73106 6692 73118
rect 6636 73054 6638 73106
rect 6690 73054 6692 73106
rect 6636 72660 6692 73054
rect 6636 72594 6692 72604
rect 6636 72324 6692 72334
rect 6636 70978 6692 72268
rect 6636 70926 6638 70978
rect 6690 70926 6692 70978
rect 6636 70914 6692 70926
rect 6748 69970 6804 74620
rect 6860 74114 6916 74126
rect 6860 74062 6862 74114
rect 6914 74062 6916 74114
rect 6860 74004 6916 74062
rect 6860 73938 6916 73948
rect 6972 73108 7028 76524
rect 7196 77810 7252 77822
rect 7196 77758 7198 77810
rect 7250 77758 7252 77810
rect 7084 76468 7140 76478
rect 7196 76468 7252 77758
rect 7420 77812 7476 81340
rect 7420 77746 7476 77756
rect 7532 77140 7588 81902
rect 7868 80946 7924 80958
rect 7868 80894 7870 80946
rect 7922 80894 7924 80946
rect 7868 79604 7924 80894
rect 7868 79538 7924 79548
rect 7756 79378 7812 79390
rect 7756 79326 7758 79378
rect 7810 79326 7812 79378
rect 7756 77588 7812 79326
rect 7980 78484 8036 82014
rect 8092 81284 8148 83470
rect 8092 80386 8148 81228
rect 8092 80334 8094 80386
rect 8146 80334 8148 80386
rect 8092 80322 8148 80334
rect 8092 79378 8148 79390
rect 8092 79326 8094 79378
rect 8146 79326 8148 79378
rect 8092 79268 8148 79326
rect 8092 79202 8148 79212
rect 7980 78418 8036 78428
rect 8092 78594 8148 78606
rect 8092 78542 8094 78594
rect 8146 78542 8148 78594
rect 7868 78036 7924 78074
rect 7868 77970 7924 77980
rect 7756 77522 7812 77532
rect 7868 77812 7924 77822
rect 7532 77074 7588 77084
rect 7756 77026 7812 77038
rect 7756 76974 7758 77026
rect 7810 76974 7812 77026
rect 7084 76466 7252 76468
rect 7084 76414 7086 76466
rect 7138 76414 7252 76466
rect 7084 76412 7252 76414
rect 7420 76466 7476 76478
rect 7420 76414 7422 76466
rect 7474 76414 7476 76466
rect 7084 76402 7140 76412
rect 7084 75908 7140 75918
rect 7084 75814 7140 75852
rect 7196 74228 7252 74238
rect 7084 74226 7252 74228
rect 7084 74174 7198 74226
rect 7250 74174 7252 74226
rect 7084 74172 7252 74174
rect 7084 73892 7140 74172
rect 7196 74162 7252 74172
rect 7420 74228 7476 76414
rect 7644 76356 7700 76366
rect 7644 76262 7700 76300
rect 7644 74674 7700 74686
rect 7644 74622 7646 74674
rect 7698 74622 7700 74674
rect 7532 74340 7588 74350
rect 7532 74246 7588 74284
rect 7084 73826 7140 73836
rect 7196 73780 7252 73790
rect 7196 73330 7252 73724
rect 7420 73668 7476 74172
rect 7420 73602 7476 73612
rect 7196 73278 7198 73330
rect 7250 73278 7252 73330
rect 7196 73266 7252 73278
rect 6972 73052 7364 73108
rect 7196 72884 7252 72894
rect 6972 71762 7028 71774
rect 6972 71710 6974 71762
rect 7026 71710 7028 71762
rect 6748 69918 6750 69970
rect 6802 69918 6804 69970
rect 6748 69636 6804 69918
rect 6748 69570 6804 69580
rect 6860 70868 6916 70878
rect 6524 67172 6580 68796
rect 6636 69188 6692 69198
rect 6636 67842 6692 69132
rect 6636 67790 6638 67842
rect 6690 67790 6692 67842
rect 6636 67778 6692 67790
rect 6748 68402 6804 68414
rect 6748 68350 6750 68402
rect 6802 68350 6804 68402
rect 6748 67284 6804 68350
rect 6300 65874 6356 65884
rect 6412 66276 6468 66286
rect 6300 65266 6356 65278
rect 6300 65214 6302 65266
rect 6354 65214 6356 65266
rect 6300 65156 6356 65214
rect 6300 65090 6356 65100
rect 6300 63700 6356 63710
rect 6300 63362 6356 63644
rect 6300 63310 6302 63362
rect 6354 63310 6356 63362
rect 6300 63298 6356 63310
rect 6412 62356 6468 66220
rect 6524 65604 6580 67116
rect 6636 67228 6804 67284
rect 6636 66274 6692 67228
rect 6636 66222 6638 66274
rect 6690 66222 6692 66274
rect 6636 66210 6692 66222
rect 6524 65538 6580 65548
rect 6524 64706 6580 64718
rect 6524 64654 6526 64706
rect 6578 64654 6580 64706
rect 6524 63922 6580 64654
rect 6524 63870 6526 63922
rect 6578 63870 6580 63922
rect 6524 63140 6580 63870
rect 6524 63074 6580 63084
rect 6412 60786 6468 62300
rect 6524 62916 6580 62926
rect 6524 61682 6580 62860
rect 6636 62244 6692 62282
rect 6636 62178 6692 62188
rect 6524 61630 6526 61682
rect 6578 61630 6580 61682
rect 6524 61618 6580 61630
rect 6412 60734 6414 60786
rect 6466 60734 6468 60786
rect 6412 60722 6468 60734
rect 6636 60676 6692 60686
rect 6636 60582 6692 60620
rect 6300 60116 6356 60126
rect 6300 60022 6356 60060
rect 6636 56868 6692 56878
rect 5740 56812 6468 56868
rect 5740 55636 5796 56812
rect 5964 56642 6020 56654
rect 5964 56590 5966 56642
rect 6018 56590 6020 56642
rect 5852 56196 5908 56206
rect 5852 56102 5908 56140
rect 5740 55580 5908 55636
rect 5628 54674 5684 54684
rect 5740 55412 5796 55422
rect 5740 54626 5796 55356
rect 5740 54574 5742 54626
rect 5794 54574 5796 54626
rect 5740 54562 5796 54574
rect 5852 55298 5908 55580
rect 5852 55246 5854 55298
rect 5906 55246 5908 55298
rect 5516 53218 5572 53228
rect 5292 51326 5294 51378
rect 5346 51326 5348 51378
rect 5292 51314 5348 51326
rect 5628 52052 5684 52062
rect 5516 51156 5572 51166
rect 5516 50706 5572 51100
rect 5516 50654 5518 50706
rect 5570 50654 5572 50706
rect 5516 50642 5572 50654
rect 5628 50484 5684 51996
rect 5852 51380 5908 55246
rect 5964 54516 6020 56590
rect 6300 55858 6356 55870
rect 6300 55806 6302 55858
rect 6354 55806 6356 55858
rect 6076 55412 6132 55422
rect 6076 55410 6244 55412
rect 6076 55358 6078 55410
rect 6130 55358 6244 55410
rect 6076 55356 6244 55358
rect 6076 55346 6132 55356
rect 6076 54516 6132 54526
rect 5964 54514 6132 54516
rect 5964 54462 6078 54514
rect 6130 54462 6132 54514
rect 5964 54460 6132 54462
rect 6076 54450 6132 54460
rect 5852 51378 6132 51380
rect 5852 51326 5854 51378
rect 5906 51326 6132 51378
rect 5852 51324 6132 51326
rect 5852 51314 5908 51324
rect 5180 50372 5572 50428
rect 3804 50204 4068 50214
rect 3860 50148 3908 50204
rect 3964 50148 4012 50204
rect 3804 50138 4068 50148
rect 4956 49924 5012 49934
rect 4464 49420 4728 49430
rect 4520 49364 4568 49420
rect 4624 49364 4672 49420
rect 4464 49354 4728 49364
rect 3724 49138 3780 49150
rect 3724 49086 3726 49138
rect 3778 49086 3780 49138
rect 3612 49026 3668 49038
rect 3612 48974 3614 49026
rect 3666 48974 3668 49026
rect 3612 48804 3668 48974
rect 3724 49028 3780 49086
rect 3724 48962 3780 48972
rect 4172 49026 4228 49038
rect 4172 48974 4174 49026
rect 4226 48974 4228 49026
rect 3612 48738 3668 48748
rect 3804 48636 4068 48646
rect 3860 48580 3908 48636
rect 3964 48580 4012 48636
rect 3804 48570 4068 48580
rect 3612 48356 3668 48366
rect 3388 48078 3390 48130
rect 3442 48078 3444 48130
rect 3388 48066 3444 48078
rect 3500 48244 3556 48254
rect 3276 47630 3278 47682
rect 3330 47630 3332 47682
rect 3276 47618 3332 47630
rect 3052 47406 3054 47458
rect 3106 47406 3108 47458
rect 3052 47394 3108 47406
rect 3164 47236 3220 47246
rect 2828 46844 3108 46900
rect 2268 45724 2436 45780
rect 2940 46676 2996 46686
rect 1932 44210 2100 44212
rect 1932 44158 1934 44210
rect 1986 44158 2100 44210
rect 1932 44156 2100 44158
rect 2156 45668 2212 45678
rect 1932 42644 1988 44156
rect 1932 42550 1988 42588
rect 2044 43540 2100 43550
rect 1932 41972 1988 41982
rect 2044 41972 2100 43484
rect 2156 43426 2212 45612
rect 2156 43374 2158 43426
rect 2210 43374 2212 43426
rect 2156 43362 2212 43374
rect 1708 40462 1710 40514
rect 1762 40462 1764 40514
rect 1596 39732 1652 39742
rect 1484 39730 1652 39732
rect 1484 39678 1598 39730
rect 1650 39678 1652 39730
rect 1484 39676 1652 39678
rect 1596 39666 1652 39676
rect 1708 39508 1764 40462
rect 1708 39442 1764 39452
rect 1820 41970 2100 41972
rect 1820 41918 1934 41970
rect 1986 41918 2100 41970
rect 1820 41916 2100 41918
rect 1372 37998 1374 38050
rect 1426 37998 1428 38050
rect 1372 37986 1428 37998
rect 1596 39396 1652 39406
rect 1596 38722 1652 39340
rect 1596 38670 1598 38722
rect 1650 38670 1652 38722
rect 1484 37938 1540 37950
rect 1484 37886 1486 37938
rect 1538 37886 1540 37938
rect 1484 37380 1540 37886
rect 1484 37314 1540 37324
rect 1484 36484 1540 36494
rect 1484 36390 1540 36428
rect 1148 35812 1204 35822
rect 1148 35718 1204 35756
rect 1484 35700 1540 35710
rect 1036 35186 1092 35196
rect 1260 35698 1540 35700
rect 1260 35646 1486 35698
rect 1538 35646 1540 35698
rect 1260 35644 1540 35646
rect 1148 32788 1204 32798
rect 1148 32694 1204 32732
rect 1148 29652 1204 29662
rect 1260 29652 1316 35644
rect 1484 35634 1540 35644
rect 1148 29650 1316 29652
rect 1148 29598 1150 29650
rect 1202 29598 1316 29650
rect 1148 29596 1316 29598
rect 1372 32228 1428 32238
rect 1148 29586 1204 29596
rect 1260 28644 1316 28654
rect 1148 27972 1204 27982
rect 1148 27878 1204 27916
rect 1260 26402 1316 28588
rect 1260 26350 1262 26402
rect 1314 26350 1316 26402
rect 1260 26338 1316 26350
rect 812 25116 980 25172
rect 1148 25284 1204 25294
rect 812 23380 868 25116
rect 1036 24052 1092 24062
rect 812 23314 868 23324
rect 924 24050 1092 24052
rect 924 23998 1038 24050
rect 1090 23998 1092 24050
rect 924 23996 1092 23998
rect 700 17378 756 17388
rect 812 23044 868 23054
rect 812 15204 868 22988
rect 924 20468 980 23996
rect 1036 23986 1092 23996
rect 1036 22930 1092 22942
rect 1036 22878 1038 22930
rect 1090 22878 1092 22930
rect 1036 21364 1092 22878
rect 1036 21298 1092 21308
rect 924 20402 980 20412
rect 1148 20356 1204 25228
rect 1260 24724 1316 24734
rect 1260 23716 1316 24668
rect 1372 24162 1428 32172
rect 1596 31332 1652 38670
rect 1820 37044 1876 41916
rect 1932 41906 1988 41916
rect 2268 41860 2324 45724
rect 2828 45668 2884 45678
rect 2380 45666 2884 45668
rect 2380 45614 2830 45666
rect 2882 45614 2884 45666
rect 2380 45612 2884 45614
rect 2380 44324 2436 45612
rect 2828 45602 2884 45612
rect 2828 44884 2884 44894
rect 2828 44790 2884 44828
rect 2940 44546 2996 46620
rect 2940 44494 2942 44546
rect 2994 44494 2996 44546
rect 2940 44482 2996 44494
rect 2380 44322 2660 44324
rect 2380 44270 2382 44322
rect 2434 44270 2660 44322
rect 2380 44268 2660 44270
rect 2380 44258 2436 44268
rect 2604 43538 2660 44268
rect 2604 43486 2606 43538
rect 2658 43486 2660 43538
rect 2604 43474 2660 43486
rect 2828 44322 2884 44334
rect 2828 44270 2830 44322
rect 2882 44270 2884 44322
rect 2380 42754 2436 42766
rect 2380 42702 2382 42754
rect 2434 42702 2436 42754
rect 2380 41972 2436 42702
rect 2828 42754 2884 44270
rect 2828 42702 2830 42754
rect 2882 42702 2884 42754
rect 2716 41972 2772 41982
rect 2380 41970 2772 41972
rect 2380 41918 2718 41970
rect 2770 41918 2772 41970
rect 2380 41916 2772 41918
rect 2268 41804 2436 41860
rect 2156 41748 2212 41758
rect 2156 41654 2212 41692
rect 2380 41636 2436 41804
rect 2268 41580 2436 41636
rect 2604 41636 2660 41646
rect 2044 40292 2100 40302
rect 2044 40198 2100 40236
rect 1932 38164 1988 38174
rect 1932 38070 1988 38108
rect 2268 37380 2324 41580
rect 2380 40628 2436 40638
rect 2380 38668 2436 40572
rect 2604 39060 2660 41580
rect 2716 39844 2772 41916
rect 2828 41860 2884 42702
rect 2940 42866 2996 42878
rect 2940 42814 2942 42866
rect 2994 42814 2996 42866
rect 2940 42084 2996 42814
rect 2940 42018 2996 42028
rect 2828 41804 2996 41860
rect 2828 41074 2884 41086
rect 2828 41022 2830 41074
rect 2882 41022 2884 41074
rect 2828 40292 2884 41022
rect 2940 41076 2996 41804
rect 2940 41010 2996 41020
rect 2828 40226 2884 40236
rect 2828 39844 2884 39854
rect 2716 39842 2884 39844
rect 2716 39790 2830 39842
rect 2882 39790 2884 39842
rect 2716 39788 2884 39790
rect 2828 39778 2884 39788
rect 2828 39060 2884 39070
rect 2604 39058 2884 39060
rect 2604 39006 2830 39058
rect 2882 39006 2884 39058
rect 2604 39004 2884 39006
rect 2828 38994 2884 39004
rect 2828 38724 2884 38734
rect 3052 38668 3108 46844
rect 3164 46898 3220 47180
rect 3164 46846 3166 46898
rect 3218 46846 3220 46898
rect 3164 46834 3220 46846
rect 3500 46788 3556 48188
rect 3500 46722 3556 46732
rect 3612 47348 3668 48300
rect 3724 48244 3780 48254
rect 3724 48150 3780 48188
rect 4060 48020 4116 48030
rect 3724 47572 3780 47582
rect 3724 47478 3780 47516
rect 3388 44884 3444 44894
rect 3388 44434 3444 44828
rect 3388 44382 3390 44434
rect 3442 44382 3444 44434
rect 3388 44370 3444 44382
rect 3164 43538 3220 43550
rect 3164 43486 3166 43538
rect 3218 43486 3220 43538
rect 3164 41970 3220 43486
rect 3164 41918 3166 41970
rect 3218 41918 3220 41970
rect 3164 41860 3220 41918
rect 3164 41794 3220 41804
rect 3388 42754 3444 42766
rect 3388 42702 3390 42754
rect 3442 42702 3444 42754
rect 3388 41636 3444 42702
rect 3388 41570 3444 41580
rect 3276 41524 3332 41534
rect 3276 41410 3332 41468
rect 3276 41358 3278 41410
rect 3330 41358 3332 41410
rect 3276 41346 3332 41358
rect 3388 41188 3444 41198
rect 3276 40404 3332 40414
rect 3276 40310 3332 40348
rect 2380 38612 2660 38668
rect 2268 37324 2436 37380
rect 1932 37268 1988 37278
rect 1932 37174 1988 37212
rect 2156 37044 2212 37054
rect 1820 36978 1876 36988
rect 1932 37042 2212 37044
rect 1932 36990 2158 37042
rect 2210 36990 2212 37042
rect 1932 36988 2212 36990
rect 1820 36482 1876 36494
rect 1820 36430 1822 36482
rect 1874 36430 1876 36482
rect 1708 34914 1764 34926
rect 1708 34862 1710 34914
rect 1762 34862 1764 34914
rect 1708 34804 1764 34862
rect 1708 34738 1764 34748
rect 1820 33684 1876 36430
rect 1708 33628 1876 33684
rect 1708 32788 1764 33628
rect 1708 32722 1764 32732
rect 1820 33458 1876 33470
rect 1820 33406 1822 33458
rect 1874 33406 1876 33458
rect 1820 32228 1876 33406
rect 1820 32162 1876 32172
rect 1484 31276 1652 31332
rect 1708 31892 1764 31902
rect 1932 31892 1988 36988
rect 2156 36978 2212 36988
rect 2268 36482 2324 36494
rect 2268 36430 2270 36482
rect 2322 36430 2324 36482
rect 2268 36372 2324 36430
rect 2044 35698 2100 35710
rect 2044 35646 2046 35698
rect 2098 35646 2100 35698
rect 2044 34580 2100 35646
rect 2044 34514 2100 34524
rect 2156 35474 2212 35486
rect 2156 35422 2158 35474
rect 2210 35422 2212 35474
rect 1484 28868 1540 31276
rect 1708 31220 1764 31836
rect 1596 31164 1764 31220
rect 1820 31836 1988 31892
rect 2044 33796 2100 33806
rect 1596 30994 1652 31164
rect 1596 30942 1598 30994
rect 1650 30942 1652 30994
rect 1596 30436 1652 30942
rect 1596 30370 1652 30380
rect 1708 30996 1764 31006
rect 1484 28802 1540 28812
rect 1708 28644 1764 30940
rect 1820 29204 1876 31836
rect 1932 31668 1988 31678
rect 1932 31574 1988 31612
rect 2044 31108 2100 33740
rect 2156 33684 2212 35422
rect 2156 33618 2212 33628
rect 2156 33460 2212 33470
rect 2156 33366 2212 33404
rect 2268 33236 2324 36316
rect 2380 34468 2436 37324
rect 2492 37268 2548 37278
rect 2492 36706 2548 37212
rect 2492 36654 2494 36706
rect 2546 36654 2548 36706
rect 2492 36642 2548 36654
rect 2604 36372 2660 38612
rect 2716 37380 2772 37390
rect 2716 37286 2772 37324
rect 2604 36306 2660 36316
rect 2716 35698 2772 35710
rect 2716 35646 2718 35698
rect 2770 35646 2772 35698
rect 2716 35252 2772 35646
rect 2716 35186 2772 35196
rect 2716 34916 2772 34926
rect 2828 34916 2884 38668
rect 2940 38612 3108 38668
rect 2940 36708 2996 38612
rect 3052 37828 3108 37838
rect 3052 37734 3108 37772
rect 3164 37044 3220 37054
rect 3164 36950 3220 36988
rect 2940 36652 3108 36708
rect 2716 34914 2884 34916
rect 2716 34862 2718 34914
rect 2770 34862 2884 34914
rect 2716 34860 2884 34862
rect 2940 36482 2996 36494
rect 2940 36430 2942 36482
rect 2994 36430 2996 36482
rect 2380 34412 2660 34468
rect 2380 34244 2436 34254
rect 2380 34150 2436 34188
rect 2156 33180 2324 33236
rect 2380 33796 2436 33806
rect 2156 31668 2212 33180
rect 2380 32450 2436 33740
rect 2604 33684 2660 34412
rect 2380 32398 2382 32450
rect 2434 32398 2436 32450
rect 2380 32386 2436 32398
rect 2492 33628 2660 33684
rect 2492 31892 2548 33628
rect 2604 33460 2660 33470
rect 2716 33460 2772 34860
rect 2940 34244 2996 36430
rect 2940 34178 2996 34188
rect 2604 33458 2772 33460
rect 2604 33406 2606 33458
rect 2658 33406 2772 33458
rect 2604 33404 2772 33406
rect 2604 33394 2660 33404
rect 2940 33346 2996 33358
rect 2940 33294 2942 33346
rect 2994 33294 2996 33346
rect 2828 32562 2884 32574
rect 2828 32510 2830 32562
rect 2882 32510 2884 32562
rect 2828 32452 2884 32510
rect 2828 32386 2884 32396
rect 2940 32116 2996 33294
rect 2492 31826 2548 31836
rect 2828 32060 2996 32116
rect 2156 31602 2212 31612
rect 2268 31780 2324 31790
rect 2268 31220 2324 31724
rect 2380 31778 2436 31790
rect 2380 31726 2382 31778
rect 2434 31726 2436 31778
rect 2380 31332 2436 31726
rect 2716 31780 2772 31818
rect 2716 31714 2772 31724
rect 2716 31556 2772 31566
rect 2380 31276 2660 31332
rect 2268 31164 2436 31220
rect 2044 30882 2100 31052
rect 2044 30830 2046 30882
rect 2098 30830 2100 30882
rect 2044 30818 2100 30830
rect 1820 29138 1876 29148
rect 2044 29988 2100 29998
rect 1708 28550 1764 28588
rect 1484 27972 1540 27982
rect 1484 27186 1540 27916
rect 1484 27134 1486 27186
rect 1538 27134 1540 27186
rect 1484 27122 1540 27134
rect 1596 27858 1652 27870
rect 1596 27806 1598 27858
rect 1650 27806 1652 27858
rect 1596 26908 1652 27806
rect 2044 27858 2100 29932
rect 2268 29316 2324 29326
rect 2268 29222 2324 29260
rect 2156 28868 2212 28878
rect 2156 28774 2212 28812
rect 2044 27806 2046 27858
rect 2098 27806 2100 27858
rect 2044 27794 2100 27806
rect 1932 27748 1988 27758
rect 1372 24110 1374 24162
rect 1426 24110 1428 24162
rect 1372 24098 1428 24110
rect 1484 26852 1652 26908
rect 1820 27074 1876 27086
rect 1820 27022 1822 27074
rect 1874 27022 1876 27074
rect 1260 23650 1316 23660
rect 1036 20300 1204 20356
rect 1260 23154 1316 23166
rect 1260 23102 1262 23154
rect 1314 23102 1316 23154
rect 1260 20356 1316 23102
rect 1372 21700 1428 21710
rect 1372 21606 1428 21644
rect 1036 20244 1092 20300
rect 1260 20290 1316 20300
rect 924 20188 1092 20244
rect 1484 20188 1540 26852
rect 1708 26516 1764 26526
rect 1596 26180 1652 26190
rect 1596 24610 1652 26124
rect 1708 24724 1764 26460
rect 1820 25284 1876 27022
rect 1932 26516 1988 27692
rect 2156 27634 2212 27646
rect 2156 27582 2158 27634
rect 2210 27582 2212 27634
rect 2156 27412 2212 27582
rect 2156 27346 2212 27356
rect 1932 26450 1988 26460
rect 2380 27074 2436 31164
rect 2492 30436 2548 30446
rect 2492 30100 2548 30380
rect 2492 29540 2548 30044
rect 2492 27748 2548 29484
rect 2492 27682 2548 27692
rect 2380 27022 2382 27074
rect 2434 27022 2436 27074
rect 1820 25218 1876 25228
rect 1932 26292 1988 26302
rect 1708 24658 1764 24668
rect 1596 24558 1598 24610
rect 1650 24558 1652 24610
rect 1596 23044 1652 24558
rect 1932 24052 1988 26236
rect 2156 25508 2212 25518
rect 2156 25414 2212 25452
rect 2380 24276 2436 27022
rect 2492 27186 2548 27198
rect 2492 27134 2494 27186
rect 2546 27134 2548 27186
rect 2492 26964 2548 27134
rect 2492 26898 2548 26908
rect 2604 24948 2660 31276
rect 2716 30322 2772 31500
rect 2716 30270 2718 30322
rect 2770 30270 2772 30322
rect 2716 30258 2772 30270
rect 2716 29540 2772 29550
rect 2716 29446 2772 29484
rect 2716 27858 2772 27870
rect 2716 27806 2718 27858
rect 2770 27806 2772 27858
rect 2716 25172 2772 27806
rect 2828 26514 2884 32060
rect 2940 31892 2996 31902
rect 2940 31798 2996 31836
rect 3052 31780 3108 36652
rect 3388 36484 3444 41132
rect 3276 35700 3332 35710
rect 3388 35700 3444 36428
rect 3500 41076 3556 41086
rect 3500 36482 3556 41020
rect 3500 36430 3502 36482
rect 3554 36430 3556 36482
rect 3500 36418 3556 36430
rect 3612 35924 3668 47292
rect 4060 47236 4116 47964
rect 4172 47460 4228 48974
rect 4844 49026 4900 49038
rect 4844 48974 4846 49026
rect 4898 48974 4900 49026
rect 4464 47852 4728 47862
rect 4520 47796 4568 47852
rect 4624 47796 4672 47852
rect 4464 47786 4728 47796
rect 4172 47394 4228 47404
rect 4284 47458 4340 47470
rect 4284 47406 4286 47458
rect 4338 47406 4340 47458
rect 4060 47180 4228 47236
rect 3804 47068 4068 47078
rect 3860 47012 3908 47068
rect 3964 47012 4012 47068
rect 3804 47002 4068 47012
rect 3804 45500 4068 45510
rect 3860 45444 3908 45500
rect 3964 45444 4012 45500
rect 3804 45434 4068 45444
rect 4172 44322 4228 47180
rect 4172 44270 4174 44322
rect 4226 44270 4228 44322
rect 3804 43932 4068 43942
rect 3860 43876 3908 43932
rect 3964 43876 4012 43932
rect 3804 43866 4068 43876
rect 4172 43764 4228 44270
rect 4060 43708 4228 43764
rect 4060 42756 4116 43708
rect 4172 43538 4228 43550
rect 4172 43486 4174 43538
rect 4226 43486 4228 43538
rect 4172 42868 4228 43486
rect 4284 43540 4340 47406
rect 4844 47124 4900 48974
rect 4956 48804 5012 49868
rect 5292 49588 5348 49598
rect 4956 48738 5012 48748
rect 5068 48916 5124 48926
rect 4844 47058 4900 47068
rect 5068 47012 5124 48860
rect 5068 46946 5124 46956
rect 4956 46788 5012 46798
rect 4464 46284 4728 46294
rect 4520 46228 4568 46284
rect 4624 46228 4672 46284
rect 4464 46218 4728 46228
rect 4844 46002 4900 46014
rect 4844 45950 4846 46002
rect 4898 45950 4900 46002
rect 4844 45892 4900 45950
rect 4844 45826 4900 45836
rect 4396 45778 4452 45790
rect 4396 45726 4398 45778
rect 4450 45726 4452 45778
rect 4396 45556 4452 45726
rect 4396 45490 4452 45500
rect 4956 45444 5012 46732
rect 5180 46674 5236 46686
rect 5180 46622 5182 46674
rect 5234 46622 5236 46674
rect 5068 46562 5124 46574
rect 5068 46510 5070 46562
rect 5122 46510 5124 46562
rect 5068 45668 5124 46510
rect 5068 45602 5124 45612
rect 4956 45378 5012 45388
rect 4464 44716 4728 44726
rect 4520 44660 4568 44716
rect 4624 44660 4672 44716
rect 4464 44650 4728 44660
rect 4284 43474 4340 43484
rect 4956 44322 5012 44334
rect 4956 44270 4958 44322
rect 5010 44270 5012 44322
rect 4956 43764 5012 44270
rect 4464 43148 4728 43158
rect 4520 43092 4568 43148
rect 4624 43092 4672 43148
rect 4464 43082 4728 43092
rect 4172 42812 4452 42868
rect 4060 42754 4340 42756
rect 4060 42702 4062 42754
rect 4114 42702 4340 42754
rect 4060 42700 4340 42702
rect 4060 42690 4116 42700
rect 3804 42364 4068 42374
rect 3860 42308 3908 42364
rect 3964 42308 4012 42364
rect 3804 42298 4068 42308
rect 4172 41972 4228 41982
rect 4172 41412 4228 41916
rect 4172 41346 4228 41356
rect 4284 41860 4340 42700
rect 4396 41972 4452 42812
rect 4956 42756 5012 43708
rect 4396 41906 4452 41916
rect 4844 42754 5012 42756
rect 4844 42702 4958 42754
rect 5010 42702 5012 42754
rect 4844 42700 5012 42702
rect 3804 40796 4068 40806
rect 3860 40740 3908 40796
rect 3964 40740 4012 40796
rect 3804 40730 4068 40740
rect 3804 39228 4068 39238
rect 3860 39172 3908 39228
rect 3964 39172 4012 39228
rect 3804 39162 4068 39172
rect 4284 38724 4340 41804
rect 4844 41748 4900 42700
rect 4956 42690 5012 42700
rect 4956 41972 5012 41982
rect 4956 41878 5012 41916
rect 5068 41748 5124 41758
rect 4844 41692 5012 41748
rect 4464 41580 4728 41590
rect 4520 41524 4568 41580
rect 4624 41524 4672 41580
rect 4464 41514 4728 41524
rect 4396 41412 4452 41422
rect 4396 41318 4452 41356
rect 4844 41188 4900 41198
rect 4844 41094 4900 41132
rect 4956 40964 5012 41692
rect 4844 40908 5012 40964
rect 4464 40012 4728 40022
rect 4520 39956 4568 40012
rect 4624 39956 4672 40012
rect 4464 39946 4728 39956
rect 4844 38836 4900 40908
rect 4956 40292 5012 40302
rect 4956 39620 5012 40236
rect 5068 40290 5124 41692
rect 5180 40964 5236 46622
rect 5292 45892 5348 49532
rect 5404 47460 5460 47470
rect 5404 47366 5460 47404
rect 5292 45556 5348 45836
rect 5292 43650 5348 45500
rect 5516 44996 5572 50372
rect 5628 45108 5684 50428
rect 5964 51154 6020 51166
rect 5964 51102 5966 51154
rect 6018 51102 6020 51154
rect 5852 49028 5908 49038
rect 5852 48934 5908 48972
rect 5964 48244 6020 51102
rect 6076 50596 6132 51324
rect 6076 50502 6132 50540
rect 6188 48916 6244 55356
rect 6300 54404 6356 55806
rect 6412 54516 6468 56812
rect 6636 56196 6692 56812
rect 6860 56308 6916 70812
rect 6972 70756 7028 71710
rect 6972 67842 7028 70700
rect 6972 67790 6974 67842
rect 7026 67790 7028 67842
rect 6972 67778 7028 67790
rect 7084 71538 7140 71550
rect 7084 71486 7086 71538
rect 7138 71486 7140 71538
rect 7084 67284 7140 71486
rect 7196 70306 7252 72828
rect 7308 70978 7364 73052
rect 7420 72324 7476 72334
rect 7420 72230 7476 72268
rect 7644 71762 7700 74622
rect 7756 73332 7812 76974
rect 7868 73332 7924 77756
rect 8092 76466 8148 78542
rect 8204 77588 8260 84028
rect 8428 84018 8484 84028
rect 8428 83860 8484 83870
rect 8316 82740 8372 82750
rect 8316 82516 8372 82684
rect 8316 82450 8372 82460
rect 8316 82292 8372 82302
rect 8316 82178 8372 82236
rect 8316 82126 8318 82178
rect 8370 82126 8372 82178
rect 8316 82114 8372 82126
rect 8428 81508 8484 83804
rect 8540 82180 8596 91868
rect 8540 82114 8596 82124
rect 8316 81452 8484 81508
rect 8316 80500 8372 81452
rect 8540 81170 8596 81182
rect 8540 81118 8542 81170
rect 8594 81118 8596 81170
rect 8540 81060 8596 81118
rect 8540 80994 8596 81004
rect 8316 80444 8484 80500
rect 8428 79714 8484 80444
rect 8652 79828 8708 97580
rect 8988 97522 9044 97534
rect 8988 97470 8990 97522
rect 9042 97470 9044 97522
rect 8988 97468 9044 97470
rect 8764 97412 9044 97468
rect 9100 97468 9156 98142
rect 9212 97636 9268 104636
rect 9660 104468 9716 105310
rect 9660 104374 9716 104412
rect 9996 105812 10164 105868
rect 9772 103796 9828 103806
rect 9324 103124 9380 103134
rect 9324 103030 9380 103068
rect 9660 102564 9716 102574
rect 9436 102114 9492 102126
rect 9436 102062 9438 102114
rect 9490 102062 9492 102114
rect 9436 100212 9492 102062
rect 9548 101554 9604 101566
rect 9548 101502 9550 101554
rect 9602 101502 9604 101554
rect 9548 100884 9604 101502
rect 9660 101442 9716 102508
rect 9660 101390 9662 101442
rect 9714 101390 9716 101442
rect 9660 101378 9716 101390
rect 9548 100818 9604 100828
rect 9436 100146 9492 100156
rect 9548 100658 9604 100670
rect 9548 100606 9550 100658
rect 9602 100606 9604 100658
rect 9548 100548 9604 100606
rect 9324 99988 9380 99998
rect 9324 99894 9380 99932
rect 9548 99876 9604 100492
rect 9548 99810 9604 99820
rect 9660 99652 9716 99662
rect 9660 99316 9716 99596
rect 9212 97570 9268 97580
rect 9548 98196 9604 98206
rect 9100 97412 9268 97468
rect 8764 94836 8820 97412
rect 8764 94770 8820 94780
rect 8876 95732 8932 95742
rect 8876 95282 8932 95676
rect 8876 95230 8878 95282
rect 8930 95230 8932 95282
rect 8876 94052 8932 95230
rect 8764 93492 8820 93502
rect 8876 93492 8932 93996
rect 8988 95284 9044 95294
rect 8988 93714 9044 95228
rect 9100 95058 9156 95070
rect 9100 95006 9102 95058
rect 9154 95006 9156 95058
rect 9100 94948 9156 95006
rect 9100 94882 9156 94892
rect 9212 94836 9268 97412
rect 9324 96628 9380 96638
rect 9324 96626 9492 96628
rect 9324 96574 9326 96626
rect 9378 96574 9492 96626
rect 9324 96572 9492 96574
rect 9324 96562 9380 96572
rect 9212 94780 9380 94836
rect 8988 93662 8990 93714
rect 9042 93662 9044 93714
rect 8988 93650 9044 93662
rect 9212 94610 9268 94622
rect 9212 94558 9214 94610
rect 9266 94558 9268 94610
rect 8876 93436 9044 93492
rect 8764 92932 8820 93436
rect 8876 93044 8932 93054
rect 8876 92950 8932 92988
rect 8764 91924 8820 92876
rect 8988 92146 9044 93436
rect 9212 93156 9268 94558
rect 9324 93940 9380 94780
rect 9324 93874 9380 93884
rect 9324 93714 9380 93726
rect 9324 93662 9326 93714
rect 9378 93662 9380 93714
rect 9324 93492 9380 93662
rect 9324 93426 9380 93436
rect 8988 92094 8990 92146
rect 9042 92094 9044 92146
rect 8988 92082 9044 92094
rect 9100 93100 9268 93156
rect 9100 92036 9156 93100
rect 9324 92932 9380 92942
rect 9436 92932 9492 96572
rect 9548 95284 9604 98140
rect 9548 95190 9604 95228
rect 9660 94836 9716 99260
rect 9772 98530 9828 103740
rect 9884 100772 9940 100782
rect 9884 100678 9940 100716
rect 9996 100436 10052 105812
rect 10108 103684 10164 103694
rect 10332 103684 10388 103694
rect 10108 103234 10164 103628
rect 10108 103182 10110 103234
rect 10162 103182 10164 103234
rect 10108 103170 10164 103182
rect 10220 103682 10388 103684
rect 10220 103630 10334 103682
rect 10386 103630 10388 103682
rect 10220 103628 10388 103630
rect 10108 102450 10164 102462
rect 10108 102398 10110 102450
rect 10162 102398 10164 102450
rect 10108 101668 10164 102398
rect 10220 102338 10276 103628
rect 10332 103618 10388 103628
rect 10220 102286 10222 102338
rect 10274 102286 10276 102338
rect 10220 102274 10276 102286
rect 10444 101892 10500 105980
rect 10668 106034 10724 106046
rect 10668 105982 10670 106034
rect 10722 105982 10724 106034
rect 10556 102900 10612 102910
rect 10556 102806 10612 102844
rect 10668 102564 10724 105982
rect 10668 102498 10724 102508
rect 10780 106036 10836 106046
rect 10780 103684 10836 105980
rect 11004 105700 11060 106204
rect 11116 106036 11172 106046
rect 11116 106034 11284 106036
rect 11116 105982 11118 106034
rect 11170 105982 11284 106034
rect 11116 105980 11284 105982
rect 11116 105970 11172 105980
rect 11116 105700 11172 105710
rect 11004 105698 11172 105700
rect 11004 105646 11118 105698
rect 11170 105646 11172 105698
rect 11004 105644 11172 105646
rect 11116 105634 11172 105644
rect 11228 105476 11284 105980
rect 11340 105476 11396 105486
rect 11228 105474 11396 105476
rect 11228 105422 11342 105474
rect 11394 105422 11396 105474
rect 11228 105420 11396 105422
rect 10444 101826 10500 101836
rect 10108 101612 10500 101668
rect 10108 101444 10164 101454
rect 10108 101350 10164 101388
rect 9884 100380 10052 100436
rect 10108 101108 10164 101118
rect 9884 99986 9940 100380
rect 9884 99934 9886 99986
rect 9938 99934 9940 99986
rect 9884 99764 9940 99934
rect 9996 100212 10052 100222
rect 9996 99874 10052 100156
rect 9996 99822 9998 99874
rect 10050 99822 10052 99874
rect 9996 99810 10052 99822
rect 9884 99698 9940 99708
rect 10108 99204 10164 101052
rect 10332 100884 10388 100894
rect 10332 100770 10388 100828
rect 10332 100718 10334 100770
rect 10386 100718 10388 100770
rect 10332 100706 10388 100718
rect 10332 100212 10388 100222
rect 9996 99148 10164 99204
rect 10220 99988 10276 99998
rect 10220 99208 10276 99932
rect 10220 99156 10222 99208
rect 10274 99156 10276 99208
rect 9772 98478 9774 98530
rect 9826 98478 9828 98530
rect 9772 98466 9828 98478
rect 9884 99090 9940 99102
rect 9884 99038 9886 99090
rect 9938 99038 9940 99090
rect 9884 95284 9940 99038
rect 9996 98868 10052 99148
rect 10220 99144 10276 99156
rect 9996 98812 10276 98868
rect 10108 98532 10164 98542
rect 10108 98306 10164 98476
rect 10108 98254 10110 98306
rect 10162 98254 10164 98306
rect 10108 98242 10164 98254
rect 10220 97746 10276 98812
rect 10220 97694 10222 97746
rect 10274 97694 10276 97746
rect 9996 97412 10052 97422
rect 9996 96964 10052 97356
rect 9996 96962 10164 96964
rect 9996 96910 9998 96962
rect 10050 96910 10164 96962
rect 9996 96908 10164 96910
rect 9996 96898 10052 96908
rect 9884 95218 9940 95228
rect 9996 95620 10052 95630
rect 9548 94780 9716 94836
rect 9548 93828 9604 94780
rect 9660 94612 9716 94622
rect 9660 94610 9828 94612
rect 9660 94558 9662 94610
rect 9714 94558 9828 94610
rect 9660 94556 9828 94558
rect 9660 94546 9716 94556
rect 9548 93772 9716 93828
rect 9548 93604 9604 93614
rect 9548 93510 9604 93548
rect 9660 93156 9716 93772
rect 9324 92930 9492 92932
rect 9324 92878 9326 92930
rect 9378 92878 9492 92930
rect 9324 92876 9492 92878
rect 9324 92866 9380 92876
rect 9324 92372 9380 92382
rect 9212 92036 9268 92046
rect 9100 92034 9268 92036
rect 9100 91982 9214 92034
rect 9266 91982 9268 92034
rect 9100 91980 9268 91982
rect 9212 91970 9268 91980
rect 8764 91858 8820 91868
rect 9212 90578 9268 90590
rect 9212 90526 9214 90578
rect 9266 90526 9268 90578
rect 8988 89012 9044 89022
rect 8988 88918 9044 88956
rect 8988 88788 9044 88798
rect 8876 85874 8932 85886
rect 8876 85822 8878 85874
rect 8930 85822 8932 85874
rect 8876 85764 8932 85822
rect 8876 85698 8932 85708
rect 8988 85762 9044 88732
rect 8988 85710 8990 85762
rect 9042 85710 9044 85762
rect 8988 85698 9044 85710
rect 9100 87442 9156 87454
rect 9100 87390 9102 87442
rect 9154 87390 9156 87442
rect 8988 85092 9044 85102
rect 8876 84308 8932 84318
rect 8876 84214 8932 84252
rect 8876 83636 8932 83646
rect 8876 83542 8932 83580
rect 8876 83412 8932 83422
rect 8764 82852 8820 82862
rect 8764 82626 8820 82796
rect 8764 82574 8766 82626
rect 8818 82574 8820 82626
rect 8764 82562 8820 82574
rect 8652 79762 8708 79772
rect 8876 81058 8932 83356
rect 8988 82178 9044 85036
rect 9100 84644 9156 87390
rect 9100 84578 9156 84588
rect 9212 83748 9268 90526
rect 9324 89908 9380 92316
rect 9436 92260 9492 92876
rect 9436 92194 9492 92204
rect 9548 93100 9716 93156
rect 9324 89842 9380 89852
rect 8988 82126 8990 82178
rect 9042 82126 9044 82178
rect 8988 82114 9044 82126
rect 9100 83692 9268 83748
rect 9324 89012 9380 89022
rect 9100 81396 9156 83692
rect 9212 83524 9268 83534
rect 9212 83430 9268 83468
rect 9100 81330 9156 81340
rect 9212 83300 9268 83310
rect 8876 81006 8878 81058
rect 8930 81006 8932 81058
rect 8428 79662 8430 79714
rect 8482 79662 8484 79714
rect 8428 79492 8484 79662
rect 8764 79604 8820 79614
rect 8764 79510 8820 79548
rect 8428 79426 8484 79436
rect 8876 79380 8932 81006
rect 8764 79324 8932 79380
rect 9100 79828 9156 79838
rect 9100 79380 9156 79772
rect 9212 79602 9268 83244
rect 9324 81956 9380 88956
rect 9436 87332 9492 87342
rect 9436 86658 9492 87276
rect 9436 86606 9438 86658
rect 9490 86606 9492 86658
rect 9436 86594 9492 86606
rect 9436 85988 9492 85998
rect 9436 85874 9492 85932
rect 9436 85822 9438 85874
rect 9490 85822 9492 85874
rect 9436 85810 9492 85822
rect 9548 82348 9604 93100
rect 9660 92932 9716 92942
rect 9660 92838 9716 92876
rect 9660 92260 9716 92270
rect 9660 92146 9716 92204
rect 9660 92094 9662 92146
rect 9714 92094 9716 92146
rect 9660 92082 9716 92094
rect 9772 90804 9828 94556
rect 9884 94274 9940 94286
rect 9884 94222 9886 94274
rect 9938 94222 9940 94274
rect 9884 93154 9940 94222
rect 9996 94164 10052 95564
rect 10108 95396 10164 96908
rect 10108 95330 10164 95340
rect 10220 94500 10276 97694
rect 10332 97300 10388 100156
rect 10444 99540 10500 101612
rect 10668 101554 10724 101566
rect 10668 101502 10670 101554
rect 10722 101502 10724 101554
rect 10556 100882 10612 100894
rect 10556 100830 10558 100882
rect 10610 100830 10612 100882
rect 10556 99764 10612 100830
rect 10668 100212 10724 101502
rect 10668 100146 10724 100156
rect 10668 99988 10724 99998
rect 10668 99894 10724 99932
rect 10556 99698 10612 99708
rect 10780 99652 10836 103628
rect 11004 104804 11060 104814
rect 10892 102228 10948 102238
rect 10892 102134 10948 102172
rect 11004 102116 11060 104748
rect 11116 104468 11172 104478
rect 11116 104374 11172 104412
rect 11340 104468 11396 105420
rect 11452 104804 11508 108780
rect 11676 108610 11732 109116
rect 11676 108558 11678 108610
rect 11730 108558 11732 108610
rect 11676 108546 11732 108558
rect 11900 108722 11956 108734
rect 11900 108670 11902 108722
rect 11954 108670 11956 108722
rect 11788 107380 11844 107390
rect 11564 106818 11620 106830
rect 11564 106766 11566 106818
rect 11618 106766 11620 106818
rect 11564 106484 11620 106766
rect 11564 106418 11620 106428
rect 11788 106596 11844 107324
rect 11452 104738 11508 104748
rect 11676 104914 11732 104926
rect 11676 104862 11678 104914
rect 11730 104862 11732 104914
rect 11564 104690 11620 104702
rect 11564 104638 11566 104690
rect 11618 104638 11620 104690
rect 11340 104402 11396 104412
rect 11452 104466 11508 104478
rect 11452 104414 11454 104466
rect 11506 104414 11508 104466
rect 11452 104244 11508 104414
rect 11004 101108 11060 102060
rect 11004 101042 11060 101052
rect 11116 104188 11508 104244
rect 11116 100884 11172 104188
rect 11452 104018 11508 104030
rect 11452 103966 11454 104018
rect 11506 103966 11508 104018
rect 11452 103908 11508 103966
rect 11116 100818 11172 100828
rect 11228 103684 11284 103694
rect 11228 100770 11284 103628
rect 11452 103124 11508 103852
rect 11564 103236 11620 104638
rect 11676 104468 11732 104862
rect 11676 104402 11732 104412
rect 11788 104244 11844 106540
rect 11676 104188 11844 104244
rect 11676 103908 11732 104188
rect 11900 104132 11956 108670
rect 12012 107826 12068 107838
rect 12012 107774 12014 107826
rect 12066 107774 12068 107826
rect 12012 107604 12068 107774
rect 12012 107538 12068 107548
rect 12124 105250 12180 105262
rect 12124 105198 12126 105250
rect 12178 105198 12180 105250
rect 11900 104066 11956 104076
rect 12012 104580 12068 104590
rect 12124 104580 12180 105198
rect 12012 104578 12180 104580
rect 12012 104526 12014 104578
rect 12066 104526 12180 104578
rect 12012 104524 12180 104526
rect 12236 104578 12292 104590
rect 12236 104526 12238 104578
rect 12290 104526 12292 104578
rect 11676 103842 11732 103852
rect 12012 103908 12068 104524
rect 12236 104132 12292 104526
rect 12348 104580 12404 110908
rect 12460 110516 12516 111806
rect 12908 111076 12964 112254
rect 13468 112084 13524 114800
rect 13692 113652 13748 114800
rect 13692 113596 13860 113652
rect 13692 113428 13748 113438
rect 13692 113334 13748 113372
rect 13468 112018 13524 112028
rect 12908 111010 12964 111020
rect 13132 111860 13188 111870
rect 12460 110450 12516 110460
rect 13020 110740 13076 110750
rect 12908 110068 12964 110078
rect 12908 109974 12964 110012
rect 12460 109954 12516 109966
rect 12460 109902 12462 109954
rect 12514 109902 12516 109954
rect 12460 108610 12516 109902
rect 12460 108558 12462 108610
rect 12514 108558 12516 108610
rect 12460 108546 12516 108558
rect 12908 109732 12964 109742
rect 12908 109060 12964 109676
rect 13020 109508 13076 110684
rect 13020 109442 13076 109452
rect 12908 108610 12964 109004
rect 12908 108558 12910 108610
rect 12962 108558 12964 108610
rect 12908 108546 12964 108558
rect 12796 107604 12852 107614
rect 12684 107268 12740 107278
rect 12684 107174 12740 107212
rect 12348 104514 12404 104524
rect 12796 104802 12852 107548
rect 13132 107380 13188 111804
rect 13692 111860 13748 111870
rect 13692 111636 13748 111804
rect 13692 111570 13748 111580
rect 13580 111524 13636 111534
rect 13468 111522 13636 111524
rect 13468 111470 13582 111522
rect 13634 111470 13636 111522
rect 13468 111468 13636 111470
rect 13244 111412 13300 111422
rect 13244 110180 13300 111356
rect 13244 110114 13300 110124
rect 13356 110180 13412 110190
rect 13468 110180 13524 111468
rect 13580 111458 13636 111468
rect 13580 110964 13636 111002
rect 13580 110898 13636 110908
rect 13692 110852 13748 110862
rect 13356 110178 13524 110180
rect 13356 110126 13358 110178
rect 13410 110126 13524 110178
rect 13356 110124 13524 110126
rect 13580 110740 13636 110750
rect 13356 110114 13412 110124
rect 13244 109620 13300 109630
rect 13244 109060 13300 109564
rect 13468 109508 13524 109518
rect 13468 109414 13524 109452
rect 13244 108994 13300 109004
rect 13580 108724 13636 110684
rect 13692 110178 13748 110796
rect 13692 110126 13694 110178
rect 13746 110126 13748 110178
rect 13692 110114 13748 110126
rect 13468 108668 13636 108724
rect 13468 108052 13524 108668
rect 13356 107996 13524 108052
rect 13580 108276 13636 108286
rect 13356 107492 13412 107996
rect 13468 107828 13524 107838
rect 13468 107734 13524 107772
rect 13356 107426 13412 107436
rect 13132 107314 13188 107324
rect 13132 106930 13188 106942
rect 13132 106878 13134 106930
rect 13186 106878 13188 106930
rect 12796 104750 12798 104802
rect 12850 104750 12852 104802
rect 12348 104132 12404 104142
rect 12236 104130 12404 104132
rect 12236 104078 12350 104130
rect 12402 104078 12404 104130
rect 12236 104076 12404 104078
rect 12348 104066 12404 104076
rect 12012 103842 12068 103852
rect 12572 104018 12628 104030
rect 12572 103966 12574 104018
rect 12626 103966 12628 104018
rect 11900 103796 11956 103806
rect 11900 103702 11956 103740
rect 11676 103684 11732 103694
rect 11676 103346 11732 103628
rect 11676 103294 11678 103346
rect 11730 103294 11732 103346
rect 11676 103282 11732 103294
rect 12124 103684 12180 103694
rect 11564 103170 11620 103180
rect 12124 103234 12180 103628
rect 12236 103348 12292 103358
rect 12572 103348 12628 103966
rect 12684 104020 12740 104030
rect 12796 104020 12852 104750
rect 12684 104018 12852 104020
rect 12684 103966 12686 104018
rect 12738 103966 12852 104018
rect 12684 103964 12852 103966
rect 12684 103954 12740 103964
rect 12796 103572 12852 103964
rect 12908 106820 12964 106830
rect 12908 103796 12964 106764
rect 13020 106484 13076 106494
rect 13020 106260 13076 106428
rect 13020 106166 13076 106204
rect 13132 106260 13188 106878
rect 13356 106596 13412 106606
rect 13244 106260 13300 106270
rect 13132 106204 13244 106260
rect 13132 106036 13188 106204
rect 13244 106194 13300 106204
rect 13132 105970 13188 105980
rect 13356 106146 13412 106540
rect 13356 106094 13358 106146
rect 13410 106094 13412 106146
rect 13356 106036 13412 106094
rect 13468 106036 13524 106046
rect 13356 105980 13468 106036
rect 13132 105812 13188 105822
rect 13132 104690 13188 105756
rect 13356 105586 13412 105980
rect 13468 105970 13524 105980
rect 13356 105534 13358 105586
rect 13410 105534 13412 105586
rect 13356 105522 13412 105534
rect 13468 105588 13524 105598
rect 13132 104638 13134 104690
rect 13186 104638 13188 104690
rect 13132 104626 13188 104638
rect 13468 104692 13524 105532
rect 13468 104626 13524 104636
rect 13580 104690 13636 108220
rect 13692 107716 13748 107726
rect 13692 107622 13748 107660
rect 13804 107604 13860 113596
rect 13916 110740 13972 114800
rect 14140 113428 14196 114800
rect 14140 113362 14196 113372
rect 14140 113202 14196 113214
rect 14140 113150 14142 113202
rect 14194 113150 14196 113202
rect 14140 112756 14196 113150
rect 14140 112690 14196 112700
rect 14364 112644 14420 114800
rect 14588 113428 14644 114800
rect 14700 113540 14756 113550
rect 14700 113446 14756 113484
rect 14588 113362 14644 113372
rect 14588 113204 14644 113214
rect 14364 112578 14420 112588
rect 14476 112756 14532 112766
rect 14476 112530 14532 112700
rect 14476 112478 14478 112530
rect 14530 112478 14532 112530
rect 14028 112306 14084 112318
rect 14028 112254 14030 112306
rect 14082 112254 14084 112306
rect 14028 111300 14084 112254
rect 14364 111748 14420 111758
rect 14028 111234 14084 111244
rect 14252 111746 14420 111748
rect 14252 111694 14366 111746
rect 14418 111694 14420 111746
rect 14252 111692 14420 111694
rect 14252 110964 14308 111692
rect 14364 111682 14420 111692
rect 14476 111636 14532 112478
rect 14476 111570 14532 111580
rect 14588 111188 14644 113148
rect 14812 112644 14868 114800
rect 15036 113540 15092 114800
rect 15036 113474 15092 113484
rect 14812 112578 14868 112588
rect 15036 113314 15092 113326
rect 15036 113262 15038 113314
rect 15090 113262 15092 113314
rect 14924 111860 14980 111898
rect 14924 111794 14980 111804
rect 14252 110898 14308 110908
rect 14364 111132 14644 111188
rect 14924 111636 14980 111646
rect 13916 110674 13972 110684
rect 14028 110738 14084 110750
rect 14028 110686 14030 110738
rect 14082 110686 14084 110738
rect 13916 110516 13972 110526
rect 13916 110402 13972 110460
rect 13916 110350 13918 110402
rect 13970 110350 13972 110402
rect 13916 110338 13972 110350
rect 14028 110068 14084 110686
rect 14028 110002 14084 110012
rect 14252 109956 14308 109966
rect 13916 109396 13972 109406
rect 13916 109282 13972 109340
rect 13916 109230 13918 109282
rect 13970 109230 13972 109282
rect 13916 109218 13972 109230
rect 13916 108612 13972 108622
rect 13916 108518 13972 108556
rect 14028 108164 14084 108174
rect 13804 107538 13860 107548
rect 13916 107940 13972 107950
rect 13916 107380 13972 107884
rect 14028 107714 14084 108108
rect 14028 107662 14030 107714
rect 14082 107662 14084 107714
rect 14028 107650 14084 107662
rect 14140 107828 14196 107838
rect 13692 107324 13972 107380
rect 14028 107492 14084 107502
rect 13692 105700 13748 107324
rect 14028 107266 14084 107436
rect 14028 107214 14030 107266
rect 14082 107214 14084 107266
rect 14028 107202 14084 107214
rect 13804 107044 13860 107054
rect 13804 107042 13972 107044
rect 13804 106990 13806 107042
rect 13858 106990 13972 107042
rect 13804 106988 13972 106990
rect 13804 106978 13860 106988
rect 13804 105700 13860 105710
rect 13692 105644 13804 105700
rect 13580 104638 13582 104690
rect 13634 104638 13636 104690
rect 12908 103730 12964 103740
rect 13132 103684 13188 103694
rect 13132 103590 13188 103628
rect 12796 103516 13076 103572
rect 12796 103348 12852 103358
rect 12236 103346 12852 103348
rect 12236 103294 12238 103346
rect 12290 103294 12798 103346
rect 12850 103294 12852 103346
rect 12236 103292 12852 103294
rect 12236 103282 12292 103292
rect 12796 103282 12852 103292
rect 12124 103182 12126 103234
rect 12178 103182 12180 103234
rect 12124 103170 12180 103182
rect 12908 103236 12964 103246
rect 12908 103142 12964 103180
rect 11452 103058 11508 103068
rect 11676 103124 11732 103134
rect 11732 103068 11788 103124
rect 11676 103058 11788 103068
rect 11732 103012 11788 103058
rect 11732 102956 12068 103012
rect 11228 100718 11230 100770
rect 11282 100718 11284 100770
rect 11228 100706 11284 100718
rect 11340 102450 11396 102462
rect 11340 102398 11342 102450
rect 11394 102398 11396 102450
rect 11340 101108 11396 102398
rect 11228 99986 11284 99998
rect 11228 99934 11230 99986
rect 11282 99934 11284 99986
rect 11228 99876 11284 99934
rect 11228 99810 11284 99820
rect 11340 99764 11396 101052
rect 11676 101554 11732 101566
rect 11676 101502 11678 101554
rect 11730 101502 11732 101554
rect 11564 100770 11620 100782
rect 11564 100718 11566 100770
rect 11618 100718 11620 100770
rect 11340 99698 11396 99708
rect 11452 99988 11508 99998
rect 10780 99596 11060 99652
rect 10444 99484 10836 99540
rect 10780 99428 10836 99484
rect 10780 99372 10948 99428
rect 10892 99314 10948 99372
rect 10892 99262 10894 99314
rect 10946 99262 10948 99314
rect 10892 99250 10948 99262
rect 10780 99202 10836 99214
rect 10780 99150 10782 99202
rect 10834 99150 10836 99202
rect 10780 98308 10836 99150
rect 11004 98644 11060 99596
rect 11452 99202 11508 99932
rect 11564 99428 11620 100718
rect 11564 99362 11620 99372
rect 11452 99150 11454 99202
rect 11506 99150 11508 99202
rect 11004 98578 11060 98588
rect 11228 98644 11284 98654
rect 11228 98420 11284 98588
rect 11340 98644 11396 98654
rect 11452 98644 11508 99150
rect 11340 98642 11508 98644
rect 11340 98590 11342 98642
rect 11394 98590 11508 98642
rect 11340 98588 11508 98590
rect 11676 99204 11732 101502
rect 11340 98578 11396 98588
rect 11228 98364 11396 98420
rect 10780 98252 11284 98308
rect 10332 96068 10388 97244
rect 10556 97748 10612 97758
rect 10556 97634 10612 97692
rect 10556 97582 10558 97634
rect 10610 97582 10612 97634
rect 10444 96628 10500 96638
rect 10444 96534 10500 96572
rect 10332 96002 10388 96012
rect 10444 95954 10500 95966
rect 10444 95902 10446 95954
rect 10498 95902 10500 95954
rect 10444 95732 10500 95902
rect 10444 95666 10500 95676
rect 10332 95282 10388 95294
rect 10332 95230 10334 95282
rect 10386 95230 10388 95282
rect 10332 95060 10388 95230
rect 10556 95172 10612 97582
rect 10892 96852 10948 96862
rect 10892 96066 10948 96796
rect 10892 96014 10894 96066
rect 10946 96014 10948 96066
rect 10892 96002 10948 96014
rect 11228 96066 11284 98252
rect 11340 97634 11396 98364
rect 11340 97582 11342 97634
rect 11394 97582 11396 97634
rect 11340 97412 11396 97582
rect 11340 97346 11396 97356
rect 11564 96852 11620 96862
rect 11452 96292 11508 96302
rect 11452 96198 11508 96236
rect 11228 96014 11230 96066
rect 11282 96014 11284 96066
rect 10780 95396 10836 95406
rect 10556 95116 10724 95172
rect 10332 95004 10612 95060
rect 9996 94098 10052 94108
rect 10108 94444 10276 94500
rect 10332 94836 10388 94846
rect 9884 93102 9886 93154
rect 9938 93102 9940 93154
rect 9884 93090 9940 93102
rect 9996 90804 10052 90814
rect 9772 90802 10052 90804
rect 9772 90750 9998 90802
rect 10050 90750 10052 90802
rect 9772 90748 10052 90750
rect 9996 90738 10052 90748
rect 10108 90580 10164 94444
rect 10220 94276 10276 94286
rect 10220 94182 10276 94220
rect 10220 93716 10276 93726
rect 10332 93716 10388 94780
rect 10220 93714 10388 93716
rect 10220 93662 10222 93714
rect 10274 93662 10388 93714
rect 10220 93660 10388 93662
rect 10444 93940 10500 93950
rect 10220 93650 10276 93660
rect 10332 93044 10388 93054
rect 9996 90524 10164 90580
rect 10220 92146 10276 92158
rect 10220 92094 10222 92146
rect 10274 92094 10276 92146
rect 9660 90244 9716 90254
rect 9660 89682 9716 90188
rect 9660 89630 9662 89682
rect 9714 89630 9716 89682
rect 9660 89124 9716 89630
rect 9660 89030 9716 89068
rect 9996 88898 10052 90524
rect 10220 90468 10276 92094
rect 10220 90402 10276 90412
rect 10108 89908 10164 89918
rect 10108 89814 10164 89852
rect 9996 88846 9998 88898
rect 10050 88846 10052 88898
rect 9996 88788 10052 88846
rect 9772 88732 10052 88788
rect 9660 84308 9716 84318
rect 9660 84214 9716 84252
rect 9660 84084 9716 84094
rect 9660 83522 9716 84028
rect 9660 83470 9662 83522
rect 9714 83470 9716 83522
rect 9660 83458 9716 83470
rect 9772 83412 9828 88732
rect 9884 88340 9940 88350
rect 9884 86882 9940 88284
rect 9884 86830 9886 86882
rect 9938 86830 9940 86882
rect 9884 84196 9940 86830
rect 10108 87442 10164 87454
rect 10108 87390 10110 87442
rect 10162 87390 10164 87442
rect 9884 84130 9940 84140
rect 9996 86772 10052 86782
rect 9884 83748 9940 83758
rect 9884 83654 9940 83692
rect 9772 83346 9828 83356
rect 9884 83524 9940 83534
rect 9884 82962 9940 83468
rect 9884 82910 9886 82962
rect 9938 82910 9940 82962
rect 9884 82898 9940 82910
rect 9548 82292 9940 82348
rect 9324 81508 9380 81900
rect 9324 81442 9380 81452
rect 9660 81060 9716 81070
rect 9660 80500 9716 81004
rect 9212 79550 9214 79602
rect 9266 79550 9268 79602
rect 9212 79538 9268 79550
rect 9436 80444 9716 80500
rect 9884 80498 9940 82292
rect 9884 80446 9886 80498
rect 9938 80446 9940 80498
rect 9436 79604 9492 80444
rect 9548 80276 9604 80286
rect 9548 80274 9716 80276
rect 9548 80222 9550 80274
rect 9602 80222 9716 80274
rect 9548 80220 9716 80222
rect 9548 80210 9604 80220
rect 9436 79548 9604 79604
rect 9436 79380 9492 79390
rect 9100 79324 9268 79380
rect 8428 79156 8484 79166
rect 8316 78932 8372 78942
rect 8316 78148 8372 78876
rect 8316 77922 8372 78092
rect 8316 77870 8318 77922
rect 8370 77870 8372 77922
rect 8316 77858 8372 77870
rect 8428 77588 8484 79100
rect 8540 79044 8596 79054
rect 8540 77812 8596 78988
rect 8540 77746 8596 77756
rect 8204 77532 8372 77588
rect 8092 76414 8094 76466
rect 8146 76414 8148 76466
rect 8092 76402 8148 76414
rect 8092 76244 8148 76254
rect 8092 74786 8148 76188
rect 8204 75684 8260 75694
rect 8204 75590 8260 75628
rect 8092 74734 8094 74786
rect 8146 74734 8148 74786
rect 8092 74722 8148 74734
rect 8204 75236 8260 75246
rect 8204 74338 8260 75180
rect 8316 74898 8372 77532
rect 8316 74846 8318 74898
rect 8370 74846 8372 74898
rect 8316 74834 8372 74846
rect 8204 74286 8206 74338
rect 8258 74286 8260 74338
rect 7980 74116 8036 74126
rect 7980 74022 8036 74060
rect 8204 73444 8260 74286
rect 8204 73378 8260 73388
rect 8316 74114 8372 74126
rect 8316 74062 8318 74114
rect 8370 74062 8372 74114
rect 8092 73332 8148 73342
rect 7868 73330 8148 73332
rect 7868 73278 8094 73330
rect 8146 73278 8148 73330
rect 7868 73276 8148 73278
rect 7756 73266 7812 73276
rect 7868 72658 7924 72670
rect 7868 72606 7870 72658
rect 7922 72606 7924 72658
rect 7644 71710 7646 71762
rect 7698 71710 7700 71762
rect 7644 71698 7700 71710
rect 7756 72548 7812 72558
rect 7756 71540 7812 72492
rect 7756 71474 7812 71484
rect 7308 70926 7310 70978
rect 7362 70926 7364 70978
rect 7308 70914 7364 70926
rect 7756 71092 7812 71102
rect 7196 70254 7198 70306
rect 7250 70254 7252 70306
rect 7196 70242 7252 70254
rect 7308 70194 7364 70206
rect 7308 70142 7310 70194
rect 7362 70142 7364 70194
rect 7308 69748 7364 70142
rect 7756 70082 7812 71036
rect 7756 70030 7758 70082
rect 7810 70030 7812 70082
rect 7756 70018 7812 70030
rect 7868 69972 7924 72606
rect 8092 72324 8148 73276
rect 8316 73220 8372 74062
rect 8316 73154 8372 73164
rect 8092 72258 8148 72268
rect 8204 72546 8260 72558
rect 8204 72494 8206 72546
rect 8258 72494 8260 72546
rect 8092 71764 8148 71774
rect 7868 69906 7924 69916
rect 7980 71762 8148 71764
rect 7980 71710 8094 71762
rect 8146 71710 8148 71762
rect 7980 71708 8148 71710
rect 7980 69748 8036 71708
rect 8092 71698 8148 71708
rect 8092 71540 8148 71550
rect 8092 70978 8148 71484
rect 8092 70926 8094 70978
rect 8146 70926 8148 70978
rect 8092 70914 8148 70926
rect 8092 70084 8148 70094
rect 8092 69990 8148 70028
rect 7308 69692 7924 69748
rect 7980 69692 8148 69748
rect 7308 69188 7364 69198
rect 7308 69094 7364 69132
rect 7308 68852 7364 68862
rect 7308 68626 7364 68796
rect 7308 68574 7310 68626
rect 7362 68574 7364 68626
rect 7308 68562 7364 68574
rect 7756 68516 7812 68526
rect 7756 68422 7812 68460
rect 7196 67842 7252 67854
rect 7196 67790 7198 67842
rect 7250 67790 7252 67842
rect 7196 67732 7252 67790
rect 7196 67676 7812 67732
rect 7084 67218 7140 67228
rect 7644 67396 7700 67406
rect 6972 67172 7028 67182
rect 6972 66836 7028 67116
rect 6972 66770 7028 66780
rect 7308 67060 7364 67070
rect 7308 66946 7364 67004
rect 7308 66894 7310 66946
rect 7362 66894 7364 66946
rect 7308 66724 7364 66894
rect 7308 66658 7364 66668
rect 7308 66274 7364 66286
rect 7308 66222 7310 66274
rect 7362 66222 7364 66274
rect 7308 65828 7364 66222
rect 7308 65772 7588 65828
rect 7420 65268 7476 65278
rect 7308 65266 7476 65268
rect 7308 65214 7422 65266
rect 7474 65214 7476 65266
rect 7308 65212 7476 65214
rect 6972 64818 7028 64830
rect 6972 64766 6974 64818
rect 7026 64766 7028 64818
rect 6972 61572 7028 64766
rect 7084 63700 7140 63710
rect 7084 63698 7252 63700
rect 7084 63646 7086 63698
rect 7138 63646 7252 63698
rect 7084 63644 7252 63646
rect 7084 63634 7140 63644
rect 6972 61506 7028 61516
rect 7196 58548 7252 63644
rect 7308 62354 7364 65212
rect 7420 65202 7476 65212
rect 7532 64596 7588 65772
rect 7420 62916 7476 62926
rect 7420 62822 7476 62860
rect 7308 62302 7310 62354
rect 7362 62302 7364 62354
rect 7308 62290 7364 62302
rect 7532 62188 7588 64540
rect 7644 63812 7700 67340
rect 7644 63746 7700 63756
rect 7644 62354 7700 62366
rect 7644 62302 7646 62354
rect 7698 62302 7700 62354
rect 7644 62188 7700 62302
rect 7420 62132 7700 62188
rect 7308 61572 7364 61582
rect 7420 61572 7476 62132
rect 7308 61570 7476 61572
rect 7308 61518 7310 61570
rect 7362 61518 7476 61570
rect 7308 61516 7476 61518
rect 7308 61506 7364 61516
rect 7308 60786 7364 60798
rect 7308 60734 7310 60786
rect 7362 60734 7364 60786
rect 7308 60228 7364 60734
rect 7420 60788 7476 61516
rect 7644 60788 7700 60798
rect 7420 60786 7700 60788
rect 7420 60734 7646 60786
rect 7698 60734 7700 60786
rect 7420 60732 7700 60734
rect 7644 60722 7700 60732
rect 7420 60228 7476 60238
rect 7308 60226 7476 60228
rect 7308 60174 7422 60226
rect 7474 60174 7476 60226
rect 7308 60172 7476 60174
rect 7420 60162 7476 60172
rect 7196 58482 7252 58492
rect 7756 57876 7812 67676
rect 7756 57810 7812 57820
rect 7084 56980 7140 56990
rect 7084 56978 7252 56980
rect 7084 56926 7086 56978
rect 7138 56926 7252 56978
rect 7084 56924 7252 56926
rect 7084 56914 7140 56924
rect 6916 56252 7140 56308
rect 6860 56242 6916 56252
rect 6636 56130 6692 56140
rect 6524 55300 6580 55310
rect 6524 55206 6580 55244
rect 6636 54852 6692 54862
rect 6524 54516 6580 54526
rect 6412 54514 6580 54516
rect 6412 54462 6526 54514
rect 6578 54462 6580 54514
rect 6412 54460 6580 54462
rect 6524 54450 6580 54460
rect 6300 53956 6356 54348
rect 6300 53890 6356 53900
rect 6636 53844 6692 54796
rect 6748 54292 6804 54302
rect 6748 54290 6916 54292
rect 6748 54238 6750 54290
rect 6802 54238 6916 54290
rect 6748 54236 6916 54238
rect 6748 54226 6804 54236
rect 6524 53788 6636 53844
rect 6300 53172 6356 53182
rect 6300 50428 6356 53116
rect 6412 52724 6468 52734
rect 6412 51378 6468 52668
rect 6412 51326 6414 51378
rect 6466 51326 6468 51378
rect 6412 51314 6468 51326
rect 6300 50372 6468 50428
rect 6188 48850 6244 48860
rect 5964 48178 6020 48188
rect 6412 48020 6468 50372
rect 6412 47954 6468 47964
rect 6524 47796 6580 53788
rect 6636 53778 6692 53788
rect 6748 53732 6804 53742
rect 6748 53638 6804 53676
rect 6636 52612 6692 52622
rect 6636 52164 6692 52556
rect 6860 52388 6916 54236
rect 6972 53732 7028 53742
rect 6972 52948 7028 53676
rect 6972 52854 7028 52892
rect 6636 52098 6692 52108
rect 6748 52332 6916 52388
rect 6636 49588 6692 49598
rect 6636 49026 6692 49532
rect 6636 48974 6638 49026
rect 6690 48974 6692 49026
rect 6636 48962 6692 48974
rect 6748 49028 6804 52332
rect 6860 52164 6916 52174
rect 6860 52070 6916 52108
rect 7084 51598 7140 56252
rect 6972 51542 7140 51598
rect 6748 48962 6804 48972
rect 6860 51268 6916 51278
rect 6860 50932 6916 51212
rect 6300 47740 6580 47796
rect 6636 48244 6692 48254
rect 6076 47348 6132 47358
rect 6076 47254 6132 47292
rect 5852 46676 5908 46686
rect 5852 46582 5908 46620
rect 6188 46450 6244 46462
rect 6188 46398 6190 46450
rect 6242 46398 6244 46450
rect 5964 45666 6020 45678
rect 5964 45614 5966 45666
rect 6018 45614 6020 45666
rect 5852 45444 5908 45454
rect 5628 45052 5796 45108
rect 5516 44902 5572 44940
rect 5628 44884 5684 44894
rect 5628 44790 5684 44828
rect 5292 43598 5294 43650
rect 5346 43598 5348 43650
rect 5292 43586 5348 43598
rect 5740 43540 5796 45052
rect 5852 45106 5908 45388
rect 5964 45220 6020 45614
rect 6188 45556 6244 46398
rect 6188 45490 6244 45500
rect 5964 45154 6020 45164
rect 5852 45054 5854 45106
rect 5906 45054 5908 45106
rect 5852 45042 5908 45054
rect 6076 44996 6132 45006
rect 6076 44902 6132 44940
rect 5628 43484 5796 43540
rect 5292 41970 5348 41982
rect 5292 41918 5294 41970
rect 5346 41918 5348 41970
rect 5292 41412 5348 41918
rect 5628 41748 5684 43484
rect 5740 43316 5796 43326
rect 5740 43314 5908 43316
rect 5740 43262 5742 43314
rect 5794 43262 5908 43314
rect 5740 43260 5908 43262
rect 5740 43250 5796 43260
rect 5740 43092 5796 43102
rect 5740 42754 5796 43036
rect 5852 42980 5908 43260
rect 5852 42914 5908 42924
rect 6188 42980 6244 42990
rect 6300 42980 6356 47740
rect 6524 47572 6580 47582
rect 6524 47478 6580 47516
rect 6636 47348 6692 48188
rect 6636 47282 6692 47292
rect 6748 47012 6804 47022
rect 6748 46562 6804 46956
rect 6748 46510 6750 46562
rect 6802 46510 6804 46562
rect 6748 46116 6804 46510
rect 6188 42978 6356 42980
rect 6188 42926 6190 42978
rect 6242 42926 6356 42978
rect 6188 42924 6356 42926
rect 6188 42914 6244 42924
rect 5740 42702 5742 42754
rect 5794 42702 5796 42754
rect 5740 42690 5796 42702
rect 6076 42196 6132 42206
rect 5852 42084 5908 42094
rect 5740 41972 5796 41982
rect 5740 41878 5796 41916
rect 5628 41692 5796 41748
rect 5292 41186 5348 41356
rect 5292 41134 5294 41186
rect 5346 41134 5348 41186
rect 5292 41122 5348 41134
rect 5628 41188 5684 41198
rect 5628 41094 5684 41132
rect 5180 40908 5348 40964
rect 5180 40404 5236 40414
rect 5180 40310 5236 40348
rect 5068 40238 5070 40290
rect 5122 40238 5124 40290
rect 5068 40226 5124 40238
rect 4956 39526 5012 39564
rect 4844 38770 4900 38780
rect 4284 38658 4340 38668
rect 4464 38444 4728 38454
rect 4520 38388 4568 38444
rect 4624 38388 4672 38444
rect 4464 38378 4728 38388
rect 5180 38276 5236 38286
rect 3804 37660 4068 37670
rect 3860 37604 3908 37660
rect 3964 37604 4012 37660
rect 3804 37594 4068 37604
rect 5180 37268 5236 38220
rect 5292 37828 5348 40908
rect 5404 39730 5460 39742
rect 5404 39678 5406 39730
rect 5458 39678 5460 39730
rect 5404 39284 5460 39678
rect 5404 39218 5460 39228
rect 5516 38834 5572 38846
rect 5516 38782 5518 38834
rect 5570 38782 5572 38834
rect 5516 38612 5572 38782
rect 5740 38668 5796 41692
rect 5852 41410 5908 42028
rect 5964 41748 6020 41758
rect 5964 41654 6020 41692
rect 5852 41358 5854 41410
rect 5906 41358 5908 41410
rect 5852 41346 5908 41358
rect 6076 41188 6132 42140
rect 5852 41132 6132 41188
rect 5852 40626 5908 41132
rect 5852 40574 5854 40626
rect 5906 40574 5908 40626
rect 5852 40562 5908 40574
rect 6188 40178 6244 40190
rect 6188 40126 6190 40178
rect 6242 40126 6244 40178
rect 6188 39844 6244 40126
rect 6188 39778 6244 39788
rect 6076 39508 6132 39518
rect 6132 39452 6244 39508
rect 6076 39442 6132 39452
rect 6188 38836 6244 39452
rect 5516 38546 5572 38556
rect 5628 38612 5796 38668
rect 6076 38724 6132 38762
rect 6076 38658 6132 38668
rect 5628 38388 5684 38612
rect 5292 37762 5348 37772
rect 5404 38332 5684 38388
rect 5740 38500 5796 38510
rect 4284 37042 4340 37054
rect 4284 36990 4286 37042
rect 4338 36990 4340 37042
rect 4284 36708 4340 36990
rect 4464 36876 4728 36886
rect 4520 36820 4568 36876
rect 4624 36820 4672 36876
rect 4464 36810 4728 36820
rect 4284 36642 4340 36652
rect 3724 36484 3780 36494
rect 3724 36482 4340 36484
rect 3724 36430 3726 36482
rect 3778 36430 4340 36482
rect 3724 36428 4340 36430
rect 3724 36418 3780 36428
rect 3804 36092 4068 36102
rect 3860 36036 3908 36092
rect 3964 36036 4012 36092
rect 3804 36026 4068 36036
rect 3612 35868 4004 35924
rect 3276 35698 3444 35700
rect 3276 35646 3278 35698
rect 3330 35646 3444 35698
rect 3276 35644 3444 35646
rect 3500 35812 3556 35822
rect 3276 35634 3332 35644
rect 3500 35308 3556 35756
rect 3052 31714 3108 31724
rect 3164 35252 3220 35262
rect 2828 26462 2830 26514
rect 2882 26462 2884 26514
rect 2828 26450 2884 26462
rect 2940 31668 2996 31678
rect 2940 25506 2996 31612
rect 3164 31218 3220 35196
rect 3388 35252 3556 35308
rect 3948 35252 4004 35868
rect 3388 35028 3444 35252
rect 3948 35186 4004 35196
rect 4172 35698 4228 35710
rect 4172 35646 4174 35698
rect 4226 35646 4228 35698
rect 3724 35140 3780 35150
rect 3724 35138 3892 35140
rect 3724 35086 3726 35138
rect 3778 35086 3892 35138
rect 3724 35084 3892 35086
rect 3724 35074 3780 35084
rect 3836 35028 3892 35084
rect 3948 35028 4004 35038
rect 3836 34972 3948 35028
rect 3388 34962 3444 34972
rect 3948 34962 4004 34972
rect 3164 31166 3166 31218
rect 3218 31166 3220 31218
rect 3164 31154 3220 31166
rect 3276 34914 3332 34926
rect 3276 34862 3278 34914
rect 3330 34862 3332 34914
rect 2940 25454 2942 25506
rect 2994 25454 2996 25506
rect 2940 25442 2996 25454
rect 3052 30210 3108 30222
rect 3052 30158 3054 30210
rect 3106 30158 3108 30210
rect 2716 25116 2996 25172
rect 2828 24948 2884 24958
rect 2604 24946 2884 24948
rect 2604 24894 2830 24946
rect 2882 24894 2884 24946
rect 2604 24892 2884 24894
rect 2828 24882 2884 24892
rect 2380 24210 2436 24220
rect 2716 24276 2772 24286
rect 2940 24276 2996 25116
rect 1596 22978 1652 22988
rect 1820 23996 1988 24052
rect 2268 24164 2324 24174
rect 1708 22930 1764 22942
rect 1708 22878 1710 22930
rect 1762 22878 1764 22930
rect 1708 21252 1764 22878
rect 1596 21196 1764 21252
rect 1820 21474 1876 23996
rect 1820 21422 1822 21474
rect 1874 21422 1876 21474
rect 1596 20916 1652 21196
rect 1596 20850 1652 20860
rect 1708 21028 1764 21038
rect 1708 20802 1764 20972
rect 1708 20750 1710 20802
rect 1762 20750 1764 20802
rect 1708 20738 1764 20750
rect 1708 20468 1764 20478
rect 924 17668 980 20188
rect 1148 20132 1204 20142
rect 1148 20038 1204 20076
rect 1260 20132 1540 20188
rect 1596 20356 1652 20366
rect 1260 19684 1316 20132
rect 1484 20020 1540 20030
rect 1148 19628 1316 19684
rect 1372 20018 1540 20020
rect 1372 19966 1486 20018
rect 1538 19966 1540 20018
rect 1372 19964 1540 19966
rect 1148 17890 1204 19628
rect 1260 19348 1316 19358
rect 1260 19254 1316 19292
rect 1148 17838 1150 17890
rect 1202 17838 1204 17890
rect 1148 17826 1204 17838
rect 924 17612 1204 17668
rect 1148 17106 1204 17612
rect 1148 17054 1150 17106
rect 1202 17054 1204 17106
rect 1148 17042 1204 17054
rect 1372 16436 1428 19964
rect 1484 19954 1540 19964
rect 1596 19572 1652 20300
rect 1484 19516 1652 19572
rect 1484 16772 1540 19516
rect 1596 19346 1652 19358
rect 1596 19294 1598 19346
rect 1650 19294 1652 19346
rect 1596 18452 1652 19294
rect 1708 18788 1764 20412
rect 1820 18900 1876 21422
rect 1932 23828 1988 23838
rect 1932 20132 1988 23772
rect 2044 22930 2100 22942
rect 2044 22878 2046 22930
rect 2098 22878 2100 22930
rect 2044 21476 2100 22878
rect 2044 21410 2100 21420
rect 2156 22258 2212 22270
rect 2156 22206 2158 22258
rect 2210 22206 2212 22258
rect 2156 21700 2212 22206
rect 2156 20468 2212 21644
rect 2156 20402 2212 20412
rect 1932 19460 1988 20076
rect 1932 19346 1988 19404
rect 1932 19294 1934 19346
rect 1986 19294 1988 19346
rect 1932 19282 1988 19294
rect 2044 20018 2100 20030
rect 2044 19966 2046 20018
rect 2098 19966 2100 20018
rect 2044 19236 2100 19966
rect 2156 19796 2212 19806
rect 2156 19702 2212 19740
rect 2268 19460 2324 24108
rect 2380 23940 2436 23950
rect 2380 23938 2548 23940
rect 2380 23886 2382 23938
rect 2434 23886 2548 23938
rect 2380 23884 2548 23886
rect 2380 23874 2436 23884
rect 2492 20132 2548 23884
rect 2716 23938 2772 24220
rect 2716 23886 2718 23938
rect 2770 23886 2772 23938
rect 2716 23874 2772 23886
rect 2828 24220 2996 24276
rect 2716 23716 2772 23726
rect 2716 23154 2772 23660
rect 2716 23102 2718 23154
rect 2770 23102 2772 23154
rect 2604 22484 2660 22494
rect 2604 22390 2660 22428
rect 2604 21700 2660 21710
rect 2604 20802 2660 21644
rect 2716 21588 2772 23102
rect 2716 21522 2772 21532
rect 2828 21364 2884 24220
rect 2940 24052 2996 24062
rect 2940 23958 2996 23996
rect 2940 21812 2996 21822
rect 3052 21812 3108 30158
rect 3276 28866 3332 34862
rect 3836 34902 3892 34914
rect 3836 34850 3838 34902
rect 3890 34850 3892 34902
rect 3836 34804 3892 34850
rect 3836 34738 3892 34748
rect 4172 34692 4228 35646
rect 4284 35140 4340 36428
rect 4508 36482 4564 36494
rect 4508 36430 4510 36482
rect 4562 36430 4564 36482
rect 4508 35812 4564 36430
rect 5180 36482 5236 37212
rect 5180 36430 5182 36482
rect 5234 36430 5236 36482
rect 5180 36418 5236 36430
rect 5404 36148 5460 38332
rect 5628 37938 5684 37950
rect 5628 37886 5630 37938
rect 5682 37886 5684 37938
rect 5628 37828 5684 37886
rect 5628 37762 5684 37772
rect 5740 37604 5796 38444
rect 6076 38500 6132 38510
rect 6076 38274 6132 38444
rect 6076 38222 6078 38274
rect 6130 38222 6132 38274
rect 5628 37548 5796 37604
rect 5852 37716 5908 37726
rect 5628 37380 5684 37548
rect 4508 35746 4564 35756
rect 5180 36092 5460 36148
rect 5516 37044 5572 37054
rect 5180 35812 5236 36092
rect 4464 35308 4728 35318
rect 4520 35252 4568 35308
rect 4624 35252 4672 35308
rect 4464 35242 4728 35252
rect 4284 35084 4900 35140
rect 3804 34524 4068 34534
rect 3612 34468 3668 34478
rect 3860 34468 3908 34524
rect 3964 34468 4012 34524
rect 3804 34458 4068 34468
rect 3500 34132 3556 34142
rect 3612 34132 3668 34412
rect 3724 34132 3780 34142
rect 3612 34076 3724 34132
rect 3500 34018 3556 34076
rect 3724 34066 3780 34076
rect 3948 34130 4004 34142
rect 3948 34078 3950 34130
rect 4002 34078 4004 34130
rect 3500 33966 3502 34018
rect 3554 33966 3556 34018
rect 3500 33954 3556 33966
rect 3948 33796 4004 34078
rect 4172 33908 4228 34636
rect 4172 33842 4228 33852
rect 4284 34914 4340 34926
rect 4284 34862 4286 34914
rect 4338 34862 4340 34914
rect 3948 33730 4004 33740
rect 4284 33572 4340 34862
rect 4732 34916 4788 34926
rect 4732 34822 4788 34860
rect 4464 33740 4728 33750
rect 4520 33684 4568 33740
rect 4624 33684 4672 33740
rect 4464 33674 4728 33684
rect 4284 33506 4340 33516
rect 3612 33460 3668 33470
rect 3612 33366 3668 33404
rect 3276 28814 3278 28866
rect 3330 28814 3332 28866
rect 3276 28802 3332 28814
rect 3388 33348 3444 33358
rect 3388 30212 3444 33292
rect 4284 33348 4340 33358
rect 4620 33348 4676 33358
rect 4284 33254 4340 33292
rect 4396 33346 4676 33348
rect 4396 33294 4622 33346
rect 4674 33294 4676 33346
rect 4396 33292 4676 33294
rect 4396 33124 4452 33292
rect 4620 33282 4676 33292
rect 4844 33346 4900 35084
rect 5068 34804 5124 34814
rect 5068 34132 5124 34748
rect 5180 34580 5236 35756
rect 5404 35588 5460 35598
rect 5292 35586 5460 35588
rect 5292 35534 5406 35586
rect 5458 35534 5460 35586
rect 5292 35532 5460 35534
rect 5292 34804 5348 35532
rect 5404 35522 5460 35532
rect 5516 35364 5572 36988
rect 5292 34738 5348 34748
rect 5404 35308 5572 35364
rect 5404 34692 5460 35308
rect 5516 34916 5572 34926
rect 5516 34822 5572 34860
rect 5404 34626 5460 34636
rect 5180 34524 5348 34580
rect 5068 34066 5124 34076
rect 4844 33294 4846 33346
rect 4898 33294 4900 33346
rect 4844 33282 4900 33294
rect 4956 33908 5012 33918
rect 4172 33068 4452 33124
rect 3804 32956 4068 32966
rect 3860 32900 3908 32956
rect 3964 32900 4012 32956
rect 3804 32890 4068 32900
rect 3612 31778 3668 31790
rect 3612 31726 3614 31778
rect 3666 31726 3668 31778
rect 3612 30436 3668 31726
rect 4172 31778 4228 33068
rect 4464 32172 4728 32182
rect 4520 32116 4568 32172
rect 4624 32116 4672 32172
rect 4464 32106 4728 32116
rect 4172 31726 4174 31778
rect 4226 31726 4228 31778
rect 4172 31714 4228 31726
rect 4844 31892 4900 31902
rect 3804 31388 4068 31398
rect 3860 31332 3908 31388
rect 3964 31332 4012 31388
rect 3804 31322 4068 31332
rect 4464 30604 4728 30614
rect 4520 30548 4568 30604
rect 4624 30548 4672 30604
rect 4464 30538 4728 30548
rect 3612 30370 3668 30380
rect 3724 30322 3780 30334
rect 3724 30270 3726 30322
rect 3778 30270 3780 30322
rect 3500 30212 3556 30222
rect 3388 30210 3556 30212
rect 3388 30158 3502 30210
rect 3554 30158 3556 30210
rect 3388 30156 3556 30158
rect 3388 29988 3444 30156
rect 3500 30146 3556 30156
rect 3724 29988 3780 30270
rect 3276 27860 3332 27870
rect 3164 27074 3220 27086
rect 3164 27022 3166 27074
rect 3218 27022 3220 27074
rect 3164 26068 3220 27022
rect 3164 26002 3220 26012
rect 3164 25506 3220 25518
rect 3164 25454 3166 25506
rect 3218 25454 3220 25506
rect 3164 25284 3220 25454
rect 3164 25218 3220 25228
rect 3164 22932 3220 22942
rect 3164 22838 3220 22876
rect 2940 21810 3108 21812
rect 2940 21758 2942 21810
rect 2994 21758 3108 21810
rect 2940 21756 3108 21758
rect 2940 21746 2996 21756
rect 3276 21700 3332 27804
rect 3388 24388 3444 29932
rect 3612 29932 3780 29988
rect 4172 30212 4228 30222
rect 3612 25284 3668 29932
rect 3804 29820 4068 29830
rect 3860 29764 3908 29820
rect 3964 29764 4012 29820
rect 3804 29754 4068 29764
rect 3804 28252 4068 28262
rect 3860 28196 3908 28252
rect 3964 28196 4012 28252
rect 3804 28186 4068 28196
rect 3948 27860 4004 27870
rect 3724 27300 3780 27310
rect 3724 27074 3780 27244
rect 3724 27022 3726 27074
rect 3778 27022 3780 27074
rect 3724 27010 3780 27022
rect 3948 27076 4004 27804
rect 3948 27010 4004 27020
rect 4172 27858 4228 30156
rect 4172 27806 4174 27858
rect 4226 27806 4228 27858
rect 4172 27076 4228 27806
rect 4172 27010 4228 27020
rect 4284 30210 4340 30222
rect 4284 30158 4286 30210
rect 4338 30158 4340 30210
rect 3804 26684 4068 26694
rect 3860 26628 3908 26684
rect 3964 26628 4012 26684
rect 3804 26618 4068 26628
rect 4172 26404 4228 26414
rect 3724 25732 3780 25742
rect 3724 25618 3780 25676
rect 4172 25730 4228 26348
rect 4172 25678 4174 25730
rect 4226 25678 4228 25730
rect 4172 25666 4228 25678
rect 4284 25732 4340 30158
rect 4844 30210 4900 31836
rect 4844 30158 4846 30210
rect 4898 30158 4900 30210
rect 4844 30146 4900 30158
rect 4956 31778 5012 33852
rect 4956 31726 4958 31778
rect 5010 31726 5012 31778
rect 4956 30212 5012 31726
rect 5068 33348 5124 33358
rect 5068 31218 5124 33292
rect 5068 31166 5070 31218
rect 5122 31166 5124 31218
rect 5068 31154 5124 31166
rect 4956 30146 5012 30156
rect 5068 30436 5124 30446
rect 5068 29650 5124 30380
rect 5068 29598 5070 29650
rect 5122 29598 5124 29650
rect 5068 29586 5124 29598
rect 4464 29036 4728 29046
rect 4520 28980 4568 29036
rect 4624 28980 4672 29036
rect 4464 28970 4728 28980
rect 5180 28642 5236 28654
rect 5180 28590 5182 28642
rect 5234 28590 5236 28642
rect 4464 27468 4728 27478
rect 4520 27412 4568 27468
rect 4624 27412 4672 27468
rect 4464 27402 4728 27412
rect 4508 27076 4564 27086
rect 4508 26982 4564 27020
rect 5180 27074 5236 28590
rect 5180 27022 5182 27074
rect 5234 27022 5236 27074
rect 5180 26852 5236 27022
rect 5180 26786 5236 26796
rect 5292 25956 5348 34524
rect 5628 34132 5684 37324
rect 5740 37156 5796 37166
rect 5740 35698 5796 37100
rect 5740 35646 5742 35698
rect 5794 35646 5796 35698
rect 5740 35634 5796 35646
rect 5852 35308 5908 37660
rect 6076 37716 6132 38222
rect 6076 37650 6132 37660
rect 6188 37828 6244 38780
rect 5628 34066 5684 34076
rect 5740 35252 5908 35308
rect 5964 37604 6020 37614
rect 5628 33908 5684 33918
rect 5516 33572 5572 33582
rect 5516 31892 5572 33516
rect 5628 33346 5684 33852
rect 5628 33294 5630 33346
rect 5682 33294 5684 33346
rect 5628 33282 5684 33294
rect 5628 31892 5684 31902
rect 5516 31890 5684 31892
rect 5516 31838 5630 31890
rect 5682 31838 5684 31890
rect 5516 31836 5684 31838
rect 5628 31826 5684 31836
rect 5740 31668 5796 35252
rect 5852 35140 5908 35150
rect 5852 34914 5908 35084
rect 5852 34862 5854 34914
rect 5906 34862 5908 34914
rect 5852 34850 5908 34862
rect 5852 34692 5908 34702
rect 5852 33012 5908 34636
rect 5964 33124 6020 37548
rect 6188 37380 6244 37772
rect 6300 37716 6356 42924
rect 6412 46060 6804 46116
rect 6412 41300 6468 46060
rect 6524 45892 6580 45902
rect 6524 45798 6580 45836
rect 6636 45778 6692 45790
rect 6636 45726 6638 45778
rect 6690 45726 6692 45778
rect 6636 45668 6692 45726
rect 6524 45106 6580 45118
rect 6524 45054 6526 45106
rect 6578 45054 6580 45106
rect 6524 43764 6580 45054
rect 6636 44322 6692 45612
rect 6860 45332 6916 50876
rect 6972 50428 7028 51542
rect 7084 51378 7140 51390
rect 7084 51326 7086 51378
rect 7138 51326 7140 51378
rect 7084 50596 7140 51326
rect 7084 50530 7140 50540
rect 6972 50372 7140 50428
rect 6972 49810 7028 49822
rect 6972 49758 6974 49810
rect 7026 49758 7028 49810
rect 6972 49700 7028 49758
rect 6972 49634 7028 49644
rect 7084 49364 7140 50372
rect 6972 49308 7140 49364
rect 6972 47348 7028 49308
rect 6972 47282 7028 47292
rect 7084 49138 7140 49150
rect 7084 49086 7086 49138
rect 7138 49086 7140 49138
rect 7084 48692 7140 49086
rect 7084 48132 7140 48636
rect 6972 47124 7028 47134
rect 6972 45444 7028 47068
rect 7084 46452 7140 48076
rect 7196 48356 7252 56924
rect 7420 55858 7476 55870
rect 7420 55806 7422 55858
rect 7474 55806 7476 55858
rect 7308 55298 7364 55310
rect 7308 55246 7310 55298
rect 7362 55246 7364 55298
rect 7308 54292 7364 55246
rect 7420 54514 7476 55806
rect 7756 54516 7812 54526
rect 7420 54462 7422 54514
rect 7474 54462 7476 54514
rect 7420 54450 7476 54462
rect 7644 54514 7812 54516
rect 7644 54462 7758 54514
rect 7810 54462 7812 54514
rect 7644 54460 7812 54462
rect 7644 54292 7700 54460
rect 7756 54450 7812 54460
rect 7308 54236 7700 54292
rect 7532 53620 7588 53630
rect 7420 49588 7476 49598
rect 7420 49494 7476 49532
rect 7532 48692 7588 53564
rect 7644 50596 7700 54236
rect 7868 53172 7924 69692
rect 7980 69522 8036 69534
rect 7980 69470 7982 69522
rect 8034 69470 8036 69522
rect 7980 68404 8036 69470
rect 7980 68338 8036 68348
rect 8092 68068 8148 69692
rect 8204 69636 8260 72494
rect 8204 69570 8260 69580
rect 8316 72436 8372 72446
rect 8316 69634 8372 72380
rect 8316 69582 8318 69634
rect 8370 69582 8372 69634
rect 8316 69570 8372 69582
rect 8092 67842 8148 68012
rect 8092 67790 8094 67842
rect 8146 67790 8148 67842
rect 8092 66274 8148 67790
rect 8092 66222 8094 66274
rect 8146 66222 8148 66274
rect 7980 63364 8036 63374
rect 7980 63270 8036 63308
rect 8092 62188 8148 66222
rect 8316 64820 8372 64830
rect 8204 64708 8260 64718
rect 8204 64614 8260 64652
rect 8204 64148 8260 64158
rect 8204 64054 8260 64092
rect 8316 63362 8372 64764
rect 8428 63812 8484 77532
rect 8540 75684 8596 75694
rect 8540 73330 8596 75628
rect 8764 73948 8820 79324
rect 9100 78706 9156 78718
rect 9100 78654 9102 78706
rect 9154 78654 9156 78706
rect 9100 78260 9156 78654
rect 9100 78194 9156 78204
rect 9212 78036 9268 79324
rect 9436 79286 9492 79324
rect 9548 78932 9604 79548
rect 9548 78838 9604 78876
rect 9100 77980 9268 78036
rect 9324 78596 9380 78606
rect 8988 77700 9044 77710
rect 8876 76468 8932 76478
rect 8876 76374 8932 76412
rect 8540 73278 8542 73330
rect 8594 73278 8596 73330
rect 8540 73266 8596 73278
rect 8652 73892 8820 73948
rect 8988 74114 9044 77644
rect 8988 74062 8990 74114
rect 9042 74062 9044 74114
rect 8652 67172 8708 73892
rect 8876 72884 8932 72894
rect 8876 71428 8932 72828
rect 8988 71876 9044 74062
rect 9100 72548 9156 77980
rect 9324 77476 9380 78540
rect 9660 78484 9716 80220
rect 9884 80052 9940 80446
rect 9884 79986 9940 79996
rect 9996 79858 10052 86716
rect 10108 84756 10164 87390
rect 10220 86436 10276 86446
rect 10220 85874 10276 86380
rect 10220 85822 10222 85874
rect 10274 85822 10276 85874
rect 10220 85810 10276 85822
rect 10108 84420 10164 84700
rect 10108 84354 10164 84364
rect 10332 83748 10388 92988
rect 10444 92930 10500 93884
rect 10444 92878 10446 92930
rect 10498 92878 10500 92930
rect 10444 92866 10500 92878
rect 10444 92148 10500 92158
rect 10556 92148 10612 95004
rect 10668 93268 10724 95116
rect 10780 94052 10836 95340
rect 11116 95284 11172 95294
rect 10780 93986 10836 93996
rect 10892 94612 10948 94622
rect 10892 93828 10948 94556
rect 11004 94386 11060 94398
rect 11004 94334 11006 94386
rect 11058 94334 11060 94386
rect 11004 94164 11060 94334
rect 11004 94098 11060 94108
rect 10892 93772 11060 93828
rect 10780 93716 10836 93726
rect 10780 93604 10836 93660
rect 10780 93548 10948 93604
rect 10668 93202 10724 93212
rect 10780 93380 10836 93390
rect 10444 92146 10612 92148
rect 10444 92094 10446 92146
rect 10498 92094 10612 92146
rect 10444 92092 10612 92094
rect 10444 92082 10500 92092
rect 10780 91476 10836 93324
rect 10892 92932 10948 93548
rect 10892 92838 10948 92876
rect 10668 91420 10836 91476
rect 10892 91476 10948 91486
rect 10556 91250 10612 91262
rect 10556 91198 10558 91250
rect 10610 91198 10612 91250
rect 10556 89124 10612 91198
rect 10556 89058 10612 89068
rect 10556 84420 10612 84430
rect 10556 84306 10612 84364
rect 10556 84254 10558 84306
rect 10610 84254 10612 84306
rect 10556 84242 10612 84254
rect 10332 83692 10500 83748
rect 10332 83524 10388 83534
rect 10332 83430 10388 83468
rect 10220 82740 10276 82750
rect 10108 82516 10164 82526
rect 10108 82180 10164 82460
rect 10108 81844 10164 82124
rect 10220 82066 10276 82684
rect 10220 82014 10222 82066
rect 10274 82014 10276 82066
rect 10220 82002 10276 82014
rect 10332 82516 10388 82526
rect 10108 81788 10276 81844
rect 9828 79802 10052 79858
rect 10108 80946 10164 80958
rect 10108 80894 10110 80946
rect 10162 80894 10164 80946
rect 9828 79716 9884 79802
rect 9828 79660 9940 79716
rect 9436 78148 9492 78158
rect 9436 78054 9492 78092
rect 9548 78036 9604 78046
rect 9548 77588 9604 77980
rect 9660 77700 9716 78428
rect 9660 77634 9716 77644
rect 9772 77924 9828 77934
rect 9548 77522 9604 77532
rect 9436 77476 9492 77486
rect 9324 77420 9436 77476
rect 9212 77362 9268 77374
rect 9212 77310 9214 77362
rect 9266 77310 9268 77362
rect 9212 77252 9268 77310
rect 9324 77252 9380 77262
rect 9212 77196 9324 77252
rect 9324 77186 9380 77196
rect 9436 74226 9492 77420
rect 9548 77252 9604 77262
rect 9548 77158 9604 77196
rect 9772 76466 9828 77868
rect 9772 76414 9774 76466
rect 9826 76414 9828 76466
rect 9772 76402 9828 76414
rect 9884 77362 9940 79660
rect 9996 79604 10052 79614
rect 10108 79604 10164 80894
rect 10220 80724 10276 81788
rect 10332 80948 10388 82460
rect 10332 80882 10388 80892
rect 10220 80668 10388 80724
rect 9996 79602 10164 79604
rect 9996 79550 9998 79602
rect 10050 79550 10164 79602
rect 9996 79548 10164 79550
rect 10220 80500 10276 80510
rect 9996 79538 10052 79548
rect 10108 79380 10164 79390
rect 10108 78484 10164 79324
rect 9996 78428 10164 78484
rect 9996 77924 10052 78428
rect 10108 78260 10164 78270
rect 10108 78146 10164 78204
rect 10108 78094 10110 78146
rect 10162 78094 10164 78146
rect 10108 78082 10164 78094
rect 9996 77868 10164 77924
rect 9884 77310 9886 77362
rect 9938 77310 9940 77362
rect 9884 76468 9940 77310
rect 9884 76402 9940 76412
rect 9436 74174 9438 74226
rect 9490 74174 9492 74226
rect 9436 74162 9492 74174
rect 9884 74116 9940 74126
rect 9548 73892 9604 73902
rect 9324 73556 9380 73566
rect 9324 73330 9380 73500
rect 9324 73278 9326 73330
rect 9378 73278 9380 73330
rect 9212 73106 9268 73118
rect 9212 73054 9214 73106
rect 9266 73054 9268 73106
rect 9212 72884 9268 73054
rect 9324 73108 9380 73278
rect 9324 73042 9380 73052
rect 9212 72818 9268 72828
rect 9436 72770 9492 72782
rect 9436 72718 9438 72770
rect 9490 72718 9492 72770
rect 9436 72548 9492 72718
rect 9100 72492 9268 72548
rect 9100 72324 9156 72334
rect 9100 72230 9156 72268
rect 8988 71810 9044 71820
rect 8876 71362 8932 71372
rect 9212 71762 9268 72492
rect 9436 72482 9492 72492
rect 9548 72546 9604 73836
rect 9772 73332 9828 73342
rect 9772 73238 9828 73276
rect 9884 72658 9940 74060
rect 10108 72772 10164 77868
rect 10220 76356 10276 80444
rect 10332 79380 10388 80668
rect 10444 79828 10500 83692
rect 10556 82738 10612 82750
rect 10556 82686 10558 82738
rect 10610 82686 10612 82738
rect 10556 82516 10612 82686
rect 10668 82628 10724 91420
rect 10892 91382 10948 91420
rect 11004 90356 11060 93772
rect 11116 92148 11172 95228
rect 11228 93716 11284 96014
rect 11452 94500 11508 94510
rect 11564 94500 11620 96796
rect 11452 94498 11620 94500
rect 11452 94446 11454 94498
rect 11506 94446 11620 94498
rect 11452 94444 11620 94446
rect 11676 96180 11732 99148
rect 11900 99428 11956 99438
rect 11900 99202 11956 99372
rect 11900 99150 11902 99202
rect 11954 99150 11956 99202
rect 11900 99138 11956 99150
rect 11788 97972 11844 97982
rect 11788 97858 11844 97916
rect 11788 97806 11790 97858
rect 11842 97806 11844 97858
rect 11788 97794 11844 97806
rect 12012 97468 12068 102956
rect 12684 102452 12740 102462
rect 12460 102114 12516 102126
rect 12460 102062 12462 102114
rect 12514 102062 12516 102114
rect 12460 101892 12516 102062
rect 12460 101826 12516 101836
rect 12348 100884 12404 100894
rect 12124 99988 12180 99998
rect 12124 99894 12180 99932
rect 12012 97412 12292 97468
rect 12124 97300 12180 97310
rect 11452 94434 11508 94444
rect 11228 93650 11284 93660
rect 11564 93716 11620 93726
rect 11564 93622 11620 93660
rect 11676 93044 11732 96124
rect 12012 96852 12068 96862
rect 12012 94722 12068 96796
rect 12124 96066 12180 97244
rect 12124 96014 12126 96066
rect 12178 96014 12180 96066
rect 12124 96002 12180 96014
rect 12012 94670 12014 94722
rect 12066 94670 12068 94722
rect 12012 94658 12068 94670
rect 12236 94724 12292 97412
rect 11900 94612 11956 94622
rect 11900 94498 11956 94556
rect 11900 94446 11902 94498
rect 11954 94446 11956 94498
rect 11900 94108 11956 94446
rect 11676 92978 11732 92988
rect 11788 94052 11956 94108
rect 11788 92708 11844 94052
rect 11788 92642 11844 92652
rect 11900 93716 11956 93726
rect 11900 92930 11956 93660
rect 11900 92878 11902 92930
rect 11954 92878 11956 92930
rect 11900 92484 11956 92878
rect 11900 92418 11956 92428
rect 11228 92148 11284 92158
rect 11116 92146 11284 92148
rect 11116 92094 11230 92146
rect 11282 92094 11284 92146
rect 11116 92092 11284 92094
rect 11116 90356 11172 90366
rect 11004 90300 11116 90356
rect 11116 90262 11172 90300
rect 11228 90132 11284 92092
rect 12124 91364 12180 91374
rect 12124 91270 12180 91308
rect 11900 90916 11956 90926
rect 11676 90578 11732 90590
rect 11676 90526 11678 90578
rect 11730 90526 11732 90578
rect 11676 90244 11732 90526
rect 11676 90178 11732 90188
rect 11116 90076 11284 90132
rect 11116 89012 11172 90076
rect 11228 89572 11284 89582
rect 11228 89478 11284 89516
rect 11788 89572 11844 89582
rect 11116 88946 11172 88956
rect 11228 88788 11284 88798
rect 10780 88786 11284 88788
rect 10780 88734 11230 88786
rect 11282 88734 11284 88786
rect 10780 88732 11284 88734
rect 10780 87442 10836 88732
rect 11228 88722 11284 88732
rect 11452 88340 11508 88350
rect 11452 88246 11508 88284
rect 10780 87390 10782 87442
rect 10834 87390 10836 87442
rect 10780 87378 10836 87390
rect 11004 88114 11060 88126
rect 11004 88062 11006 88114
rect 11058 88062 11060 88114
rect 11004 87332 11060 88062
rect 11452 87556 11508 87566
rect 11004 87266 11060 87276
rect 11228 87444 11284 87454
rect 11228 87330 11284 87388
rect 11452 87442 11508 87500
rect 11452 87390 11454 87442
rect 11506 87390 11508 87442
rect 11452 87378 11508 87390
rect 11564 87444 11620 87454
rect 11228 87278 11230 87330
rect 11282 87278 11284 87330
rect 11228 87266 11284 87278
rect 11340 86884 11396 86894
rect 11004 86660 11060 86670
rect 11004 86566 11060 86604
rect 11340 86324 11396 86828
rect 11452 86772 11508 86782
rect 11564 86772 11620 87388
rect 11788 87442 11844 89516
rect 11788 87390 11790 87442
rect 11842 87390 11844 87442
rect 11788 87378 11844 87390
rect 11452 86770 11620 86772
rect 11452 86718 11454 86770
rect 11506 86718 11620 86770
rect 11452 86716 11620 86718
rect 11452 86706 11508 86716
rect 11004 86100 11060 86110
rect 11004 85874 11060 86044
rect 11004 85822 11006 85874
rect 11058 85822 11060 85874
rect 10892 85316 10948 85326
rect 10892 85090 10948 85260
rect 10892 85038 10894 85090
rect 10946 85038 10948 85090
rect 10892 85026 10948 85038
rect 11004 82964 11060 85822
rect 11004 82898 11060 82908
rect 11116 85988 11172 85998
rect 11116 83522 11172 85932
rect 11228 85204 11284 85214
rect 11228 85110 11284 85148
rect 11116 83470 11118 83522
rect 11170 83470 11172 83522
rect 10892 82628 10948 82638
rect 10668 82626 10948 82628
rect 10668 82574 10894 82626
rect 10946 82574 10948 82626
rect 10668 82572 10948 82574
rect 10892 82562 10948 82572
rect 10556 82450 10612 82460
rect 11004 82404 11060 82414
rect 10668 81956 10724 81966
rect 11004 81956 11060 82348
rect 10668 81954 11060 81956
rect 10668 81902 10670 81954
rect 10722 81902 11060 81954
rect 10668 81900 11060 81902
rect 11116 81956 11172 83470
rect 10668 81890 10724 81900
rect 11116 81890 11172 81900
rect 11228 84644 11284 84654
rect 10668 81508 10724 81518
rect 10556 81058 10612 81070
rect 10556 81006 10558 81058
rect 10610 81006 10612 81058
rect 10556 80164 10612 81006
rect 10556 80098 10612 80108
rect 10444 79762 10500 79772
rect 10668 79604 10724 81452
rect 10892 81284 10948 81294
rect 10892 81282 11060 81284
rect 10892 81230 10894 81282
rect 10946 81230 11060 81282
rect 10892 81228 11060 81230
rect 10892 81218 10948 81228
rect 10780 80948 10836 80958
rect 10780 80854 10836 80892
rect 10892 79940 10948 79950
rect 10668 79602 10836 79604
rect 10668 79550 10670 79602
rect 10722 79550 10836 79602
rect 10668 79548 10836 79550
rect 10668 79538 10724 79548
rect 10332 79314 10388 79324
rect 10780 78708 10836 79548
rect 10780 78642 10836 78652
rect 10668 78594 10724 78606
rect 10668 78542 10670 78594
rect 10722 78542 10724 78594
rect 10668 78484 10724 78542
rect 10332 78428 10724 78484
rect 10332 77250 10388 78428
rect 10892 78372 10948 79884
rect 11004 78932 11060 81228
rect 11228 80612 11284 84588
rect 11340 84420 11396 86268
rect 11340 84326 11396 84364
rect 11452 84980 11508 84990
rect 11228 80546 11284 80556
rect 11340 83188 11396 83198
rect 11116 80164 11172 80174
rect 11116 80162 11284 80164
rect 11116 80110 11118 80162
rect 11170 80110 11284 80162
rect 11116 80108 11284 80110
rect 11116 80098 11172 80108
rect 11228 78932 11284 80108
rect 11004 78876 11172 78932
rect 11116 78818 11172 78876
rect 11228 78866 11284 78876
rect 11116 78766 11118 78818
rect 11170 78766 11172 78818
rect 11116 78754 11172 78766
rect 10892 78306 10948 78316
rect 11228 78708 11284 78718
rect 11228 78372 11284 78652
rect 11228 78306 11284 78316
rect 10332 77198 10334 77250
rect 10386 77198 10388 77250
rect 10332 77186 10388 77198
rect 10444 78260 10500 78270
rect 10220 76290 10276 76300
rect 10444 76466 10500 78204
rect 11340 78260 11396 83132
rect 11452 79940 11508 84924
rect 11452 79874 11508 79884
rect 11452 79716 11508 79726
rect 11452 79602 11508 79660
rect 11452 79550 11454 79602
rect 11506 79550 11508 79602
rect 11452 79538 11508 79550
rect 11452 79044 11508 79054
rect 11452 78950 11508 78988
rect 11452 78596 11508 78606
rect 11452 78502 11508 78540
rect 11340 78194 11396 78204
rect 10444 76414 10446 76466
rect 10498 76414 10500 76466
rect 10444 73948 10500 76414
rect 10556 77924 10612 77934
rect 11564 77924 11620 86716
rect 11788 86660 11844 86670
rect 11788 86566 11844 86604
rect 11900 85708 11956 90860
rect 12236 90804 12292 94668
rect 12012 90748 12292 90804
rect 12012 85876 12068 90748
rect 12124 90580 12180 90590
rect 12124 87556 12180 90524
rect 12236 90132 12292 90142
rect 12236 90018 12292 90076
rect 12236 89966 12238 90018
rect 12290 89966 12292 90018
rect 12236 89954 12292 89966
rect 12236 87556 12292 87566
rect 12124 87554 12292 87556
rect 12124 87502 12238 87554
rect 12290 87502 12292 87554
rect 12124 87500 12292 87502
rect 12236 87490 12292 87500
rect 12012 85810 12068 85820
rect 12348 86658 12404 100828
rect 12572 100770 12628 100782
rect 12572 100718 12574 100770
rect 12626 100718 12628 100770
rect 12572 99204 12628 100718
rect 12572 99138 12628 99148
rect 12684 97468 12740 102396
rect 12908 102452 12964 102462
rect 13020 102452 13076 103516
rect 13132 103124 13188 103134
rect 13132 103122 13412 103124
rect 13132 103070 13134 103122
rect 13186 103070 13412 103122
rect 13132 103068 13412 103070
rect 13132 103058 13188 103068
rect 12908 102450 13188 102452
rect 12908 102398 12910 102450
rect 12962 102398 13188 102450
rect 12908 102396 13188 102398
rect 12908 102386 12964 102396
rect 13132 101668 13188 102396
rect 13244 102338 13300 102350
rect 13244 102286 13246 102338
rect 13298 102286 13300 102338
rect 13244 101892 13300 102286
rect 13244 101826 13300 101836
rect 13244 101668 13300 101678
rect 13132 101666 13300 101668
rect 13132 101614 13246 101666
rect 13298 101614 13300 101666
rect 13132 101612 13300 101614
rect 12908 101556 12964 101566
rect 12908 100210 12964 101500
rect 12908 100158 12910 100210
rect 12962 100158 12964 100210
rect 12908 100146 12964 100158
rect 13132 100212 13188 100222
rect 12908 99204 12964 99214
rect 12908 99110 12964 99148
rect 12572 97412 12740 97468
rect 13020 98644 13076 98654
rect 13020 98418 13076 98588
rect 13020 98366 13022 98418
rect 13074 98366 13076 98418
rect 13020 97524 13076 98366
rect 13020 97458 13076 97468
rect 12460 96068 12516 96078
rect 12460 95974 12516 96012
rect 12460 90804 12516 90814
rect 12460 87780 12516 90748
rect 12572 90132 12628 97412
rect 12908 97410 12964 97422
rect 12908 97358 12910 97410
rect 12962 97358 12964 97410
rect 12684 97300 12740 97310
rect 12684 94498 12740 97244
rect 12908 97300 12964 97358
rect 12908 97234 12964 97244
rect 12684 94446 12686 94498
rect 12738 94446 12740 94498
rect 12684 94434 12740 94446
rect 12796 97076 12852 97086
rect 12684 92930 12740 92942
rect 12684 92878 12686 92930
rect 12738 92878 12740 92930
rect 12684 91588 12740 92878
rect 12684 91522 12740 91532
rect 12796 91476 12852 97020
rect 13020 96850 13076 96862
rect 13020 96798 13022 96850
rect 13074 96798 13076 96850
rect 12908 96738 12964 96750
rect 12908 96686 12910 96738
rect 12962 96686 12964 96738
rect 12908 96292 12964 96686
rect 12908 96226 12964 96236
rect 12908 95508 12964 95518
rect 13020 95508 13076 96798
rect 12908 95506 13076 95508
rect 12908 95454 12910 95506
rect 12962 95454 13076 95506
rect 12908 95452 13076 95454
rect 12908 95442 12964 95452
rect 13020 94498 13076 94510
rect 13020 94446 13022 94498
rect 13074 94446 13076 94498
rect 12908 93042 12964 93054
rect 12908 92990 12910 93042
rect 12962 92990 12964 93042
rect 12908 92484 12964 92990
rect 12908 92418 12964 92428
rect 12908 91476 12964 91486
rect 12796 91474 12964 91476
rect 12796 91422 12910 91474
rect 12962 91422 12964 91474
rect 12796 91420 12964 91422
rect 12908 91410 12964 91420
rect 13020 90692 13076 94446
rect 13132 93716 13188 100156
rect 13244 95844 13300 101612
rect 13356 100212 13412 103068
rect 13356 100146 13412 100156
rect 13468 102452 13524 102462
rect 13468 99876 13524 102396
rect 13580 102340 13636 104638
rect 13692 105362 13748 105374
rect 13692 105310 13694 105362
rect 13746 105310 13748 105362
rect 13692 105252 13748 105310
rect 13804 105364 13860 105644
rect 13804 105298 13860 105308
rect 13692 103796 13748 105196
rect 13692 103122 13748 103740
rect 13804 104466 13860 104478
rect 13804 104414 13806 104466
rect 13858 104414 13860 104466
rect 13804 103348 13860 104414
rect 13804 103282 13860 103292
rect 13692 103070 13694 103122
rect 13746 103070 13748 103122
rect 13692 102564 13748 103070
rect 13916 102676 13972 106988
rect 13692 102498 13748 102508
rect 13804 102620 13972 102676
rect 14028 106484 14084 106494
rect 13692 102340 13748 102350
rect 13580 102338 13748 102340
rect 13580 102286 13694 102338
rect 13746 102286 13748 102338
rect 13580 102284 13748 102286
rect 13580 101556 13636 101566
rect 13580 101462 13636 101500
rect 13468 98084 13524 99820
rect 13244 95778 13300 95788
rect 13356 98028 13524 98084
rect 13580 101332 13636 101342
rect 13580 98306 13636 101276
rect 13692 100884 13748 102284
rect 13692 100818 13748 100828
rect 13580 98254 13582 98306
rect 13634 98254 13636 98306
rect 13244 94500 13300 94510
rect 13356 94500 13412 98028
rect 13468 96180 13524 96190
rect 13468 96066 13524 96124
rect 13468 96014 13470 96066
rect 13522 96014 13524 96066
rect 13468 96002 13524 96014
rect 13244 94498 13412 94500
rect 13244 94446 13246 94498
rect 13298 94446 13412 94498
rect 13244 94444 13412 94446
rect 13244 94434 13300 94444
rect 13132 93650 13188 93660
rect 13468 94052 13524 94062
rect 13468 93492 13524 93996
rect 13580 93940 13636 98254
rect 13804 97524 13860 102620
rect 13916 102452 13972 102462
rect 13916 102358 13972 102396
rect 14028 102228 14084 106428
rect 14140 103460 14196 107772
rect 14252 107826 14308 109900
rect 14252 107774 14254 107826
rect 14306 107774 14308 107826
rect 14252 107762 14308 107774
rect 14364 107492 14420 111132
rect 14588 110964 14644 110974
rect 14476 110740 14532 110750
rect 14476 109396 14532 110684
rect 14588 110178 14644 110908
rect 14588 110126 14590 110178
rect 14642 110126 14644 110178
rect 14588 110114 14644 110126
rect 14476 109330 14532 109340
rect 14812 108836 14868 108846
rect 14924 108836 14980 111580
rect 15036 111412 15092 113262
rect 15148 113316 15204 113326
rect 15148 112530 15204 113260
rect 15260 112644 15316 114800
rect 15372 114212 15428 114222
rect 15372 113538 15428 114156
rect 15372 113486 15374 113538
rect 15426 113486 15428 113538
rect 15372 113474 15428 113486
rect 15260 112578 15316 112588
rect 15372 113316 15428 113326
rect 15148 112478 15150 112530
rect 15202 112478 15204 112530
rect 15148 112466 15204 112478
rect 15036 111346 15092 111356
rect 15148 110964 15204 110974
rect 15148 110870 15204 110908
rect 15036 110178 15092 110190
rect 15036 110126 15038 110178
rect 15090 110126 15092 110178
rect 15036 109620 15092 110126
rect 15036 109554 15092 109564
rect 15036 109284 15092 109294
rect 15036 109282 15316 109284
rect 15036 109230 15038 109282
rect 15090 109230 15316 109282
rect 15036 109228 15316 109230
rect 15036 109218 15092 109228
rect 14812 108834 14980 108836
rect 14812 108782 14814 108834
rect 14866 108782 14980 108834
rect 14812 108780 14980 108782
rect 15148 109172 15316 109228
rect 14812 108770 14868 108780
rect 15036 108610 15092 108622
rect 15036 108558 15038 108610
rect 15090 108558 15092 108610
rect 14700 107714 14756 107726
rect 14700 107662 14702 107714
rect 14754 107662 14756 107714
rect 14700 107604 14756 107662
rect 15036 107716 15092 108558
rect 15148 107826 15204 109172
rect 15148 107774 15150 107826
rect 15202 107774 15204 107826
rect 15148 107762 15204 107774
rect 15260 108948 15316 108958
rect 15036 107650 15092 107660
rect 14700 107538 14756 107548
rect 14364 107426 14420 107436
rect 14812 107492 14868 107502
rect 14588 106932 14644 106942
rect 14588 106838 14644 106876
rect 14588 106034 14644 106046
rect 14588 105982 14590 106034
rect 14642 105982 14644 106034
rect 14364 105474 14420 105486
rect 14364 105422 14366 105474
rect 14418 105422 14420 105474
rect 14364 105252 14420 105422
rect 14364 105186 14420 105196
rect 14252 105028 14308 105038
rect 14252 104130 14308 104972
rect 14476 104692 14532 104702
rect 14588 104692 14644 105982
rect 14476 104690 14644 104692
rect 14476 104638 14478 104690
rect 14530 104638 14644 104690
rect 14476 104636 14644 104638
rect 14476 104626 14532 104636
rect 14252 104078 14254 104130
rect 14306 104078 14308 104130
rect 14252 104066 14308 104078
rect 14700 103796 14756 103806
rect 14700 103702 14756 103740
rect 14140 103404 14420 103460
rect 13916 102172 14084 102228
rect 14140 103236 14196 103246
rect 14140 102898 14196 103180
rect 14140 102846 14142 102898
rect 14194 102846 14196 102898
rect 13916 100770 13972 102172
rect 14140 101668 14196 102846
rect 14140 101602 14196 101612
rect 14028 101554 14084 101566
rect 14028 101502 14030 101554
rect 14082 101502 14084 101554
rect 14028 100884 14084 101502
rect 14252 101332 14308 101342
rect 14028 100818 14084 100828
rect 14140 101330 14308 101332
rect 14140 101278 14254 101330
rect 14306 101278 14308 101330
rect 14140 101276 14308 101278
rect 13916 100718 13918 100770
rect 13970 100718 13972 100770
rect 13916 100212 13972 100718
rect 13916 100146 13972 100156
rect 14140 99988 14196 101276
rect 14252 101266 14308 101276
rect 14028 99762 14084 99774
rect 14028 99710 14030 99762
rect 14082 99710 14084 99762
rect 14028 99428 14084 99710
rect 14028 99362 14084 99372
rect 14140 97748 14196 99932
rect 14252 100882 14308 100894
rect 14252 100830 14254 100882
rect 14306 100830 14308 100882
rect 14252 100772 14308 100830
rect 14252 97860 14308 100716
rect 14364 99316 14420 103404
rect 14588 102340 14644 102350
rect 14588 102246 14644 102284
rect 14476 100212 14532 100222
rect 14476 100100 14532 100156
rect 14476 100098 14644 100100
rect 14476 100046 14478 100098
rect 14530 100046 14644 100098
rect 14476 100044 14644 100046
rect 14476 100034 14532 100044
rect 14364 99260 14532 99316
rect 14364 99090 14420 99102
rect 14364 99038 14366 99090
rect 14418 99038 14420 99090
rect 14364 98084 14420 99038
rect 14364 98018 14420 98028
rect 14476 97860 14532 99260
rect 14252 97804 14420 97860
rect 14140 97692 14308 97748
rect 13748 97468 13860 97524
rect 13748 97412 13804 97468
rect 13748 97356 13860 97412
rect 13692 96852 13748 96862
rect 13692 96758 13748 96796
rect 13580 93884 13748 93940
rect 13468 93426 13524 93436
rect 13580 93714 13636 93726
rect 13580 93662 13582 93714
rect 13634 93662 13636 93714
rect 13580 93268 13636 93662
rect 13580 92932 13636 93212
rect 13468 92706 13524 92718
rect 13468 92654 13470 92706
rect 13522 92654 13524 92706
rect 13020 90626 13076 90636
rect 13244 91364 13300 91374
rect 12796 90468 12852 90478
rect 12796 90374 12852 90412
rect 13132 90468 13188 90478
rect 13132 90374 13188 90412
rect 12572 90076 12740 90132
rect 12572 89908 12628 89918
rect 12572 89814 12628 89852
rect 12684 88228 12740 90076
rect 13244 89794 13300 91308
rect 13356 91362 13412 91374
rect 13356 91310 13358 91362
rect 13410 91310 13412 91362
rect 13356 90132 13412 91310
rect 13468 90356 13524 92654
rect 13468 90290 13524 90300
rect 13580 92146 13636 92876
rect 13580 92094 13582 92146
rect 13634 92094 13636 92146
rect 13580 90578 13636 92094
rect 13580 90526 13582 90578
rect 13634 90526 13636 90578
rect 13580 90244 13636 90526
rect 13580 90178 13636 90188
rect 13356 90066 13412 90076
rect 13244 89742 13246 89794
rect 13298 89742 13300 89794
rect 13244 89730 13300 89742
rect 13692 89796 13748 93884
rect 13804 93154 13860 97356
rect 13916 96964 13972 96974
rect 13916 96292 13972 96908
rect 13916 96226 13972 96236
rect 14028 96626 14084 96638
rect 14028 96574 14030 96626
rect 14082 96574 14084 96626
rect 14028 95844 14084 96574
rect 14028 95778 14084 95788
rect 14252 95396 14308 97692
rect 14028 95340 14308 95396
rect 14028 94500 14084 95340
rect 14140 95172 14196 95182
rect 14196 95116 14308 95172
rect 14140 95078 14196 95116
rect 14140 94500 14196 94510
rect 14028 94498 14196 94500
rect 14028 94446 14142 94498
rect 14194 94446 14196 94498
rect 14028 94444 14196 94446
rect 13916 94388 13972 94398
rect 13972 94332 14084 94388
rect 13916 94322 13972 94332
rect 13804 93102 13806 93154
rect 13858 93102 13860 93154
rect 13804 93090 13860 93102
rect 13916 94164 13972 94174
rect 13916 93156 13972 94108
rect 14028 93828 14084 94332
rect 14140 94052 14196 94444
rect 14140 93986 14196 93996
rect 14028 93772 14196 93828
rect 14028 93490 14084 93502
rect 14028 93438 14030 93490
rect 14082 93438 14084 93490
rect 14028 93380 14084 93438
rect 14028 93314 14084 93324
rect 13916 93100 14084 93156
rect 13916 92484 13972 92494
rect 13916 91586 13972 92428
rect 13916 91534 13918 91586
rect 13970 91534 13972 91586
rect 13916 91522 13972 91534
rect 14028 92034 14084 93100
rect 14028 91982 14030 92034
rect 14082 91982 14084 92034
rect 13804 91362 13860 91374
rect 13804 91310 13806 91362
rect 13858 91310 13860 91362
rect 13804 91140 13860 91310
rect 14028 91252 14084 91982
rect 14028 91186 14084 91196
rect 13804 91074 13860 91084
rect 13916 90356 13972 90366
rect 13916 90018 13972 90300
rect 14140 90354 14196 93772
rect 14140 90302 14142 90354
rect 14194 90302 14196 90354
rect 14140 90020 14196 90302
rect 13916 89966 13918 90018
rect 13970 89966 13972 90018
rect 13916 89954 13972 89966
rect 14028 89964 14196 90020
rect 13692 89730 13748 89740
rect 13804 89794 13860 89806
rect 14028 89796 14084 89964
rect 13804 89742 13806 89794
rect 13858 89742 13860 89794
rect 12908 89684 12964 89694
rect 12908 89682 13188 89684
rect 12908 89630 12910 89682
rect 12962 89630 13188 89682
rect 12908 89628 13188 89630
rect 12908 89618 12964 89628
rect 13020 89124 13076 89134
rect 13020 89030 13076 89068
rect 13132 88452 13188 89628
rect 13356 88898 13412 88910
rect 13356 88846 13358 88898
rect 13410 88846 13412 88898
rect 13356 88676 13412 88846
rect 13356 88610 13412 88620
rect 13132 88396 13412 88452
rect 12684 88162 12740 88172
rect 13244 88228 13300 88238
rect 12572 88004 12628 88014
rect 12572 88002 12964 88004
rect 12572 87950 12574 88002
rect 12626 87950 12964 88002
rect 12572 87948 12964 87950
rect 12572 87938 12628 87948
rect 12796 87780 12852 87790
rect 12460 87724 12740 87780
rect 12460 86772 12516 86782
rect 12460 86678 12516 86716
rect 12348 86606 12350 86658
rect 12402 86606 12404 86658
rect 11788 85652 11956 85708
rect 11676 78932 11732 78942
rect 11676 78708 11732 78876
rect 11676 78642 11732 78652
rect 10556 77810 10612 77868
rect 10556 77758 10558 77810
rect 10610 77758 10612 77810
rect 10556 76132 10612 77758
rect 11452 77868 11620 77924
rect 10892 77362 10948 77374
rect 10892 77310 10894 77362
rect 10946 77310 10948 77362
rect 10556 76066 10612 76076
rect 10780 77250 10836 77262
rect 10780 77198 10782 77250
rect 10834 77198 10836 77250
rect 10556 74900 10612 74910
rect 10556 74898 10724 74900
rect 10556 74846 10558 74898
rect 10610 74846 10724 74898
rect 10556 74844 10724 74846
rect 10556 74834 10612 74844
rect 10668 74116 10724 74844
rect 10668 74050 10724 74060
rect 10332 73892 10500 73948
rect 10668 73892 10724 73902
rect 10220 73444 10276 73454
rect 10220 73350 10276 73388
rect 10332 72996 10388 73892
rect 10668 73798 10724 73836
rect 10556 73668 10612 73678
rect 10556 73554 10612 73612
rect 10556 73502 10558 73554
rect 10610 73502 10612 73554
rect 10556 73490 10612 73502
rect 10780 73556 10836 77198
rect 10892 77252 10948 77310
rect 10892 77186 10948 77196
rect 11452 77028 11508 77868
rect 11676 77812 11732 77822
rect 11564 77810 11732 77812
rect 11564 77758 11678 77810
rect 11730 77758 11732 77810
rect 11564 77756 11732 77758
rect 11564 77250 11620 77756
rect 11676 77746 11732 77756
rect 11564 77198 11566 77250
rect 11618 77198 11620 77250
rect 11564 77186 11620 77198
rect 11676 77364 11732 77374
rect 11452 76972 11620 77028
rect 10892 76356 10948 76366
rect 10892 76262 10948 76300
rect 11228 76356 11284 76366
rect 11004 75124 11060 75134
rect 11004 74786 11060 75068
rect 11004 74734 11006 74786
rect 11058 74734 11060 74786
rect 11004 74722 11060 74734
rect 11228 73948 11284 76300
rect 10780 73490 10836 73500
rect 11004 73892 11284 73948
rect 11452 74116 11508 74126
rect 11452 74002 11508 74060
rect 11452 73950 11454 74002
rect 11506 73950 11508 74002
rect 11340 73892 11396 73902
rect 10780 73220 10836 73230
rect 10780 73126 10836 73164
rect 10668 73106 10724 73118
rect 10668 73054 10670 73106
rect 10722 73054 10724 73106
rect 10332 72940 10500 72996
rect 10332 72772 10388 72810
rect 10108 72716 10276 72772
rect 9884 72606 9886 72658
rect 9938 72606 9940 72658
rect 9884 72594 9940 72606
rect 9548 72494 9550 72546
rect 9602 72494 9604 72546
rect 9548 72482 9604 72494
rect 10108 72546 10164 72558
rect 10108 72494 10110 72546
rect 10162 72494 10164 72546
rect 9324 72436 9380 72446
rect 9324 72342 9380 72380
rect 9772 72436 9828 72446
rect 9772 71986 9828 72380
rect 10108 72436 10164 72494
rect 10108 72370 10164 72380
rect 9772 71934 9774 71986
rect 9826 71934 9828 71986
rect 9772 71922 9828 71934
rect 10108 72212 10164 72222
rect 9212 71710 9214 71762
rect 9266 71710 9268 71762
rect 9212 71204 9268 71710
rect 9212 71148 9604 71204
rect 8876 71090 8932 71102
rect 8876 71038 8878 71090
rect 8930 71038 8932 71090
rect 8876 69300 8932 71038
rect 9100 70978 9156 70990
rect 9100 70926 9102 70978
rect 9154 70926 9156 70978
rect 9100 70532 9156 70926
rect 9100 70466 9156 70476
rect 9212 70364 9492 70420
rect 8988 70308 9044 70318
rect 9212 70308 9268 70364
rect 8988 70306 9268 70308
rect 8988 70254 8990 70306
rect 9042 70254 9268 70306
rect 8988 70252 9268 70254
rect 8988 70242 9044 70252
rect 9324 70196 9380 70206
rect 9212 70194 9380 70196
rect 9212 70142 9326 70194
rect 9378 70142 9380 70194
rect 9212 70140 9380 70142
rect 8988 69636 9044 69646
rect 9212 69636 9268 70140
rect 9324 70130 9380 70140
rect 8988 69634 9268 69636
rect 8988 69582 8990 69634
rect 9042 69582 9268 69634
rect 8988 69580 9268 69582
rect 8988 69570 9044 69580
rect 9436 69524 9492 70364
rect 8876 69234 8932 69244
rect 9324 69468 9492 69524
rect 8652 67106 8708 67116
rect 8988 68402 9044 68414
rect 8988 68350 8990 68402
rect 9042 68350 9044 68402
rect 8988 67060 9044 68350
rect 8988 66994 9044 67004
rect 9324 67620 9380 69468
rect 9436 68404 9492 68414
rect 9436 68310 9492 68348
rect 9548 68180 9604 71148
rect 9772 70756 9828 70766
rect 9772 70662 9828 70700
rect 9884 70194 9940 70206
rect 9884 70142 9886 70194
rect 9938 70142 9940 70194
rect 9772 69972 9828 69982
rect 9772 68626 9828 69916
rect 9772 68574 9774 68626
rect 9826 68574 9828 68626
rect 9772 68562 9828 68574
rect 8540 66834 8596 66846
rect 8540 66782 8542 66834
rect 8594 66782 8596 66834
rect 8540 65492 8596 66782
rect 9324 66164 9380 67564
rect 9212 66162 9380 66164
rect 9212 66110 9326 66162
rect 9378 66110 9380 66162
rect 9212 66108 9380 66110
rect 8540 65426 8596 65436
rect 8876 65604 8932 65614
rect 8428 63746 8484 63756
rect 8764 64036 8820 64046
rect 8316 63310 8318 63362
rect 8370 63310 8372 63362
rect 8316 63298 8372 63310
rect 8764 63364 8820 63980
rect 8876 64036 8932 65548
rect 8988 65380 9044 65390
rect 9212 65380 9268 66108
rect 9324 66098 9380 66108
rect 9436 68124 9604 68180
rect 9324 65492 9380 65502
rect 9324 65398 9380 65436
rect 8988 65378 9268 65380
rect 8988 65326 8990 65378
rect 9042 65326 9268 65378
rect 8988 65324 9268 65326
rect 8988 64818 9044 65324
rect 9436 65268 9492 68124
rect 9548 67732 9604 67742
rect 9548 67730 9716 67732
rect 9548 67678 9550 67730
rect 9602 67678 9716 67730
rect 9548 67676 9716 67678
rect 9548 67666 9604 67676
rect 9548 67060 9604 67070
rect 9548 66276 9604 67004
rect 9660 67058 9716 67676
rect 9660 67006 9662 67058
rect 9714 67006 9716 67058
rect 9660 66836 9716 67006
rect 9660 66770 9716 66780
rect 9884 67060 9940 70142
rect 9996 69972 10052 69982
rect 9996 69878 10052 69916
rect 10108 69634 10164 72156
rect 10108 69582 10110 69634
rect 10162 69582 10164 69634
rect 10108 69570 10164 69582
rect 9996 69524 10052 69534
rect 9996 68964 10052 69468
rect 9996 68066 10052 68908
rect 9996 68014 9998 68066
rect 10050 68014 10052 68066
rect 9996 68002 10052 68014
rect 9660 66276 9716 66286
rect 9548 66274 9716 66276
rect 9548 66222 9662 66274
rect 9714 66222 9716 66274
rect 9548 66220 9716 66222
rect 9660 66210 9716 66220
rect 9884 66276 9940 67004
rect 9996 67172 10052 67182
rect 9996 66946 10052 67116
rect 9996 66894 9998 66946
rect 10050 66894 10052 66946
rect 9996 66882 10052 66894
rect 10108 66276 10164 66286
rect 9884 66274 10164 66276
rect 9884 66222 10110 66274
rect 10162 66222 10164 66274
rect 9884 66220 10164 66222
rect 8988 64766 8990 64818
rect 9042 64766 9044 64818
rect 8988 64754 9044 64766
rect 9100 65212 9492 65268
rect 9884 65490 9940 66220
rect 10108 66210 10164 66220
rect 9884 65438 9886 65490
rect 9938 65438 9940 65490
rect 8876 64034 9044 64036
rect 8876 63982 8878 64034
rect 8930 63982 9044 64034
rect 8876 63980 9044 63982
rect 8876 63970 8932 63980
rect 8876 63364 8932 63374
rect 8764 63362 8932 63364
rect 8764 63310 8878 63362
rect 8930 63310 8932 63362
rect 8764 63308 8932 63310
rect 8876 63298 8932 63308
rect 8652 62354 8708 62366
rect 8652 62302 8654 62354
rect 8706 62302 8708 62354
rect 8092 62132 8260 62188
rect 8204 61570 8260 62132
rect 8204 61518 8206 61570
rect 8258 61518 8260 61570
rect 8204 60788 8260 61518
rect 8652 60788 8708 62302
rect 8988 61796 9044 63980
rect 8988 61730 9044 61740
rect 8204 60786 8708 60788
rect 8204 60734 8654 60786
rect 8706 60734 8708 60786
rect 8204 60732 8708 60734
rect 8652 60722 8708 60732
rect 8764 59780 8820 59790
rect 8316 59218 8372 59230
rect 8316 59166 8318 59218
rect 8370 59166 8372 59218
rect 8316 58772 8372 59166
rect 8764 59106 8820 59724
rect 8764 59054 8766 59106
rect 8818 59054 8820 59106
rect 8764 59042 8820 59054
rect 8092 58716 8316 58772
rect 8092 57762 8148 58716
rect 8316 58706 8372 58716
rect 8092 57710 8094 57762
rect 8146 57710 8148 57762
rect 8092 56868 8148 57710
rect 8540 57764 8596 57774
rect 8540 57538 8596 57708
rect 8540 57486 8542 57538
rect 8594 57486 8596 57538
rect 8540 57474 8596 57486
rect 8092 56802 8148 56812
rect 8988 56980 9044 56990
rect 8204 56642 8260 56654
rect 8204 56590 8206 56642
rect 8258 56590 8260 56642
rect 8092 55300 8148 55310
rect 7644 50530 7700 50540
rect 7756 53116 7924 53172
rect 7980 55298 8148 55300
rect 7980 55246 8094 55298
rect 8146 55246 8148 55298
rect 7980 55244 8148 55246
rect 7980 54516 8036 55244
rect 8092 55234 8148 55244
rect 7756 50428 7812 53116
rect 7980 51378 8036 54460
rect 8204 53844 8260 56590
rect 8988 56194 9044 56924
rect 8988 56142 8990 56194
rect 9042 56142 9044 56194
rect 8988 56130 9044 56142
rect 9100 54964 9156 65212
rect 9212 65044 9268 65054
rect 9212 63362 9268 64988
rect 9324 64708 9380 64718
rect 9324 64614 9380 64652
rect 9884 64706 9940 65438
rect 9996 65266 10052 65278
rect 9996 65214 9998 65266
rect 10050 65214 10052 65266
rect 9996 65044 10052 65214
rect 9996 64978 10052 64988
rect 9996 64820 10052 64830
rect 9996 64726 10052 64764
rect 9884 64654 9886 64706
rect 9938 64654 9940 64706
rect 9884 64642 9940 64654
rect 9548 63924 9604 63934
rect 9324 63812 9380 63822
rect 9324 63718 9380 63756
rect 9212 63310 9214 63362
rect 9266 63310 9268 63362
rect 9212 63298 9268 63310
rect 9548 62354 9604 63868
rect 9548 62302 9550 62354
rect 9602 62302 9604 62354
rect 9548 62290 9604 62302
rect 9884 63812 9940 63822
rect 9884 63476 9940 63756
rect 9212 62130 9268 62142
rect 9212 62078 9214 62130
rect 9266 62078 9268 62130
rect 9212 61460 9268 62078
rect 9212 61394 9268 61404
rect 9436 61796 9492 61806
rect 9436 61570 9492 61740
rect 9436 61518 9438 61570
rect 9490 61518 9492 61570
rect 9436 59892 9492 61518
rect 9548 61124 9604 61134
rect 9548 60002 9604 61068
rect 9548 59950 9550 60002
rect 9602 59950 9604 60002
rect 9548 59938 9604 59950
rect 9884 60114 9940 63420
rect 9996 62580 10052 62590
rect 9996 61908 10052 62524
rect 9996 61794 10052 61852
rect 9996 61742 9998 61794
rect 10050 61742 10052 61794
rect 9996 61730 10052 61742
rect 9884 60062 9886 60114
rect 9938 60062 9940 60114
rect 9884 60004 9940 60062
rect 9884 59938 9940 59948
rect 9436 59220 9492 59836
rect 9436 59154 9492 59164
rect 10108 59892 10164 59902
rect 9884 58996 9940 59006
rect 9436 58994 9940 58996
rect 9436 58942 9886 58994
rect 9938 58942 9940 58994
rect 9436 58940 9940 58942
rect 9324 58772 9380 58782
rect 9324 55298 9380 58716
rect 9436 56082 9492 58940
rect 9884 58930 9940 58940
rect 10108 58772 10164 59836
rect 9660 58716 10108 58772
rect 9660 58434 9716 58716
rect 10108 58706 10164 58716
rect 9660 58382 9662 58434
rect 9714 58382 9716 58434
rect 9660 58370 9716 58382
rect 9996 58546 10052 58558
rect 9996 58494 9998 58546
rect 10050 58494 10052 58546
rect 9996 58212 10052 58494
rect 9996 58146 10052 58156
rect 9660 57426 9716 57438
rect 9660 57374 9662 57426
rect 9714 57374 9716 57426
rect 9436 56030 9438 56082
rect 9490 56030 9492 56082
rect 9436 56018 9492 56030
rect 9548 56980 9604 56990
rect 9324 55246 9326 55298
rect 9378 55246 9380 55298
rect 9324 55234 9380 55246
rect 9100 54908 9492 54964
rect 8764 54516 8820 54526
rect 8764 54422 8820 54460
rect 8204 53778 8260 53788
rect 8092 52948 8148 52958
rect 8092 52854 8148 52892
rect 8428 52946 8484 52958
rect 8428 52894 8430 52946
rect 8482 52894 8484 52946
rect 7980 51326 7982 51378
rect 8034 51326 8036 51378
rect 7756 50372 7924 50428
rect 7532 48626 7588 48636
rect 7756 49028 7812 49038
rect 7196 47572 7252 48300
rect 7196 47506 7252 47516
rect 7644 47236 7700 47246
rect 7196 47234 7700 47236
rect 7196 47182 7646 47234
rect 7698 47182 7700 47234
rect 7196 47180 7700 47182
rect 7196 46674 7252 47180
rect 7644 47170 7700 47180
rect 7196 46622 7198 46674
rect 7250 46622 7252 46674
rect 7196 46610 7252 46622
rect 7532 47012 7588 47022
rect 7532 46674 7588 46956
rect 7756 46788 7812 48972
rect 7868 48244 7924 50372
rect 7868 48178 7924 48188
rect 7756 46732 7924 46788
rect 7532 46622 7534 46674
rect 7586 46622 7588 46674
rect 7532 46610 7588 46622
rect 7756 46564 7812 46574
rect 7756 46470 7812 46508
rect 7084 46396 7364 46452
rect 7084 46004 7140 46014
rect 7084 45910 7140 45948
rect 6972 45388 7140 45444
rect 6860 45276 7028 45332
rect 6860 45108 6916 45118
rect 6860 45014 6916 45052
rect 6972 44436 7028 45276
rect 7084 44996 7140 45388
rect 7084 44994 7252 44996
rect 7084 44942 7086 44994
rect 7138 44942 7252 44994
rect 7084 44940 7252 44942
rect 7084 44930 7140 44940
rect 7084 44436 7140 44446
rect 6972 44380 7084 44436
rect 7084 44342 7140 44380
rect 6636 44270 6638 44322
rect 6690 44270 6692 44322
rect 6636 44258 6692 44270
rect 6524 43708 6692 43764
rect 6636 43652 6692 43708
rect 6860 43652 6916 43662
rect 6636 43650 6916 43652
rect 6636 43598 6862 43650
rect 6914 43598 6916 43650
rect 6636 43596 6916 43598
rect 6860 43586 6916 43596
rect 6860 43092 6916 43102
rect 6412 41234 6468 41244
rect 6524 41970 6580 41982
rect 6524 41918 6526 41970
rect 6578 41918 6580 41970
rect 6524 41186 6580 41918
rect 6524 41134 6526 41186
rect 6578 41134 6580 41186
rect 6300 37650 6356 37660
rect 6412 40180 6468 40190
rect 6188 37324 6356 37380
rect 6188 36596 6244 36606
rect 6076 36482 6132 36494
rect 6076 36430 6078 36482
rect 6130 36430 6132 36482
rect 6076 35476 6132 36430
rect 6076 35410 6132 35420
rect 6188 35700 6244 36540
rect 6188 35140 6244 35644
rect 6188 35074 6244 35084
rect 6076 35028 6132 35038
rect 6076 34934 6132 34972
rect 6188 34916 6244 34926
rect 6188 33572 6244 34860
rect 6300 34242 6356 37324
rect 6412 37154 6468 40124
rect 6524 39842 6580 41134
rect 6524 39790 6526 39842
rect 6578 39790 6580 39842
rect 6524 39778 6580 39790
rect 6860 40514 6916 43036
rect 7196 42980 7252 44940
rect 7308 44884 7364 46396
rect 7532 45220 7588 45230
rect 7532 45106 7588 45164
rect 7532 45054 7534 45106
rect 7586 45054 7588 45106
rect 7532 45042 7588 45054
rect 7308 44828 7588 44884
rect 7084 42924 7196 42980
rect 7084 41188 7140 42924
rect 7196 42914 7252 42924
rect 7196 42756 7252 42766
rect 7196 42532 7252 42700
rect 7196 41970 7252 42476
rect 7196 41918 7198 41970
rect 7250 41918 7252 41970
rect 7196 41906 7252 41918
rect 7308 42530 7364 42542
rect 7308 42478 7310 42530
rect 7362 42478 7364 42530
rect 7308 41860 7364 42478
rect 7308 41794 7364 41804
rect 6860 40462 6862 40514
rect 6914 40462 6916 40514
rect 6860 39620 6916 40462
rect 6412 37102 6414 37154
rect 6466 37102 6468 37154
rect 6412 36484 6468 37102
rect 6412 36418 6468 36428
rect 6524 39172 6580 39182
rect 6412 35588 6468 35598
rect 6524 35588 6580 39116
rect 6860 38724 6916 39564
rect 6860 38658 6916 38668
rect 6972 41186 7140 41188
rect 6972 41134 7086 41186
rect 7138 41134 7140 41186
rect 6972 41132 7140 41134
rect 6860 37828 6916 37838
rect 6860 37266 6916 37772
rect 6860 37214 6862 37266
rect 6914 37214 6916 37266
rect 6412 35586 6580 35588
rect 6412 35534 6414 35586
rect 6466 35534 6580 35586
rect 6412 35532 6580 35534
rect 6636 36708 6692 36718
rect 6412 35522 6468 35532
rect 6636 35476 6692 36652
rect 6524 35420 6692 35476
rect 6748 36482 6804 36494
rect 6748 36430 6750 36482
rect 6802 36430 6804 36482
rect 6524 35026 6580 35420
rect 6748 35140 6804 36430
rect 6860 35698 6916 37214
rect 6860 35646 6862 35698
rect 6914 35646 6916 35698
rect 6860 35634 6916 35646
rect 6524 34974 6526 35026
rect 6578 34974 6580 35026
rect 6524 34962 6580 34974
rect 6636 35084 6804 35140
rect 6636 34916 6692 35084
rect 6636 34850 6692 34860
rect 6972 34580 7028 41132
rect 7084 41122 7140 41132
rect 7308 40178 7364 40190
rect 7308 40126 7310 40178
rect 7362 40126 7364 40178
rect 7308 40068 7364 40126
rect 7308 40002 7364 40012
rect 7084 39730 7140 39742
rect 7084 39678 7086 39730
rect 7138 39678 7140 39730
rect 7084 39172 7140 39678
rect 7084 39106 7140 39116
rect 7196 38612 7252 38622
rect 7196 38610 7364 38612
rect 7196 38558 7198 38610
rect 7250 38558 7364 38610
rect 7196 38556 7364 38558
rect 7196 38546 7252 38556
rect 7196 37828 7252 37838
rect 7196 37734 7252 37772
rect 7196 37266 7252 37278
rect 7196 37214 7198 37266
rect 7250 37214 7252 37266
rect 7196 37044 7252 37214
rect 7308 37156 7364 38556
rect 7308 37090 7364 37100
rect 7420 37604 7476 37614
rect 7420 37154 7476 37548
rect 7532 37380 7588 44828
rect 7756 43538 7812 43550
rect 7756 43486 7758 43538
rect 7810 43486 7812 43538
rect 7756 43316 7812 43486
rect 7756 43250 7812 43260
rect 7756 42196 7812 42206
rect 7532 37314 7588 37324
rect 7644 39730 7700 39742
rect 7644 39678 7646 39730
rect 7698 39678 7700 39730
rect 7420 37102 7422 37154
rect 7474 37102 7476 37154
rect 7420 37090 7476 37102
rect 7196 36978 7252 36988
rect 7532 37044 7588 37054
rect 7308 36596 7364 36606
rect 7308 36502 7364 36540
rect 7532 36482 7588 36988
rect 7532 36430 7534 36482
rect 7586 36430 7588 36482
rect 7532 36418 7588 36430
rect 7196 35924 7252 35934
rect 6300 34190 6302 34242
rect 6354 34190 6356 34242
rect 6300 34178 6356 34190
rect 6748 34524 7028 34580
rect 7084 34914 7140 34926
rect 7084 34862 7086 34914
rect 7138 34862 7140 34914
rect 6636 34018 6692 34030
rect 6636 33966 6638 34018
rect 6690 33966 6692 34018
rect 6300 33572 6356 33582
rect 6188 33570 6356 33572
rect 6188 33518 6302 33570
rect 6354 33518 6356 33570
rect 6188 33516 6356 33518
rect 6300 33506 6356 33516
rect 6636 33124 6692 33966
rect 5964 33068 6692 33124
rect 5852 32956 6020 33012
rect 5516 31612 5796 31668
rect 4464 25900 4728 25910
rect 4520 25844 4568 25900
rect 4624 25844 4672 25900
rect 4464 25834 4728 25844
rect 5068 25900 5348 25956
rect 5404 29316 5460 29326
rect 4508 25732 4564 25742
rect 4284 25676 4452 25732
rect 3724 25566 3726 25618
rect 3778 25566 3780 25618
rect 3724 25554 3780 25566
rect 3612 25218 3668 25228
rect 4284 25506 4340 25518
rect 4284 25454 4286 25506
rect 4338 25454 4340 25506
rect 4284 25172 4340 25454
rect 3804 25116 4068 25126
rect 3612 25060 3668 25070
rect 3860 25060 3908 25116
rect 3964 25060 4012 25116
rect 4284 25106 4340 25116
rect 3804 25050 4068 25060
rect 3612 24836 3668 25004
rect 4396 24948 4452 25676
rect 4508 25508 4564 25676
rect 4956 25620 5012 25630
rect 4508 25442 4564 25452
rect 4844 25506 4900 25518
rect 4844 25454 4846 25506
rect 4898 25454 4900 25506
rect 4284 24892 4452 24948
rect 3612 24780 3780 24836
rect 3612 24612 3668 24622
rect 3388 24332 3556 24388
rect 3388 24164 3444 24174
rect 3388 24050 3444 24108
rect 3388 23998 3390 24050
rect 3442 23998 3444 24050
rect 3388 23986 3444 23998
rect 3388 21700 3444 21710
rect 3276 21644 3388 21700
rect 3388 21634 3444 21644
rect 3500 21588 3556 24332
rect 3612 22596 3668 24556
rect 3724 23940 3780 24780
rect 4060 23940 4116 23950
rect 3724 23938 4116 23940
rect 3724 23886 4062 23938
rect 4114 23886 4116 23938
rect 3724 23884 4116 23886
rect 4060 23828 4116 23884
rect 4060 23762 4116 23772
rect 4172 23940 4228 23950
rect 3804 23548 4068 23558
rect 3860 23492 3908 23548
rect 3964 23492 4012 23548
rect 3804 23482 4068 23492
rect 4060 22708 4116 22718
rect 3724 22596 3780 22606
rect 3612 22594 3780 22596
rect 3612 22542 3726 22594
rect 3778 22542 3780 22594
rect 3612 22540 3780 22542
rect 3724 22530 3780 22540
rect 4060 22260 4116 22652
rect 4060 22194 4116 22204
rect 3804 21980 4068 21990
rect 3860 21924 3908 21980
rect 3964 21924 4012 21980
rect 3804 21914 4068 21924
rect 3500 21532 3892 21588
rect 2828 21308 3332 21364
rect 3052 20804 3108 20814
rect 2604 20750 2606 20802
rect 2658 20750 2660 20802
rect 2604 20692 2660 20750
rect 2604 20626 2660 20636
rect 2940 20802 3108 20804
rect 2940 20750 3054 20802
rect 3106 20750 3108 20802
rect 2940 20748 3108 20750
rect 2492 20076 2884 20132
rect 2604 19906 2660 19918
rect 2604 19854 2606 19906
rect 2658 19854 2660 19906
rect 2268 19404 2548 19460
rect 2044 19170 2100 19180
rect 2380 19234 2436 19246
rect 2380 19182 2382 19234
rect 2434 19182 2436 19234
rect 1820 18844 2324 18900
rect 1708 18732 1876 18788
rect 1596 18386 1652 18396
rect 1708 18450 1764 18462
rect 1708 18398 1710 18450
rect 1762 18398 1764 18450
rect 1484 16706 1540 16716
rect 1708 18116 1764 18398
rect 1148 16380 1428 16436
rect 812 15138 868 15148
rect 1036 15540 1092 15550
rect 924 14644 980 14654
rect 700 13300 756 13310
rect 700 8260 756 13244
rect 812 12180 868 12190
rect 812 10388 868 12124
rect 812 10322 868 10332
rect 812 10164 868 10174
rect 812 8260 868 10108
rect 924 8372 980 14588
rect 1036 8930 1092 15484
rect 1148 10050 1204 16380
rect 1708 16100 1764 18060
rect 1820 17892 1876 18732
rect 2156 18340 2212 18350
rect 2156 18246 2212 18284
rect 1820 17826 1876 17836
rect 2268 17890 2324 18844
rect 2268 17838 2270 17890
rect 2322 17838 2324 17890
rect 2268 17826 2324 17838
rect 2268 17668 2324 17678
rect 2156 17556 2212 17566
rect 2156 16322 2212 17500
rect 2268 16770 2324 17612
rect 2268 16718 2270 16770
rect 2322 16718 2324 16770
rect 2268 16706 2324 16718
rect 2156 16270 2158 16322
rect 2210 16270 2212 16322
rect 2156 16258 2212 16270
rect 1708 16098 1988 16100
rect 1708 16046 1710 16098
rect 1762 16046 1988 16098
rect 1708 16044 1988 16046
rect 1708 16034 1764 16044
rect 1260 15428 1316 15438
rect 1260 15334 1316 15372
rect 1932 15428 1988 16044
rect 1372 15316 1428 15326
rect 1260 14756 1316 14766
rect 1260 13746 1316 14700
rect 1260 13694 1262 13746
rect 1314 13694 1316 13746
rect 1260 13682 1316 13694
rect 1260 11282 1316 11294
rect 1260 11230 1262 11282
rect 1314 11230 1316 11282
rect 1260 10836 1316 11230
rect 1260 10722 1316 10780
rect 1260 10670 1262 10722
rect 1314 10670 1316 10722
rect 1260 10658 1316 10670
rect 1148 9998 1150 10050
rect 1202 9998 1204 10050
rect 1148 9986 1204 9998
rect 1260 10388 1316 10398
rect 1036 8878 1038 8930
rect 1090 8878 1092 8930
rect 1036 8866 1092 8878
rect 1260 8820 1316 10332
rect 1372 9042 1428 15260
rect 1596 15204 1652 15242
rect 1596 15138 1652 15148
rect 1820 14980 1876 14990
rect 1484 14868 1540 14878
rect 1484 10500 1540 14812
rect 1708 14756 1764 14766
rect 1708 14530 1764 14700
rect 1708 14478 1710 14530
rect 1762 14478 1764 14530
rect 1708 12962 1764 14478
rect 1708 12910 1710 12962
rect 1762 12910 1764 12962
rect 1708 12898 1764 12910
rect 1820 12404 1876 14924
rect 1708 12348 1876 12404
rect 1596 11620 1652 11630
rect 1596 11506 1652 11564
rect 1596 11454 1598 11506
rect 1650 11454 1652 11506
rect 1596 11442 1652 11454
rect 1596 10500 1652 10510
rect 1484 10498 1652 10500
rect 1484 10446 1598 10498
rect 1650 10446 1652 10498
rect 1484 10444 1652 10446
rect 1596 10434 1652 10444
rect 1372 8990 1374 9042
rect 1426 8990 1428 9042
rect 1372 8978 1428 8990
rect 1708 8930 1764 12348
rect 1820 12180 1876 12190
rect 1932 12180 1988 15372
rect 1820 12178 1988 12180
rect 1820 12126 1822 12178
rect 1874 12126 1988 12178
rect 1820 12124 1988 12126
rect 2044 14644 2100 14654
rect 1820 11788 1876 12124
rect 2044 11844 2100 14588
rect 2268 14532 2324 14542
rect 2268 13748 2324 14476
rect 2268 13654 2324 13692
rect 2268 12964 2324 12974
rect 2268 12066 2324 12908
rect 2268 12014 2270 12066
rect 2322 12014 2324 12066
rect 2268 12002 2324 12014
rect 2044 11788 2324 11844
rect 1820 11732 1988 11788
rect 1820 11060 1876 11070
rect 1820 10164 1876 11004
rect 1932 10948 1988 11732
rect 1932 10882 1988 10892
rect 2044 11172 2100 11182
rect 1820 10098 1876 10108
rect 1932 10724 1988 10734
rect 1708 8878 1710 8930
rect 1762 8878 1764 8930
rect 1708 8866 1764 8878
rect 1820 9268 1876 9278
rect 1148 8764 1316 8820
rect 1036 8372 1092 8382
rect 924 8370 1092 8372
rect 924 8318 1038 8370
rect 1090 8318 1092 8370
rect 924 8316 1092 8318
rect 1036 8306 1092 8316
rect 812 8204 980 8260
rect 700 8194 756 8204
rect 924 3780 980 8204
rect 1036 8148 1092 8158
rect 1036 5794 1092 8092
rect 1036 5742 1038 5794
rect 1090 5742 1092 5794
rect 1036 5730 1092 5742
rect 1036 5348 1092 5358
rect 1036 5254 1092 5292
rect 1036 4228 1092 4238
rect 1036 4134 1092 4172
rect 1036 3780 1092 3790
rect 924 3778 1092 3780
rect 924 3726 1038 3778
rect 1090 3726 1092 3778
rect 924 3724 1092 3726
rect 1036 3714 1092 3724
rect 1148 3388 1204 8764
rect 1260 8596 1316 8606
rect 1820 8596 1876 9212
rect 1260 5906 1316 8540
rect 1708 8540 1876 8596
rect 1484 8484 1540 8494
rect 1372 8260 1428 8270
rect 1372 8166 1428 8204
rect 1372 6692 1428 6702
rect 1372 6598 1428 6636
rect 1260 5854 1262 5906
rect 1314 5854 1316 5906
rect 1260 5842 1316 5854
rect 1372 5348 1428 5358
rect 1372 5254 1428 5292
rect 1372 4340 1428 4350
rect 1372 4246 1428 4284
rect 1372 3780 1428 3790
rect 1484 3780 1540 8428
rect 1708 7028 1764 8540
rect 1932 8484 1988 10668
rect 2044 9042 2100 11116
rect 2268 11060 2324 11788
rect 2380 11284 2436 19182
rect 2492 16324 2548 19404
rect 2492 16258 2548 16268
rect 2492 13748 2548 13758
rect 2492 12962 2548 13692
rect 2492 12910 2494 12962
rect 2546 12910 2548 12962
rect 2492 12898 2548 12910
rect 2380 11218 2436 11228
rect 2492 12516 2548 12526
rect 2268 11004 2436 11060
rect 2268 10052 2324 10062
rect 2268 9958 2324 9996
rect 2044 8990 2046 9042
rect 2098 8990 2100 9042
rect 2044 8978 2100 8990
rect 1932 8428 2100 8484
rect 1820 8372 1876 8382
rect 1820 8370 1988 8372
rect 1820 8318 1822 8370
rect 1874 8318 1988 8370
rect 1820 8316 1988 8318
rect 1820 8306 1876 8316
rect 1596 6972 1764 7028
rect 1820 7474 1876 7486
rect 1820 7422 1822 7474
rect 1874 7422 1876 7474
rect 1596 6244 1652 6972
rect 1708 6802 1764 6814
rect 1708 6750 1710 6802
rect 1762 6750 1764 6802
rect 1708 6468 1764 6750
rect 1708 6402 1764 6412
rect 1820 6356 1876 7422
rect 1820 6290 1876 6300
rect 1596 6188 1764 6244
rect 1708 5460 1764 6188
rect 1708 5404 1876 5460
rect 1708 5234 1764 5246
rect 1708 5182 1710 5234
rect 1762 5182 1764 5234
rect 1708 5124 1764 5182
rect 1708 5058 1764 5068
rect 1708 4228 1764 4238
rect 1708 4134 1764 4172
rect 1372 3778 1540 3780
rect 1372 3726 1374 3778
rect 1426 3726 1540 3778
rect 1372 3724 1540 3726
rect 1708 3780 1764 3790
rect 1820 3780 1876 5404
rect 1932 4340 1988 8316
rect 2044 6468 2100 8428
rect 2156 8260 2212 8270
rect 2380 8260 2436 11004
rect 2156 8258 2436 8260
rect 2156 8206 2158 8258
rect 2210 8206 2436 8258
rect 2156 8204 2436 8206
rect 2156 8194 2212 8204
rect 2268 7364 2324 7374
rect 2268 7270 2324 7308
rect 2380 6802 2436 6814
rect 2380 6750 2382 6802
rect 2434 6750 2436 6802
rect 2156 6692 2212 6702
rect 2156 6598 2212 6636
rect 2380 6692 2436 6750
rect 2380 6626 2436 6636
rect 2044 6412 2436 6468
rect 2268 6244 2324 6254
rect 2268 5906 2324 6188
rect 2268 5854 2270 5906
rect 2322 5854 2324 5906
rect 2156 5684 2212 5694
rect 2044 5348 2100 5358
rect 2044 5254 2100 5292
rect 1932 4274 1988 4284
rect 2044 4452 2100 4462
rect 2044 4338 2100 4396
rect 2044 4286 2046 4338
rect 2098 4286 2100 4338
rect 2044 4274 2100 4286
rect 1708 3778 1876 3780
rect 1708 3726 1710 3778
rect 1762 3726 1876 3778
rect 1708 3724 1876 3726
rect 2044 3780 2100 3790
rect 1372 3714 1428 3724
rect 1708 3714 1764 3724
rect 2044 3686 2100 3724
rect 1148 3332 1540 3388
rect 1148 2212 1204 2222
rect 588 2210 1204 2212
rect 588 2158 1150 2210
rect 1202 2158 1204 2210
rect 588 2156 1204 2158
rect 1148 2146 1204 2156
rect 1484 2210 1540 3332
rect 1484 2158 1486 2210
rect 1538 2158 1540 2210
rect 1484 2146 1540 2158
rect 1596 3332 1652 3342
rect 924 1876 980 1886
rect 924 756 980 1820
rect 924 690 980 700
rect 1596 308 1652 3276
rect 1708 2770 1764 2782
rect 1708 2718 1710 2770
rect 1762 2718 1764 2770
rect 1708 2212 1764 2718
rect 2156 2658 2212 5628
rect 2268 3556 2324 5854
rect 2380 5346 2436 6412
rect 2380 5294 2382 5346
rect 2434 5294 2436 5346
rect 2380 5282 2436 5294
rect 2492 5124 2548 12460
rect 2604 11732 2660 19854
rect 2716 19796 2772 19806
rect 2716 19236 2772 19740
rect 2716 19142 2772 19180
rect 2716 18340 2772 18350
rect 2716 18116 2772 18284
rect 2716 17666 2772 18060
rect 2716 17614 2718 17666
rect 2770 17614 2772 17666
rect 2716 17602 2772 17614
rect 2716 17220 2772 17230
rect 2716 16994 2772 17164
rect 2716 16942 2718 16994
rect 2770 16942 2772 16994
rect 2716 16930 2772 16942
rect 2716 15540 2772 15550
rect 2716 14530 2772 15484
rect 2828 15538 2884 20076
rect 2940 19572 2996 20748
rect 3052 20738 3108 20748
rect 3164 20692 3220 20702
rect 3164 20018 3220 20636
rect 3164 19966 3166 20018
rect 3218 19966 3220 20018
rect 3164 19954 3220 19966
rect 2940 19516 3108 19572
rect 2828 15486 2830 15538
rect 2882 15486 2884 15538
rect 2828 15474 2884 15486
rect 2940 19346 2996 19358
rect 2940 19294 2942 19346
rect 2994 19294 2996 19346
rect 2716 14478 2718 14530
rect 2770 14478 2772 14530
rect 2716 14466 2772 14478
rect 2940 13860 2996 19294
rect 2828 13804 2996 13860
rect 2828 12852 2884 13804
rect 2940 13636 2996 13646
rect 2940 13542 2996 13580
rect 3052 13188 3108 19516
rect 3276 18450 3332 21308
rect 3388 20018 3444 20030
rect 3388 19966 3390 20018
rect 3442 19966 3444 20018
rect 3388 19236 3444 19966
rect 3500 19796 3556 21532
rect 3724 21364 3780 21374
rect 3612 21362 3780 21364
rect 3612 21310 3726 21362
rect 3778 21310 3780 21362
rect 3612 21308 3780 21310
rect 3612 20244 3668 21308
rect 3724 21298 3780 21308
rect 3724 20914 3780 20926
rect 3724 20862 3726 20914
rect 3778 20862 3780 20914
rect 3724 20580 3780 20862
rect 3836 20802 3892 21532
rect 4060 21364 4116 21374
rect 4060 21270 4116 21308
rect 4172 21028 4228 23884
rect 4284 23378 4340 24892
rect 4464 24332 4728 24342
rect 4520 24276 4568 24332
rect 4624 24276 4672 24332
rect 4464 24266 4728 24276
rect 4284 23326 4286 23378
rect 4338 23326 4340 23378
rect 4284 23314 4340 23326
rect 4396 23828 4452 23838
rect 4396 23044 4452 23772
rect 4396 22978 4452 22988
rect 4464 22764 4728 22774
rect 4520 22708 4568 22764
rect 4624 22708 4672 22764
rect 4464 22698 4728 22708
rect 4284 22596 4340 22606
rect 4844 22596 4900 25454
rect 4956 23940 5012 25564
rect 4956 23846 5012 23884
rect 4284 22594 4900 22596
rect 4284 22542 4286 22594
rect 4338 22542 4900 22594
rect 4284 22540 4900 22542
rect 4956 23380 5012 23390
rect 4284 22530 4340 22540
rect 4844 22148 4900 22158
rect 4464 21196 4728 21206
rect 4520 21140 4568 21196
rect 4624 21140 4672 21196
rect 4464 21130 4728 21140
rect 4172 20962 4228 20972
rect 4396 21028 4452 21038
rect 3836 20750 3838 20802
rect 3890 20750 3892 20802
rect 3836 20738 3892 20750
rect 4284 20802 4340 20814
rect 4284 20750 4286 20802
rect 4338 20750 4340 20802
rect 3724 20524 4228 20580
rect 3804 20412 4068 20422
rect 3860 20356 3908 20412
rect 3964 20356 4012 20412
rect 3804 20346 4068 20356
rect 4172 20244 4228 20524
rect 3612 20178 3668 20188
rect 4060 20188 4228 20244
rect 3500 19730 3556 19740
rect 3388 19170 3444 19180
rect 3500 19234 3556 19246
rect 3500 19182 3502 19234
rect 3554 19182 3556 19234
rect 3276 18398 3278 18450
rect 3330 18398 3332 18450
rect 3276 18386 3332 18398
rect 3276 17892 3332 17902
rect 3164 17332 3220 17342
rect 3164 15204 3220 17276
rect 3276 17220 3332 17836
rect 3276 17154 3332 17164
rect 3388 17444 3444 17454
rect 3276 16996 3332 17006
rect 3276 16770 3332 16940
rect 3276 16718 3278 16770
rect 3330 16718 3332 16770
rect 3276 16706 3332 16718
rect 3276 16324 3332 16334
rect 3276 16230 3332 16268
rect 3388 15316 3444 17388
rect 3500 15540 3556 19182
rect 3948 19236 4004 19246
rect 3948 19142 4004 19180
rect 3612 19124 3668 19134
rect 3612 18676 3668 19068
rect 4060 19012 4116 20188
rect 4172 20020 4228 20030
rect 4172 19926 4228 19964
rect 4060 18946 4116 18956
rect 3804 18844 4068 18854
rect 3860 18788 3908 18844
rect 3964 18788 4012 18844
rect 3804 18778 4068 18788
rect 3612 18620 4004 18676
rect 3948 18338 4004 18620
rect 4172 18452 4228 18462
rect 4172 18358 4228 18396
rect 3948 18286 3950 18338
rect 4002 18286 4004 18338
rect 3948 18274 4004 18286
rect 4284 18004 4340 20750
rect 4396 20244 4452 20972
rect 4732 20690 4788 20702
rect 4732 20638 4734 20690
rect 4786 20638 4788 20690
rect 4732 20580 4788 20638
rect 4732 20514 4788 20524
rect 4396 20178 4452 20188
rect 4464 19628 4728 19638
rect 4520 19572 4568 19628
rect 4624 19572 4672 19628
rect 4464 19562 4728 19572
rect 4172 17948 4340 18004
rect 4464 18060 4728 18070
rect 4520 18004 4568 18060
rect 4624 18004 4672 18060
rect 4464 17994 4728 18004
rect 4844 18004 4900 22092
rect 4956 21140 5012 23324
rect 4956 21074 5012 21084
rect 5068 20690 5124 25900
rect 5292 25732 5348 25742
rect 5180 25620 5236 25630
rect 5180 25526 5236 25564
rect 5180 25172 5236 25182
rect 5180 24834 5236 25116
rect 5180 24782 5182 24834
rect 5234 24782 5236 24834
rect 5180 24770 5236 24782
rect 5180 23828 5236 23838
rect 5180 23266 5236 23772
rect 5180 23214 5182 23266
rect 5234 23214 5236 23266
rect 5180 23202 5236 23214
rect 5068 20638 5070 20690
rect 5122 20638 5124 20690
rect 5068 20580 5124 20638
rect 5068 20514 5124 20524
rect 5180 23044 5236 23054
rect 4956 20244 5012 20254
rect 4956 19234 5012 20188
rect 5068 19908 5124 19918
rect 5180 19908 5236 22988
rect 5292 22484 5348 25676
rect 5404 22708 5460 29260
rect 5516 24610 5572 31612
rect 5740 30212 5796 30222
rect 5740 30118 5796 30156
rect 5628 28308 5684 28318
rect 5628 25732 5684 28252
rect 5628 25666 5684 25676
rect 5740 25620 5796 25630
rect 5628 25508 5684 25518
rect 5628 25284 5684 25452
rect 5740 25508 5796 25564
rect 5740 25506 5908 25508
rect 5740 25454 5742 25506
rect 5794 25454 5908 25506
rect 5740 25452 5908 25454
rect 5740 25442 5796 25452
rect 5852 25284 5908 25452
rect 5628 25228 5796 25284
rect 5516 24558 5518 24610
rect 5570 24558 5572 24610
rect 5516 24546 5572 24558
rect 5628 22932 5684 22942
rect 5628 22838 5684 22876
rect 5404 22652 5684 22708
rect 5404 22484 5460 22494
rect 5292 22482 5460 22484
rect 5292 22430 5406 22482
rect 5458 22430 5460 22482
rect 5292 22428 5460 22430
rect 5404 21700 5460 22428
rect 5404 21634 5460 21644
rect 5516 20802 5572 20814
rect 5516 20750 5518 20802
rect 5570 20750 5572 20802
rect 5404 20020 5460 20030
rect 5404 19926 5460 19964
rect 5068 19906 5236 19908
rect 5068 19854 5070 19906
rect 5122 19854 5236 19906
rect 5068 19852 5236 19854
rect 5068 19684 5124 19852
rect 5068 19618 5124 19628
rect 5516 19572 5572 20750
rect 4956 19182 4958 19234
rect 5010 19182 5012 19234
rect 4956 19170 5012 19182
rect 5404 19516 5572 19572
rect 4956 18228 5012 18238
rect 4956 18134 5012 18172
rect 5292 18226 5348 18238
rect 5292 18174 5294 18226
rect 5346 18174 5348 18226
rect 4844 17948 5012 18004
rect 3612 17780 3668 17790
rect 3612 17108 3668 17724
rect 3948 17556 4004 17566
rect 3948 17462 4004 17500
rect 3804 17276 4068 17286
rect 3860 17220 3908 17276
rect 3964 17220 4012 17276
rect 3804 17210 4068 17220
rect 3612 17052 4004 17108
rect 3948 16770 4004 17052
rect 3948 16718 3950 16770
rect 4002 16718 4004 16770
rect 3948 16706 4004 16718
rect 3612 16658 3668 16670
rect 3612 16606 3614 16658
rect 3666 16606 3668 16658
rect 3612 16212 3668 16606
rect 4172 16324 4228 17948
rect 4284 17780 4340 17790
rect 4284 17686 4340 17724
rect 4284 17220 4340 17230
rect 4284 16882 4340 17164
rect 4284 16830 4286 16882
rect 4338 16830 4340 16882
rect 4284 16818 4340 16830
rect 4844 16884 4900 16894
rect 4464 16492 4728 16502
rect 4520 16436 4568 16492
rect 4624 16436 4672 16492
rect 4464 16426 4728 16436
rect 4620 16324 4676 16334
rect 4844 16324 4900 16828
rect 4172 16268 4452 16324
rect 3612 16146 3668 16156
rect 3948 16212 4004 16222
rect 3948 16210 4228 16212
rect 3948 16158 3950 16210
rect 4002 16158 4228 16210
rect 3948 16156 4228 16158
rect 3948 16146 4004 16156
rect 3804 15708 4068 15718
rect 3860 15652 3908 15708
rect 3964 15652 4012 15708
rect 3804 15642 4068 15652
rect 4172 15652 4228 16156
rect 4284 16100 4340 16110
rect 4284 16006 4340 16044
rect 4172 15596 4340 15652
rect 3500 15484 3780 15540
rect 3612 15316 3668 15326
rect 3388 15314 3668 15316
rect 3388 15262 3614 15314
rect 3666 15262 3668 15314
rect 3388 15260 3668 15262
rect 3612 15250 3668 15260
rect 3276 15204 3332 15214
rect 3164 15202 3332 15204
rect 3164 15150 3278 15202
rect 3330 15150 3332 15202
rect 3164 15148 3332 15150
rect 3724 15148 3780 15484
rect 4172 15428 4228 15438
rect 3276 15138 3332 15148
rect 3612 15092 3780 15148
rect 4060 15316 4116 15326
rect 4060 15202 4116 15260
rect 4060 15150 4062 15202
rect 4114 15150 4116 15202
rect 4060 15138 4116 15150
rect 3276 14530 3332 14542
rect 3276 14478 3278 14530
rect 3330 14478 3332 14530
rect 2828 12786 2884 12796
rect 2940 13132 3108 13188
rect 3164 13860 3220 13870
rect 2604 11676 2884 11732
rect 2828 11618 2884 11676
rect 2828 11566 2830 11618
rect 2882 11566 2884 11618
rect 2828 11554 2884 11566
rect 2828 11284 2884 11294
rect 2716 10836 2772 10846
rect 2716 10276 2772 10780
rect 2828 10834 2884 11228
rect 2828 10782 2830 10834
rect 2882 10782 2884 10834
rect 2828 10770 2884 10782
rect 2940 10612 2996 13132
rect 2492 5058 2548 5068
rect 2604 10164 2660 10174
rect 2604 4228 2660 10108
rect 2716 9714 2772 10220
rect 2716 9662 2718 9714
rect 2770 9662 2772 9714
rect 2716 9044 2772 9662
rect 2716 8950 2772 8988
rect 2828 10556 2996 10612
rect 3052 12962 3108 12974
rect 3052 12910 3054 12962
rect 3106 12910 3108 12962
rect 2828 7700 2884 10556
rect 2828 7634 2884 7644
rect 2940 8708 2996 8718
rect 2716 5684 2772 5694
rect 2716 5590 2772 5628
rect 2716 5348 2772 5358
rect 2716 5254 2772 5292
rect 2716 4676 2772 4686
rect 2716 4338 2772 4620
rect 2716 4286 2718 4338
rect 2770 4286 2772 4338
rect 2716 4274 2772 4286
rect 2604 4162 2660 4172
rect 2716 3780 2772 3790
rect 2940 3780 2996 8652
rect 3052 8372 3108 12910
rect 3164 10500 3220 13804
rect 3276 10948 3332 14478
rect 3500 13748 3556 13758
rect 3500 13654 3556 13692
rect 3388 13524 3444 13534
rect 3388 13430 3444 13468
rect 3612 13188 3668 15092
rect 3724 14644 3780 14654
rect 3724 14550 3780 14588
rect 3836 14532 3892 14542
rect 3836 14438 3892 14476
rect 3804 14140 4068 14150
rect 3860 14084 3908 14140
rect 3964 14084 4012 14140
rect 3804 14074 4068 14084
rect 4060 13860 4116 13870
rect 3388 13132 3668 13188
rect 3948 13748 4004 13758
rect 3388 12402 3444 13132
rect 3724 13076 3780 13086
rect 3388 12350 3390 12402
rect 3442 12350 3444 12402
rect 3388 12338 3444 12350
rect 3612 13074 3780 13076
rect 3612 13022 3726 13074
rect 3778 13022 3780 13074
rect 3612 13020 3780 13022
rect 3500 12180 3556 12190
rect 3388 11620 3444 11630
rect 3500 11620 3556 12124
rect 3388 11618 3556 11620
rect 3388 11566 3390 11618
rect 3442 11566 3556 11618
rect 3388 11564 3556 11566
rect 3388 11554 3444 11564
rect 3276 10882 3332 10892
rect 3500 10836 3556 10846
rect 3500 10610 3556 10780
rect 3612 10724 3668 13020
rect 3724 13010 3780 13020
rect 3948 12962 4004 13692
rect 4060 13746 4116 13804
rect 4060 13694 4062 13746
rect 4114 13694 4116 13746
rect 4060 13682 4116 13694
rect 3948 12910 3950 12962
rect 4002 12910 4004 12962
rect 3948 12898 4004 12910
rect 3804 12572 4068 12582
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 3804 12506 4068 12516
rect 4172 12180 4228 15372
rect 4284 14084 4340 15596
rect 4396 15428 4452 16268
rect 4620 16322 4900 16324
rect 4620 16270 4622 16322
rect 4674 16270 4900 16322
rect 4620 16268 4900 16270
rect 4956 16322 5012 17948
rect 5292 17444 5348 18174
rect 5404 17892 5460 19516
rect 5516 19346 5572 19358
rect 5516 19294 5518 19346
rect 5570 19294 5572 19346
rect 5516 18676 5572 19294
rect 5628 19236 5684 22652
rect 5740 21810 5796 25228
rect 5852 25218 5908 25228
rect 5852 23828 5908 23838
rect 5852 23734 5908 23772
rect 5964 22484 6020 32956
rect 6188 31108 6244 31118
rect 6188 30882 6244 31052
rect 6188 30830 6190 30882
rect 6242 30830 6244 30882
rect 6076 30772 6132 30782
rect 6076 28642 6132 30716
rect 6188 29316 6244 30830
rect 6188 29222 6244 29260
rect 6300 29092 6356 33068
rect 6412 32788 6468 32798
rect 6412 32676 6468 32732
rect 6412 32674 6580 32676
rect 6412 32622 6414 32674
rect 6466 32622 6580 32674
rect 6412 32620 6580 32622
rect 6412 32610 6468 32620
rect 6524 30548 6580 32620
rect 6748 32116 6804 34524
rect 6972 34356 7028 34366
rect 6860 32340 6916 32350
rect 6860 32246 6916 32284
rect 6748 32060 6916 32116
rect 6636 32004 6692 32014
rect 6636 31892 6692 31948
rect 6748 31892 6804 31902
rect 6636 31890 6804 31892
rect 6636 31838 6750 31890
rect 6802 31838 6804 31890
rect 6636 31836 6804 31838
rect 6748 31826 6804 31836
rect 6748 30996 6804 31006
rect 6748 30902 6804 30940
rect 6524 30492 6692 30548
rect 6524 30324 6580 30334
rect 6524 29540 6580 30268
rect 6636 30212 6692 30492
rect 6636 30118 6692 30156
rect 6636 29540 6692 29550
rect 6524 29538 6692 29540
rect 6524 29486 6638 29538
rect 6690 29486 6692 29538
rect 6524 29484 6692 29486
rect 6636 29474 6692 29484
rect 6076 28590 6078 28642
rect 6130 28590 6132 28642
rect 6076 27074 6132 28590
rect 6076 27022 6078 27074
rect 6130 27022 6132 27074
rect 6076 27010 6132 27022
rect 6188 29036 6356 29092
rect 6188 26516 6244 29036
rect 6188 25730 6244 26460
rect 6300 28868 6356 28878
rect 6860 28868 6916 32060
rect 6300 27970 6356 28812
rect 6300 27918 6302 27970
rect 6354 27918 6356 27970
rect 6300 26292 6356 27918
rect 6748 28812 6916 28868
rect 6636 27748 6692 27758
rect 6636 27654 6692 27692
rect 6748 27300 6804 28812
rect 6972 28756 7028 34300
rect 7084 33124 7140 34862
rect 7084 33058 7140 33068
rect 7196 32004 7252 35868
rect 7420 35700 7476 35710
rect 7308 35698 7476 35700
rect 7308 35646 7422 35698
rect 7474 35646 7476 35698
rect 7308 35644 7476 35646
rect 7308 34914 7364 35644
rect 7420 35634 7476 35644
rect 7308 34862 7310 34914
rect 7362 34862 7364 34914
rect 7308 34850 7364 34862
rect 7420 35476 7476 35486
rect 7420 34692 7476 35420
rect 7196 31938 7252 31948
rect 7308 34636 7476 34692
rect 7532 34916 7588 34926
rect 7196 31666 7252 31678
rect 7196 31614 7198 31666
rect 7250 31614 7252 31666
rect 7196 30996 7252 31614
rect 7196 30930 7252 30940
rect 7308 30772 7364 34636
rect 7420 34468 7476 34478
rect 7420 33458 7476 34412
rect 7420 33406 7422 33458
rect 7474 33406 7476 33458
rect 7420 32116 7476 33406
rect 7420 32050 7476 32060
rect 7532 31220 7588 34860
rect 7644 34356 7700 39678
rect 7644 34290 7700 34300
rect 7532 31154 7588 31164
rect 7420 31108 7476 31118
rect 7420 31014 7476 31052
rect 7756 30772 7812 42140
rect 7868 41186 7924 46732
rect 7980 44548 8036 51326
rect 8428 50428 8484 52894
rect 9212 52948 9268 52958
rect 9212 52854 9268 52892
rect 9100 52722 9156 52734
rect 9100 52670 9102 52722
rect 9154 52670 9156 52722
rect 9100 52164 9156 52670
rect 9100 52098 9156 52108
rect 8204 50372 8484 50428
rect 8540 51492 8596 51502
rect 8204 49250 8260 50372
rect 8540 50034 8596 51436
rect 9324 51492 9380 51502
rect 9324 51378 9380 51436
rect 9324 51326 9326 51378
rect 9378 51326 9380 51378
rect 9324 51314 9380 51326
rect 8988 51268 9044 51278
rect 8540 49982 8542 50034
rect 8594 49982 8596 50034
rect 8540 49970 8596 49982
rect 8652 51266 9044 51268
rect 8652 51214 8990 51266
rect 9042 51214 9044 51266
rect 8652 51212 9044 51214
rect 8204 49198 8206 49250
rect 8258 49198 8260 49250
rect 8204 49186 8260 49198
rect 8316 48018 8372 48030
rect 8316 47966 8318 48018
rect 8370 47966 8372 48018
rect 8204 47346 8260 47358
rect 8204 47294 8206 47346
rect 8258 47294 8260 47346
rect 8092 47234 8148 47246
rect 8092 47182 8094 47234
rect 8146 47182 8148 47234
rect 8092 44884 8148 47182
rect 8204 46116 8260 47294
rect 8316 46674 8372 47966
rect 8652 47012 8708 51212
rect 8988 51202 9044 51212
rect 8316 46622 8318 46674
rect 8370 46622 8372 46674
rect 8316 46610 8372 46622
rect 8428 46956 8708 47012
rect 8764 51044 8820 51054
rect 8204 46060 8372 46116
rect 8204 45892 8260 45902
rect 8204 45798 8260 45836
rect 8204 45108 8260 45118
rect 8204 45014 8260 45052
rect 8092 44818 8148 44828
rect 7980 44482 8036 44492
rect 8204 44548 8260 44558
rect 8316 44548 8372 46060
rect 8204 44546 8372 44548
rect 8204 44494 8206 44546
rect 8258 44494 8372 44546
rect 8204 44492 8372 44494
rect 8204 44482 8260 44492
rect 8092 44436 8148 44446
rect 7980 42196 8036 42206
rect 7980 41970 8036 42140
rect 7980 41918 7982 41970
rect 8034 41918 8036 41970
rect 7980 41906 8036 41918
rect 7868 41134 7870 41186
rect 7922 41134 7924 41186
rect 7868 41076 7924 41134
rect 7868 41010 7924 41020
rect 7980 40740 8036 40750
rect 7980 40516 8036 40684
rect 7868 39394 7924 39406
rect 7868 39342 7870 39394
rect 7922 39342 7924 39394
rect 7868 37604 7924 39342
rect 7868 37538 7924 37548
rect 7868 37156 7924 37166
rect 7868 37062 7924 37100
rect 7868 36708 7924 36718
rect 7868 36482 7924 36652
rect 7868 36430 7870 36482
rect 7922 36430 7924 36482
rect 7868 36418 7924 36430
rect 7868 34356 7924 34366
rect 7868 34262 7924 34300
rect 7980 33572 8036 40460
rect 8092 38668 8148 44380
rect 8316 44324 8372 44492
rect 8316 44258 8372 44268
rect 8204 43540 8260 43550
rect 8204 43426 8260 43484
rect 8204 43374 8206 43426
rect 8258 43374 8260 43426
rect 8204 43362 8260 43374
rect 8428 41412 8484 46956
rect 8764 46900 8820 50988
rect 9436 50428 9492 54908
rect 9324 50372 9492 50428
rect 9548 53730 9604 56924
rect 9660 56868 9716 57374
rect 10108 56980 10164 56990
rect 10108 56886 10164 56924
rect 9660 56802 9716 56812
rect 10220 56308 10276 72716
rect 10332 72706 10388 72716
rect 10332 72548 10388 72558
rect 10332 72454 10388 72492
rect 10444 72324 10500 72940
rect 10668 72546 10724 73054
rect 10668 72494 10670 72546
rect 10722 72494 10724 72546
rect 10668 72482 10724 72494
rect 10780 72548 10836 72558
rect 10332 72268 10500 72324
rect 10332 68068 10388 72268
rect 10444 70756 10500 70766
rect 10444 70194 10500 70700
rect 10444 70142 10446 70194
rect 10498 70142 10500 70194
rect 10444 70130 10500 70142
rect 10556 69298 10612 69310
rect 10556 69246 10558 69298
rect 10610 69246 10612 69298
rect 10556 69076 10612 69246
rect 10556 68738 10612 69020
rect 10556 68686 10558 68738
rect 10610 68686 10612 68738
rect 10556 68674 10612 68686
rect 10332 68012 10612 68068
rect 10332 66386 10388 66398
rect 10332 66334 10334 66386
rect 10386 66334 10388 66386
rect 10332 63924 10388 66334
rect 10444 64706 10500 64718
rect 10444 64654 10446 64706
rect 10498 64654 10500 64706
rect 10444 64148 10500 64654
rect 10444 64082 10500 64092
rect 10332 63858 10388 63868
rect 10444 63698 10500 63710
rect 10444 63646 10446 63698
rect 10498 63646 10500 63698
rect 10444 62916 10500 63646
rect 10444 62850 10500 62860
rect 10556 61348 10612 68012
rect 10668 67284 10724 67294
rect 10668 65490 10724 67228
rect 10780 66724 10836 72492
rect 10892 71652 10948 71662
rect 10892 71558 10948 71596
rect 11004 71092 11060 73892
rect 11340 73442 11396 73836
rect 11340 73390 11342 73442
rect 11394 73390 11396 73442
rect 11340 73378 11396 73390
rect 11228 73220 11284 73230
rect 11452 73220 11508 73950
rect 11228 73126 11284 73164
rect 11340 73164 11508 73220
rect 11340 72996 11396 73164
rect 11004 70998 11060 71036
rect 11116 72884 11172 72894
rect 10892 68516 10948 68526
rect 11116 68516 11172 72828
rect 11228 72548 11284 72558
rect 11340 72548 11396 72940
rect 11228 72546 11396 72548
rect 11228 72494 11230 72546
rect 11282 72494 11396 72546
rect 11228 72492 11396 72494
rect 11452 72772 11508 72782
rect 11228 72482 11284 72492
rect 11340 71876 11396 71886
rect 11340 71782 11396 71820
rect 11340 70866 11396 70878
rect 11340 70814 11342 70866
rect 11394 70814 11396 70866
rect 10892 68514 11172 68516
rect 10892 68462 10894 68514
rect 10946 68462 11172 68514
rect 10892 68460 11172 68462
rect 11228 70194 11284 70206
rect 11228 70142 11230 70194
rect 11282 70142 11284 70194
rect 10892 66948 10948 68460
rect 11228 67844 11284 70142
rect 11340 69076 11396 70814
rect 11340 69010 11396 69020
rect 11116 67618 11172 67630
rect 11116 67566 11118 67618
rect 11170 67566 11172 67618
rect 11116 67284 11172 67566
rect 11116 67218 11172 67228
rect 11228 67060 11284 67788
rect 11228 67004 11396 67060
rect 10892 66882 10948 66892
rect 11228 66836 11284 66846
rect 11004 66834 11284 66836
rect 11004 66782 11230 66834
rect 11282 66782 11284 66834
rect 11004 66780 11284 66782
rect 10780 66668 10948 66724
rect 10668 65438 10670 65490
rect 10722 65438 10724 65490
rect 10668 65426 10724 65438
rect 10780 64036 10836 64046
rect 10780 63942 10836 63980
rect 10892 63700 10948 66668
rect 11004 66274 11060 66780
rect 11228 66770 11284 66780
rect 11340 66276 11396 67004
rect 11004 66222 11006 66274
rect 11058 66222 11060 66274
rect 11004 66210 11060 66222
rect 11228 66274 11396 66276
rect 11228 66222 11342 66274
rect 11394 66222 11396 66274
rect 11228 66220 11396 66222
rect 11004 65490 11060 65502
rect 11004 65438 11006 65490
rect 11058 65438 11060 65490
rect 11004 64706 11060 65438
rect 11228 65490 11284 66220
rect 11340 66210 11396 66220
rect 11228 65438 11230 65490
rect 11282 65438 11284 65490
rect 11228 65426 11284 65438
rect 11004 64654 11006 64706
rect 11058 64654 11060 64706
rect 11004 64596 11060 64654
rect 11004 64530 11060 64540
rect 10892 63634 10948 63644
rect 11228 63138 11284 63150
rect 11228 63086 11230 63138
rect 11282 63086 11284 63138
rect 10892 63028 10948 63038
rect 10556 61282 10612 61292
rect 10780 63026 10948 63028
rect 10780 62974 10894 63026
rect 10946 62974 10948 63026
rect 10780 62972 10948 62974
rect 10556 61124 10612 61134
rect 10556 60898 10612 61068
rect 10556 60846 10558 60898
rect 10610 60846 10612 60898
rect 10556 60834 10612 60846
rect 10780 60676 10836 62972
rect 10892 62962 10948 62972
rect 10892 62468 10948 62478
rect 10892 62374 10948 62412
rect 10780 60610 10836 60620
rect 11004 61908 11060 61918
rect 11004 60674 11060 61852
rect 11116 61572 11172 61582
rect 11116 61478 11172 61516
rect 11004 60622 11006 60674
rect 11058 60622 11060 60674
rect 11004 60610 11060 60622
rect 11116 60228 11172 60238
rect 11228 60228 11284 63086
rect 11116 60226 11284 60228
rect 11116 60174 11118 60226
rect 11170 60174 11284 60226
rect 11116 60172 11284 60174
rect 11116 60162 11172 60172
rect 10780 59444 10836 59454
rect 10332 58772 10388 58782
rect 10332 57762 10388 58716
rect 10332 57710 10334 57762
rect 10386 57710 10388 57762
rect 10332 57698 10388 57710
rect 10668 57988 10724 57998
rect 10444 56868 10500 56878
rect 10444 56774 10500 56812
rect 10220 56252 10500 56308
rect 9884 56084 9940 56094
rect 9884 55990 9940 56028
rect 10332 56084 10388 56094
rect 9996 55860 10052 55870
rect 9996 55858 10164 55860
rect 9996 55806 9998 55858
rect 10050 55806 10164 55858
rect 9996 55804 10164 55806
rect 9996 55794 10052 55804
rect 9548 53678 9550 53730
rect 9602 53678 9604 53730
rect 8876 50260 8932 50270
rect 8876 47236 8932 50204
rect 8988 49700 9044 49710
rect 8988 47572 9044 49644
rect 9324 48468 9380 50372
rect 9548 48580 9604 53678
rect 9772 55410 9828 55422
rect 9772 55358 9774 55410
rect 9826 55358 9828 55410
rect 9772 53620 9828 55358
rect 9884 53844 9940 53854
rect 9884 53730 9940 53788
rect 9884 53678 9886 53730
rect 9938 53678 9940 53730
rect 9884 53666 9940 53678
rect 9660 52946 9716 52958
rect 9660 52894 9662 52946
rect 9714 52894 9716 52946
rect 9660 52388 9716 52894
rect 9772 52500 9828 53564
rect 10108 53060 10164 55804
rect 10332 53730 10388 56028
rect 10332 53678 10334 53730
rect 10386 53678 10388 53730
rect 10108 53004 10276 53060
rect 10108 52836 10164 52846
rect 10108 52742 10164 52780
rect 10220 52612 10276 53004
rect 9772 52434 9828 52444
rect 10108 52556 10276 52612
rect 9660 52322 9716 52332
rect 9772 52276 9828 52286
rect 9660 50370 9716 50382
rect 9660 50318 9662 50370
rect 9714 50318 9716 50370
rect 9660 48804 9716 50318
rect 9660 48738 9716 48748
rect 9548 48514 9604 48524
rect 9324 48402 9380 48412
rect 9100 48020 9156 48030
rect 9100 48018 9604 48020
rect 9100 47966 9102 48018
rect 9154 47966 9604 48018
rect 9100 47964 9604 47966
rect 9100 47954 9156 47964
rect 9212 47684 9268 47694
rect 9212 47572 9268 47628
rect 8988 47516 9156 47572
rect 8876 47170 8932 47180
rect 8540 46844 8820 46900
rect 8540 41524 8596 46844
rect 8988 46676 9044 46686
rect 8988 46582 9044 46620
rect 9100 46228 9156 47516
rect 9212 47570 9492 47572
rect 9212 47518 9214 47570
rect 9266 47518 9492 47570
rect 9212 47516 9492 47518
rect 9212 47506 9268 47516
rect 8652 46172 9156 46228
rect 9212 47348 9268 47358
rect 8652 43316 8708 46172
rect 9212 46116 9268 47292
rect 9436 47068 9492 47516
rect 9548 47458 9604 47964
rect 9548 47406 9550 47458
rect 9602 47406 9604 47458
rect 9548 47394 9604 47406
rect 9436 47012 9604 47068
rect 8652 43250 8708 43260
rect 8764 46060 9268 46116
rect 8652 41972 8708 41982
rect 8652 41878 8708 41916
rect 8540 41468 8708 41524
rect 8428 41356 8596 41412
rect 8428 40628 8484 40638
rect 8428 40534 8484 40572
rect 8204 39396 8260 39406
rect 8204 39302 8260 39340
rect 8316 39172 8372 39182
rect 8316 38946 8372 39116
rect 8316 38894 8318 38946
rect 8370 38894 8372 38946
rect 8316 38882 8372 38894
rect 8092 38612 8260 38668
rect 8204 35308 8260 38612
rect 8316 36484 8372 36494
rect 8316 36390 8372 36428
rect 8428 35700 8484 35710
rect 8540 35700 8596 41356
rect 8428 35698 8596 35700
rect 8428 35646 8430 35698
rect 8482 35646 8596 35698
rect 8428 35644 8596 35646
rect 8652 37266 8708 41468
rect 8764 38836 8820 46060
rect 8876 45890 8932 45902
rect 9100 45892 9156 45902
rect 8876 45838 8878 45890
rect 8930 45838 8932 45890
rect 8876 45444 8932 45838
rect 8876 45378 8932 45388
rect 8988 45836 9100 45892
rect 8988 44322 9044 45836
rect 9100 45798 9156 45836
rect 9436 45666 9492 45678
rect 9436 45614 9438 45666
rect 9490 45614 9492 45666
rect 9212 45106 9268 45118
rect 9212 45054 9214 45106
rect 9266 45054 9268 45106
rect 8988 44270 8990 44322
rect 9042 44270 9044 44322
rect 8988 44258 9044 44270
rect 9100 44324 9156 44334
rect 9100 44230 9156 44268
rect 9212 44100 9268 45054
rect 9436 44434 9492 45614
rect 9548 44660 9604 47012
rect 9772 46900 9828 52220
rect 10108 52274 10164 52556
rect 10108 52222 10110 52274
rect 10162 52222 10164 52274
rect 10108 52052 10164 52222
rect 10108 51986 10164 51996
rect 10220 52388 10276 52398
rect 9884 51828 9940 51838
rect 9884 51378 9940 51772
rect 10220 51380 10276 52332
rect 9884 51326 9886 51378
rect 9938 51326 9940 51378
rect 9884 51044 9940 51326
rect 10108 51324 10276 51380
rect 10332 51380 10388 53678
rect 10444 54514 10500 56252
rect 10668 56082 10724 57932
rect 10780 57540 10836 59388
rect 11228 58210 11284 58222
rect 11228 58158 11230 58210
rect 11282 58158 11284 58210
rect 11228 57988 11284 58158
rect 11228 57922 11284 57932
rect 10780 57538 11396 57540
rect 10780 57486 10782 57538
rect 10834 57486 11396 57538
rect 10780 57484 11396 57486
rect 10780 57474 10836 57484
rect 10668 56030 10670 56082
rect 10722 56030 10724 56082
rect 10668 56018 10724 56030
rect 11004 56980 11060 56990
rect 11004 56866 11060 56924
rect 11004 56814 11006 56866
rect 11058 56814 11060 56866
rect 11004 56084 11060 56814
rect 11004 56018 11060 56028
rect 11116 56978 11172 56990
rect 11116 56926 11118 56978
rect 11170 56926 11172 56978
rect 11116 55300 11172 56926
rect 11228 56084 11284 56094
rect 11228 55990 11284 56028
rect 10444 54462 10446 54514
rect 10498 54462 10500 54514
rect 10444 53620 10500 54462
rect 10780 55244 11172 55300
rect 10556 53842 10612 53854
rect 10556 53790 10558 53842
rect 10610 53790 10612 53842
rect 10556 53732 10612 53790
rect 10556 53676 10724 53732
rect 10444 53564 10612 53620
rect 10444 52162 10500 52174
rect 10444 52110 10446 52162
rect 10498 52110 10500 52162
rect 10444 51492 10500 52110
rect 10444 51426 10500 51436
rect 9996 51268 10052 51278
rect 10108 51268 10164 51324
rect 10332 51314 10388 51324
rect 9996 51266 10164 51268
rect 9996 51214 9998 51266
rect 10050 51214 10164 51266
rect 9996 51212 10164 51214
rect 9996 51202 10052 51212
rect 9884 50978 9940 50988
rect 10332 50484 10388 50494
rect 9884 49812 9940 49822
rect 9884 49810 10164 49812
rect 9884 49758 9886 49810
rect 9938 49758 10164 49810
rect 9884 49756 10164 49758
rect 9884 49746 9940 49756
rect 9996 49586 10052 49598
rect 9996 49534 9998 49586
rect 10050 49534 10052 49586
rect 9996 49140 10052 49534
rect 9884 49084 10052 49140
rect 9884 48132 9940 49084
rect 9996 48916 10052 48926
rect 9996 48822 10052 48860
rect 10108 48692 10164 49756
rect 10220 49700 10276 49710
rect 10220 48916 10276 49644
rect 10220 48850 10276 48860
rect 10108 48626 10164 48636
rect 9884 48066 9940 48076
rect 10108 48468 10164 48478
rect 10108 47684 10164 48412
rect 10220 48020 10276 48030
rect 10220 47926 10276 47964
rect 10220 47684 10276 47694
rect 10108 47682 10276 47684
rect 10108 47630 10222 47682
rect 10274 47630 10276 47682
rect 10108 47628 10276 47630
rect 10220 47618 10276 47628
rect 9996 47458 10052 47470
rect 9996 47406 9998 47458
rect 10050 47406 10052 47458
rect 9996 47012 10052 47406
rect 9996 46956 10164 47012
rect 9772 46844 10052 46900
rect 9884 46674 9940 46686
rect 9884 46622 9886 46674
rect 9938 46622 9940 46674
rect 9884 46564 9940 46622
rect 9884 46498 9940 46508
rect 9660 46116 9716 46126
rect 9660 46022 9716 46060
rect 9660 45890 9716 45902
rect 9660 45838 9662 45890
rect 9714 45838 9716 45890
rect 9660 45220 9716 45838
rect 9772 45220 9828 45230
rect 9660 45218 9828 45220
rect 9660 45166 9774 45218
rect 9826 45166 9828 45218
rect 9660 45164 9828 45166
rect 9772 45154 9828 45164
rect 9660 44994 9716 45006
rect 9660 44942 9662 44994
rect 9714 44942 9716 44994
rect 9660 44884 9716 44942
rect 9660 44818 9716 44828
rect 9884 44884 9940 44894
rect 9884 44790 9940 44828
rect 9548 44604 9940 44660
rect 9436 44382 9438 44434
rect 9490 44382 9492 44434
rect 9436 44370 9492 44382
rect 9772 44436 9828 44446
rect 9324 44100 9380 44138
rect 9212 44044 9324 44100
rect 9324 44034 9380 44044
rect 9324 43876 9380 43886
rect 9324 43650 9380 43820
rect 9324 43598 9326 43650
rect 9378 43598 9380 43650
rect 9324 43586 9380 43598
rect 9772 43764 9828 44380
rect 9884 44434 9940 44604
rect 9884 44382 9886 44434
rect 9938 44382 9940 44434
rect 9884 44370 9940 44382
rect 9996 43988 10052 46844
rect 9324 42980 9380 42990
rect 9324 42866 9380 42924
rect 9324 42814 9326 42866
rect 9378 42814 9380 42866
rect 9324 42802 9380 42814
rect 9660 42756 9716 42766
rect 9436 42754 9716 42756
rect 9436 42702 9662 42754
rect 9714 42702 9716 42754
rect 9436 42700 9716 42702
rect 9436 42644 9492 42700
rect 9660 42690 9716 42700
rect 9100 42588 9492 42644
rect 8988 42084 9044 42094
rect 8988 41990 9044 42028
rect 8988 40628 9044 40638
rect 9100 40628 9156 42588
rect 9660 42532 9716 42542
rect 9324 42420 9380 42430
rect 9212 41860 9268 41870
rect 9212 41766 9268 41804
rect 8988 40626 9156 40628
rect 8988 40574 8990 40626
rect 9042 40574 9156 40626
rect 8988 40572 9156 40574
rect 8988 40562 9044 40572
rect 8764 38780 9156 38836
rect 8764 38722 8820 38780
rect 8764 38670 8766 38722
rect 8818 38670 8820 38722
rect 8764 38658 8820 38670
rect 8876 38500 8932 38510
rect 8652 37214 8654 37266
rect 8706 37214 8708 37266
rect 8652 36372 8708 37214
rect 8204 35252 8372 35308
rect 8092 34916 8148 34926
rect 8092 34822 8148 34860
rect 8316 33796 8372 35252
rect 8428 34916 8484 35644
rect 8652 35476 8708 36316
rect 8652 35410 8708 35420
rect 8764 37940 8820 37950
rect 8764 35252 8820 37884
rect 8428 34850 8484 34860
rect 8652 35196 8820 35252
rect 8316 33740 8484 33796
rect 7980 33506 8036 33516
rect 8316 33572 8372 33582
rect 8092 33348 8148 33358
rect 7868 33236 7924 33246
rect 7868 33142 7924 33180
rect 7980 32788 8036 32798
rect 7980 32694 8036 32732
rect 7308 30716 7476 30772
rect 7084 30436 7140 30446
rect 7084 30342 7140 30380
rect 7308 30324 7364 30334
rect 7308 28866 7364 30268
rect 7308 28814 7310 28866
rect 7362 28814 7364 28866
rect 7308 28802 7364 28814
rect 6972 28690 7028 28700
rect 6748 27234 6804 27244
rect 6860 28642 6916 28654
rect 6860 28590 6862 28642
rect 6914 28590 6916 28642
rect 6748 27074 6804 27086
rect 6748 27022 6750 27074
rect 6802 27022 6804 27074
rect 6748 26516 6804 27022
rect 6860 26908 6916 28590
rect 7308 27186 7364 27198
rect 7308 27134 7310 27186
rect 7362 27134 7364 27186
rect 6860 26852 7140 26908
rect 6972 26628 7028 26638
rect 6748 26460 6916 26516
rect 6636 26292 6692 26302
rect 6300 26290 6692 26292
rect 6300 26238 6638 26290
rect 6690 26238 6692 26290
rect 6300 26236 6692 26238
rect 6188 25678 6190 25730
rect 6242 25678 6244 25730
rect 6188 25666 6244 25678
rect 6524 25956 6580 25966
rect 6188 24050 6244 24062
rect 6188 23998 6190 24050
rect 6242 23998 6244 24050
rect 6188 23940 6244 23998
rect 6188 23874 6244 23884
rect 6412 22932 6468 22942
rect 5964 22428 6356 22484
rect 5852 22258 5908 22270
rect 5852 22206 5854 22258
rect 5906 22206 5908 22258
rect 5852 22148 5908 22206
rect 5852 22082 5908 22092
rect 6188 22260 6244 22270
rect 5740 21758 5742 21810
rect 5794 21758 5796 21810
rect 5740 21746 5796 21758
rect 6076 20914 6132 20926
rect 6076 20862 6078 20914
rect 6130 20862 6132 20914
rect 5964 20802 6020 20814
rect 5964 20750 5966 20802
rect 6018 20750 6020 20802
rect 5964 20692 6020 20750
rect 5964 20626 6020 20636
rect 5852 20018 5908 20030
rect 6076 20020 6132 20862
rect 5852 19966 5854 20018
rect 5906 19966 5908 20018
rect 5852 19796 5908 19966
rect 5852 19730 5908 19740
rect 5964 19964 6132 20020
rect 5964 19348 6020 19964
rect 5964 19282 6020 19292
rect 6076 19794 6132 19806
rect 6076 19742 6078 19794
rect 6130 19742 6132 19794
rect 5740 19236 5796 19246
rect 5628 19234 5796 19236
rect 5628 19182 5742 19234
rect 5794 19182 5796 19234
rect 5628 19180 5796 19182
rect 5740 19170 5796 19180
rect 5516 18610 5572 18620
rect 5740 19012 5796 19022
rect 5628 18228 5684 18238
rect 5628 18134 5684 18172
rect 5740 18004 5796 18956
rect 5964 18226 6020 18238
rect 5964 18174 5966 18226
rect 6018 18174 6020 18226
rect 5964 18116 6020 18174
rect 5964 18050 6020 18060
rect 5628 17948 5796 18004
rect 5516 17892 5572 17902
rect 5404 17890 5572 17892
rect 5404 17838 5518 17890
rect 5570 17838 5572 17890
rect 5404 17836 5572 17838
rect 5516 17826 5572 17836
rect 5292 17378 5348 17388
rect 5404 17668 5460 17678
rect 5404 17108 5460 17612
rect 5404 16994 5460 17052
rect 5404 16942 5406 16994
rect 5458 16942 5460 16994
rect 5404 16930 5460 16942
rect 5516 17556 5572 17566
rect 4956 16270 4958 16322
rect 5010 16270 5012 16322
rect 4620 16258 4676 16268
rect 4956 16258 5012 16270
rect 5516 16100 5572 17500
rect 5404 16044 5516 16100
rect 4396 15362 4452 15372
rect 4844 15988 4900 15998
rect 4396 15204 4452 15214
rect 4620 15204 4676 15214
rect 4396 15202 4620 15204
rect 4396 15150 4398 15202
rect 4450 15150 4620 15202
rect 4396 15148 4620 15150
rect 4396 15138 4452 15148
rect 4620 15138 4676 15148
rect 4464 14924 4728 14934
rect 4520 14868 4568 14924
rect 4624 14868 4672 14924
rect 4464 14858 4728 14868
rect 4396 14532 4452 14542
rect 4396 14438 4452 14476
rect 4732 14418 4788 14430
rect 4732 14366 4734 14418
rect 4786 14366 4788 14418
rect 4284 14018 4340 14028
rect 4396 14196 4452 14206
rect 4396 13634 4452 14140
rect 4732 14196 4788 14366
rect 4844 14308 4900 15932
rect 5068 15652 5124 15662
rect 5068 15538 5124 15596
rect 5068 15486 5070 15538
rect 5122 15486 5124 15538
rect 5068 15474 5124 15486
rect 5180 14980 5236 14990
rect 5068 14644 5124 14654
rect 5068 14550 5124 14588
rect 4844 14252 5012 14308
rect 4732 14130 4788 14140
rect 4396 13582 4398 13634
rect 4450 13582 4452 13634
rect 4396 13570 4452 13582
rect 4844 14084 4900 14094
rect 4172 12114 4228 12124
rect 4284 13524 4340 13534
rect 3836 11954 3892 11966
rect 3836 11902 3838 11954
rect 3890 11902 3892 11954
rect 3836 11172 3892 11902
rect 4172 11956 4228 11966
rect 4284 11956 4340 13468
rect 4464 13356 4728 13366
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4464 13290 4728 13300
rect 4396 12962 4452 12974
rect 4396 12910 4398 12962
rect 4450 12910 4452 12962
rect 4396 12516 4452 12910
rect 4732 12850 4788 12862
rect 4732 12798 4734 12850
rect 4786 12798 4788 12850
rect 4732 12628 4788 12798
rect 4732 12562 4788 12572
rect 4396 12450 4452 12460
rect 4172 11954 4340 11956
rect 4172 11902 4174 11954
rect 4226 11902 4340 11954
rect 4172 11900 4340 11902
rect 4172 11890 4228 11900
rect 4464 11788 4728 11798
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4464 11722 4728 11732
rect 4284 11620 4340 11630
rect 3836 11116 4228 11172
rect 3804 11004 4068 11014
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 3804 10938 4068 10948
rect 3612 10658 3668 10668
rect 3500 10558 3502 10610
rect 3554 10558 3556 10610
rect 3500 10546 3556 10558
rect 4172 10610 4228 11116
rect 4172 10558 4174 10610
rect 4226 10558 4228 10610
rect 4172 10546 4228 10558
rect 3164 10434 3220 10444
rect 3948 10500 4004 10510
rect 3948 10406 4004 10444
rect 3276 10386 3332 10398
rect 3276 10334 3278 10386
rect 3330 10334 3332 10386
rect 3164 10052 3220 10062
rect 3164 8930 3220 9996
rect 3164 8878 3166 8930
rect 3218 8878 3220 8930
rect 3164 8866 3220 8878
rect 3276 8596 3332 10334
rect 3804 9436 4068 9446
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 3804 9370 4068 9380
rect 4284 9266 4340 11564
rect 4620 11506 4676 11518
rect 4620 11454 4622 11506
rect 4674 11454 4676 11506
rect 4620 11060 4676 11454
rect 4844 11172 4900 14028
rect 4956 13634 5012 14252
rect 4956 13582 4958 13634
rect 5010 13582 5012 13634
rect 4956 13570 5012 13582
rect 5068 13076 5124 13086
rect 5068 12982 5124 13020
rect 4956 12292 5012 12302
rect 4956 12066 5012 12236
rect 4956 12014 4958 12066
rect 5010 12014 5012 12066
rect 4956 12002 5012 12014
rect 5180 11788 5236 14924
rect 5292 13972 5348 13982
rect 5292 13746 5348 13916
rect 5292 13694 5294 13746
rect 5346 13694 5348 13746
rect 5292 13682 5348 13694
rect 5404 13636 5460 16044
rect 5516 16006 5572 16044
rect 5404 13570 5460 13580
rect 5516 14530 5572 14542
rect 5516 14478 5518 14530
rect 5570 14478 5572 14530
rect 5404 12962 5460 12974
rect 5404 12910 5406 12962
rect 5458 12910 5460 12962
rect 5292 11956 5348 11966
rect 5292 11862 5348 11900
rect 5068 11732 5236 11788
rect 4956 11396 5012 11406
rect 4956 11302 5012 11340
rect 4844 11106 4900 11116
rect 4620 10994 4676 11004
rect 4464 10220 4728 10230
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4464 10154 4728 10164
rect 4732 10052 4788 10062
rect 4732 9938 4788 9996
rect 4732 9886 4734 9938
rect 4786 9886 4788 9938
rect 4284 9214 4286 9266
rect 4338 9214 4340 9266
rect 4284 9202 4340 9214
rect 4396 9714 4452 9726
rect 4396 9662 4398 9714
rect 4450 9662 4452 9714
rect 4396 9156 4452 9662
rect 4732 9492 4788 9886
rect 4732 9426 4788 9436
rect 4844 9716 4900 9726
rect 4396 9090 4452 9100
rect 3276 8530 3332 8540
rect 3948 9044 4004 9054
rect 3052 8316 3332 8372
rect 3052 8146 3108 8158
rect 3052 8094 3054 8146
rect 3106 8094 3108 8146
rect 3052 6802 3108 8094
rect 3276 6916 3332 8316
rect 3500 8260 3556 8270
rect 3500 8166 3556 8204
rect 3948 8258 4004 8988
rect 4284 8932 4340 8942
rect 3948 8206 3950 8258
rect 4002 8206 4004 8258
rect 3948 8194 4004 8206
rect 4060 8370 4116 8382
rect 4060 8318 4062 8370
rect 4114 8318 4116 8370
rect 4060 8036 4116 8318
rect 3612 7980 4116 8036
rect 3388 7700 3444 7710
rect 3388 7606 3444 7644
rect 3276 6860 3556 6916
rect 3052 6750 3054 6802
rect 3106 6750 3108 6802
rect 3052 5684 3108 6750
rect 3388 6692 3444 6702
rect 3388 6598 3444 6636
rect 3052 5618 3108 5628
rect 3388 6020 3444 6030
rect 3388 5122 3444 5964
rect 3388 5070 3390 5122
rect 3442 5070 3444 5122
rect 3164 5012 3220 5022
rect 3164 4226 3220 4956
rect 3164 4174 3166 4226
rect 3218 4174 3220 4226
rect 3164 4162 3220 4174
rect 2716 3778 2996 3780
rect 2716 3726 2718 3778
rect 2770 3726 2996 3778
rect 2716 3724 2996 3726
rect 2716 3714 2772 3724
rect 2268 3490 2324 3500
rect 2380 3666 2436 3678
rect 2380 3614 2382 3666
rect 2434 3614 2436 3666
rect 2156 2606 2158 2658
rect 2210 2606 2212 2658
rect 2156 2594 2212 2606
rect 1708 2146 1764 2156
rect 1820 2548 1876 2558
rect 1820 2210 1876 2492
rect 1820 2158 1822 2210
rect 1874 2158 1876 2210
rect 1820 2146 1876 2158
rect 2156 2098 2212 2110
rect 2156 2046 2158 2098
rect 2210 2046 2212 2098
rect 2156 1988 2212 2046
rect 2380 1988 2436 3614
rect 3164 3556 3220 3566
rect 3164 3388 3220 3500
rect 3388 3554 3444 5070
rect 3388 3502 3390 3554
rect 3442 3502 3444 3554
rect 3388 3490 3444 3502
rect 3164 3332 3332 3388
rect 3276 2660 3332 3332
rect 3388 2996 3444 3006
rect 3388 2902 3444 2940
rect 3388 2660 3444 2670
rect 3276 2604 3388 2660
rect 2492 2324 2548 2334
rect 2492 2210 2548 2268
rect 2492 2158 2494 2210
rect 2546 2158 2548 2210
rect 2492 2146 2548 2158
rect 2716 1988 2772 1998
rect 2380 1986 2772 1988
rect 2380 1934 2718 1986
rect 2770 1934 2772 1986
rect 2380 1932 2772 1934
rect 2156 1922 2212 1932
rect 2716 1922 2772 1932
rect 3388 1986 3444 2604
rect 3388 1934 3390 1986
rect 3442 1934 3444 1986
rect 1820 1764 1876 1774
rect 1820 1314 1876 1708
rect 3388 1764 3444 1934
rect 3388 1698 3444 1708
rect 1820 1262 1822 1314
rect 1874 1262 1876 1314
rect 1820 1250 1876 1262
rect 2268 1428 2324 1438
rect 2268 1090 2324 1372
rect 3388 1428 3444 1438
rect 3500 1428 3556 6860
rect 3388 1426 3556 1428
rect 3388 1374 3390 1426
rect 3442 1374 3556 1426
rect 3388 1372 3556 1374
rect 3612 1428 3668 7980
rect 3804 7868 4068 7878
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 3804 7802 4068 7812
rect 3948 6804 4004 6814
rect 3948 6690 4004 6748
rect 3948 6638 3950 6690
rect 4002 6638 4004 6690
rect 3948 6626 4004 6638
rect 4060 6802 4116 6814
rect 4060 6750 4062 6802
rect 4114 6750 4116 6802
rect 4060 6692 4116 6750
rect 4060 6626 4116 6636
rect 3804 6300 4068 6310
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 3804 6234 4068 6244
rect 3836 5908 3892 5918
rect 3836 5814 3892 5852
rect 4172 5124 4228 5134
rect 3804 4732 4068 4742
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 3804 4666 4068 4676
rect 4172 3554 4228 5068
rect 4284 4562 4340 8876
rect 4464 8652 4728 8662
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4464 8586 4728 8596
rect 4732 8258 4788 8270
rect 4732 8206 4734 8258
rect 4786 8206 4788 8258
rect 4732 7812 4788 8206
rect 4732 7746 4788 7756
rect 4844 7364 4900 9660
rect 5068 9044 5124 11732
rect 5404 11620 5460 12910
rect 5404 11554 5460 11564
rect 5516 10052 5572 14478
rect 5628 11060 5684 17948
rect 5740 17668 5796 17678
rect 5740 16770 5796 17612
rect 5740 16718 5742 16770
rect 5794 16718 5796 16770
rect 5740 12964 5796 16718
rect 5964 16548 6020 16558
rect 5852 16436 5908 16446
rect 5852 14530 5908 16380
rect 5964 16322 6020 16492
rect 5964 16270 5966 16322
rect 6018 16270 6020 16322
rect 5964 16258 6020 16270
rect 6076 15988 6132 19742
rect 6188 19124 6244 22204
rect 6188 19058 6244 19068
rect 6188 18004 6244 18014
rect 6188 17666 6244 17948
rect 6188 17614 6190 17666
rect 6242 17614 6244 17666
rect 6188 17556 6244 17614
rect 6188 17490 6244 17500
rect 5852 14478 5854 14530
rect 5906 14478 5908 14530
rect 5852 14420 5908 14478
rect 5852 14354 5908 14364
rect 5964 15932 6132 15988
rect 5964 13524 6020 15932
rect 6076 15204 6132 15214
rect 6076 14754 6132 15148
rect 6188 15092 6244 15102
rect 6188 14998 6244 15036
rect 6076 14702 6078 14754
rect 6130 14702 6132 14754
rect 6076 14690 6132 14702
rect 6300 13972 6356 22428
rect 5964 13458 6020 13468
rect 6188 13916 6356 13972
rect 6076 13076 6132 13086
rect 5964 13074 6132 13076
rect 5964 13022 6078 13074
rect 6130 13022 6132 13074
rect 5964 13020 6132 13022
rect 5740 12898 5796 12908
rect 5852 12962 5908 12974
rect 5852 12910 5854 12962
rect 5906 12910 5908 12962
rect 5852 12628 5908 12910
rect 5852 12562 5908 12572
rect 5964 11620 6020 13020
rect 6076 13010 6132 13020
rect 6188 12852 6244 13916
rect 6076 12796 6244 12852
rect 6300 13746 6356 13758
rect 6300 13694 6302 13746
rect 6354 13694 6356 13746
rect 6300 13636 6356 13694
rect 6076 11956 6132 12796
rect 6076 11890 6132 11900
rect 6188 12292 6244 12302
rect 5852 11564 6020 11620
rect 6076 11620 6132 11630
rect 5740 11284 5796 11294
rect 5740 11190 5796 11228
rect 5628 11004 5796 11060
rect 5628 10610 5684 10622
rect 5628 10558 5630 10610
rect 5682 10558 5684 10610
rect 5628 10500 5684 10558
rect 5628 10434 5684 10444
rect 5516 9986 5572 9996
rect 5068 8978 5124 8988
rect 5292 9044 5348 9054
rect 5292 8950 5348 8988
rect 4956 8818 5012 8830
rect 5628 8820 5684 8830
rect 4956 8766 4958 8818
rect 5010 8766 5012 8818
rect 4956 8484 5012 8766
rect 4956 8418 5012 8428
rect 5404 8818 5684 8820
rect 5404 8766 5630 8818
rect 5682 8766 5684 8818
rect 5404 8764 5684 8766
rect 4956 8260 5012 8270
rect 4956 7924 5012 8204
rect 4956 7858 5012 7868
rect 5068 8258 5124 8270
rect 5068 8206 5070 8258
rect 5122 8206 5124 8258
rect 4956 7364 5012 7374
rect 4844 7362 5012 7364
rect 4844 7310 4958 7362
rect 5010 7310 5012 7362
rect 4844 7308 5012 7310
rect 4956 7298 5012 7308
rect 4464 7084 4728 7094
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4464 7018 4728 7028
rect 4732 6916 4788 6926
rect 4732 6690 4788 6860
rect 4732 6638 4734 6690
rect 4786 6638 4788 6690
rect 4732 6626 4788 6638
rect 5068 6690 5124 8206
rect 5292 7476 5348 7486
rect 5404 7476 5460 8764
rect 5628 8754 5684 8764
rect 5292 7474 5460 7476
rect 5292 7422 5294 7474
rect 5346 7422 5460 7474
rect 5292 7420 5460 7422
rect 5740 7474 5796 11004
rect 5740 7422 5742 7474
rect 5794 7422 5796 7474
rect 5292 7410 5348 7420
rect 5740 7410 5796 7422
rect 5852 7252 5908 11564
rect 6076 11508 6132 11564
rect 5964 11506 6132 11508
rect 5964 11454 6078 11506
rect 6130 11454 6132 11506
rect 5964 11452 6132 11454
rect 5964 10500 6020 11452
rect 6076 11442 6132 11452
rect 5964 10406 6020 10444
rect 6076 11284 6132 11294
rect 5964 10052 6020 10062
rect 5964 9958 6020 9996
rect 6076 9156 6132 11228
rect 6188 10276 6244 12236
rect 6300 12180 6356 13580
rect 6300 11284 6356 12124
rect 6412 11620 6468 22876
rect 6524 21028 6580 25900
rect 6636 25508 6692 26236
rect 6636 25442 6692 25452
rect 6748 24948 6804 24958
rect 6748 24854 6804 24892
rect 6860 24164 6916 26460
rect 6860 24098 6916 24108
rect 6972 23548 7028 26572
rect 7084 25732 7140 26852
rect 7196 26066 7252 26078
rect 7196 26014 7198 26066
rect 7250 26014 7252 26066
rect 7196 25956 7252 26014
rect 7308 25956 7364 27134
rect 7420 26628 7476 30716
rect 7644 30716 7812 30772
rect 7868 32116 7924 32126
rect 7868 30770 7924 32060
rect 7868 30718 7870 30770
rect 7922 30718 7924 30770
rect 7532 30212 7588 30222
rect 7532 29538 7588 30156
rect 7532 29486 7534 29538
rect 7586 29486 7588 29538
rect 7532 28868 7588 29486
rect 7532 28802 7588 28812
rect 7532 28642 7588 28654
rect 7532 28590 7534 28642
rect 7586 28590 7588 28642
rect 7532 27074 7588 28590
rect 7532 27022 7534 27074
rect 7586 27022 7588 27074
rect 7532 26964 7588 27022
rect 7532 26898 7588 26908
rect 7420 26562 7476 26572
rect 7308 25900 7476 25956
rect 7196 25890 7252 25900
rect 7308 25732 7364 25742
rect 7084 25730 7364 25732
rect 7084 25678 7310 25730
rect 7362 25678 7364 25730
rect 7084 25676 7364 25678
rect 7308 25666 7364 25676
rect 7308 24722 7364 24734
rect 7308 24670 7310 24722
rect 7362 24670 7364 24722
rect 7308 24612 7364 24670
rect 7308 24546 7364 24556
rect 7420 24388 7476 25900
rect 7532 24724 7588 24734
rect 7532 24610 7588 24668
rect 7532 24558 7534 24610
rect 7586 24558 7588 24610
rect 7532 24546 7588 24558
rect 7420 24332 7588 24388
rect 7420 24164 7476 24174
rect 7420 24070 7476 24108
rect 6972 23492 7252 23548
rect 6748 23380 6804 23390
rect 6748 23286 6804 23324
rect 7196 23042 7252 23492
rect 7196 22990 7198 23042
rect 7250 22990 7252 23042
rect 6860 22484 6916 22494
rect 6636 22260 6692 22270
rect 6636 22166 6692 22204
rect 6860 21474 6916 22428
rect 7084 22482 7140 22494
rect 7084 22430 7086 22482
rect 7138 22430 7140 22482
rect 7084 22372 7140 22430
rect 7084 22306 7140 22316
rect 6860 21422 6862 21474
rect 6914 21422 6916 21474
rect 6860 21410 6916 21422
rect 6524 20972 6692 21028
rect 6524 20802 6580 20814
rect 6524 20750 6526 20802
rect 6578 20750 6580 20802
rect 6524 16324 6580 20750
rect 6636 19348 6692 20972
rect 6748 20020 6804 20030
rect 6748 19926 6804 19964
rect 7196 19796 7252 22990
rect 7308 22148 7364 22158
rect 7308 21586 7364 22092
rect 7308 21534 7310 21586
rect 7362 21534 7364 21586
rect 7308 21252 7364 21534
rect 7308 21186 7364 21196
rect 7308 20804 7364 20814
rect 7308 20018 7364 20748
rect 7532 20580 7588 24332
rect 7644 23604 7700 30716
rect 7868 28308 7924 30718
rect 7980 29316 8036 29326
rect 8092 29316 8148 33292
rect 8204 29988 8260 29998
rect 8204 29894 8260 29932
rect 7980 29314 8260 29316
rect 7980 29262 7982 29314
rect 8034 29262 8260 29314
rect 7980 29260 8260 29262
rect 7980 29250 8036 29260
rect 7868 28242 7924 28252
rect 7980 28642 8036 28654
rect 7980 28590 7982 28642
rect 8034 28590 8036 28642
rect 7868 27636 7924 27646
rect 7756 27634 7924 27636
rect 7756 27582 7870 27634
rect 7922 27582 7924 27634
rect 7756 27580 7924 27582
rect 7756 27076 7812 27580
rect 7868 27570 7924 27580
rect 7756 27010 7812 27020
rect 7868 27074 7924 27086
rect 7868 27022 7870 27074
rect 7922 27022 7924 27074
rect 7868 26908 7924 27022
rect 7644 23538 7700 23548
rect 7756 26852 7924 26908
rect 7756 23380 7812 26852
rect 7980 24948 8036 28590
rect 7980 24882 8036 24892
rect 8092 26068 8148 26078
rect 8092 24946 8148 26012
rect 8092 24894 8094 24946
rect 8146 24894 8148 24946
rect 8092 24882 8148 24894
rect 8204 23548 8260 29260
rect 8316 28754 8372 33516
rect 8428 33348 8484 33740
rect 8428 33282 8484 33292
rect 8428 33124 8484 33134
rect 8428 29316 8484 33068
rect 8652 31108 8708 35196
rect 8652 31042 8708 31052
rect 8764 34018 8820 34030
rect 8764 33966 8766 34018
rect 8818 33966 8820 34018
rect 8764 30212 8820 33966
rect 8428 29250 8484 29260
rect 8540 30156 8820 30212
rect 8316 28702 8318 28754
rect 8370 28702 8372 28754
rect 8316 28690 8372 28702
rect 8428 28756 8484 28766
rect 8428 28532 8484 28700
rect 8316 28476 8484 28532
rect 8316 27970 8372 28476
rect 8316 27918 8318 27970
rect 8370 27918 8372 27970
rect 8316 27906 8372 27918
rect 8540 27972 8596 30156
rect 8540 27906 8596 27916
rect 8652 29988 8708 29998
rect 8652 28644 8708 29932
rect 8876 28756 8932 38444
rect 9100 35308 9156 38780
rect 9212 37044 9268 37054
rect 9212 35698 9268 36988
rect 9212 35646 9214 35698
rect 9266 35646 9268 35698
rect 9212 35476 9268 35646
rect 9212 35410 9268 35420
rect 8988 35252 9156 35308
rect 8988 34356 9044 35252
rect 9100 35028 9156 35038
rect 9100 34934 9156 34972
rect 8988 34290 9044 34300
rect 9212 34914 9268 34926
rect 9212 34862 9214 34914
rect 9266 34862 9268 34914
rect 9100 34132 9156 34142
rect 8988 34130 9156 34132
rect 8988 34078 9102 34130
rect 9154 34078 9156 34130
rect 8988 34076 9156 34078
rect 8988 31218 9044 34076
rect 9100 34066 9156 34076
rect 9212 32788 9268 34862
rect 9212 32722 9268 32732
rect 8988 31166 8990 31218
rect 9042 31166 9044 31218
rect 8988 31154 9044 31166
rect 9100 31666 9156 31678
rect 9100 31614 9102 31666
rect 9154 31614 9156 31666
rect 9100 31108 9156 31614
rect 8988 30324 9044 30334
rect 9100 30324 9156 31052
rect 9044 30268 9156 30324
rect 8988 28980 9044 30268
rect 9324 30100 9380 42364
rect 9548 41858 9604 41870
rect 9548 41806 9550 41858
rect 9602 41806 9604 41858
rect 9548 41748 9604 41806
rect 9548 41682 9604 41692
rect 9436 38612 9492 38622
rect 9436 37940 9492 38556
rect 9436 37846 9492 37884
rect 9436 37268 9492 37278
rect 9660 37268 9716 42476
rect 9492 37212 9716 37268
rect 9436 37174 9492 37212
rect 9772 36820 9828 43708
rect 9884 43932 10052 43988
rect 10108 46116 10164 46956
rect 10220 46788 10276 46798
rect 10220 46228 10276 46732
rect 10220 46162 10276 46172
rect 9884 40852 9940 43932
rect 9996 43538 10052 43550
rect 9996 43486 9998 43538
rect 10050 43486 10052 43538
rect 9996 43316 10052 43486
rect 9996 43250 10052 43260
rect 10108 42754 10164 46060
rect 10332 46004 10388 50428
rect 10556 49810 10612 53564
rect 10668 51828 10724 53676
rect 10780 52276 10836 55244
rect 11004 55076 11060 55086
rect 11004 55074 11172 55076
rect 11004 55022 11006 55074
rect 11058 55022 11172 55074
rect 11004 55020 11172 55022
rect 11004 55010 11060 55020
rect 10892 54404 10948 54414
rect 10892 53844 10948 54348
rect 10892 53778 10948 53788
rect 11116 53730 11172 55020
rect 11116 53678 11118 53730
rect 11170 53678 11172 53730
rect 11116 53666 11172 53678
rect 10892 53284 10948 53294
rect 10892 53170 10948 53228
rect 10892 53118 10894 53170
rect 10946 53118 10948 53170
rect 10892 53106 10948 53118
rect 11228 52946 11284 52958
rect 11228 52894 11230 52946
rect 11282 52894 11284 52946
rect 11116 52388 11172 52398
rect 11228 52388 11284 52894
rect 11116 52386 11284 52388
rect 11116 52334 11118 52386
rect 11170 52334 11284 52386
rect 11116 52332 11284 52334
rect 11116 52322 11172 52332
rect 10780 52210 10836 52220
rect 10668 51762 10724 51772
rect 10892 52164 10948 52174
rect 10668 51378 10724 51390
rect 10668 51326 10670 51378
rect 10722 51326 10724 51378
rect 10668 51268 10724 51326
rect 10668 51202 10724 51212
rect 10780 51044 10836 51054
rect 10780 50818 10836 50988
rect 10780 50766 10782 50818
rect 10834 50766 10836 50818
rect 10780 50754 10836 50766
rect 10556 49758 10558 49810
rect 10610 49758 10612 49810
rect 10556 49700 10612 49758
rect 10556 49634 10612 49644
rect 10444 49364 10500 49374
rect 10444 49250 10500 49308
rect 10444 49198 10446 49250
rect 10498 49198 10500 49250
rect 10444 49186 10500 49198
rect 10668 48804 10724 48814
rect 10444 48020 10500 48030
rect 10444 46788 10500 47964
rect 10668 47570 10724 48748
rect 10780 48244 10836 48254
rect 10780 48150 10836 48188
rect 10668 47518 10670 47570
rect 10722 47518 10724 47570
rect 10668 47506 10724 47518
rect 10892 47124 10948 52108
rect 11116 51380 11172 51390
rect 11004 50932 11060 50942
rect 11004 50596 11060 50876
rect 11004 50530 11060 50540
rect 11004 49812 11060 49822
rect 11004 49698 11060 49756
rect 11004 49646 11006 49698
rect 11058 49646 11060 49698
rect 11004 49634 11060 49646
rect 10444 46722 10500 46732
rect 10780 47068 10948 47124
rect 11004 48468 11060 48478
rect 10444 46452 10500 46462
rect 10444 46450 10724 46452
rect 10444 46398 10446 46450
rect 10498 46398 10724 46450
rect 10444 46396 10724 46398
rect 10444 46386 10500 46396
rect 10220 45948 10388 46004
rect 10220 45108 10276 45948
rect 10668 45890 10724 46396
rect 10668 45838 10670 45890
rect 10722 45838 10724 45890
rect 10668 45826 10724 45838
rect 10332 45780 10388 45790
rect 10332 45686 10388 45724
rect 10220 45042 10276 45052
rect 10444 45444 10500 45454
rect 10444 45106 10500 45388
rect 10444 45054 10446 45106
rect 10498 45054 10500 45106
rect 10444 45042 10500 45054
rect 10220 44322 10276 44334
rect 10220 44270 10222 44322
rect 10274 44270 10276 44322
rect 10220 43876 10276 44270
rect 10780 44324 10836 47068
rect 10892 46900 10948 46910
rect 10892 45780 10948 46844
rect 11004 46564 11060 48412
rect 11004 46498 11060 46508
rect 11116 46676 11172 51324
rect 11228 51378 11284 51390
rect 11228 51326 11230 51378
rect 11282 51326 11284 51378
rect 11228 50820 11284 51326
rect 11228 50754 11284 50764
rect 11228 50596 11284 50606
rect 11228 48244 11284 50540
rect 11340 49364 11396 57484
rect 11452 56420 11508 72716
rect 11564 61682 11620 76972
rect 11676 75906 11732 77308
rect 11676 75854 11678 75906
rect 11730 75854 11732 75906
rect 11676 75842 11732 75854
rect 11676 75124 11732 75134
rect 11676 72884 11732 75068
rect 11788 74228 11844 85652
rect 11900 84532 11956 84542
rect 11900 82404 11956 84476
rect 12348 84308 12404 86606
rect 12684 85708 12740 87724
rect 12572 85652 12740 85708
rect 12460 85092 12516 85102
rect 12460 84998 12516 85036
rect 12348 84242 12404 84252
rect 12460 84868 12516 84878
rect 11900 82338 11956 82348
rect 12012 83522 12068 83534
rect 12012 83470 12014 83522
rect 12066 83470 12068 83522
rect 12012 83300 12068 83470
rect 12012 82628 12068 83244
rect 12460 83188 12516 84812
rect 12460 83122 12516 83132
rect 12012 82066 12068 82572
rect 12124 82516 12180 82526
rect 12124 82514 12404 82516
rect 12124 82462 12126 82514
rect 12178 82462 12404 82514
rect 12124 82460 12404 82462
rect 12124 82450 12180 82460
rect 12012 82014 12014 82066
rect 12066 82014 12068 82066
rect 12012 82002 12068 82014
rect 12348 81954 12404 82460
rect 12348 81902 12350 81954
rect 12402 81902 12404 81954
rect 12348 81890 12404 81902
rect 12348 81172 12404 81182
rect 12236 80948 12292 80958
rect 12236 79602 12292 80892
rect 12236 79550 12238 79602
rect 12290 79550 12292 79602
rect 12124 79492 12180 79502
rect 12124 79398 12180 79436
rect 11900 79378 11956 79390
rect 11900 79326 11902 79378
rect 11954 79326 11956 79378
rect 11900 78930 11956 79326
rect 12236 79156 12292 79550
rect 12124 79100 12292 79156
rect 12348 80386 12404 81116
rect 12348 80334 12350 80386
rect 12402 80334 12404 80386
rect 11900 78878 11902 78930
rect 11954 78878 11956 78930
rect 11900 78866 11956 78878
rect 12012 78932 12068 78942
rect 12012 78484 12068 78876
rect 12012 78418 12068 78428
rect 12124 78258 12180 79100
rect 12348 78932 12404 80334
rect 12572 79044 12628 85652
rect 12796 85428 12852 87724
rect 12908 86770 12964 87948
rect 12908 86718 12910 86770
rect 12962 86718 12964 86770
rect 12908 86706 12964 86718
rect 13132 87668 13188 87678
rect 13132 87554 13188 87612
rect 13132 87502 13134 87554
rect 13186 87502 13188 87554
rect 13020 85988 13076 85998
rect 13132 85988 13188 87502
rect 13020 85986 13188 85988
rect 13020 85934 13022 85986
rect 13074 85934 13188 85986
rect 13020 85932 13188 85934
rect 13020 85708 13076 85932
rect 13020 85652 13188 85708
rect 12796 85362 12852 85372
rect 12908 84978 12964 84990
rect 12908 84926 12910 84978
rect 12962 84926 12964 84978
rect 12796 84084 12852 84094
rect 12908 84084 12964 84926
rect 13132 84868 13188 85652
rect 13244 85316 13300 88172
rect 13356 85540 13412 88396
rect 13692 88340 13748 88350
rect 13692 88246 13748 88284
rect 13804 88116 13860 89742
rect 13580 87218 13636 87230
rect 13580 87166 13582 87218
rect 13634 87166 13636 87218
rect 13468 86660 13524 86670
rect 13468 86566 13524 86604
rect 13580 86212 13636 87166
rect 13580 86146 13636 86156
rect 13580 85988 13636 85998
rect 13468 85876 13524 85886
rect 13468 85762 13524 85820
rect 13468 85710 13470 85762
rect 13522 85710 13524 85762
rect 13468 85698 13524 85710
rect 13356 85484 13524 85540
rect 13244 85250 13300 85260
rect 13244 85092 13300 85102
rect 13244 84998 13300 85036
rect 13132 84812 13300 84868
rect 13132 84420 13188 84430
rect 13020 84196 13076 84206
rect 13020 84102 13076 84140
rect 12684 84082 12964 84084
rect 12684 84030 12798 84082
rect 12850 84030 12964 84082
rect 12684 84028 12964 84030
rect 12684 79044 12740 84028
rect 12796 84018 12852 84028
rect 12796 83860 12852 83870
rect 12796 81954 12852 83804
rect 13020 83748 13076 83758
rect 12908 82514 12964 82526
rect 12908 82462 12910 82514
rect 12962 82462 12964 82514
rect 12908 82068 12964 82462
rect 13020 82516 13076 83692
rect 13020 82450 13076 82460
rect 12908 82002 12964 82012
rect 13020 82066 13076 82078
rect 13020 82014 13022 82066
rect 13074 82014 13076 82066
rect 12796 81902 12798 81954
rect 12850 81902 12852 81954
rect 12796 81890 12852 81902
rect 13020 81396 13076 82014
rect 13020 81330 13076 81340
rect 12908 81172 12964 81182
rect 12908 81078 12964 81116
rect 12908 80612 12964 80622
rect 12908 80518 12964 80556
rect 12908 79492 12964 79502
rect 12684 78988 12852 79044
rect 12572 78978 12628 78988
rect 12348 78866 12404 78876
rect 12684 78820 12740 78830
rect 12460 78818 12740 78820
rect 12460 78766 12686 78818
rect 12738 78766 12740 78818
rect 12460 78764 12740 78766
rect 12236 78596 12292 78606
rect 12236 78502 12292 78540
rect 12348 78594 12404 78606
rect 12348 78542 12350 78594
rect 12402 78542 12404 78594
rect 12348 78372 12404 78542
rect 12348 78306 12404 78316
rect 12124 78206 12126 78258
rect 12178 78206 12180 78258
rect 12124 78194 12180 78206
rect 12236 78148 12292 78158
rect 12460 78148 12516 78764
rect 12684 78754 12740 78764
rect 12572 78596 12628 78606
rect 12572 78502 12628 78540
rect 12796 78372 12852 78988
rect 12292 78092 12516 78148
rect 12684 78316 12852 78372
rect 12236 78054 12292 78092
rect 11900 77250 11956 77262
rect 11900 77198 11902 77250
rect 11954 77198 11956 77250
rect 11900 76580 11956 77198
rect 11900 76514 11956 76524
rect 12124 76468 12180 76478
rect 12124 76374 12180 76412
rect 12348 75796 12404 75806
rect 12012 75682 12068 75694
rect 12012 75630 12014 75682
rect 12066 75630 12068 75682
rect 12012 74788 12068 75630
rect 12236 75572 12292 75582
rect 12124 74900 12180 74910
rect 12124 74806 12180 74844
rect 12012 74722 12068 74732
rect 11788 74226 12180 74228
rect 11788 74174 11790 74226
rect 11842 74174 12180 74226
rect 11788 74172 12180 74174
rect 11788 74162 11844 74172
rect 11788 74004 11844 74014
rect 11788 73220 11844 73948
rect 11900 73220 11956 73230
rect 11788 73218 11956 73220
rect 11788 73166 11902 73218
rect 11954 73166 11956 73218
rect 11788 73164 11956 73166
rect 11900 73154 11956 73164
rect 11676 72818 11732 72828
rect 11676 72660 11732 72670
rect 11676 72658 11844 72660
rect 11676 72606 11678 72658
rect 11730 72606 11844 72658
rect 11676 72604 11844 72606
rect 11676 72594 11732 72604
rect 11788 72548 11844 72604
rect 11788 72482 11844 72492
rect 11676 72436 11732 72446
rect 11676 63138 11732 72380
rect 12012 70194 12068 70206
rect 12012 70142 12014 70194
rect 12066 70142 12068 70194
rect 11900 69636 11956 69646
rect 11900 69542 11956 69580
rect 11788 68628 11844 68638
rect 11788 63924 11844 68572
rect 12012 68068 12068 70142
rect 12124 69188 12180 74172
rect 12236 74116 12292 75516
rect 12348 75236 12404 75740
rect 12572 75572 12628 75582
rect 12572 75478 12628 75516
rect 12684 75348 12740 78316
rect 12908 78260 12964 79436
rect 13132 79492 13188 84364
rect 13244 83748 13300 84812
rect 13468 84420 13524 85484
rect 13468 84354 13524 84364
rect 13244 83682 13300 83692
rect 13356 83298 13412 83310
rect 13356 83246 13358 83298
rect 13410 83246 13412 83298
rect 13356 80724 13412 83246
rect 13468 83300 13524 83310
rect 13468 83206 13524 83244
rect 13468 82068 13524 82078
rect 13468 81974 13524 82012
rect 13356 80658 13412 80668
rect 13468 80946 13524 80958
rect 13468 80894 13470 80946
rect 13522 80894 13524 80946
rect 13468 80836 13524 80894
rect 13468 80500 13524 80780
rect 13132 79426 13188 79436
rect 13356 80444 13524 80500
rect 13132 79044 13188 79054
rect 12572 75292 12740 75348
rect 12796 78204 12964 78260
rect 13020 78260 13076 78270
rect 12348 75180 12516 75236
rect 12236 74050 12292 74060
rect 12348 74676 12404 74686
rect 12236 73108 12292 73118
rect 12236 73014 12292 73052
rect 12236 69412 12292 69422
rect 12236 69318 12292 69356
rect 12124 69132 12292 69188
rect 12236 68516 12292 69132
rect 12348 68740 12404 74620
rect 12460 70644 12516 75180
rect 12460 70578 12516 70588
rect 12348 68674 12404 68684
rect 12572 68628 12628 75292
rect 12796 74788 12852 78204
rect 13020 78146 13076 78204
rect 13020 78094 13022 78146
rect 13074 78094 13076 78146
rect 13020 78082 13076 78094
rect 12908 77250 12964 77262
rect 12908 77198 12910 77250
rect 12962 77198 12964 77250
rect 12908 76804 12964 77198
rect 12908 76738 12964 76748
rect 12908 76580 12964 76590
rect 12908 76486 12964 76524
rect 13020 75908 13076 75918
rect 13132 75908 13188 78988
rect 13356 77922 13412 80444
rect 13356 77870 13358 77922
rect 13410 77870 13412 77922
rect 13356 76804 13412 77870
rect 13468 77362 13524 77374
rect 13468 77310 13470 77362
rect 13522 77310 13524 77362
rect 13468 77140 13524 77310
rect 13468 77074 13524 77084
rect 13356 76748 13524 76804
rect 13244 76468 13300 76478
rect 13244 76374 13300 76412
rect 13468 76132 13524 76748
rect 13580 76244 13636 85932
rect 13804 85988 13860 88060
rect 13916 89740 14084 89796
rect 14140 89796 14196 89806
rect 13916 86548 13972 89740
rect 13916 86482 13972 86492
rect 14028 88340 14084 88350
rect 13804 85922 13860 85932
rect 14028 85708 14084 88284
rect 14140 85876 14196 89740
rect 14252 86212 14308 95116
rect 14364 94108 14420 97804
rect 14476 97794 14532 97804
rect 14476 97524 14532 97534
rect 14476 95396 14532 97468
rect 14588 97188 14644 100044
rect 14812 99426 14868 107436
rect 15148 106372 15204 106382
rect 15148 106278 15204 106316
rect 15260 105700 15316 108892
rect 15372 108724 15428 113260
rect 15484 109732 15540 114800
rect 15596 113314 15652 113326
rect 15596 113262 15598 113314
rect 15650 113262 15652 113314
rect 15596 112868 15652 113262
rect 15596 112802 15652 112812
rect 15708 110180 15764 114800
rect 15820 111076 15876 111086
rect 15820 110962 15876 111020
rect 15820 110910 15822 110962
rect 15874 110910 15876 110962
rect 15820 110516 15876 110910
rect 15932 110628 15988 114800
rect 16156 112644 16212 114800
rect 16380 113316 16436 114800
rect 16380 113250 16436 113260
rect 16380 113092 16436 113102
rect 16380 112998 16436 113036
rect 16604 112644 16660 114800
rect 16156 112578 16212 112588
rect 16268 112588 16660 112644
rect 16716 112756 16772 112766
rect 16716 112642 16772 112700
rect 16716 112590 16718 112642
rect 16770 112590 16772 112642
rect 16268 112420 16324 112588
rect 16716 112578 16772 112590
rect 16156 112364 16324 112420
rect 16380 112418 16436 112430
rect 16380 112366 16382 112418
rect 16434 112366 16436 112418
rect 15932 110562 15988 110572
rect 16044 111522 16100 111534
rect 16044 111470 16046 111522
rect 16098 111470 16100 111522
rect 15820 110450 15876 110460
rect 15708 110114 15764 110124
rect 15932 110178 15988 110190
rect 15932 110126 15934 110178
rect 15986 110126 15988 110178
rect 15932 110068 15988 110126
rect 15932 110002 15988 110012
rect 15484 109666 15540 109676
rect 15932 109396 15988 109406
rect 16044 109396 16100 111470
rect 15932 109394 16100 109396
rect 15932 109342 15934 109394
rect 15986 109342 16100 109394
rect 15932 109340 16100 109342
rect 15932 109330 15988 109340
rect 15372 108658 15428 108668
rect 15484 109282 15540 109294
rect 15484 109230 15486 109282
rect 15538 109230 15540 109282
rect 15372 108500 15428 108510
rect 15484 108500 15540 109230
rect 16156 109228 16212 112364
rect 16380 111412 16436 112366
rect 16828 112308 16884 114800
rect 16940 113428 16996 113438
rect 16940 112420 16996 113372
rect 17052 112644 17108 114800
rect 17276 113204 17332 114800
rect 17500 113428 17556 114800
rect 17500 113362 17556 113372
rect 17612 113426 17668 113438
rect 17612 113374 17614 113426
rect 17666 113374 17668 113426
rect 17276 113148 17556 113204
rect 17052 112578 17108 112588
rect 16940 112364 17108 112420
rect 16828 112252 16996 112308
rect 16828 111524 16884 111534
rect 16828 111430 16884 111468
rect 16268 110738 16324 110750
rect 16268 110686 16270 110738
rect 16322 110686 16324 110738
rect 16268 110628 16324 110686
rect 16268 109844 16324 110572
rect 16268 109778 16324 109788
rect 16380 109620 16436 111356
rect 15428 108444 15540 108500
rect 15596 109172 16212 109228
rect 16268 109564 16436 109620
rect 16828 109954 16884 109966
rect 16828 109902 16830 109954
rect 16882 109902 16884 109954
rect 16268 109228 16324 109564
rect 16380 109396 16436 109406
rect 16380 109302 16436 109340
rect 16268 109172 16436 109228
rect 15372 108406 15428 108444
rect 15596 107826 15652 109172
rect 16156 108724 16212 108734
rect 16156 108630 16212 108668
rect 15820 108610 15876 108622
rect 15820 108558 15822 108610
rect 15874 108558 15876 108610
rect 15596 107774 15598 107826
rect 15650 107774 15652 107826
rect 15596 107762 15652 107774
rect 15708 108052 15764 108062
rect 15708 107714 15764 107996
rect 15708 107662 15710 107714
rect 15762 107662 15764 107714
rect 15708 107650 15764 107662
rect 15260 105644 15540 105700
rect 14924 105588 14980 105598
rect 14924 105494 14980 105532
rect 15036 104690 15092 104702
rect 15036 104638 15038 104690
rect 15090 104638 15092 104690
rect 15036 102508 15092 104638
rect 15260 104020 15316 104030
rect 15260 103926 15316 103964
rect 15372 103684 15428 103694
rect 15372 103590 15428 103628
rect 15260 102898 15316 102910
rect 15260 102846 15262 102898
rect 15314 102846 15316 102898
rect 15036 102452 15204 102508
rect 15148 102338 15204 102452
rect 15148 102286 15150 102338
rect 15202 102286 15204 102338
rect 14924 101556 14980 101566
rect 15148 101556 15204 102286
rect 15260 102340 15316 102846
rect 15484 102452 15540 105644
rect 15820 105028 15876 108558
rect 16156 107714 16212 107726
rect 16156 107662 16158 107714
rect 16210 107662 16212 107714
rect 15820 104962 15876 104972
rect 15932 107604 15988 107614
rect 15820 104690 15876 104702
rect 15820 104638 15822 104690
rect 15874 104638 15876 104690
rect 15596 103908 15652 103918
rect 15596 103814 15652 103852
rect 15820 103906 15876 104638
rect 15820 103854 15822 103906
rect 15874 103854 15876 103906
rect 15260 102274 15316 102284
rect 15372 102396 15540 102452
rect 15260 101556 15316 101566
rect 15148 101554 15316 101556
rect 15148 101502 15262 101554
rect 15314 101502 15316 101554
rect 15148 101500 15316 101502
rect 14924 101462 14980 101500
rect 15260 101444 15316 101500
rect 15260 101378 15316 101388
rect 14812 99374 14814 99426
rect 14866 99374 14868 99426
rect 14700 98194 14756 98206
rect 14700 98142 14702 98194
rect 14754 98142 14756 98194
rect 14700 97524 14756 98142
rect 14812 98084 14868 99374
rect 14812 98018 14868 98028
rect 14924 101108 14980 101118
rect 14924 97858 14980 101052
rect 14924 97806 14926 97858
rect 14978 97806 14980 97858
rect 14924 97794 14980 97806
rect 15148 98306 15204 98318
rect 15148 98254 15150 98306
rect 15202 98254 15204 98306
rect 14700 97468 15092 97524
rect 14588 97122 14644 97132
rect 14924 97188 14980 97198
rect 14700 97076 14756 97086
rect 14700 96962 14756 97020
rect 14700 96910 14702 96962
rect 14754 96910 14756 96962
rect 14700 96898 14756 96910
rect 14476 95394 14756 95396
rect 14476 95342 14478 95394
rect 14530 95342 14756 95394
rect 14476 95340 14756 95342
rect 14476 95330 14532 95340
rect 14700 95060 14756 95340
rect 14588 95004 14756 95060
rect 14364 94052 14532 94108
rect 14476 93380 14532 94052
rect 14476 93314 14532 93324
rect 14476 92932 14532 92942
rect 14476 92838 14532 92876
rect 14364 91364 14420 91374
rect 14364 91270 14420 91308
rect 14476 91252 14532 91262
rect 14364 90132 14420 90142
rect 14364 89906 14420 90076
rect 14364 89854 14366 89906
rect 14418 89854 14420 89906
rect 14364 89842 14420 89854
rect 14476 89012 14532 91196
rect 14588 90356 14644 95004
rect 14812 94948 14868 94958
rect 14812 94610 14868 94892
rect 14812 94558 14814 94610
rect 14866 94558 14868 94610
rect 14812 94546 14868 94558
rect 14700 94500 14756 94510
rect 14700 94406 14756 94444
rect 14812 93044 14868 93054
rect 14812 92950 14868 92988
rect 14588 90290 14644 90300
rect 14700 92708 14756 92718
rect 14588 89794 14644 89806
rect 14588 89742 14590 89794
rect 14642 89742 14644 89794
rect 14588 89234 14644 89742
rect 14588 89182 14590 89234
rect 14642 89182 14644 89234
rect 14588 89170 14644 89182
rect 14476 88946 14532 88956
rect 14700 88340 14756 92652
rect 14812 91588 14868 91598
rect 14924 91588 14980 97132
rect 15036 96850 15092 97468
rect 15148 97468 15204 98254
rect 15148 97412 15316 97468
rect 15036 96798 15038 96850
rect 15090 96798 15092 96850
rect 15036 96786 15092 96798
rect 15036 96404 15092 96414
rect 15036 93044 15092 96348
rect 15260 95956 15316 97412
rect 15372 96180 15428 102396
rect 15820 102340 15876 103854
rect 15932 103796 15988 107548
rect 16044 105700 16100 105710
rect 16156 105700 16212 107662
rect 16044 105698 16212 105700
rect 16044 105646 16046 105698
rect 16098 105646 16212 105698
rect 16044 105644 16212 105646
rect 16268 106034 16324 106046
rect 16268 105982 16270 106034
rect 16322 105982 16324 106034
rect 16044 105634 16100 105644
rect 16268 104468 16324 105982
rect 16268 104402 16324 104412
rect 15932 103730 15988 103740
rect 16044 102340 16100 102350
rect 15820 102338 16100 102340
rect 15820 102286 16046 102338
rect 16098 102286 16100 102338
rect 15820 102284 16100 102286
rect 15484 101556 15540 101566
rect 16044 101556 16100 102284
rect 16268 101556 16324 101566
rect 16044 101554 16324 101556
rect 16044 101502 16270 101554
rect 16322 101502 16324 101554
rect 16044 101500 16324 101502
rect 15484 100770 15540 101500
rect 15484 100718 15486 100770
rect 15538 100718 15540 100770
rect 15484 100706 15540 100718
rect 15932 98980 15988 98990
rect 15596 98978 15988 98980
rect 15596 98926 15934 98978
rect 15986 98926 15988 98978
rect 15596 98924 15988 98926
rect 15484 98532 15540 98542
rect 15484 96850 15540 98476
rect 15596 98418 15652 98924
rect 15932 98914 15988 98924
rect 15596 98366 15598 98418
rect 15650 98366 15652 98418
rect 15596 98354 15652 98366
rect 15708 98756 15764 98766
rect 16268 98756 16324 101500
rect 15708 97468 15764 98700
rect 15484 96798 15486 96850
rect 15538 96798 15540 96850
rect 15484 96786 15540 96798
rect 15596 97412 15764 97468
rect 15932 98700 16324 98756
rect 15932 97524 15988 98700
rect 16044 98532 16100 98542
rect 16044 98418 16100 98476
rect 16044 98366 16046 98418
rect 16098 98366 16100 98418
rect 16044 98354 16100 98366
rect 16156 98308 16212 98318
rect 16156 98214 16212 98252
rect 16380 97972 16436 109172
rect 16380 97906 16436 97916
rect 16492 109170 16548 109182
rect 16492 109118 16494 109170
rect 16546 109118 16548 109170
rect 15932 97458 15988 97468
rect 16380 97524 16436 97534
rect 15372 96114 15428 96124
rect 15484 96404 15540 96414
rect 15260 95890 15316 95900
rect 15484 94500 15540 96348
rect 15372 94444 15540 94500
rect 15148 93716 15204 93726
rect 15148 93622 15204 93660
rect 15036 92596 15092 92988
rect 15036 92530 15092 92540
rect 15148 91924 15204 91934
rect 15148 91830 15204 91868
rect 14924 91532 15092 91588
rect 14812 91364 14868 91532
rect 14924 91364 14980 91374
rect 14812 91362 14980 91364
rect 14812 91310 14926 91362
rect 14978 91310 14980 91362
rect 14812 91308 14980 91310
rect 14812 88452 14868 91308
rect 14924 91298 14980 91308
rect 15036 90020 15092 91532
rect 15260 91364 15316 91374
rect 15260 90802 15316 91308
rect 15260 90750 15262 90802
rect 15314 90750 15316 90802
rect 15260 90738 15316 90750
rect 14812 88386 14868 88396
rect 14924 89964 15092 90020
rect 15148 90356 15204 90366
rect 14588 88284 14756 88340
rect 14252 86146 14308 86156
rect 14364 87108 14420 87118
rect 14140 85810 14196 85820
rect 14252 85988 14308 85998
rect 13804 85652 13860 85662
rect 14028 85652 14196 85708
rect 13804 85090 13860 85596
rect 14028 85540 14084 85550
rect 13804 85038 13806 85090
rect 13858 85038 13860 85090
rect 13804 85026 13860 85038
rect 13916 85202 13972 85214
rect 13916 85150 13918 85202
rect 13970 85150 13972 85202
rect 13916 84308 13972 85150
rect 13916 84084 13972 84252
rect 13916 84018 13972 84028
rect 14028 83748 14084 85484
rect 13804 83692 14084 83748
rect 13692 83298 13748 83310
rect 13692 83246 13694 83298
rect 13746 83246 13748 83298
rect 13692 81172 13748 83246
rect 13692 81106 13748 81116
rect 13804 79492 13860 83692
rect 14140 83636 14196 85652
rect 14028 83580 14196 83636
rect 13916 83522 13972 83534
rect 13916 83470 13918 83522
rect 13970 83470 13972 83522
rect 13916 81396 13972 83470
rect 14028 82740 14084 83580
rect 14028 82674 14084 82684
rect 14140 82628 14196 82638
rect 14252 82628 14308 85932
rect 14364 85764 14420 87052
rect 14588 86660 14644 88284
rect 14924 88228 14980 89964
rect 15036 89796 15092 89806
rect 15036 89702 15092 89740
rect 15148 89572 15204 90300
rect 14812 88002 14868 88014
rect 14812 87950 14814 88002
rect 14866 87950 14868 88002
rect 14700 87444 14756 87454
rect 14700 87350 14756 87388
rect 14364 85698 14420 85708
rect 14476 86658 14644 86660
rect 14476 86606 14590 86658
rect 14642 86606 14644 86658
rect 14476 86604 14644 86606
rect 14476 83636 14532 86604
rect 14588 86594 14644 86604
rect 14700 86548 14756 86558
rect 14700 85988 14756 86492
rect 14700 85922 14756 85932
rect 14588 85764 14644 85802
rect 14588 85698 14644 85708
rect 14588 85092 14644 85102
rect 14812 85092 14868 87950
rect 14924 87332 14980 88172
rect 15036 89516 15204 89572
rect 15036 87668 15092 89516
rect 15036 87602 15092 87612
rect 15372 87556 15428 94444
rect 15484 94274 15540 94286
rect 15484 94222 15486 94274
rect 15538 94222 15540 94274
rect 15484 93604 15540 94222
rect 15596 93828 15652 97412
rect 16044 97410 16100 97422
rect 16044 97358 16046 97410
rect 16098 97358 16100 97410
rect 16044 96852 16100 97358
rect 16156 96852 16212 96862
rect 16044 96850 16212 96852
rect 16044 96798 16158 96850
rect 16210 96798 16212 96850
rect 16044 96796 16212 96798
rect 16156 96786 16212 96796
rect 15708 96628 15764 96638
rect 15708 96534 15764 96572
rect 15932 96292 15988 96302
rect 15708 95956 15764 95966
rect 15708 94164 15764 95900
rect 15820 94388 15876 94398
rect 15820 94294 15876 94332
rect 15708 94108 15876 94164
rect 15596 93772 15764 93828
rect 15484 93538 15540 93548
rect 15596 93602 15652 93614
rect 15596 93550 15598 93602
rect 15650 93550 15652 93602
rect 15484 93380 15540 93390
rect 15484 90692 15540 93324
rect 15596 92260 15652 93550
rect 15596 92166 15652 92204
rect 15708 91588 15764 93772
rect 15484 90626 15540 90636
rect 15596 91532 15764 91588
rect 15372 87490 15428 87500
rect 14924 87266 14980 87276
rect 15484 87444 15540 87454
rect 15148 85988 15204 85998
rect 15148 85894 15204 85932
rect 15484 85874 15540 87388
rect 15484 85822 15486 85874
rect 15538 85822 15540 85874
rect 15484 85810 15540 85822
rect 15372 85764 15428 85774
rect 14588 85090 14868 85092
rect 14588 85038 14590 85090
rect 14642 85038 14868 85090
rect 14588 85036 14868 85038
rect 14924 85092 14980 85102
rect 14588 85026 14644 85036
rect 14924 84196 14980 85036
rect 15148 84980 15204 84990
rect 15036 84420 15092 84430
rect 15036 84326 15092 84364
rect 14924 84130 14980 84140
rect 15036 83972 15092 83982
rect 14140 82626 14308 82628
rect 14140 82574 14142 82626
rect 14194 82574 14308 82626
rect 14140 82572 14308 82574
rect 14364 83580 14532 83636
rect 14924 83634 14980 83646
rect 14924 83582 14926 83634
rect 14978 83582 14980 83634
rect 14140 82562 14196 82572
rect 14364 82348 14420 83580
rect 14476 83412 14532 83422
rect 14476 83318 14532 83356
rect 14812 83412 14868 83422
rect 14588 83188 14644 83198
rect 14476 82964 14532 82974
rect 14476 82738 14532 82908
rect 14476 82686 14478 82738
rect 14530 82686 14532 82738
rect 14476 82516 14532 82686
rect 14476 82450 14532 82460
rect 14028 82292 14084 82302
rect 14028 81732 14084 82236
rect 14028 81666 14084 81676
rect 14140 82292 14420 82348
rect 13916 80612 13972 81340
rect 14028 80612 14084 80622
rect 13916 80610 14084 80612
rect 13916 80558 14030 80610
rect 14082 80558 14084 80610
rect 13916 80556 14084 80558
rect 14028 80546 14084 80556
rect 14028 79492 14084 79502
rect 13804 79490 14084 79492
rect 13804 79438 14030 79490
rect 14082 79438 14084 79490
rect 13804 79436 14084 79438
rect 13692 78148 13748 78158
rect 13692 76466 13748 78092
rect 13692 76414 13694 76466
rect 13746 76414 13748 76466
rect 13692 76402 13748 76414
rect 13804 77250 13860 77262
rect 13804 77198 13806 77250
rect 13858 77198 13860 77250
rect 13804 76356 13860 77198
rect 13916 76356 13972 76366
rect 13804 76354 13972 76356
rect 13804 76302 13918 76354
rect 13970 76302 13972 76354
rect 13804 76300 13972 76302
rect 13916 76290 13972 76300
rect 13580 76188 13748 76244
rect 13020 75906 13188 75908
rect 13020 75854 13022 75906
rect 13074 75854 13188 75906
rect 13020 75852 13188 75854
rect 13356 76076 13524 76132
rect 12796 74786 12964 74788
rect 12796 74734 12798 74786
rect 12850 74734 12964 74786
rect 12796 74732 12964 74734
rect 12796 74722 12852 74732
rect 12796 73444 12852 73454
rect 12796 73350 12852 73388
rect 12796 72772 12852 72782
rect 12796 72678 12852 72716
rect 12908 68964 12964 74732
rect 13020 74676 13076 75852
rect 13132 74900 13188 74910
rect 13132 74806 13188 74844
rect 13020 74610 13076 74620
rect 13020 73892 13076 73902
rect 13020 73890 13188 73892
rect 13020 73838 13022 73890
rect 13074 73838 13188 73890
rect 13020 73836 13188 73838
rect 13020 73826 13076 73836
rect 13132 73330 13188 73836
rect 13132 73278 13134 73330
rect 13186 73278 13188 73330
rect 13132 73266 13188 73278
rect 13244 73332 13300 73342
rect 12796 68908 12964 68964
rect 13020 70644 13076 70654
rect 12796 68628 12852 68908
rect 12572 68572 12740 68628
rect 12236 68460 12628 68516
rect 12124 68404 12180 68414
rect 12124 68402 12516 68404
rect 12124 68350 12126 68402
rect 12178 68350 12516 68402
rect 12124 68348 12516 68350
rect 12124 68338 12180 68348
rect 12012 68002 12068 68012
rect 12348 68068 12404 68078
rect 12124 67956 12180 67966
rect 12124 67862 12180 67900
rect 12348 66276 12404 68012
rect 12460 67842 12516 68348
rect 12460 67790 12462 67842
rect 12514 67790 12516 67842
rect 12460 67778 12516 67790
rect 12124 66274 12404 66276
rect 12124 66222 12350 66274
rect 12402 66222 12404 66274
rect 12124 66220 12404 66222
rect 12124 65490 12180 66220
rect 12348 66210 12404 66220
rect 12124 65438 12126 65490
rect 12178 65438 12180 65490
rect 12124 64706 12180 65438
rect 12124 64654 12126 64706
rect 12178 64654 12180 64706
rect 12124 64642 12180 64654
rect 11788 63858 11844 63868
rect 11900 63364 11956 63374
rect 11900 63270 11956 63308
rect 12348 63140 12404 63150
rect 11676 63086 11678 63138
rect 11730 63086 11732 63138
rect 11676 62468 11732 63086
rect 12236 63138 12404 63140
rect 12236 63086 12350 63138
rect 12402 63086 12404 63138
rect 12236 63084 12404 63086
rect 11676 62402 11732 62412
rect 11900 62916 11956 62926
rect 11564 61630 11566 61682
rect 11618 61630 11620 61682
rect 11564 61618 11620 61630
rect 11900 61570 11956 62860
rect 11900 61518 11902 61570
rect 11954 61518 11956 61570
rect 11900 61506 11956 61518
rect 12124 61012 12180 61022
rect 12236 61012 12292 63084
rect 12348 63074 12404 63084
rect 12572 62188 12628 68460
rect 12348 62132 12628 62188
rect 12348 61684 12404 62132
rect 12348 61236 12404 61628
rect 12572 61682 12628 61694
rect 12572 61630 12574 61682
rect 12626 61630 12628 61682
rect 12348 61170 12404 61180
rect 12460 61570 12516 61582
rect 12460 61518 12462 61570
rect 12514 61518 12516 61570
rect 12124 61010 12292 61012
rect 12124 60958 12126 61010
rect 12178 60958 12292 61010
rect 12124 60956 12292 60958
rect 12124 60946 12180 60956
rect 12460 60900 12516 61518
rect 12460 60834 12516 60844
rect 11900 60228 11956 60238
rect 12572 60228 12628 61630
rect 11900 60226 12628 60228
rect 11900 60174 11902 60226
rect 11954 60174 12628 60226
rect 11900 60172 12628 60174
rect 11900 60162 11956 60172
rect 11564 60114 11620 60126
rect 11564 60062 11566 60114
rect 11618 60062 11620 60114
rect 11564 58660 11620 60062
rect 11564 58594 11620 58604
rect 11900 57428 11956 57438
rect 11676 57426 11956 57428
rect 11676 57374 11902 57426
rect 11954 57374 11956 57426
rect 11676 57372 11956 57374
rect 11676 56866 11732 57372
rect 11900 57362 11956 57372
rect 11676 56814 11678 56866
rect 11730 56814 11732 56866
rect 11676 56802 11732 56814
rect 12236 56868 12292 56878
rect 11452 56354 11508 56364
rect 11676 56084 11732 56094
rect 11676 53730 11732 56028
rect 12124 56084 12180 56094
rect 12236 56084 12292 56812
rect 12124 56082 12292 56084
rect 12124 56030 12126 56082
rect 12178 56030 12292 56082
rect 12124 56028 12292 56030
rect 12124 56018 12180 56028
rect 12124 54292 12180 54302
rect 11676 53678 11678 53730
rect 11730 53678 11732 53730
rect 11564 52162 11620 52174
rect 11564 52110 11566 52162
rect 11618 52110 11620 52162
rect 11340 49298 11396 49308
rect 11452 51828 11508 51838
rect 11452 50708 11508 51772
rect 11228 48178 11284 48188
rect 11340 48580 11396 48590
rect 11340 48130 11396 48524
rect 11452 48356 11508 50652
rect 11564 51268 11620 52110
rect 11564 49250 11620 51212
rect 11564 49198 11566 49250
rect 11618 49198 11620 49250
rect 11564 49186 11620 49198
rect 11676 48468 11732 53678
rect 12012 54290 12180 54292
rect 12012 54238 12126 54290
rect 12178 54238 12180 54290
rect 12012 54236 12180 54238
rect 12012 52946 12068 54236
rect 12124 54226 12180 54236
rect 12236 53732 12292 56028
rect 12348 56866 12404 56878
rect 12348 56814 12350 56866
rect 12402 56814 12404 56866
rect 12348 56084 12404 56814
rect 12348 56018 12404 56028
rect 12572 53732 12628 53742
rect 12236 53730 12628 53732
rect 12236 53678 12574 53730
rect 12626 53678 12628 53730
rect 12236 53676 12628 53678
rect 12012 52894 12014 52946
rect 12066 52894 12068 52946
rect 12012 52882 12068 52894
rect 12236 52948 12292 52958
rect 11788 52834 11844 52846
rect 11788 52782 11790 52834
rect 11842 52782 11844 52834
rect 11788 52388 11844 52782
rect 11788 52322 11844 52332
rect 12236 52612 12292 52892
rect 12124 52164 12180 52174
rect 11900 52162 12180 52164
rect 11900 52110 12126 52162
rect 12178 52110 12180 52162
rect 11900 52108 12180 52110
rect 11900 51380 11956 52108
rect 12124 52098 12180 52108
rect 11788 50484 11844 50522
rect 11900 50484 11956 51324
rect 11844 50428 11956 50484
rect 12012 51378 12068 51390
rect 12012 51326 12014 51378
rect 12066 51326 12068 51378
rect 12012 50484 12068 51326
rect 11788 50418 11844 50428
rect 12012 50418 12068 50428
rect 12124 50594 12180 50606
rect 12124 50542 12126 50594
rect 12178 50542 12180 50594
rect 12124 50034 12180 50542
rect 12124 49982 12126 50034
rect 12178 49982 12180 50034
rect 12124 49970 12180 49982
rect 11676 48402 11732 48412
rect 11788 49476 11844 49486
rect 11452 48300 11620 48356
rect 11340 48078 11342 48130
rect 11394 48078 11396 48130
rect 11228 47458 11284 47470
rect 11228 47406 11230 47458
rect 11282 47406 11284 47458
rect 11228 47124 11284 47406
rect 11228 47058 11284 47068
rect 11116 45890 11172 46620
rect 11340 46228 11396 48078
rect 11452 48132 11508 48142
rect 11452 48038 11508 48076
rect 11564 47068 11620 48300
rect 11676 48132 11732 48142
rect 11676 48038 11732 48076
rect 11564 47012 11732 47068
rect 11564 46452 11620 46462
rect 11116 45838 11118 45890
rect 11170 45838 11172 45890
rect 11116 45826 11172 45838
rect 11228 46172 11396 46228
rect 11452 46450 11620 46452
rect 11452 46398 11566 46450
rect 11618 46398 11620 46450
rect 11452 46396 11620 46398
rect 11228 45892 11284 46172
rect 11228 45826 11284 45836
rect 11340 46002 11396 46014
rect 11340 45950 11342 46002
rect 11394 45950 11396 46002
rect 10892 45724 11060 45780
rect 11004 45108 11060 45724
rect 11228 45444 11284 45454
rect 11004 45052 11172 45108
rect 11004 44882 11060 44894
rect 11004 44830 11006 44882
rect 11058 44830 11060 44882
rect 10892 44548 10948 44558
rect 10892 44454 10948 44492
rect 10780 44322 10948 44324
rect 10780 44270 10782 44322
rect 10834 44270 10948 44322
rect 10780 44268 10948 44270
rect 10780 44258 10836 44268
rect 10220 43810 10276 43820
rect 10332 43988 10388 43998
rect 10332 43426 10388 43932
rect 10332 43374 10334 43426
rect 10386 43374 10388 43426
rect 10332 43362 10388 43374
rect 10892 43092 10948 44268
rect 11004 43988 11060 44830
rect 11004 43922 11060 43932
rect 10332 42868 10388 42878
rect 10108 42702 10110 42754
rect 10162 42702 10164 42754
rect 10108 42690 10164 42702
rect 10220 42866 10388 42868
rect 10220 42814 10334 42866
rect 10386 42814 10388 42866
rect 10220 42812 10388 42814
rect 9996 41076 10052 41086
rect 9996 40982 10052 41020
rect 9884 40796 10052 40852
rect 9884 39060 9940 39070
rect 9884 38966 9940 39004
rect 9884 38276 9940 38286
rect 9884 36932 9940 38220
rect 9996 37156 10052 40796
rect 10220 40516 10276 42812
rect 10332 42802 10388 42812
rect 10780 42754 10836 42766
rect 10780 42702 10782 42754
rect 10834 42702 10836 42754
rect 10332 42196 10388 42206
rect 10780 42196 10836 42702
rect 10332 42194 10836 42196
rect 10332 42142 10334 42194
rect 10386 42142 10836 42194
rect 10332 42140 10836 42142
rect 10332 42130 10388 42140
rect 10892 42084 10948 43036
rect 10668 42028 10948 42084
rect 10556 41972 10612 41982
rect 10332 41186 10388 41198
rect 10332 41134 10334 41186
rect 10386 41134 10388 41186
rect 10332 40628 10388 41134
rect 10332 40562 10388 40572
rect 10220 40450 10276 40460
rect 10556 40514 10612 41916
rect 10668 40852 10724 42028
rect 11004 41412 11060 41422
rect 11004 41318 11060 41356
rect 10668 40786 10724 40796
rect 10780 41188 10836 41198
rect 10556 40462 10558 40514
rect 10610 40462 10612 40514
rect 10108 40404 10164 40414
rect 10108 40290 10164 40348
rect 10108 40238 10110 40290
rect 10162 40238 10164 40290
rect 10108 40180 10164 40238
rect 10108 40114 10164 40124
rect 10220 39956 10276 39966
rect 10108 39172 10164 39182
rect 10108 37266 10164 39116
rect 10108 37214 10110 37266
rect 10162 37214 10164 37266
rect 10108 37202 10164 37214
rect 10220 38164 10276 39900
rect 9996 37090 10052 37100
rect 10220 37044 10276 38108
rect 10108 36988 10276 37044
rect 10444 39508 10500 39518
rect 9884 36876 10052 36932
rect 9772 36764 9940 36820
rect 9772 36596 9828 36606
rect 9324 30034 9380 30044
rect 9436 35476 9492 35486
rect 9100 29204 9156 29214
rect 9100 29202 9268 29204
rect 9100 29150 9102 29202
rect 9154 29150 9268 29202
rect 9100 29148 9268 29150
rect 9100 29138 9156 29148
rect 8988 28924 9156 28980
rect 8652 27858 8708 28588
rect 8652 27806 8654 27858
rect 8706 27806 8708 27858
rect 8652 27794 8708 27806
rect 8764 28700 8932 28756
rect 8988 28756 9044 28766
rect 8316 27748 8372 27758
rect 8316 27186 8372 27692
rect 8316 27134 8318 27186
rect 8370 27134 8372 27186
rect 8316 27122 8372 27134
rect 8764 26908 8820 28700
rect 8988 28644 9044 28700
rect 8876 28588 9044 28644
rect 8876 28530 8932 28588
rect 9100 28532 9156 28924
rect 8876 28478 8878 28530
rect 8930 28478 8932 28530
rect 8876 28466 8932 28478
rect 8988 28476 9156 28532
rect 9212 28642 9268 29148
rect 9212 28590 9214 28642
rect 9266 28590 9268 28642
rect 8652 26852 8820 26908
rect 8876 26962 8932 26974
rect 8876 26910 8878 26962
rect 8930 26910 8932 26962
rect 8876 26852 8932 26910
rect 8316 26292 8372 26302
rect 8316 26198 8372 26236
rect 7756 23314 7812 23324
rect 7868 23492 8260 23548
rect 8316 25172 8372 25182
rect 7532 20514 7588 20524
rect 7644 23154 7700 23166
rect 7868 23156 7924 23492
rect 8092 23156 8148 23166
rect 8316 23156 8372 25116
rect 8652 25172 8708 26852
rect 8764 26404 8820 26414
rect 8876 26404 8932 26796
rect 8764 26402 8932 26404
rect 8764 26350 8766 26402
rect 8818 26350 8932 26402
rect 8764 26348 8932 26350
rect 8764 26338 8820 26348
rect 8988 25620 9044 28476
rect 9100 28308 9156 28318
rect 9100 27858 9156 28252
rect 9100 27806 9102 27858
rect 9154 27806 9156 27858
rect 9100 27794 9156 27806
rect 9212 27636 9268 28590
rect 9212 27570 9268 27580
rect 9324 27634 9380 27646
rect 9324 27582 9326 27634
rect 9378 27582 9380 27634
rect 9100 27300 9156 27310
rect 9100 26292 9156 27244
rect 9212 27076 9268 27086
rect 9212 26982 9268 27020
rect 9100 26198 9156 26236
rect 8988 25554 9044 25564
rect 9100 25508 9156 25518
rect 9100 25414 9156 25452
rect 8652 25106 8708 25116
rect 9324 24724 9380 27582
rect 9324 24658 9380 24668
rect 8988 24612 9044 24622
rect 8988 24518 9044 24556
rect 8428 24500 8484 24510
rect 8428 24498 8932 24500
rect 8428 24446 8430 24498
rect 8482 24446 8932 24498
rect 8428 24444 8932 24446
rect 8428 24434 8484 24444
rect 7644 23102 7646 23154
rect 7698 23102 7700 23154
rect 7308 19966 7310 20018
rect 7362 19966 7364 20018
rect 7308 19954 7364 19966
rect 7196 19740 7476 19796
rect 6860 19460 6916 19470
rect 6636 19292 6804 19348
rect 6636 19124 6692 19134
rect 6636 19030 6692 19068
rect 6748 18900 6804 19292
rect 6636 18844 6804 18900
rect 6636 18562 6692 18844
rect 6636 18510 6638 18562
rect 6690 18510 6692 18562
rect 6636 18004 6692 18510
rect 6636 17938 6692 17948
rect 6860 18340 6916 19404
rect 7084 19346 7140 19358
rect 7084 19294 7086 19346
rect 7138 19294 7140 19346
rect 7084 18564 7140 19294
rect 7084 18498 7140 18508
rect 6972 18340 7028 18350
rect 6860 18338 7028 18340
rect 6860 18286 6974 18338
rect 7026 18286 7028 18338
rect 6860 18284 7028 18286
rect 6636 17780 6692 17790
rect 6748 17780 6804 17790
rect 6636 17778 6748 17780
rect 6636 17726 6638 17778
rect 6690 17726 6748 17778
rect 6636 17724 6748 17726
rect 6636 17714 6692 17724
rect 6524 16258 6580 16268
rect 6636 17332 6692 17342
rect 6636 17108 6692 17276
rect 6636 15426 6692 17052
rect 6636 15374 6638 15426
rect 6690 15374 6692 15426
rect 6636 15148 6692 15374
rect 6412 11554 6468 11564
rect 6524 15092 6692 15148
rect 6748 15092 6804 17724
rect 6860 17668 6916 18284
rect 6972 18274 7028 18284
rect 6860 17602 6916 17612
rect 6972 17108 7028 17118
rect 6972 17014 7028 17052
rect 7084 16324 7140 16334
rect 7084 16230 7140 16268
rect 6300 11218 6356 11228
rect 6524 11396 6580 15092
rect 6748 15026 6804 15036
rect 6636 14530 6692 14542
rect 6636 14478 6638 14530
rect 6690 14478 6692 14530
rect 6636 11620 6692 14478
rect 7308 14532 7364 14542
rect 7420 14532 7476 19740
rect 7308 14530 7476 14532
rect 7308 14478 7310 14530
rect 7362 14478 7476 14530
rect 7308 14476 7476 14478
rect 7532 19572 7588 19582
rect 7308 14466 7364 14476
rect 7532 13748 7588 19516
rect 7644 17892 7700 23102
rect 7756 23100 7924 23156
rect 7980 23154 8372 23156
rect 7980 23102 8094 23154
rect 8146 23102 8372 23154
rect 7980 23100 8372 23102
rect 7756 22148 7812 23100
rect 7756 19460 7812 22092
rect 7868 21476 7924 21486
rect 7868 21382 7924 21420
rect 7756 19394 7812 19404
rect 7868 21252 7924 21262
rect 7868 18340 7924 21196
rect 7980 19572 8036 23100
rect 8092 23090 8148 23100
rect 8652 23044 8708 23054
rect 8316 23042 8708 23044
rect 8316 22990 8654 23042
rect 8706 22990 8708 23042
rect 8316 22988 8708 22990
rect 8204 22932 8260 22942
rect 8092 22930 8260 22932
rect 8092 22878 8206 22930
rect 8258 22878 8260 22930
rect 8092 22876 8260 22878
rect 8092 21586 8148 22876
rect 8204 22866 8260 22876
rect 8092 21534 8094 21586
rect 8146 21534 8148 21586
rect 8092 21522 8148 21534
rect 8204 22146 8260 22158
rect 8204 22094 8206 22146
rect 8258 22094 8260 22146
rect 7980 19506 8036 19516
rect 8092 20802 8148 20814
rect 8092 20750 8094 20802
rect 8146 20750 8148 20802
rect 8092 20244 8148 20750
rect 8092 20018 8148 20188
rect 8092 19966 8094 20018
rect 8146 19966 8148 20018
rect 7756 17892 7812 17902
rect 7644 17890 7812 17892
rect 7644 17838 7758 17890
rect 7810 17838 7812 17890
rect 7644 17836 7812 17838
rect 7756 17826 7812 17836
rect 7868 17668 7924 18284
rect 7868 16994 7924 17612
rect 7868 16942 7870 16994
rect 7922 16942 7924 16994
rect 7868 16930 7924 16942
rect 7980 16772 8036 16782
rect 7980 16322 8036 16716
rect 7980 16270 7982 16322
rect 8034 16270 8036 16322
rect 7980 16258 8036 16270
rect 8092 16100 8148 19966
rect 8204 20020 8260 22094
rect 8204 19954 8260 19964
rect 8204 19460 8260 19470
rect 8204 19366 8260 19404
rect 8204 18452 8260 18462
rect 8316 18452 8372 22988
rect 8652 22978 8708 22988
rect 8540 21362 8596 21374
rect 8540 21310 8542 21362
rect 8594 21310 8596 21362
rect 8540 20132 8596 21310
rect 8540 20066 8596 20076
rect 8764 20132 8820 20142
rect 8652 19908 8708 19918
rect 8652 19814 8708 19852
rect 8652 18564 8708 18574
rect 8764 18564 8820 20076
rect 8876 18900 8932 24444
rect 8988 23268 9044 23278
rect 9044 23212 9380 23268
rect 8988 23202 9044 23212
rect 9324 22260 9380 23212
rect 9212 21140 9268 21150
rect 8988 20018 9044 20030
rect 8988 19966 8990 20018
rect 9042 19966 9044 20018
rect 8988 19460 9044 19966
rect 8988 19394 9044 19404
rect 8876 18834 8932 18844
rect 8652 18562 8820 18564
rect 8652 18510 8654 18562
rect 8706 18510 8820 18562
rect 8652 18508 8820 18510
rect 8652 18498 8708 18508
rect 8204 18450 8372 18452
rect 8204 18398 8206 18450
rect 8258 18398 8372 18450
rect 8204 18396 8372 18398
rect 8988 18452 9044 18462
rect 8204 18386 8260 18396
rect 8988 18358 9044 18396
rect 9100 17668 9156 17678
rect 9100 17574 9156 17612
rect 9212 17332 9268 21084
rect 9324 19796 9380 22204
rect 9436 23154 9492 35420
rect 9660 35364 9716 35374
rect 9548 34916 9604 34926
rect 9548 31890 9604 34860
rect 9660 34130 9716 35308
rect 9772 34914 9828 36540
rect 9772 34862 9774 34914
rect 9826 34862 9828 34914
rect 9772 34850 9828 34862
rect 9660 34078 9662 34130
rect 9714 34078 9716 34130
rect 9660 33460 9716 34078
rect 9772 34692 9828 34702
rect 9772 34018 9828 34636
rect 9884 34132 9940 36764
rect 9996 36708 10052 36876
rect 9996 36642 10052 36652
rect 10108 34916 10164 36988
rect 10444 36932 10500 39452
rect 10556 39172 10612 40462
rect 10556 38946 10612 39116
rect 10556 38894 10558 38946
rect 10610 38894 10612 38946
rect 10556 38882 10612 38894
rect 10668 40516 10724 40526
rect 10556 37716 10612 37726
rect 10556 37044 10612 37660
rect 10668 37268 10724 40460
rect 10780 40404 10836 41132
rect 10780 40338 10836 40348
rect 10892 41076 10948 41086
rect 10892 39730 10948 41020
rect 11116 40068 11172 45052
rect 11228 40516 11284 45388
rect 11340 45108 11396 45950
rect 11340 45042 11396 45052
rect 11452 43764 11508 46396
rect 11564 46386 11620 46396
rect 11452 43698 11508 43708
rect 11564 44322 11620 44334
rect 11564 44270 11566 44322
rect 11618 44270 11620 44322
rect 11564 43762 11620 44270
rect 11564 43710 11566 43762
rect 11618 43710 11620 43762
rect 11564 43698 11620 43710
rect 11452 42756 11508 42766
rect 11452 42662 11508 42700
rect 11340 42644 11396 42654
rect 11340 41860 11396 42588
rect 11452 41860 11508 41870
rect 11340 41858 11508 41860
rect 11340 41806 11454 41858
rect 11506 41806 11508 41858
rect 11340 41804 11508 41806
rect 11340 40628 11396 41804
rect 11452 41794 11508 41804
rect 11340 40562 11396 40572
rect 11452 41186 11508 41198
rect 11452 41134 11454 41186
rect 11506 41134 11508 41186
rect 11228 40450 11284 40460
rect 11452 40180 11508 41134
rect 10892 39678 10894 39730
rect 10946 39678 10948 39730
rect 10892 39396 10948 39678
rect 10780 39340 10948 39396
rect 11004 40012 11172 40068
rect 11340 40124 11508 40180
rect 10780 38948 10836 39340
rect 11004 39284 11060 40012
rect 11340 39956 11396 40124
rect 10780 38882 10836 38892
rect 10892 39228 11060 39284
rect 11116 39900 11396 39956
rect 11676 39956 11732 47012
rect 11788 41972 11844 49420
rect 12124 49028 12180 49038
rect 12012 49026 12180 49028
rect 12012 48974 12126 49026
rect 12178 48974 12180 49026
rect 12012 48972 12180 48974
rect 11900 48244 11956 48254
rect 11900 48150 11956 48188
rect 12012 46674 12068 48972
rect 12124 48962 12180 48972
rect 12236 48580 12292 52556
rect 12236 48514 12292 48524
rect 12348 48916 12404 48926
rect 12236 48354 12292 48366
rect 12236 48302 12238 48354
rect 12290 48302 12292 48354
rect 12236 48244 12292 48302
rect 12236 48178 12292 48188
rect 12012 46622 12014 46674
rect 12066 46622 12068 46674
rect 12012 46564 12068 46622
rect 12012 46498 12068 46508
rect 12124 48018 12180 48030
rect 12124 47966 12126 48018
rect 12178 47966 12180 48018
rect 12124 46116 12180 47966
rect 12236 47460 12292 47470
rect 12236 47366 12292 47404
rect 12348 46116 12404 48860
rect 11900 46060 12180 46116
rect 12236 46060 12404 46116
rect 12460 47012 12516 53676
rect 12572 53666 12628 53676
rect 12572 50596 12628 50606
rect 12572 50502 12628 50540
rect 12684 49476 12740 68572
rect 12796 67956 12852 68572
rect 12908 68404 12964 68414
rect 12908 68310 12964 68348
rect 12796 67890 12852 67900
rect 12908 67842 12964 67854
rect 12908 67790 12910 67842
rect 12962 67790 12964 67842
rect 12908 67732 12964 67790
rect 12908 63364 12964 67676
rect 13020 66612 13076 70588
rect 13132 69412 13188 69422
rect 13132 68066 13188 69356
rect 13132 68014 13134 68066
rect 13186 68014 13188 68066
rect 13132 68002 13188 68014
rect 13244 67732 13300 73276
rect 13356 72324 13412 76076
rect 13580 76020 13636 76030
rect 13580 74898 13636 75964
rect 13580 74846 13582 74898
rect 13634 74846 13636 74898
rect 13468 74116 13524 74126
rect 13468 72546 13524 74060
rect 13580 72884 13636 74846
rect 13692 74228 13748 76188
rect 14028 76020 14084 79436
rect 14028 75954 14084 75964
rect 14140 75908 14196 82292
rect 14476 82180 14532 82190
rect 14252 81956 14308 81994
rect 14476 81956 14532 82124
rect 14308 81900 14532 81956
rect 14252 81890 14308 81900
rect 14476 81732 14532 81742
rect 14476 80948 14532 81676
rect 14588 81508 14644 83132
rect 14812 81732 14868 83356
rect 14924 82740 14980 83582
rect 14924 82674 14980 82684
rect 15036 82516 15092 83916
rect 14924 82460 15092 82516
rect 14924 81844 14980 82460
rect 15036 82292 15092 82302
rect 15036 81954 15092 82236
rect 15036 81902 15038 81954
rect 15090 81902 15092 81954
rect 15036 81890 15092 81902
rect 14924 81778 14980 81788
rect 14812 81666 14868 81676
rect 14588 81442 14644 81452
rect 14700 81396 14756 81406
rect 14756 81340 14980 81396
rect 14700 81330 14756 81340
rect 14588 81172 14644 81182
rect 14924 81172 14980 81340
rect 15148 81284 15204 84924
rect 15372 84306 15428 85708
rect 15596 85708 15652 91532
rect 15708 91028 15764 91038
rect 15820 91028 15876 94108
rect 15932 93380 15988 96236
rect 16380 94164 16436 97468
rect 16492 96404 16548 109118
rect 16828 108612 16884 109902
rect 16940 109228 16996 112252
rect 17052 110852 17108 112364
rect 17388 112308 17444 112318
rect 17388 112214 17444 112252
rect 17052 110786 17108 110796
rect 17388 110740 17444 110750
rect 17164 110738 17444 110740
rect 17164 110686 17390 110738
rect 17442 110686 17444 110738
rect 17164 110684 17444 110686
rect 17164 109394 17220 110684
rect 17388 110674 17444 110684
rect 17500 110516 17556 113148
rect 17612 112196 17668 113374
rect 17612 112130 17668 112140
rect 17164 109342 17166 109394
rect 17218 109342 17220 109394
rect 17164 109330 17220 109342
rect 17388 110460 17556 110516
rect 16940 109172 17220 109228
rect 16828 108546 16884 108556
rect 16828 108388 16884 108398
rect 16828 108386 17108 108388
rect 16828 108334 16830 108386
rect 16882 108334 17108 108386
rect 16828 108332 17108 108334
rect 16828 108322 16884 108332
rect 16828 107828 16884 107838
rect 16828 107734 16884 107772
rect 16828 107044 16884 107054
rect 16828 106950 16884 106988
rect 16716 106260 16772 106270
rect 16716 106166 16772 106204
rect 16604 105252 16660 105262
rect 16604 104802 16660 105196
rect 16604 104750 16606 104802
rect 16658 104750 16660 104802
rect 16604 103124 16660 104750
rect 16940 104578 16996 104590
rect 16940 104526 16942 104578
rect 16994 104526 16996 104578
rect 16604 103058 16660 103068
rect 16716 104468 16772 104478
rect 16940 104468 16996 104526
rect 16772 104412 16996 104468
rect 16604 102900 16660 102910
rect 16604 102806 16660 102844
rect 16716 97076 16772 104412
rect 16828 104132 16884 104142
rect 16828 103906 16884 104076
rect 16828 103854 16830 103906
rect 16882 103854 16884 103906
rect 16828 103842 16884 103854
rect 17052 103348 17108 108332
rect 17164 105252 17220 109172
rect 17388 109172 17444 110460
rect 17612 110068 17668 110078
rect 17500 109508 17556 109518
rect 17500 109394 17556 109452
rect 17500 109342 17502 109394
rect 17554 109342 17556 109394
rect 17500 109330 17556 109342
rect 17388 109106 17444 109116
rect 17164 105186 17220 105196
rect 17276 108948 17332 108958
rect 16940 103292 17108 103348
rect 16940 100660 16996 103292
rect 17276 103236 17332 108892
rect 17276 103170 17332 103180
rect 17388 108612 17444 108622
rect 17052 103124 17108 103134
rect 17108 103068 17220 103124
rect 17052 103030 17108 103068
rect 16940 100594 16996 100604
rect 17164 99988 17220 103068
rect 17276 102338 17332 102350
rect 17276 102286 17278 102338
rect 17330 102286 17332 102338
rect 17276 102116 17332 102286
rect 17276 102050 17332 102060
rect 17388 102004 17444 108556
rect 17500 107156 17556 107166
rect 17500 104468 17556 107100
rect 17612 106484 17668 110012
rect 17724 109396 17780 114800
rect 17948 113428 18004 114800
rect 17948 113372 18116 113428
rect 17948 113204 18004 113214
rect 17836 113202 18004 113204
rect 17836 113150 17950 113202
rect 18002 113150 18004 113202
rect 17836 113148 18004 113150
rect 17836 110068 17892 113148
rect 17948 113138 18004 113148
rect 17948 111860 18004 111870
rect 17948 111766 18004 111804
rect 17948 110964 18004 110974
rect 17948 110870 18004 110908
rect 17836 110002 17892 110012
rect 17948 110290 18004 110302
rect 17948 110238 17950 110290
rect 18002 110238 18004 110290
rect 17724 109330 17780 109340
rect 17948 108948 18004 110238
rect 17948 108882 18004 108892
rect 17948 108724 18004 108734
rect 17836 108722 18004 108724
rect 17836 108670 17950 108722
rect 18002 108670 18004 108722
rect 17836 108668 18004 108670
rect 17724 108388 17780 108398
rect 17724 107826 17780 108332
rect 17724 107774 17726 107826
rect 17778 107774 17780 107826
rect 17724 107762 17780 107774
rect 17612 106418 17668 106428
rect 17500 104412 17668 104468
rect 17612 103010 17668 104412
rect 17612 102958 17614 103010
rect 17666 102958 17668 103010
rect 17612 102676 17668 102958
rect 17724 103906 17780 103918
rect 17724 103854 17726 103906
rect 17778 103854 17780 103906
rect 17724 102900 17780 103854
rect 17836 103572 17892 108668
rect 17948 108658 18004 108668
rect 17948 107154 18004 107166
rect 17948 107102 17950 107154
rect 18002 107102 18004 107154
rect 17948 106708 18004 107102
rect 17948 106642 18004 106652
rect 17836 103506 17892 103516
rect 17948 105700 18004 105710
rect 17724 102834 17780 102844
rect 17388 101938 17444 101948
rect 17500 102620 17668 102676
rect 17276 100772 17332 100810
rect 17276 100706 17332 100716
rect 16940 99986 17220 99988
rect 16940 99934 17166 99986
rect 17218 99934 17220 99986
rect 16940 99932 17220 99934
rect 16940 99202 16996 99932
rect 17164 99922 17220 99932
rect 17276 100548 17332 100558
rect 16940 99150 16942 99202
rect 16994 99150 16996 99202
rect 16940 99138 16996 99150
rect 16828 98418 16884 98430
rect 17164 98420 17220 98430
rect 16828 98366 16830 98418
rect 16882 98366 16884 98418
rect 16828 97858 16884 98366
rect 16828 97806 16830 97858
rect 16882 97806 16884 97858
rect 16828 97794 16884 97806
rect 16940 98418 17220 98420
rect 16940 98366 17166 98418
rect 17218 98366 17220 98418
rect 16940 98364 17220 98366
rect 16716 97010 16772 97020
rect 16828 97524 16884 97534
rect 16492 96338 16548 96348
rect 16828 96290 16884 97468
rect 16828 96238 16830 96290
rect 16882 96238 16884 96290
rect 16828 96226 16884 96238
rect 16940 96850 16996 98364
rect 17164 98354 17220 98364
rect 16940 96798 16942 96850
rect 16994 96798 16996 96850
rect 16268 94108 16436 94164
rect 16492 96180 16548 96190
rect 16044 93716 16100 93726
rect 16044 93714 16212 93716
rect 16044 93662 16046 93714
rect 16098 93662 16212 93714
rect 16044 93660 16212 93662
rect 16044 93650 16100 93660
rect 15932 93314 15988 93324
rect 16044 92706 16100 92718
rect 16044 92654 16046 92706
rect 16098 92654 16100 92706
rect 15932 92146 15988 92158
rect 15932 92094 15934 92146
rect 15986 92094 15988 92146
rect 15932 92036 15988 92094
rect 15932 91970 15988 91980
rect 16044 92148 16100 92654
rect 15932 91362 15988 91374
rect 15932 91310 15934 91362
rect 15986 91310 15988 91362
rect 15932 91252 15988 91310
rect 15932 91186 15988 91196
rect 15764 90972 15876 91028
rect 15708 90466 15764 90972
rect 15708 90414 15710 90466
rect 15762 90414 15764 90466
rect 15708 85988 15764 90414
rect 15708 85922 15764 85932
rect 15820 90692 15876 90702
rect 15596 85652 15764 85708
rect 15372 84254 15374 84306
rect 15426 84254 15428 84306
rect 15372 84242 15428 84254
rect 15596 84756 15652 84766
rect 15484 81956 15540 81966
rect 15148 81218 15204 81228
rect 15372 81954 15540 81956
rect 15372 81902 15486 81954
rect 15538 81902 15540 81954
rect 15372 81900 15540 81902
rect 15036 81172 15092 81182
rect 14924 81170 15092 81172
rect 14924 81118 15038 81170
rect 15090 81118 15092 81170
rect 14924 81116 15092 81118
rect 14588 81078 14644 81116
rect 15036 81106 15092 81116
rect 14476 80892 14644 80948
rect 14476 80386 14532 80398
rect 14476 80334 14478 80386
rect 14530 80334 14532 80386
rect 14364 79828 14420 79838
rect 14476 79828 14532 80334
rect 14364 79826 14532 79828
rect 14364 79774 14366 79826
rect 14418 79774 14532 79826
rect 14364 79772 14532 79774
rect 14364 79762 14420 79772
rect 14364 79604 14420 79614
rect 14364 79510 14420 79548
rect 14252 78932 14308 78942
rect 14252 78818 14308 78876
rect 14252 78766 14254 78818
rect 14306 78766 14308 78818
rect 14252 78754 14308 78766
rect 14364 78706 14420 78718
rect 14364 78654 14366 78706
rect 14418 78654 14420 78706
rect 14364 77250 14420 78654
rect 14588 78372 14644 80892
rect 15148 80946 15204 80958
rect 15148 80894 15150 80946
rect 15202 80894 15204 80946
rect 14812 80724 14868 80734
rect 14812 80386 14868 80668
rect 15036 80724 15092 80734
rect 14812 80334 14814 80386
rect 14866 80334 14868 80386
rect 14812 80322 14868 80334
rect 14924 80610 14980 80622
rect 14924 80558 14926 80610
rect 14978 80558 14980 80610
rect 14700 80276 14756 80286
rect 14700 78932 14756 80220
rect 14924 80164 14980 80558
rect 15036 80498 15092 80668
rect 15036 80446 15038 80498
rect 15090 80446 15092 80498
rect 15036 80434 15092 80446
rect 15148 80612 15204 80894
rect 14924 80098 14980 80108
rect 15148 79604 15204 80556
rect 15260 80500 15316 80510
rect 15372 80500 15428 81900
rect 15484 81890 15540 81900
rect 15484 81732 15540 81742
rect 15484 81284 15540 81676
rect 15484 80948 15540 81228
rect 15596 80948 15652 84700
rect 15708 82292 15764 85652
rect 15820 84756 15876 90636
rect 16044 90578 16100 92092
rect 16156 91364 16212 93660
rect 16268 92708 16324 94108
rect 16268 92642 16324 92652
rect 16380 93828 16436 93838
rect 16380 93714 16436 93772
rect 16380 93662 16382 93714
rect 16434 93662 16436 93714
rect 16156 91298 16212 91308
rect 16268 92372 16324 92382
rect 16044 90526 16046 90578
rect 16098 90526 16100 90578
rect 16044 90514 16100 90526
rect 16044 90244 16100 90254
rect 16044 89794 16100 90188
rect 16044 89742 16046 89794
rect 16098 89742 16100 89794
rect 16044 89730 16100 89742
rect 16044 85988 16100 85998
rect 16044 85874 16100 85932
rect 16044 85822 16046 85874
rect 16098 85822 16100 85874
rect 16044 85810 16100 85822
rect 16156 85762 16212 85774
rect 16156 85710 16158 85762
rect 16210 85710 16212 85762
rect 16044 85540 16100 85550
rect 16044 85092 16100 85484
rect 16044 84998 16100 85036
rect 16156 84980 16212 85710
rect 16268 85708 16324 92316
rect 16380 92146 16436 93662
rect 16492 92372 16548 96124
rect 16828 95844 16884 95854
rect 16828 94722 16884 95788
rect 16828 94670 16830 94722
rect 16882 94670 16884 94722
rect 16828 94658 16884 94670
rect 16940 93828 16996 96798
rect 17164 97636 17220 97646
rect 17052 96180 17108 96190
rect 17052 96086 17108 96124
rect 17164 96178 17220 97580
rect 17164 96126 17166 96178
rect 17218 96126 17220 96178
rect 17164 96114 17220 96126
rect 17164 94610 17220 94622
rect 17164 94558 17166 94610
rect 17218 94558 17220 94610
rect 17164 94164 17220 94558
rect 17164 94098 17220 94108
rect 16828 93772 16996 93828
rect 16604 93490 16660 93502
rect 16604 93438 16606 93490
rect 16658 93438 16660 93490
rect 16604 92484 16660 93438
rect 16604 92418 16660 92428
rect 16492 92306 16548 92316
rect 16380 92094 16382 92146
rect 16434 92094 16436 92146
rect 16380 85876 16436 92094
rect 16604 91922 16660 91934
rect 16604 91870 16606 91922
rect 16658 91870 16660 91922
rect 16492 90578 16548 90590
rect 16492 90526 16494 90578
rect 16546 90526 16548 90578
rect 16492 90244 16548 90526
rect 16492 90178 16548 90188
rect 16604 88900 16660 91870
rect 16828 91364 16884 93772
rect 17052 93716 17108 93726
rect 16940 93660 17052 93716
rect 16940 91924 16996 93660
rect 17052 93622 17108 93660
rect 17052 92932 17108 92942
rect 17052 92838 17108 92876
rect 17052 92148 17108 92158
rect 17052 92054 17108 92092
rect 17164 92036 17220 92046
rect 16940 91868 17108 91924
rect 16828 91308 16996 91364
rect 16716 91250 16772 91262
rect 16716 91198 16718 91250
rect 16770 91198 16772 91250
rect 16716 91028 16772 91198
rect 16716 90962 16772 90972
rect 16828 91140 16884 91150
rect 16716 90356 16772 90366
rect 16716 90262 16772 90300
rect 16604 88834 16660 88844
rect 16716 87556 16772 87566
rect 16380 85810 16436 85820
rect 16492 87444 16548 87454
rect 16268 85652 16436 85708
rect 16156 84914 16212 84924
rect 15820 84700 16324 84756
rect 15932 84308 15988 84318
rect 15932 82516 15988 84252
rect 16044 84196 16100 84206
rect 16044 84102 16100 84140
rect 16156 84084 16212 84094
rect 16044 83524 16100 83534
rect 16044 83430 16100 83468
rect 16044 82964 16100 82974
rect 16044 82738 16100 82908
rect 16044 82686 16046 82738
rect 16098 82686 16100 82738
rect 16044 82674 16100 82686
rect 15932 82450 15988 82460
rect 15708 82236 16100 82292
rect 15708 82068 15764 82078
rect 15708 81974 15764 82012
rect 15820 81954 15876 81966
rect 15820 81902 15822 81954
rect 15874 81902 15876 81954
rect 15708 81284 15764 81294
rect 15708 81190 15764 81228
rect 15596 80892 15764 80948
rect 15484 80882 15540 80892
rect 15260 80498 15428 80500
rect 15260 80446 15262 80498
rect 15314 80446 15428 80498
rect 15260 80444 15428 80446
rect 15260 80434 15316 80444
rect 15148 79538 15204 79548
rect 15596 79604 15652 79614
rect 15596 79510 15652 79548
rect 14924 79156 14980 79166
rect 14812 78932 14868 78942
rect 14700 78930 14868 78932
rect 14700 78878 14814 78930
rect 14866 78878 14868 78930
rect 14700 78876 14868 78878
rect 14812 78596 14868 78876
rect 14588 78306 14644 78316
rect 14700 78540 14868 78596
rect 14364 77198 14366 77250
rect 14418 77198 14420 77250
rect 14364 77186 14420 77198
rect 14588 77810 14644 77822
rect 14588 77758 14590 77810
rect 14642 77758 14644 77810
rect 14588 76466 14644 77758
rect 14588 76414 14590 76466
rect 14642 76414 14644 76466
rect 14588 76402 14644 76414
rect 14700 76132 14756 78540
rect 14812 78372 14868 78382
rect 14812 77362 14868 78316
rect 14812 77310 14814 77362
rect 14866 77310 14868 77362
rect 14812 77298 14868 77310
rect 14364 76076 14756 76132
rect 14924 76466 14980 79100
rect 15148 78708 15204 78718
rect 15148 77364 15204 78652
rect 15484 78036 15540 78046
rect 15484 77942 15540 77980
rect 14924 76414 14926 76466
rect 14978 76414 14980 76466
rect 14140 75852 14308 75908
rect 14252 75684 14308 75852
rect 14028 75628 14308 75684
rect 13804 74788 13860 74798
rect 13804 74694 13860 74732
rect 13692 73332 13748 74172
rect 13692 73238 13748 73276
rect 13804 73108 13860 73118
rect 13804 73014 13860 73052
rect 13580 72818 13636 72828
rect 13468 72494 13470 72546
rect 13522 72494 13524 72546
rect 13468 72482 13524 72494
rect 13804 72660 13860 72670
rect 13356 72258 13412 72268
rect 13804 71652 13860 72604
rect 13916 72658 13972 72670
rect 13916 72606 13918 72658
rect 13970 72606 13972 72658
rect 13916 72324 13972 72606
rect 13916 72258 13972 72268
rect 13916 71652 13972 71662
rect 13804 71650 13972 71652
rect 13804 71598 13918 71650
rect 13970 71598 13972 71650
rect 13804 71596 13972 71598
rect 13916 71586 13972 71596
rect 14028 69748 14084 75628
rect 14140 75458 14196 75470
rect 14140 75406 14142 75458
rect 14194 75406 14196 75458
rect 14140 74900 14196 75406
rect 14252 74900 14308 74910
rect 14140 74898 14308 74900
rect 14140 74846 14254 74898
rect 14306 74846 14308 74898
rect 14140 74844 14308 74846
rect 14252 74834 14308 74844
rect 14252 73218 14308 73230
rect 14252 73166 14254 73218
rect 14306 73166 14308 73218
rect 14252 72772 14308 73166
rect 14252 72706 14308 72716
rect 14252 71540 14308 71550
rect 14252 71446 14308 71484
rect 14364 71204 14420 76076
rect 14924 74898 14980 76414
rect 14924 74846 14926 74898
rect 14978 74846 14980 74898
rect 14812 74788 14868 74798
rect 14812 74226 14868 74732
rect 14812 74174 14814 74226
rect 14866 74174 14868 74226
rect 14476 74116 14532 74126
rect 14476 74022 14532 74060
rect 14588 72996 14644 73006
rect 14812 72996 14868 74174
rect 13692 69692 14084 69748
rect 14252 71148 14420 71204
rect 14476 71988 14532 71998
rect 13244 67666 13300 67676
rect 13356 68852 13412 68862
rect 13020 66556 13188 66612
rect 13020 65604 13076 65614
rect 13020 65510 13076 65548
rect 13132 64706 13188 66556
rect 13356 65378 13412 68796
rect 13580 68404 13636 68414
rect 13580 67954 13636 68348
rect 13580 67902 13582 67954
rect 13634 67902 13636 67954
rect 13580 67890 13636 67902
rect 13468 66834 13524 66846
rect 13468 66782 13470 66834
rect 13522 66782 13524 66834
rect 13468 65716 13524 66782
rect 13692 66612 13748 69692
rect 14252 69636 14308 71148
rect 13916 69580 14308 69636
rect 14364 70978 14420 70990
rect 14364 70926 14366 70978
rect 14418 70926 14420 70978
rect 14364 70532 14420 70926
rect 13804 66836 13860 66846
rect 13804 66742 13860 66780
rect 13692 66556 13860 66612
rect 13468 65650 13524 65660
rect 13580 65828 13636 65838
rect 13356 65326 13358 65378
rect 13410 65326 13412 65378
rect 13356 65314 13412 65326
rect 13580 64930 13636 65772
rect 13580 64878 13582 64930
rect 13634 64878 13636 64930
rect 13580 64866 13636 64878
rect 13692 65156 13748 65166
rect 13132 64654 13134 64706
rect 13186 64654 13188 64706
rect 13132 64036 13188 64654
rect 13132 63970 13188 63980
rect 13580 64372 13636 64382
rect 12908 63298 12964 63308
rect 13468 63364 13524 63374
rect 12908 63138 12964 63150
rect 12908 63086 12910 63138
rect 12962 63086 12964 63138
rect 12908 62916 12964 63086
rect 12908 62850 12964 62860
rect 13468 62804 13524 63308
rect 13468 62738 13524 62748
rect 13020 61572 13076 61582
rect 13020 61478 13076 61516
rect 13580 61570 13636 64316
rect 13580 61518 13582 61570
rect 13634 61518 13636 61570
rect 13132 61348 13188 61358
rect 13132 60786 13188 61292
rect 13132 60734 13134 60786
rect 13186 60734 13188 60786
rect 13132 60676 13188 60734
rect 13132 60610 13188 60620
rect 13580 60228 13636 61518
rect 13692 60674 13748 65100
rect 13804 61572 13860 66556
rect 13916 66164 13972 69580
rect 14140 69300 14196 69310
rect 14364 69300 14420 70476
rect 14476 70082 14532 71932
rect 14588 71874 14644 72940
rect 14588 71822 14590 71874
rect 14642 71822 14644 71874
rect 14588 71810 14644 71822
rect 14700 72940 14868 72996
rect 14924 72996 14980 74846
rect 15036 77308 15204 77364
rect 15036 73556 15092 77308
rect 15484 76916 15540 76926
rect 15036 73500 15204 73556
rect 15036 73332 15092 73342
rect 15036 73238 15092 73276
rect 14476 70030 14478 70082
rect 14530 70030 14532 70082
rect 14476 70018 14532 70030
rect 14588 69522 14644 69534
rect 14588 69470 14590 69522
rect 14642 69470 14644 69522
rect 14140 69298 14420 69300
rect 14140 69246 14142 69298
rect 14194 69246 14420 69298
rect 14140 69244 14420 69246
rect 14476 69412 14532 69422
rect 14140 69234 14196 69244
rect 14476 69076 14532 69356
rect 14140 68740 14196 68750
rect 14476 68740 14532 69020
rect 14588 68852 14644 69470
rect 14588 68786 14644 68796
rect 14140 68514 14196 68684
rect 14140 68462 14142 68514
rect 14194 68462 14196 68514
rect 14140 68450 14196 68462
rect 14252 68738 14532 68740
rect 14252 68686 14478 68738
rect 14530 68686 14532 68738
rect 14252 68684 14532 68686
rect 14140 67844 14196 67854
rect 14140 67750 14196 67788
rect 14140 67396 14196 67406
rect 14140 67170 14196 67340
rect 14140 67118 14142 67170
rect 14194 67118 14196 67170
rect 14140 67106 14196 67118
rect 13916 65828 13972 66108
rect 13916 65762 13972 65772
rect 14252 66274 14308 68684
rect 14476 68674 14532 68684
rect 14700 68516 14756 72940
rect 14924 72930 14980 72940
rect 14924 72660 14980 72670
rect 14812 71092 14868 71102
rect 14812 70998 14868 71036
rect 14252 66222 14254 66274
rect 14306 66222 14308 66274
rect 14252 65604 14308 66222
rect 14252 65538 14308 65548
rect 14476 68460 14756 68516
rect 14812 69970 14868 69982
rect 14812 69918 14814 69970
rect 14866 69918 14868 69970
rect 14812 68516 14868 69918
rect 14252 64036 14308 64046
rect 14252 63942 14308 63980
rect 14476 63364 14532 68460
rect 14812 68450 14868 68460
rect 14924 67620 14980 72604
rect 15036 72322 15092 72334
rect 15036 72270 15038 72322
rect 15090 72270 15092 72322
rect 15036 71762 15092 72270
rect 15036 71710 15038 71762
rect 15090 71710 15092 71762
rect 15036 71698 15092 71710
rect 15148 71540 15204 73500
rect 15484 71762 15540 76860
rect 15484 71710 15486 71762
rect 15538 71710 15540 71762
rect 14924 67554 14980 67564
rect 15036 71484 15204 71540
rect 15260 71652 15316 71662
rect 14700 67172 14756 67182
rect 14588 67058 14644 67070
rect 14588 67006 14590 67058
rect 14642 67006 14644 67058
rect 14588 65714 14644 67006
rect 14700 66498 14756 67116
rect 14924 67060 14980 67070
rect 14924 66966 14980 67004
rect 14700 66446 14702 66498
rect 14754 66446 14756 66498
rect 14700 66434 14756 66446
rect 15036 66612 15092 71484
rect 15260 68852 15316 71596
rect 15372 70532 15428 70542
rect 15372 70306 15428 70476
rect 15372 70254 15374 70306
rect 15426 70254 15428 70306
rect 15372 70242 15428 70254
rect 15260 68796 15428 68852
rect 15260 68628 15316 68638
rect 15260 68534 15316 68572
rect 15260 67956 15316 67966
rect 15260 67842 15316 67900
rect 15260 67790 15262 67842
rect 15314 67790 15316 67842
rect 15260 67284 15316 67790
rect 15260 67218 15316 67228
rect 15148 66836 15204 66846
rect 15148 66742 15204 66780
rect 14588 65662 14590 65714
rect 14642 65662 14644 65714
rect 14588 65650 14644 65662
rect 14700 64484 14756 64494
rect 14476 63298 14532 63308
rect 14588 64482 14756 64484
rect 14588 64430 14702 64482
rect 14754 64430 14756 64482
rect 14588 64428 14756 64430
rect 13916 63140 13972 63150
rect 13916 63046 13972 63084
rect 14252 62468 14308 62478
rect 14252 62374 14308 62412
rect 14588 62354 14644 64428
rect 14700 64418 14756 64428
rect 14700 63812 14756 63822
rect 15036 63812 15092 66556
rect 14700 63810 15092 63812
rect 14700 63758 14702 63810
rect 14754 63758 15092 63810
rect 14700 63756 15092 63758
rect 14700 63746 14756 63756
rect 15148 63364 15204 63374
rect 15372 63364 15428 68796
rect 15484 67060 15540 71710
rect 15708 71652 15764 80892
rect 15820 80612 15876 81902
rect 15820 80546 15876 80556
rect 15932 81508 15988 81518
rect 15932 79828 15988 81452
rect 16044 81058 16100 82236
rect 16156 81508 16212 84028
rect 16156 81442 16212 81452
rect 16268 82628 16324 84700
rect 16380 83748 16436 85652
rect 16492 84306 16548 87388
rect 16604 85764 16660 85802
rect 16604 85698 16660 85708
rect 16492 84254 16494 84306
rect 16546 84254 16548 84306
rect 16492 84242 16548 84254
rect 16604 85540 16660 85550
rect 16604 84308 16660 85484
rect 16604 84242 16660 84252
rect 16716 84084 16772 87500
rect 16828 85988 16884 91084
rect 16828 85922 16884 85932
rect 16940 89796 16996 91308
rect 17052 91362 17108 91868
rect 17052 91310 17054 91362
rect 17106 91310 17108 91362
rect 17052 91298 17108 91310
rect 17164 90578 17220 91980
rect 17164 90526 17166 90578
rect 17218 90526 17220 90578
rect 17164 90514 17220 90526
rect 16940 85204 16996 89740
rect 17276 89684 17332 100492
rect 17388 99314 17444 99326
rect 17388 99262 17390 99314
rect 17442 99262 17444 99314
rect 17388 98980 17444 99262
rect 17388 98914 17444 98924
rect 17500 94500 17556 102620
rect 17612 102452 17668 102462
rect 17612 102358 17668 102396
rect 17948 101108 18004 105644
rect 17836 101052 18004 101108
rect 17612 100882 17668 100894
rect 17612 100830 17614 100882
rect 17666 100830 17668 100882
rect 17612 99764 17668 100830
rect 17836 100772 17892 101052
rect 17724 99876 17780 99886
rect 17724 99782 17780 99820
rect 17612 99698 17668 99708
rect 17836 98644 17892 100716
rect 18060 100548 18116 113372
rect 18172 108164 18228 114800
rect 18396 113204 18452 114800
rect 18508 113988 18564 113998
rect 18508 113538 18564 113932
rect 18620 113764 18676 114800
rect 18844 113988 18900 114800
rect 18844 113922 18900 113932
rect 18620 113698 18676 113708
rect 19068 113540 19124 114800
rect 18508 113486 18510 113538
rect 18562 113486 18564 113538
rect 18508 113474 18564 113486
rect 18732 113484 19124 113540
rect 19180 113652 19236 113662
rect 19180 113538 19236 113596
rect 19180 113486 19182 113538
rect 19234 113486 19236 113538
rect 18732 113316 18788 113484
rect 19180 113474 19236 113486
rect 18284 113148 18452 113204
rect 18508 113260 18788 113316
rect 18844 113314 18900 113326
rect 18844 113262 18846 113314
rect 18898 113262 18900 113314
rect 18284 111636 18340 113148
rect 18284 111570 18340 111580
rect 18396 111634 18452 111646
rect 18396 111582 18398 111634
rect 18450 111582 18452 111634
rect 18396 111300 18452 111582
rect 18284 111244 18452 111300
rect 18284 111188 18340 111244
rect 18284 109844 18340 111132
rect 18284 109778 18340 109788
rect 18396 110066 18452 110078
rect 18396 110014 18398 110066
rect 18450 110014 18452 110066
rect 18172 108098 18228 108108
rect 18396 106930 18452 110014
rect 18508 110068 18564 113260
rect 18620 112420 18676 112430
rect 18620 112418 18788 112420
rect 18620 112366 18622 112418
rect 18674 112366 18788 112418
rect 18620 112364 18788 112366
rect 18620 112354 18676 112364
rect 18732 110292 18788 112364
rect 18844 110404 18900 113262
rect 19068 113316 19124 113326
rect 18956 112756 19012 112766
rect 18956 112642 19012 112700
rect 18956 112590 18958 112642
rect 19010 112590 19012 112642
rect 18956 112578 19012 112590
rect 19068 111748 19124 113260
rect 19292 112084 19348 114800
rect 19516 113540 19572 114800
rect 19516 113474 19572 113484
rect 19628 113764 19684 113774
rect 19516 113314 19572 113326
rect 19516 113262 19518 113314
rect 19570 113262 19572 113314
rect 19516 113204 19572 113262
rect 19516 113138 19572 113148
rect 19516 112868 19572 112878
rect 19516 112418 19572 112812
rect 19516 112366 19518 112418
rect 19570 112366 19572 112418
rect 19516 112354 19572 112366
rect 19292 112028 19460 112084
rect 18956 111692 19124 111748
rect 18956 110628 19012 111692
rect 19068 111524 19124 111534
rect 19068 111522 19236 111524
rect 19068 111470 19070 111522
rect 19122 111470 19236 111522
rect 19068 111468 19236 111470
rect 19068 111458 19124 111468
rect 19068 110852 19124 110862
rect 19068 110758 19124 110796
rect 18956 110572 19124 110628
rect 18956 110404 19012 110414
rect 18844 110402 19012 110404
rect 18844 110350 18958 110402
rect 19010 110350 19012 110402
rect 18844 110348 19012 110350
rect 18956 110338 19012 110348
rect 18732 110236 18900 110292
rect 18508 110012 18788 110068
rect 18396 106878 18398 106930
rect 18450 106878 18452 106930
rect 18396 106820 18452 106878
rect 18396 106754 18452 106764
rect 18508 109844 18564 109854
rect 18508 108610 18564 109788
rect 18508 108558 18510 108610
rect 18562 108558 18564 108610
rect 18508 106260 18564 108558
rect 18620 109396 18676 109434
rect 18620 106484 18676 109340
rect 18732 106708 18788 110012
rect 18732 106642 18788 106652
rect 18620 106418 18676 106428
rect 18508 106194 18564 106204
rect 18844 105924 18900 110236
rect 18956 110180 19012 110190
rect 18956 109396 19012 110124
rect 18956 109330 19012 109340
rect 19068 109394 19124 110572
rect 19068 109342 19070 109394
rect 19122 109342 19124 109394
rect 19068 109330 19124 109342
rect 19180 109228 19236 111468
rect 19292 110180 19348 110190
rect 19292 110086 19348 110124
rect 19404 109956 19460 112028
rect 19516 111188 19572 111198
rect 19516 111074 19572 111132
rect 19516 111022 19518 111074
rect 19570 111022 19572 111074
rect 19516 111010 19572 111022
rect 19628 110852 19684 113708
rect 19740 112532 19796 114800
rect 19852 114324 19908 114334
rect 19852 112868 19908 114268
rect 19964 112868 20020 114800
rect 20188 113316 20244 114800
rect 20188 113250 20244 113260
rect 20412 113316 20468 114800
rect 20412 113250 20468 113260
rect 20524 114436 20580 114446
rect 20188 113092 20244 113102
rect 20188 113090 20468 113092
rect 20188 113038 20190 113090
rect 20242 113038 20468 113090
rect 20188 113036 20468 113038
rect 20188 113026 20244 113036
rect 19964 112812 20132 112868
rect 19852 112802 19908 112812
rect 19740 112466 19796 112476
rect 19964 112644 20020 112654
rect 19852 112306 19908 112318
rect 19852 112254 19854 112306
rect 19906 112254 19908 112306
rect 19852 111972 19908 112254
rect 19852 111906 19908 111916
rect 19964 111748 20020 112588
rect 18508 105868 18900 105924
rect 18956 109172 19236 109228
rect 19292 109900 19460 109956
rect 19516 110796 19684 110852
rect 19852 111692 20020 111748
rect 18172 104468 18228 104478
rect 18172 104374 18228 104412
rect 18508 104132 18564 105868
rect 18956 105588 19012 109172
rect 19180 108948 19236 108958
rect 18396 104076 18564 104132
rect 18844 105532 19012 105588
rect 19068 105588 19124 105626
rect 18396 103236 18452 104076
rect 18508 103906 18564 103918
rect 18508 103854 18510 103906
rect 18562 103854 18564 103906
rect 18508 103348 18564 103854
rect 18732 103348 18788 103358
rect 18508 103346 18788 103348
rect 18508 103294 18734 103346
rect 18786 103294 18788 103346
rect 18508 103292 18788 103294
rect 18732 103282 18788 103292
rect 18396 103180 18564 103236
rect 18508 101108 18564 103180
rect 18844 101780 18900 105532
rect 19068 105522 19124 105532
rect 19068 105252 19124 105262
rect 18956 104020 19012 104030
rect 18956 103926 19012 103964
rect 19068 103906 19124 105196
rect 19068 103854 19070 103906
rect 19122 103854 19124 103906
rect 19068 103842 19124 103854
rect 19180 103122 19236 108892
rect 19180 103070 19182 103122
rect 19234 103070 19236 103122
rect 19180 103058 19236 103070
rect 18844 101714 18900 101724
rect 19292 101108 19348 109900
rect 19404 109282 19460 109294
rect 19404 109230 19406 109282
rect 19458 109230 19460 109282
rect 19404 109172 19460 109230
rect 19404 109106 19460 109116
rect 19404 105588 19460 105598
rect 19404 105494 19460 105532
rect 19516 104692 19572 110796
rect 19740 110628 19796 110638
rect 19628 110290 19684 110302
rect 19628 110238 19630 110290
rect 19682 110238 19684 110290
rect 19628 109060 19684 110238
rect 19628 108994 19684 109004
rect 19740 108948 19796 110572
rect 19852 109394 19908 111692
rect 20076 110964 20132 112812
rect 20300 112532 20356 112542
rect 20076 110898 20132 110908
rect 20188 111858 20244 111870
rect 20188 111806 20190 111858
rect 20242 111806 20244 111858
rect 19964 110404 20020 110414
rect 19964 110310 20020 110348
rect 19852 109342 19854 109394
rect 19906 109342 19908 109394
rect 19852 109330 19908 109342
rect 19964 109508 20020 109518
rect 19740 108882 19796 108892
rect 19852 106484 19908 106494
rect 19516 104636 19796 104692
rect 19516 104468 19572 104478
rect 19516 103906 19572 104412
rect 19516 103854 19518 103906
rect 19570 103854 19572 103906
rect 19516 103842 19572 103854
rect 19628 104020 19684 104030
rect 19516 102900 19572 102910
rect 19516 102806 19572 102844
rect 19292 101052 19460 101108
rect 18508 101042 18564 101052
rect 18060 100482 18116 100492
rect 18844 99762 18900 99774
rect 18844 99710 18846 99762
rect 18898 99710 18900 99762
rect 18844 99204 18900 99710
rect 18956 99428 19012 99438
rect 18956 99334 19012 99372
rect 19292 99316 19348 99326
rect 19292 99222 19348 99260
rect 18844 99138 18900 99148
rect 18508 98980 18564 98990
rect 18508 98978 19012 98980
rect 18508 98926 18510 98978
rect 18562 98926 19012 98978
rect 18508 98924 19012 98926
rect 18508 98914 18564 98924
rect 17724 98588 17892 98644
rect 17724 97468 17780 98588
rect 18844 98532 18900 98542
rect 18844 98438 18900 98476
rect 18172 98420 18228 98430
rect 18172 98326 18228 98364
rect 18620 98420 18676 98430
rect 18284 98196 18340 98206
rect 18060 97972 18116 97982
rect 18060 97746 18116 97916
rect 18060 97694 18062 97746
rect 18114 97694 18116 97746
rect 18060 97682 18116 97694
rect 17500 94434 17556 94444
rect 17612 97412 17780 97468
rect 18284 97636 18340 98140
rect 17612 93154 17668 97412
rect 18284 97074 18340 97580
rect 18396 97748 18452 97758
rect 18396 97634 18452 97692
rect 18396 97582 18398 97634
rect 18450 97582 18452 97634
rect 18396 97570 18452 97582
rect 18284 97022 18286 97074
rect 18338 97022 18340 97074
rect 18284 97010 18340 97022
rect 18620 97074 18676 98364
rect 18956 98418 19012 98924
rect 18956 98366 18958 98418
rect 19010 98366 19012 98418
rect 18732 98306 18788 98318
rect 18732 98254 18734 98306
rect 18786 98254 18788 98306
rect 18732 97524 18788 98254
rect 18956 97636 19012 98366
rect 19180 98418 19236 98430
rect 19180 98366 19182 98418
rect 19234 98366 19236 98418
rect 19068 97860 19124 97870
rect 19180 97860 19236 98366
rect 19292 98420 19348 98430
rect 19292 98326 19348 98364
rect 19404 98196 19460 101052
rect 19068 97858 19236 97860
rect 19068 97806 19070 97858
rect 19122 97806 19236 97858
rect 19068 97804 19236 97806
rect 19292 98140 19460 98196
rect 19516 99204 19572 99214
rect 19068 97794 19124 97804
rect 19180 97636 19236 97646
rect 18956 97634 19236 97636
rect 18956 97582 19182 97634
rect 19234 97582 19236 97634
rect 18956 97580 19236 97582
rect 19180 97570 19236 97580
rect 18732 97458 18788 97468
rect 18620 97022 18622 97074
rect 18674 97022 18676 97074
rect 18620 97010 18676 97022
rect 19068 97410 19124 97422
rect 19068 97358 19070 97410
rect 19122 97358 19124 97410
rect 17724 96850 17780 96862
rect 17724 96798 17726 96850
rect 17778 96798 17780 96850
rect 17724 96068 17780 96798
rect 18620 96852 18676 96862
rect 18620 96850 18788 96852
rect 18620 96798 18622 96850
rect 18674 96798 18788 96850
rect 18620 96796 18788 96798
rect 18620 96786 18676 96796
rect 18284 96516 18340 96526
rect 17724 96002 17780 96012
rect 17836 96180 17892 96190
rect 17612 93102 17614 93154
rect 17666 93102 17668 93154
rect 17612 93090 17668 93102
rect 17724 94386 17780 94398
rect 17724 94334 17726 94386
rect 17778 94334 17780 94386
rect 17724 94052 17780 94334
rect 17500 93042 17556 93054
rect 17500 92990 17502 93042
rect 17554 92990 17556 93042
rect 17500 92596 17556 92990
rect 17724 92932 17780 93996
rect 17836 93940 17892 96124
rect 18060 96068 18116 96078
rect 17836 93874 17892 93884
rect 17948 95732 18004 95742
rect 17836 93716 17892 93726
rect 17836 93622 17892 93660
rect 17724 92866 17780 92876
rect 17500 92530 17556 92540
rect 17836 92372 17892 92382
rect 17836 92146 17892 92316
rect 17836 92094 17838 92146
rect 17890 92094 17892 92146
rect 17836 92082 17892 92094
rect 17948 92148 18004 95676
rect 17948 92082 18004 92092
rect 17724 91476 17780 91486
rect 17724 91382 17780 91420
rect 17500 91362 17556 91374
rect 17500 91310 17502 91362
rect 17554 91310 17556 91362
rect 17500 90244 17556 91310
rect 17948 91252 18004 91262
rect 18060 91252 18116 96012
rect 18172 94724 18228 94762
rect 18172 94658 18228 94668
rect 18172 94500 18228 94510
rect 18172 93156 18228 94444
rect 18284 93268 18340 96460
rect 18620 96068 18676 96078
rect 18508 96066 18676 96068
rect 18508 96014 18622 96066
rect 18674 96014 18676 96066
rect 18508 96012 18676 96014
rect 18396 95956 18452 95966
rect 18396 95282 18452 95900
rect 18396 95230 18398 95282
rect 18450 95230 18452 95282
rect 18396 94052 18452 95230
rect 18396 93986 18452 93996
rect 18284 93212 18452 93268
rect 18172 93100 18340 93156
rect 18172 91364 18228 91374
rect 18172 91270 18228 91308
rect 18004 91196 18116 91252
rect 17724 91140 17780 91150
rect 17724 90578 17780 91084
rect 17724 90526 17726 90578
rect 17778 90526 17780 90578
rect 17724 90514 17780 90526
rect 17500 90178 17556 90188
rect 17724 90244 17780 90254
rect 17276 89628 17668 89684
rect 17164 89572 17220 89582
rect 17164 89570 17556 89572
rect 17164 89518 17166 89570
rect 17218 89518 17556 89570
rect 17164 89516 17556 89518
rect 17164 89506 17220 89516
rect 17276 89348 17332 89358
rect 17164 85876 17220 85886
rect 17164 85782 17220 85820
rect 17164 85428 17220 85438
rect 16940 85148 17108 85204
rect 16828 85090 16884 85102
rect 16828 85038 16830 85090
rect 16882 85038 16884 85090
rect 16828 84868 16884 85038
rect 16828 84802 16884 84812
rect 16716 84018 16772 84028
rect 16940 84532 16996 84542
rect 16380 83692 16772 83748
rect 16716 83634 16772 83692
rect 16716 83582 16718 83634
rect 16770 83582 16772 83634
rect 16492 82628 16548 82638
rect 16268 82626 16548 82628
rect 16268 82574 16494 82626
rect 16546 82574 16548 82626
rect 16268 82572 16548 82574
rect 16044 81006 16046 81058
rect 16098 81006 16100 81058
rect 16044 80994 16100 81006
rect 15820 79772 15988 79828
rect 16156 80946 16212 80958
rect 16156 80894 16158 80946
rect 16210 80894 16212 80946
rect 15820 78596 15876 79772
rect 15932 79602 15988 79614
rect 15932 79550 15934 79602
rect 15986 79550 15988 79602
rect 15932 79042 15988 79550
rect 15932 78990 15934 79042
rect 15986 78990 15988 79042
rect 15932 78978 15988 78990
rect 15820 78148 15876 78540
rect 15820 78082 15876 78092
rect 16044 78820 16100 78830
rect 15932 77924 15988 77934
rect 15932 77830 15988 77868
rect 16044 77250 16100 78764
rect 16156 78708 16212 80894
rect 16156 78642 16212 78652
rect 16044 77198 16046 77250
rect 16098 77198 16100 77250
rect 16044 77186 16100 77198
rect 15932 76466 15988 76478
rect 15932 76414 15934 76466
rect 15986 76414 15988 76466
rect 15820 74898 15876 74910
rect 15820 74846 15822 74898
rect 15874 74846 15876 74898
rect 15820 73330 15876 74846
rect 15820 73278 15822 73330
rect 15874 73278 15876 73330
rect 15820 72212 15876 73278
rect 15932 73332 15988 76414
rect 16156 75572 16212 75582
rect 16044 74900 16100 74910
rect 16044 74338 16100 74844
rect 16044 74286 16046 74338
rect 16098 74286 16100 74338
rect 16044 74274 16100 74286
rect 15932 73266 15988 73276
rect 15820 72146 15876 72156
rect 15708 71586 15764 71596
rect 16044 71650 16100 71662
rect 16044 71598 16046 71650
rect 16098 71598 16100 71650
rect 15596 71540 15652 71550
rect 15596 71446 15652 71484
rect 15708 71316 15764 71326
rect 15708 69636 15764 71260
rect 16044 71202 16100 71598
rect 16044 71150 16046 71202
rect 16098 71150 16100 71202
rect 16044 71138 16100 71150
rect 15820 69972 15876 69982
rect 15820 69970 15988 69972
rect 15820 69918 15822 69970
rect 15874 69918 15988 69970
rect 15820 69916 15988 69918
rect 15820 69906 15876 69916
rect 15708 69580 15876 69636
rect 15708 69186 15764 69198
rect 15708 69134 15710 69186
rect 15762 69134 15764 69186
rect 15708 68626 15764 69134
rect 15708 68574 15710 68626
rect 15762 68574 15764 68626
rect 15708 68562 15764 68574
rect 15820 68066 15876 69580
rect 15820 68014 15822 68066
rect 15874 68014 15876 68066
rect 15820 68002 15876 68014
rect 15932 67172 15988 69916
rect 16156 68628 16212 75516
rect 16268 75124 16324 82572
rect 16492 82562 16548 82572
rect 16604 82516 16660 82526
rect 16604 79716 16660 82460
rect 16492 79660 16660 79716
rect 16380 79602 16436 79614
rect 16380 79550 16382 79602
rect 16434 79550 16436 79602
rect 16380 79044 16436 79550
rect 16380 78978 16436 78988
rect 16492 76916 16548 79660
rect 16716 79604 16772 83582
rect 16940 82852 16996 84476
rect 17052 84306 17108 85148
rect 17052 84254 17054 84306
rect 17106 84254 17108 84306
rect 17052 84242 17108 84254
rect 17052 83524 17108 83534
rect 17052 83430 17108 83468
rect 16940 82786 16996 82796
rect 16604 79492 16660 79502
rect 16604 79398 16660 79436
rect 16492 76850 16548 76860
rect 16716 78930 16772 79548
rect 16716 78878 16718 78930
rect 16770 78878 16772 78930
rect 16716 76692 16772 78878
rect 17052 78820 17108 78830
rect 17052 78726 17108 78764
rect 16268 75058 16324 75068
rect 16492 76636 16772 76692
rect 16828 78036 16884 78046
rect 16828 77250 16884 77980
rect 16828 77198 16830 77250
rect 16882 77198 16884 77250
rect 16492 76578 16548 76636
rect 16492 76526 16494 76578
rect 16546 76526 16548 76578
rect 16044 68626 16212 68628
rect 16044 68574 16158 68626
rect 16210 68574 16212 68626
rect 16044 68572 16212 68574
rect 16044 67396 16100 68572
rect 16156 68562 16212 68572
rect 16380 74452 16436 74462
rect 16268 68516 16324 68526
rect 16268 68422 16324 68460
rect 16156 67956 16212 67966
rect 16156 67862 16212 67900
rect 16044 67330 16100 67340
rect 16156 67732 16212 67742
rect 15932 67106 15988 67116
rect 15484 66994 15540 67004
rect 15820 67058 15876 67070
rect 15820 67006 15822 67058
rect 15874 67006 15876 67058
rect 15820 66498 15876 67006
rect 15820 66446 15822 66498
rect 15874 66446 15876 66498
rect 15820 66434 15876 66446
rect 16156 67058 16212 67676
rect 16156 67006 16158 67058
rect 16210 67006 16212 67058
rect 16156 65716 16212 67006
rect 16156 65650 16212 65660
rect 16268 66724 16324 66734
rect 15820 65604 15876 65614
rect 15820 65510 15876 65548
rect 16268 65378 16324 66668
rect 16268 65326 16270 65378
rect 16322 65326 16324 65378
rect 16268 65314 16324 65326
rect 15148 63362 15428 63364
rect 15148 63310 15150 63362
rect 15202 63310 15428 63362
rect 15148 63308 15428 63310
rect 15484 63812 15540 63822
rect 14588 62302 14590 62354
rect 14642 62302 14644 62354
rect 14588 62290 14644 62302
rect 14924 63138 14980 63150
rect 14924 63086 14926 63138
rect 14978 63086 14980 63138
rect 14924 61908 14980 63086
rect 15148 62468 15204 63308
rect 15260 63140 15316 63150
rect 15260 63046 15316 63084
rect 15148 62402 15204 62412
rect 15036 62354 15092 62366
rect 15036 62302 15038 62354
rect 15090 62302 15092 62354
rect 15036 62244 15092 62302
rect 15036 62178 15092 62188
rect 15260 62132 15316 62142
rect 15260 62038 15316 62076
rect 14924 61852 15428 61908
rect 15372 61682 15428 61852
rect 15372 61630 15374 61682
rect 15426 61630 15428 61682
rect 15372 61618 15428 61630
rect 14588 61572 14644 61582
rect 13804 61570 14644 61572
rect 13804 61518 14590 61570
rect 14642 61518 14644 61570
rect 13804 61516 14644 61518
rect 13692 60622 13694 60674
rect 13746 60622 13748 60674
rect 13692 60610 13748 60622
rect 13804 61124 13860 61134
rect 13580 60162 13636 60172
rect 13692 59220 13748 59230
rect 13692 58434 13748 59164
rect 13692 58382 13694 58434
rect 13746 58382 13748 58434
rect 13692 58370 13748 58382
rect 13580 57540 13636 57550
rect 13580 57446 13636 57484
rect 13244 57426 13300 57438
rect 13244 57374 13246 57426
rect 13298 57374 13300 57426
rect 13132 56868 13188 56878
rect 13132 56774 13188 56812
rect 12908 55860 12964 55870
rect 12908 55858 13076 55860
rect 12908 55806 12910 55858
rect 12962 55806 13076 55858
rect 12908 55804 13076 55806
rect 12908 55794 12964 55804
rect 13020 51380 13076 55804
rect 13132 52276 13188 52286
rect 13132 52162 13188 52220
rect 13132 52110 13134 52162
rect 13186 52110 13188 52162
rect 13132 52098 13188 52110
rect 13132 51380 13188 51390
rect 13020 51378 13188 51380
rect 13020 51326 13134 51378
rect 13186 51326 13188 51378
rect 13020 51324 13188 51326
rect 13132 51314 13188 51324
rect 12796 51268 12852 51278
rect 12796 51266 12964 51268
rect 12796 51214 12798 51266
rect 12850 51214 12964 51266
rect 12796 51212 12964 51214
rect 12796 51202 12852 51212
rect 12796 50708 12852 50718
rect 12796 50614 12852 50652
rect 12684 49410 12740 49420
rect 12796 50372 12852 50382
rect 12684 49252 12740 49262
rect 12684 49158 12740 49196
rect 11900 45220 11956 46060
rect 12012 45890 12068 45902
rect 12012 45838 12014 45890
rect 12066 45838 12068 45890
rect 12012 45332 12068 45838
rect 12124 45332 12180 45342
rect 12012 45330 12180 45332
rect 12012 45278 12126 45330
rect 12178 45278 12180 45330
rect 12012 45276 12180 45278
rect 12124 45266 12180 45276
rect 11900 45164 12068 45220
rect 11900 44322 11956 44334
rect 11900 44270 11902 44322
rect 11954 44270 11956 44322
rect 11900 43204 11956 44270
rect 11900 42420 11956 43148
rect 12012 42532 12068 45164
rect 12012 42466 12068 42476
rect 11900 42354 11956 42364
rect 11900 42084 11956 42094
rect 11900 41990 11956 42028
rect 11788 41906 11844 41916
rect 12012 41186 12068 41198
rect 12012 41134 12014 41186
rect 12066 41134 12068 41186
rect 10892 38722 10948 39228
rect 11116 39172 11172 39900
rect 11676 39890 11732 39900
rect 11788 40292 11844 40302
rect 10892 38670 10894 38722
rect 10946 38670 10948 38722
rect 10892 37380 10948 38670
rect 11004 39116 11172 39172
rect 11228 39618 11284 39630
rect 11228 39566 11230 39618
rect 11282 39566 11284 39618
rect 11004 38274 11060 39116
rect 11228 39060 11284 39566
rect 11676 39618 11732 39630
rect 11676 39566 11678 39618
rect 11730 39566 11732 39618
rect 11676 39508 11732 39566
rect 11676 39442 11732 39452
rect 11228 38994 11284 39004
rect 11004 38222 11006 38274
rect 11058 38222 11060 38274
rect 11004 38210 11060 38222
rect 11564 38948 11620 38958
rect 10892 37324 11284 37380
rect 10668 37212 10948 37268
rect 10668 37044 10724 37054
rect 10556 36988 10668 37044
rect 10668 36950 10724 36988
rect 10444 36866 10500 36876
rect 10780 36820 10836 36830
rect 10332 36484 10388 36494
rect 10668 36484 10724 36494
rect 10332 36390 10388 36428
rect 10556 36482 10724 36484
rect 10556 36430 10670 36482
rect 10722 36430 10724 36482
rect 10556 36428 10724 36430
rect 10220 35698 10276 35710
rect 10556 35700 10612 36428
rect 10668 36418 10724 36428
rect 10220 35646 10222 35698
rect 10274 35646 10276 35698
rect 10220 35476 10276 35646
rect 10220 35410 10276 35420
rect 10332 35698 10612 35700
rect 10332 35646 10558 35698
rect 10610 35646 10612 35698
rect 10332 35644 10612 35646
rect 10108 34860 10276 34916
rect 10108 34690 10164 34702
rect 10108 34638 10110 34690
rect 10162 34638 10164 34690
rect 9884 34066 9940 34076
rect 9996 34356 10052 34366
rect 9772 33966 9774 34018
rect 9826 33966 9828 34018
rect 9772 33954 9828 33966
rect 9996 33796 10052 34300
rect 9660 33394 9716 33404
rect 9772 33740 9996 33796
rect 9548 31838 9550 31890
rect 9602 31838 9604 31890
rect 9548 31668 9604 31838
rect 9548 31602 9604 31612
rect 9772 30548 9828 33740
rect 9996 33730 10052 33740
rect 10108 33348 10164 34638
rect 10108 33282 10164 33292
rect 9884 32788 9940 32798
rect 9884 32694 9940 32732
rect 9660 30492 9828 30548
rect 9884 32004 9940 32014
rect 9660 28980 9716 30492
rect 9772 30324 9828 30334
rect 9772 30210 9828 30268
rect 9772 30158 9774 30210
rect 9826 30158 9828 30210
rect 9772 30146 9828 30158
rect 9884 29876 9940 31948
rect 9604 28924 9716 28980
rect 9772 29820 9940 29876
rect 9996 31668 10052 31678
rect 9604 28756 9660 28924
rect 9548 28700 9660 28756
rect 9548 26516 9604 28700
rect 9772 28642 9828 29820
rect 9884 28756 9940 28766
rect 9884 28662 9940 28700
rect 9772 28590 9774 28642
rect 9826 28590 9828 28642
rect 9772 28308 9828 28590
rect 9772 28242 9828 28252
rect 9772 27746 9828 27758
rect 9772 27694 9774 27746
rect 9826 27694 9828 27746
rect 9772 27300 9828 27694
rect 9772 27234 9828 27244
rect 9884 27188 9940 27198
rect 9884 27094 9940 27132
rect 9772 27074 9828 27086
rect 9772 27022 9774 27074
rect 9826 27022 9828 27074
rect 9772 26758 9828 27022
rect 9772 26702 9940 26758
rect 9548 26460 9716 26516
rect 9548 26292 9604 26302
rect 9548 26198 9604 26236
rect 9660 25956 9716 26460
rect 9884 26292 9940 26702
rect 9884 26226 9940 26236
rect 9772 26068 9828 26078
rect 9772 25974 9828 26012
rect 9660 25844 9716 25900
rect 9660 25788 9828 25844
rect 9436 23102 9438 23154
rect 9490 23102 9492 23154
rect 9436 20804 9492 23102
rect 9436 20738 9492 20748
rect 9548 25618 9604 25630
rect 9548 25566 9550 25618
rect 9602 25566 9604 25618
rect 9548 25172 9604 25566
rect 9548 24276 9604 25116
rect 9548 20356 9604 24220
rect 9548 20290 9604 20300
rect 9660 20690 9716 20702
rect 9660 20638 9662 20690
rect 9714 20638 9716 20690
rect 9436 20132 9492 20142
rect 9660 20132 9716 20638
rect 9436 20018 9492 20076
rect 9436 19966 9438 20018
rect 9490 19966 9492 20018
rect 9436 19954 9492 19966
rect 9548 20076 9660 20132
rect 9324 19740 9492 19796
rect 9436 18900 9492 19740
rect 9548 19234 9604 20076
rect 9660 20066 9716 20076
rect 9660 19796 9716 19806
rect 9660 19702 9716 19740
rect 9548 19182 9550 19234
rect 9602 19182 9604 19234
rect 9548 19170 9604 19182
rect 9660 19012 9716 19022
rect 9436 18844 9604 18900
rect 9100 17276 9268 17332
rect 9436 18450 9492 18462
rect 9436 18398 9438 18450
rect 9490 18398 9492 18450
rect 7980 16044 8148 16100
rect 8204 16772 8260 16782
rect 7868 15316 7924 15326
rect 7756 15090 7812 15102
rect 7756 15038 7758 15090
rect 7810 15038 7812 15090
rect 7756 13972 7812 15038
rect 7756 13906 7812 13916
rect 7868 13970 7924 15260
rect 7980 14644 8036 16044
rect 8092 15092 8148 15102
rect 8092 14998 8148 15036
rect 7980 14532 8036 14588
rect 8092 14532 8148 14542
rect 7980 14530 8148 14532
rect 7980 14478 8094 14530
rect 8146 14478 8148 14530
rect 7980 14476 8148 14478
rect 8092 14466 8148 14476
rect 7868 13918 7870 13970
rect 7922 13918 7924 13970
rect 7868 13906 7924 13918
rect 7532 13682 7588 13692
rect 7868 13748 7924 13758
rect 6748 13636 6804 13646
rect 6748 13542 6804 13580
rect 6972 13300 7028 13310
rect 6748 12964 6804 12974
rect 6748 12870 6804 12908
rect 6748 11956 6804 11966
rect 6748 11862 6804 11900
rect 6636 11554 6692 11564
rect 6188 10220 6356 10276
rect 6076 9090 6132 9100
rect 6188 10052 6244 10062
rect 5964 9044 6020 9054
rect 5964 8950 6020 8988
rect 5964 8260 6020 8270
rect 5964 7362 6020 8204
rect 5964 7310 5966 7362
rect 6018 7310 6020 7362
rect 5964 7298 6020 7310
rect 6076 8258 6132 8270
rect 6076 8206 6078 8258
rect 6130 8206 6132 8258
rect 6076 7588 6132 8206
rect 5068 6638 5070 6690
rect 5122 6638 5124 6690
rect 5068 6580 5124 6638
rect 4844 6524 5124 6580
rect 5180 7196 5908 7252
rect 4464 5516 4728 5526
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4464 5450 4728 5460
rect 4844 5124 4900 6524
rect 4956 6244 5012 6254
rect 4956 5234 5012 6188
rect 5068 5908 5124 5918
rect 5068 5814 5124 5852
rect 4956 5182 4958 5234
rect 5010 5182 5012 5234
rect 4956 5170 5012 5182
rect 4844 5058 4900 5068
rect 4284 4510 4286 4562
rect 4338 4510 4340 4562
rect 4284 4498 4340 4510
rect 5180 4338 5236 7196
rect 5964 7028 6020 7038
rect 5852 6916 5908 6926
rect 5740 6804 5796 6814
rect 5292 5682 5348 5694
rect 5628 5684 5684 5694
rect 5292 5630 5294 5682
rect 5346 5630 5348 5682
rect 5292 5348 5348 5630
rect 5292 5282 5348 5292
rect 5404 5682 5684 5684
rect 5404 5630 5630 5682
rect 5682 5630 5684 5682
rect 5404 5628 5684 5630
rect 5404 5346 5460 5628
rect 5628 5618 5684 5628
rect 5404 5294 5406 5346
rect 5458 5294 5460 5346
rect 5404 5282 5460 5294
rect 5180 4286 5182 4338
rect 5234 4286 5236 4338
rect 5180 4274 5236 4286
rect 5628 5124 5684 5134
rect 5740 5124 5796 6748
rect 5852 5236 5908 6860
rect 5964 5794 6020 6972
rect 6076 6690 6132 7532
rect 6076 6638 6078 6690
rect 6130 6638 6132 6690
rect 6076 5908 6132 6638
rect 6076 5842 6132 5852
rect 5964 5742 5966 5794
rect 6018 5742 6020 5794
rect 5964 5730 6020 5742
rect 5852 5170 5908 5180
rect 6076 5684 6132 5694
rect 5628 5122 5796 5124
rect 5628 5070 5630 5122
rect 5682 5070 5796 5122
rect 5628 5068 5796 5070
rect 6076 5122 6132 5628
rect 6076 5070 6078 5122
rect 6130 5070 6132 5122
rect 5404 4228 5460 4238
rect 5404 4134 5460 4172
rect 4956 4004 5012 4014
rect 4464 3948 4728 3958
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4464 3882 4728 3892
rect 4956 3666 5012 3948
rect 5404 3780 5460 3790
rect 5404 3686 5460 3724
rect 4956 3614 4958 3666
rect 5010 3614 5012 3666
rect 4956 3602 5012 3614
rect 4172 3502 4174 3554
rect 4226 3502 4228 3554
rect 4172 3490 4228 3502
rect 5628 3554 5684 5068
rect 6076 5058 6132 5070
rect 6076 4228 6132 4238
rect 6188 4228 6244 9996
rect 6076 4226 6244 4228
rect 6076 4174 6078 4226
rect 6130 4174 6244 4226
rect 6076 4172 6244 4174
rect 6076 4162 6132 4172
rect 5740 4116 5796 4126
rect 5740 4022 5796 4060
rect 5628 3502 5630 3554
rect 5682 3502 5684 3554
rect 5628 3490 5684 3502
rect 6076 3892 6132 3902
rect 6076 3554 6132 3836
rect 6300 3780 6356 10220
rect 6524 9826 6580 11340
rect 6524 9774 6526 9826
rect 6578 9774 6580 9826
rect 6524 9762 6580 9774
rect 6636 10164 6692 10174
rect 6412 8930 6468 8942
rect 6412 8878 6414 8930
rect 6466 8878 6468 8930
rect 6412 7700 6468 8878
rect 6636 8820 6692 10108
rect 6972 9940 7028 13244
rect 7084 12962 7140 12974
rect 7084 12910 7086 12962
rect 7138 12910 7140 12962
rect 7084 10724 7140 12910
rect 7196 12964 7252 12974
rect 7196 10834 7252 12908
rect 7868 12402 7924 13692
rect 8092 12964 8148 12974
rect 8092 12870 8148 12908
rect 7868 12350 7870 12402
rect 7922 12350 7924 12402
rect 7868 12338 7924 12350
rect 7308 11620 7364 11630
rect 7308 11526 7364 11564
rect 7756 11508 7812 11518
rect 7756 11414 7812 11452
rect 8092 11394 8148 11406
rect 8092 11342 8094 11394
rect 8146 11342 8148 11394
rect 7196 10782 7198 10834
rect 7250 10782 7252 10834
rect 7196 10770 7252 10782
rect 7308 10836 7364 10846
rect 7084 10658 7140 10668
rect 7084 9940 7140 9950
rect 6972 9938 7140 9940
rect 6972 9886 7086 9938
rect 7138 9886 7140 9938
rect 6972 9884 7140 9886
rect 6412 7634 6468 7644
rect 6524 8764 6692 8820
rect 6860 9042 6916 9054
rect 6860 8990 6862 9042
rect 6914 8990 6916 9042
rect 6300 3714 6356 3724
rect 6412 5572 6468 5582
rect 6412 5234 6468 5516
rect 6412 5182 6414 5234
rect 6466 5182 6468 5234
rect 6412 3666 6468 5182
rect 6524 4228 6580 8764
rect 6636 8370 6692 8382
rect 6636 8318 6638 8370
rect 6690 8318 6692 8370
rect 6636 8148 6692 8318
rect 6636 8082 6692 8092
rect 6748 7700 6804 7710
rect 6748 7586 6804 7644
rect 6748 7534 6750 7586
rect 6802 7534 6804 7586
rect 6748 7522 6804 7534
rect 6636 7476 6692 7486
rect 6636 6914 6692 7420
rect 6636 6862 6638 6914
rect 6690 6862 6692 6914
rect 6636 6850 6692 6862
rect 6524 4162 6580 4172
rect 6636 6580 6692 6590
rect 6412 3614 6414 3666
rect 6466 3614 6468 3666
rect 6412 3602 6468 3614
rect 6076 3502 6078 3554
rect 6130 3502 6132 3554
rect 6076 3490 6132 3502
rect 6076 3332 6132 3342
rect 3804 3164 4068 3174
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 3804 3098 4068 3108
rect 4172 3108 4228 3118
rect 3836 2772 3892 2782
rect 3836 2678 3892 2716
rect 4172 2658 4228 3052
rect 4172 2606 4174 2658
rect 4226 2606 4228 2658
rect 4172 2594 4228 2606
rect 5292 2770 5348 2782
rect 5292 2718 5294 2770
rect 5346 2718 5348 2770
rect 5292 2436 5348 2718
rect 5740 2660 5796 2670
rect 5740 2566 5796 2604
rect 4464 2380 4728 2390
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 5292 2370 5348 2380
rect 5628 2436 5684 2446
rect 4464 2314 4728 2324
rect 4956 2212 5012 2222
rect 4956 2118 5012 2156
rect 3836 2098 3892 2110
rect 3836 2046 3838 2098
rect 3890 2046 3892 2098
rect 3836 1876 3892 2046
rect 5628 2100 5684 2380
rect 6076 2210 6132 3276
rect 6636 2660 6692 6524
rect 6748 5236 6804 5246
rect 6748 5142 6804 5180
rect 6860 2994 6916 8990
rect 6972 8258 7028 8270
rect 6972 8206 6974 8258
rect 7026 8206 7028 8258
rect 6972 7028 7028 8206
rect 6972 6962 7028 6972
rect 7084 6916 7140 9884
rect 7308 9042 7364 10780
rect 7644 10612 7700 10622
rect 7644 10498 7700 10556
rect 7644 10446 7646 10498
rect 7698 10446 7700 10498
rect 7644 10434 7700 10446
rect 7980 10388 8036 10398
rect 7980 10294 8036 10332
rect 7308 8990 7310 9042
rect 7362 8990 7364 9042
rect 7308 8596 7364 8990
rect 7532 10276 7588 10286
rect 7420 8820 7476 8830
rect 7420 8726 7476 8764
rect 7308 8540 7476 8596
rect 7308 8372 7364 8382
rect 7308 8278 7364 8316
rect 7196 7474 7252 7486
rect 7196 7422 7198 7474
rect 7250 7422 7252 7474
rect 7196 7028 7252 7422
rect 7420 7476 7476 8540
rect 7420 7410 7476 7420
rect 7196 6972 7476 7028
rect 7084 6860 7252 6916
rect 6972 6804 7028 6814
rect 6972 6690 7028 6748
rect 6972 6638 6974 6690
rect 7026 6638 7028 6690
rect 6972 6626 7028 6638
rect 6972 5908 7028 5918
rect 6972 4338 7028 5852
rect 7084 5348 7140 5358
rect 7084 5254 7140 5292
rect 6972 4286 6974 4338
rect 7026 4286 7028 4338
rect 6972 4274 7028 4286
rect 6860 2942 6862 2994
rect 6914 2942 6916 2994
rect 6860 2930 6916 2942
rect 6972 4116 7028 4126
rect 6972 2772 7028 4060
rect 7196 3332 7252 6860
rect 7308 6804 7364 6814
rect 7308 6710 7364 6748
rect 7308 5236 7364 5246
rect 7308 3778 7364 5180
rect 7308 3726 7310 3778
rect 7362 3726 7364 3778
rect 7308 3714 7364 3726
rect 7196 3266 7252 3276
rect 6076 2158 6078 2210
rect 6130 2158 6132 2210
rect 6076 2146 6132 2158
rect 6188 2604 6692 2660
rect 6860 2716 7028 2772
rect 5628 1986 5684 2044
rect 5628 1934 5630 1986
rect 5682 1934 5684 1986
rect 5628 1922 5684 1934
rect 6188 1876 6244 2604
rect 3836 1810 3892 1820
rect 5964 1820 6244 1876
rect 6412 2436 6468 2446
rect 3804 1596 4068 1606
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 3804 1530 4068 1540
rect 3612 1372 3892 1428
rect 3388 1362 3444 1372
rect 3836 1202 3892 1372
rect 5628 1316 5684 1326
rect 3836 1150 3838 1202
rect 3890 1150 3892 1202
rect 3836 1138 3892 1150
rect 4172 1204 4228 1214
rect 2268 1038 2270 1090
rect 2322 1038 2324 1090
rect 2268 1026 2324 1038
rect 4172 1090 4228 1148
rect 5628 1202 5684 1260
rect 5628 1150 5630 1202
rect 5682 1150 5684 1202
rect 5628 1138 5684 1150
rect 4172 1038 4174 1090
rect 4226 1038 4228 1090
rect 4172 1026 4228 1038
rect 4844 1092 4900 1102
rect 4844 998 4900 1036
rect 5180 978 5236 990
rect 5180 926 5182 978
rect 5234 926 5236 978
rect 4464 812 4728 822
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4464 746 4728 756
rect 5180 756 5236 926
rect 5180 690 5236 700
rect 5628 980 5684 990
rect 1596 242 1652 252
rect 5404 420 5460 430
rect 5404 112 5460 364
rect 5628 112 5684 924
rect 5852 978 5908 990
rect 5852 926 5854 978
rect 5906 926 5908 978
rect 5852 868 5908 926
rect 5852 802 5908 812
rect 5964 644 6020 1820
rect 5852 588 6020 644
rect 6076 1652 6132 1662
rect 5852 112 5908 588
rect 6076 112 6132 1596
rect 6300 1540 6356 1550
rect 6300 112 6356 1484
rect 6412 1314 6468 2380
rect 6412 1262 6414 1314
rect 6466 1262 6468 1314
rect 6412 1250 6468 1262
rect 6524 1652 6580 1662
rect 6524 112 6580 1596
rect 6748 1652 6804 1662
rect 6748 112 6804 1596
rect 6860 1090 6916 2716
rect 7196 2212 7252 2222
rect 7420 2212 7476 6972
rect 7532 3780 7588 10220
rect 7868 8932 7924 8942
rect 7868 8838 7924 8876
rect 8092 8708 8148 11342
rect 8204 11060 8260 16716
rect 8316 16098 8372 16110
rect 8316 16046 8318 16098
rect 8370 16046 8372 16098
rect 8316 15204 8372 16046
rect 8988 16100 9044 16110
rect 8988 16006 9044 16044
rect 9100 15876 9156 17276
rect 8988 15820 9156 15876
rect 9212 17108 9268 17118
rect 8764 15316 8820 15326
rect 8764 15222 8820 15260
rect 8316 15138 8372 15148
rect 8428 15202 8484 15214
rect 8428 15150 8430 15202
rect 8482 15150 8484 15202
rect 8428 14868 8484 15150
rect 8316 13860 8372 13870
rect 8428 13860 8484 14812
rect 8988 14756 9044 15820
rect 9212 15764 9268 17052
rect 9436 17106 9492 18398
rect 9548 17890 9604 18844
rect 9548 17838 9550 17890
rect 9602 17838 9604 17890
rect 9548 17826 9604 17838
rect 9436 17054 9438 17106
rect 9490 17054 9492 17106
rect 9436 17042 9492 17054
rect 9548 16324 9604 16334
rect 9660 16324 9716 18956
rect 9548 16322 9716 16324
rect 9548 16270 9550 16322
rect 9602 16270 9716 16322
rect 9548 16268 9716 16270
rect 9100 15708 9268 15764
rect 9324 15764 9380 15774
rect 9100 15148 9156 15708
rect 9324 15314 9380 15708
rect 9324 15262 9326 15314
rect 9378 15262 9380 15314
rect 9324 15250 9380 15262
rect 9436 15204 9492 15242
rect 9100 15092 9268 15148
rect 9436 15138 9492 15148
rect 8988 14690 9044 14700
rect 8316 13858 8484 13860
rect 8316 13806 8318 13858
rect 8370 13806 8484 13858
rect 8316 13804 8484 13806
rect 8876 14642 8932 14654
rect 8876 14590 8878 14642
rect 8930 14590 8932 14642
rect 8316 13794 8372 13804
rect 8652 13748 8708 13758
rect 8652 13654 8708 13692
rect 8540 13636 8596 13646
rect 8428 12852 8484 12862
rect 8428 12180 8484 12796
rect 8428 12086 8484 12124
rect 8204 10994 8260 11004
rect 8428 10612 8484 10622
rect 8316 9828 8372 9838
rect 8204 9604 8260 9614
rect 8204 9510 8260 9548
rect 7868 8652 8148 8708
rect 7644 8372 7700 8382
rect 7644 8278 7700 8316
rect 7644 7477 7700 7514
rect 7644 7476 7646 7477
rect 7698 7476 7700 7477
rect 7644 7410 7700 7420
rect 7756 7250 7812 7262
rect 7756 7198 7758 7250
rect 7810 7198 7812 7250
rect 7644 6690 7700 6702
rect 7644 6638 7646 6690
rect 7698 6638 7700 6690
rect 7644 5796 7700 6638
rect 7644 5730 7700 5740
rect 7644 3780 7700 3790
rect 7532 3778 7700 3780
rect 7532 3726 7646 3778
rect 7698 3726 7700 3778
rect 7532 3724 7700 3726
rect 7644 3714 7700 3724
rect 7756 3388 7812 7198
rect 7868 6468 7924 8652
rect 8092 8484 8148 8494
rect 7980 8370 8036 8382
rect 7980 8318 7982 8370
rect 8034 8318 8036 8370
rect 7980 8036 8036 8318
rect 7980 7970 8036 7980
rect 7980 6692 8036 6702
rect 7980 6598 8036 6636
rect 8092 6468 8148 8428
rect 8204 8260 8260 8270
rect 8204 8166 8260 8204
rect 7868 6402 7924 6412
rect 7980 6412 8148 6468
rect 8204 7362 8260 7374
rect 8204 7310 8206 7362
rect 8258 7310 8260 7362
rect 7868 5908 7924 5918
rect 7868 5124 7924 5852
rect 7980 5346 8036 6412
rect 7980 5294 7982 5346
rect 8034 5294 8036 5346
rect 7980 5282 8036 5294
rect 8092 5348 8148 5358
rect 7868 4338 7924 5068
rect 7868 4286 7870 4338
rect 7922 4286 7924 4338
rect 7868 4274 7924 4286
rect 8092 3554 8148 5292
rect 8092 3502 8094 3554
rect 8146 3502 8148 3554
rect 8092 3490 8148 3502
rect 7532 3332 7812 3388
rect 7532 2548 7588 3332
rect 8204 3108 8260 7310
rect 8316 6914 8372 9772
rect 8316 6862 8318 6914
rect 8370 6862 8372 6914
rect 8316 6850 8372 6862
rect 8428 9042 8484 10556
rect 8428 8990 8430 9042
rect 8482 8990 8484 9042
rect 8428 8372 8484 8990
rect 8540 9044 8596 13580
rect 8876 13524 8932 14590
rect 9100 14532 9156 14542
rect 8876 13458 8932 13468
rect 8988 14530 9156 14532
rect 8988 14478 9102 14530
rect 9154 14478 9156 14530
rect 8988 14476 9156 14478
rect 8876 13188 8932 13198
rect 8876 13094 8932 13132
rect 8988 12180 9044 14476
rect 9100 14466 9156 14476
rect 9100 14196 9156 14206
rect 9100 13746 9156 14140
rect 9100 13694 9102 13746
rect 9154 13694 9156 13746
rect 9100 13682 9156 13694
rect 9212 13524 9268 15092
rect 9324 15092 9380 15102
rect 9324 13634 9380 15036
rect 9548 14868 9604 16268
rect 9324 13582 9326 13634
rect 9378 13582 9380 13634
rect 9324 13570 9380 13582
rect 9436 14812 9604 14868
rect 9660 15204 9716 15214
rect 8876 12124 9044 12180
rect 9100 13468 9268 13524
rect 8764 11956 8820 11966
rect 8764 11284 8820 11900
rect 8876 11732 8932 12124
rect 8988 11956 9044 11966
rect 8988 11862 9044 11900
rect 9100 11732 9156 13468
rect 9212 13074 9268 13086
rect 9212 13022 9214 13074
rect 9266 13022 9268 13074
rect 9212 12180 9268 13022
rect 9212 12114 9268 12124
rect 9436 12964 9492 14812
rect 9548 14642 9604 14654
rect 9548 14590 9550 14642
rect 9602 14590 9604 14642
rect 9548 14084 9604 14590
rect 9548 14018 9604 14028
rect 9436 11844 9492 12908
rect 9436 11778 9492 11788
rect 8876 11676 9044 11732
rect 9100 11676 9268 11732
rect 8764 11218 8820 11228
rect 8876 11506 8932 11518
rect 8876 11454 8878 11506
rect 8930 11454 8932 11506
rect 8764 10724 8820 10734
rect 8764 10610 8820 10668
rect 8764 10558 8766 10610
rect 8818 10558 8820 10610
rect 8764 10546 8820 10558
rect 8876 10164 8932 11454
rect 8764 10108 8932 10164
rect 8540 8988 8708 9044
rect 8428 6804 8484 8316
rect 8652 8708 8708 8988
rect 8652 8036 8708 8652
rect 8764 8596 8820 10108
rect 8876 9940 8932 9950
rect 8876 9846 8932 9884
rect 8988 9716 9044 11676
rect 9100 11394 9156 11406
rect 9100 11342 9102 11394
rect 9154 11342 9156 11394
rect 9100 10052 9156 11342
rect 9100 9986 9156 9996
rect 8764 8530 8820 8540
rect 8876 9660 9044 9716
rect 9100 9826 9156 9838
rect 9100 9774 9102 9826
rect 9154 9774 9156 9826
rect 8652 7970 8708 7980
rect 8876 7812 8932 9660
rect 8428 6738 8484 6748
rect 8540 7756 8932 7812
rect 8316 6692 8372 6702
rect 8316 5908 8372 6636
rect 8316 5842 8372 5852
rect 8428 5906 8484 5918
rect 8428 5854 8430 5906
rect 8482 5854 8484 5906
rect 8316 5234 8372 5246
rect 8316 5182 8318 5234
rect 8370 5182 8372 5234
rect 8316 5012 8372 5182
rect 8316 4946 8372 4956
rect 8316 3666 8372 3678
rect 8316 3614 8318 3666
rect 8370 3614 8372 3666
rect 8316 3444 8372 3614
rect 8316 3378 8372 3388
rect 7868 3052 8260 3108
rect 7756 2772 7812 2782
rect 7756 2678 7812 2716
rect 7532 2482 7588 2492
rect 7196 2210 7476 2212
rect 7196 2158 7198 2210
rect 7250 2158 7476 2210
rect 7196 2156 7476 2158
rect 7196 2146 7252 2156
rect 7644 2100 7700 2110
rect 7644 2006 7700 2044
rect 7868 1988 7924 3052
rect 7980 2884 8036 2894
rect 7980 2210 8036 2828
rect 7980 2158 7982 2210
rect 8034 2158 8036 2210
rect 7980 2146 8036 2158
rect 8092 2772 8148 2782
rect 7868 1932 8036 1988
rect 6860 1038 6862 1090
rect 6914 1038 6916 1090
rect 6860 1026 6916 1038
rect 6972 1652 7028 1662
rect 6972 112 7028 1596
rect 7420 1652 7476 1662
rect 7196 308 7252 318
rect 7196 112 7252 252
rect 7420 112 7476 1596
rect 7644 1652 7700 1662
rect 7644 112 7700 1596
rect 7868 1652 7924 1662
rect 7868 112 7924 1596
rect 7980 1426 8036 1932
rect 7980 1374 7982 1426
rect 8034 1374 8036 1426
rect 7980 1362 8036 1374
rect 8092 112 8148 2716
rect 8316 2324 8372 2334
rect 8316 2210 8372 2268
rect 8316 2158 8318 2210
rect 8370 2158 8372 2210
rect 8316 2146 8372 2158
rect 8428 2212 8484 5854
rect 8428 2146 8484 2156
rect 8540 1988 8596 7756
rect 9100 7700 9156 9774
rect 9212 7812 9268 11676
rect 9660 10836 9716 15148
rect 9772 13748 9828 25788
rect 9884 25620 9940 25630
rect 9884 22260 9940 25564
rect 9996 24500 10052 31612
rect 10220 30436 10276 34860
rect 10332 32788 10388 35644
rect 10556 35634 10612 35644
rect 10668 35924 10724 35934
rect 10332 32722 10388 32732
rect 10444 34130 10500 34142
rect 10444 34078 10446 34130
rect 10498 34078 10500 34130
rect 10444 31892 10500 34078
rect 10668 32116 10724 35868
rect 10780 34356 10836 36764
rect 10892 34804 10948 37212
rect 11004 36932 11060 36942
rect 11004 35308 11060 36876
rect 11116 36482 11172 36494
rect 11116 36430 11118 36482
rect 11170 36430 11172 36482
rect 11116 36372 11172 36430
rect 11116 36306 11172 36316
rect 11228 35924 11284 37324
rect 11564 36820 11620 38892
rect 11676 37940 11732 37950
rect 11676 37846 11732 37884
rect 11788 37268 11844 40236
rect 11564 36754 11620 36764
rect 11676 37212 11844 37268
rect 11900 39730 11956 39742
rect 11900 39678 11902 39730
rect 11954 39678 11956 39730
rect 11340 36596 11396 36606
rect 11340 36502 11396 36540
rect 11228 35858 11284 35868
rect 11564 36260 11620 36270
rect 11340 35698 11396 35710
rect 11340 35646 11342 35698
rect 11394 35646 11396 35698
rect 11228 35474 11284 35486
rect 11228 35422 11230 35474
rect 11282 35422 11284 35474
rect 11004 35252 11172 35308
rect 11116 35140 11172 35252
rect 10892 34802 11060 34804
rect 10892 34750 10894 34802
rect 10946 34750 11060 34802
rect 10892 34748 11060 34750
rect 10892 34738 10948 34748
rect 10780 34290 10836 34300
rect 10780 34132 10836 34142
rect 10780 34038 10836 34076
rect 11004 33012 11060 34748
rect 11116 34580 11172 35084
rect 11116 34514 11172 34524
rect 11228 33684 11284 35422
rect 11340 35364 11396 35646
rect 11340 35298 11396 35308
rect 11564 35364 11620 36204
rect 11564 35298 11620 35308
rect 11676 35140 11732 37212
rect 11788 37042 11844 37054
rect 11788 36990 11790 37042
rect 11842 36990 11844 37042
rect 11788 36594 11844 36990
rect 11788 36542 11790 36594
rect 11842 36542 11844 36594
rect 11788 35698 11844 36542
rect 11788 35646 11790 35698
rect 11842 35646 11844 35698
rect 11788 35634 11844 35646
rect 11452 35084 11732 35140
rect 11788 35364 11844 35374
rect 11340 35028 11396 35038
rect 11452 35028 11508 35084
rect 11340 35026 11508 35028
rect 11340 34974 11342 35026
rect 11394 34974 11508 35026
rect 11340 34972 11508 34974
rect 11340 34962 11396 34972
rect 11228 33618 11284 33628
rect 11228 33236 11284 33246
rect 11228 33234 11396 33236
rect 11228 33182 11230 33234
rect 11282 33182 11396 33234
rect 11228 33180 11396 33182
rect 11228 33170 11284 33180
rect 11004 32956 11284 33012
rect 10780 32788 10836 32798
rect 10780 32340 10836 32732
rect 10780 32274 10836 32284
rect 11004 32676 11060 32686
rect 11004 32450 11060 32620
rect 11004 32398 11006 32450
rect 11058 32398 11060 32450
rect 11004 32340 11060 32398
rect 11004 32274 11060 32284
rect 11116 32564 11172 32574
rect 10668 32060 10836 32116
rect 10668 31892 10724 31902
rect 10444 31890 10724 31892
rect 10444 31838 10670 31890
rect 10722 31838 10724 31890
rect 10444 31836 10724 31838
rect 10668 31826 10724 31836
rect 10444 30996 10500 31006
rect 10220 30434 10388 30436
rect 10220 30382 10222 30434
rect 10274 30382 10388 30434
rect 10220 30380 10388 30382
rect 10220 30370 10276 30380
rect 10108 28756 10164 28766
rect 10108 24948 10164 28700
rect 10220 28644 10276 28654
rect 10220 26908 10276 28588
rect 10332 28084 10388 30380
rect 10444 30324 10500 30940
rect 10444 30258 10500 30268
rect 10668 30772 10724 30782
rect 10556 29428 10612 29438
rect 10556 29334 10612 29372
rect 10332 28018 10388 28028
rect 10444 28642 10500 28654
rect 10444 28590 10446 28642
rect 10498 28590 10500 28642
rect 10332 27636 10388 27646
rect 10332 27186 10388 27580
rect 10332 27134 10334 27186
rect 10386 27134 10388 27186
rect 10332 27122 10388 27134
rect 10444 27076 10500 28590
rect 10556 27860 10612 27870
rect 10556 27766 10612 27804
rect 10444 27010 10500 27020
rect 10668 26908 10724 30716
rect 10780 30436 10836 32060
rect 11004 32004 11060 32014
rect 11004 30882 11060 31948
rect 11004 30830 11006 30882
rect 11058 30830 11060 30882
rect 11004 30772 11060 30830
rect 11004 30706 11060 30716
rect 10780 30370 10836 30380
rect 11004 29316 11060 29326
rect 11004 29222 11060 29260
rect 10892 28642 10948 28654
rect 10892 28590 10894 28642
rect 10946 28590 10948 28642
rect 10892 27860 10948 28590
rect 11116 28642 11172 32508
rect 11228 31668 11284 32956
rect 11340 32564 11396 33180
rect 11452 32788 11508 34972
rect 11788 34916 11844 35308
rect 11452 32722 11508 32732
rect 11564 34860 11844 34916
rect 11452 32564 11508 32574
rect 11340 32562 11508 32564
rect 11340 32510 11454 32562
rect 11506 32510 11508 32562
rect 11340 32508 11508 32510
rect 11228 31602 11284 31612
rect 11340 32340 11396 32350
rect 11340 30212 11396 32284
rect 11116 28590 11118 28642
rect 11170 28590 11172 28642
rect 11116 28578 11172 28590
rect 11228 30156 11396 30212
rect 11228 28420 11284 30156
rect 11340 29988 11396 29998
rect 11340 29894 11396 29932
rect 11340 29540 11396 29550
rect 11340 28532 11396 29484
rect 11452 29428 11508 32508
rect 11564 32004 11620 34860
rect 11900 34356 11956 39678
rect 12012 36484 12068 41134
rect 12236 41186 12292 46060
rect 12348 45890 12404 45902
rect 12348 45838 12350 45890
rect 12402 45838 12404 45890
rect 12348 45668 12404 45838
rect 12348 45602 12404 45612
rect 12348 42980 12404 42990
rect 12348 42754 12404 42924
rect 12348 42702 12350 42754
rect 12402 42702 12404 42754
rect 12348 42196 12404 42702
rect 12348 42130 12404 42140
rect 12236 41134 12238 41186
rect 12290 41134 12292 41186
rect 12236 41122 12292 41134
rect 12460 40068 12516 46956
rect 12572 48580 12628 48590
rect 12572 40292 12628 48524
rect 12684 47460 12740 47470
rect 12684 42980 12740 47404
rect 12796 46676 12852 50316
rect 12908 48916 12964 51212
rect 13244 51044 13300 57374
rect 13692 55188 13748 55198
rect 13804 55188 13860 61068
rect 14252 60676 14308 60686
rect 14252 60002 14308 60620
rect 14252 59950 14254 60002
rect 14306 59950 14308 60002
rect 14252 59938 14308 59950
rect 14028 58548 14084 58558
rect 14028 58454 14084 58492
rect 13916 58436 13972 58446
rect 13916 57538 13972 58380
rect 14476 58324 14532 61516
rect 14588 61506 14644 61516
rect 15036 61460 15092 61470
rect 14812 61012 14868 61022
rect 14812 60918 14868 60956
rect 14812 60788 14868 60798
rect 14812 60226 14868 60732
rect 14812 60174 14814 60226
rect 14866 60174 14868 60226
rect 14812 60162 14868 60174
rect 14812 59780 14868 59790
rect 14700 59220 14756 59230
rect 14700 59126 14756 59164
rect 14364 58268 14532 58324
rect 14588 58884 14644 58894
rect 13916 57486 13918 57538
rect 13970 57486 13972 57538
rect 13916 57474 13972 57486
rect 14028 58212 14084 58222
rect 14028 55972 14084 58156
rect 14252 57428 14308 57438
rect 14252 57334 14308 57372
rect 13692 55186 13860 55188
rect 13692 55134 13694 55186
rect 13746 55134 13860 55186
rect 13692 55132 13860 55134
rect 13916 55970 14084 55972
rect 13916 55918 14030 55970
rect 14082 55918 14084 55970
rect 13916 55916 14084 55918
rect 13692 52836 13748 55132
rect 13692 52770 13748 52780
rect 13916 52164 13972 55916
rect 14028 55906 14084 55916
rect 14140 56644 14196 56654
rect 14140 55410 14196 56588
rect 14140 55358 14142 55410
rect 14194 55358 14196 55410
rect 14140 55346 14196 55358
rect 14140 54740 14196 54750
rect 14140 54626 14196 54684
rect 14140 54574 14142 54626
rect 14194 54574 14196 54626
rect 14140 54404 14196 54574
rect 14140 54338 14196 54348
rect 14028 53620 14084 53630
rect 14028 52612 14084 53564
rect 14028 52546 14084 52556
rect 13244 50978 13300 50988
rect 13580 52108 13972 52164
rect 13580 50708 13636 52108
rect 13804 51940 13860 51950
rect 13804 51938 14308 51940
rect 13804 51886 13806 51938
rect 13858 51886 14308 51938
rect 13804 51884 14308 51886
rect 13804 51874 13860 51884
rect 13580 50642 13636 50652
rect 13692 51378 13748 51390
rect 13692 51326 13694 51378
rect 13746 51326 13748 51378
rect 13244 50594 13300 50606
rect 13244 50542 13246 50594
rect 13298 50542 13300 50594
rect 13244 50034 13300 50542
rect 13692 50596 13748 51326
rect 14252 51378 14308 51884
rect 14252 51326 14254 51378
rect 14306 51326 14308 51378
rect 14252 51314 14308 51326
rect 13804 51156 13860 51166
rect 14364 51156 14420 58268
rect 14588 57762 14644 58828
rect 14588 57710 14590 57762
rect 14642 57710 14644 57762
rect 14588 57698 14644 57710
rect 14476 56196 14532 56206
rect 14476 53172 14532 56140
rect 14588 55076 14644 55086
rect 14588 54514 14644 55020
rect 14588 54462 14590 54514
rect 14642 54462 14644 54514
rect 14588 54450 14644 54462
rect 14476 53116 14644 53172
rect 14476 52946 14532 52958
rect 14476 52894 14478 52946
rect 14530 52894 14532 52946
rect 14476 52836 14532 52894
rect 14476 52770 14532 52780
rect 13804 51154 14420 51156
rect 13804 51102 13806 51154
rect 13858 51102 14420 51154
rect 13804 51100 14420 51102
rect 14476 52612 14532 52622
rect 13804 51090 13860 51100
rect 14476 50932 14532 52556
rect 14252 50876 14532 50932
rect 14588 52052 14644 53116
rect 14588 50932 14644 51996
rect 13692 50428 13748 50540
rect 13804 50820 13860 50830
rect 13804 50594 13860 50764
rect 13804 50542 13806 50594
rect 13858 50542 13860 50594
rect 13804 50530 13860 50542
rect 14028 50594 14084 50606
rect 14028 50542 14030 50594
rect 14082 50542 14084 50594
rect 14028 50428 14084 50542
rect 13692 50372 13972 50428
rect 14028 50372 14196 50428
rect 13244 49982 13246 50034
rect 13298 49982 13300 50034
rect 13244 49970 13300 49982
rect 12908 48850 12964 48860
rect 13804 48804 13860 48814
rect 13356 48802 13860 48804
rect 13356 48750 13806 48802
rect 13858 48750 13860 48802
rect 13356 48748 13860 48750
rect 12908 48692 12964 48702
rect 12908 47236 12964 48636
rect 13356 48242 13412 48748
rect 13804 48738 13860 48748
rect 13356 48190 13358 48242
rect 13410 48190 13412 48242
rect 13356 48178 13412 48190
rect 13468 48242 13524 48254
rect 13468 48190 13470 48242
rect 13522 48190 13524 48242
rect 13020 48132 13076 48142
rect 13020 48038 13076 48076
rect 13244 48130 13300 48142
rect 13244 48078 13246 48130
rect 13298 48078 13300 48130
rect 13020 47460 13076 47470
rect 13244 47460 13300 48078
rect 13468 47570 13524 48190
rect 13580 48244 13636 48254
rect 13580 48150 13636 48188
rect 13804 48020 13860 48030
rect 13916 48020 13972 50372
rect 13804 48018 13972 48020
rect 13804 47966 13806 48018
rect 13858 47966 13972 48018
rect 13804 47964 13972 47966
rect 13804 47954 13860 47964
rect 13468 47518 13470 47570
rect 13522 47518 13524 47570
rect 13468 47506 13524 47518
rect 13020 47458 13300 47460
rect 13020 47406 13022 47458
rect 13074 47406 13300 47458
rect 13020 47404 13300 47406
rect 13020 47394 13076 47404
rect 13132 47236 13188 47246
rect 12908 47234 13188 47236
rect 12908 47182 13134 47234
rect 13186 47182 13188 47234
rect 12908 47180 13188 47182
rect 12908 46898 12964 47180
rect 13132 47170 13188 47180
rect 13356 47234 13412 47246
rect 13356 47182 13358 47234
rect 13410 47182 13412 47234
rect 12908 46846 12910 46898
rect 12962 46846 12964 46898
rect 12908 46834 12964 46846
rect 13356 47012 13412 47182
rect 12796 46620 13076 46676
rect 13020 44996 13076 46620
rect 13356 45890 13412 46956
rect 14028 46450 14084 46462
rect 14028 46398 14030 46450
rect 14082 46398 14084 46450
rect 14028 46340 14084 46398
rect 14028 46274 14084 46284
rect 13356 45838 13358 45890
rect 13410 45838 13412 45890
rect 13356 45826 13412 45838
rect 13468 45220 13524 45230
rect 13020 44940 13412 44996
rect 13020 44322 13076 44334
rect 13020 44270 13022 44322
rect 13074 44270 13076 44322
rect 13020 43652 13076 44270
rect 13020 43586 13076 43596
rect 12684 42914 12740 42924
rect 12908 42756 12964 42766
rect 12572 40226 12628 40236
rect 12684 41188 12740 41198
rect 12460 40012 12628 40068
rect 12348 39618 12404 39630
rect 12348 39566 12350 39618
rect 12402 39566 12404 39618
rect 12124 39060 12180 39070
rect 12348 39060 12404 39566
rect 12124 39058 12404 39060
rect 12124 39006 12126 39058
rect 12178 39006 12404 39058
rect 12124 39004 12404 39006
rect 12124 38994 12180 39004
rect 12572 38724 12628 40012
rect 12684 39620 12740 41132
rect 12684 39554 12740 39564
rect 12908 39618 12964 42700
rect 13132 42756 13188 42766
rect 13132 42754 13300 42756
rect 13132 42702 13134 42754
rect 13186 42702 13300 42754
rect 13132 42700 13300 42702
rect 13132 42690 13188 42700
rect 13020 41188 13076 41198
rect 13020 41094 13076 41132
rect 13244 40852 13300 42700
rect 13132 40796 13300 40852
rect 13020 40516 13076 40526
rect 13020 40422 13076 40460
rect 12908 39566 12910 39618
rect 12962 39566 12964 39618
rect 12908 39554 12964 39566
rect 12460 38668 12628 38724
rect 12012 36418 12068 36428
rect 12124 38276 12180 38286
rect 11788 34300 11956 34356
rect 12124 34580 12180 38220
rect 12236 37828 12292 37838
rect 12236 37380 12292 37772
rect 12236 37314 12292 37324
rect 12348 36482 12404 36494
rect 12348 36430 12350 36482
rect 12402 36430 12404 36482
rect 12236 35812 12292 35822
rect 12236 35718 12292 35756
rect 12348 35700 12404 36430
rect 12348 35634 12404 35644
rect 12460 35252 12516 38668
rect 11676 33458 11732 33470
rect 11676 33406 11678 33458
rect 11730 33406 11732 33458
rect 11676 32116 11732 33406
rect 11676 32050 11732 32060
rect 11564 31938 11620 31948
rect 11788 31892 11844 34300
rect 11900 34132 11956 34142
rect 11900 34038 11956 34076
rect 11788 31826 11844 31836
rect 11900 31890 11956 31902
rect 11900 31838 11902 31890
rect 11954 31838 11956 31890
rect 11900 31780 11956 31838
rect 11900 31714 11956 31724
rect 11564 31666 11620 31678
rect 11564 31614 11566 31666
rect 11618 31614 11620 31666
rect 11564 31444 11620 31614
rect 12124 31556 12180 34524
rect 12124 31490 12180 31500
rect 12348 35196 12516 35252
rect 12572 37380 12628 37390
rect 11564 30996 11620 31388
rect 11564 30930 11620 30940
rect 11676 30884 11732 30894
rect 11676 30212 11732 30828
rect 12124 30772 12180 30782
rect 12124 30770 12292 30772
rect 12124 30718 12126 30770
rect 12178 30718 12292 30770
rect 12124 30716 12292 30718
rect 12124 30706 12180 30716
rect 11788 30212 11844 30222
rect 11676 30210 11844 30212
rect 11676 30158 11790 30210
rect 11842 30158 11844 30210
rect 11676 30156 11844 30158
rect 11452 29362 11508 29372
rect 11788 28647 11844 30156
rect 12236 30210 12292 30716
rect 12236 30158 12238 30210
rect 12290 30158 12292 30210
rect 11788 28644 11790 28647
rect 11340 28466 11396 28476
rect 11452 28595 11790 28644
rect 11842 28595 11844 28647
rect 11452 28588 11844 28595
rect 10892 27794 10948 27804
rect 11116 28364 11284 28420
rect 10220 26852 10388 26908
rect 10108 24882 10164 24892
rect 10220 26628 10276 26638
rect 10108 24500 10164 24510
rect 9996 24498 10164 24500
rect 9996 24446 10110 24498
rect 10162 24446 10164 24498
rect 9996 24444 10164 24446
rect 9996 22484 10052 24444
rect 10108 24434 10164 24444
rect 10220 24276 10276 26572
rect 10332 26290 10388 26852
rect 10332 26238 10334 26290
rect 10386 26238 10388 26290
rect 10332 26226 10388 26238
rect 10444 26852 10724 26908
rect 10892 27076 10948 27086
rect 10108 24220 10276 24276
rect 10108 22820 10164 24220
rect 10444 24052 10500 26852
rect 10892 26290 10948 27020
rect 11116 26404 11172 28364
rect 11228 28084 11284 28094
rect 11228 26628 11284 28028
rect 11452 27858 11508 28588
rect 11788 28583 11844 28588
rect 12124 29202 12180 29214
rect 12124 29150 12126 29202
rect 12178 29150 12180 29202
rect 12124 28644 12180 29150
rect 12124 28578 12180 28588
rect 11452 27806 11454 27858
rect 11506 27806 11508 27858
rect 11452 27794 11508 27806
rect 11564 28084 11620 28094
rect 11228 26562 11284 26572
rect 11452 27524 11508 27534
rect 11564 27524 11620 28028
rect 11508 27468 11620 27524
rect 11900 27860 11956 27870
rect 11116 26348 11396 26404
rect 10892 26238 10894 26290
rect 10946 26238 10948 26290
rect 10892 26180 10948 26238
rect 10892 26124 11172 26180
rect 10556 25396 10612 25406
rect 10556 24834 10612 25340
rect 10556 24782 10558 24834
rect 10610 24782 10612 24834
rect 10556 24770 10612 24782
rect 10668 25282 10724 25294
rect 10668 25230 10670 25282
rect 10722 25230 10724 25282
rect 10332 23996 10500 24052
rect 10220 23154 10276 23166
rect 10220 23102 10222 23154
rect 10274 23102 10276 23154
rect 10220 23044 10276 23102
rect 10220 22978 10276 22988
rect 10108 22764 10276 22820
rect 9996 22418 10052 22428
rect 10108 22260 10164 22270
rect 9884 22258 10164 22260
rect 9884 22206 10110 22258
rect 10162 22206 10164 22258
rect 9884 22204 10164 22206
rect 10108 22036 10164 22204
rect 10108 21970 10164 21980
rect 9996 21140 10052 21150
rect 9996 20914 10052 21084
rect 9996 20862 9998 20914
rect 10050 20862 10052 20914
rect 9996 20850 10052 20862
rect 9884 20356 9940 20366
rect 9884 19012 9940 20300
rect 10108 20020 10164 20030
rect 10108 19926 10164 19964
rect 9996 19348 10052 19358
rect 9996 19254 10052 19292
rect 10220 19348 10276 22764
rect 10220 19282 10276 19292
rect 9884 18946 9940 18956
rect 10332 18564 10388 23996
rect 10444 23828 10500 23838
rect 10500 23772 10612 23828
rect 10444 23734 10500 23772
rect 10444 22482 10500 22494
rect 10444 22430 10446 22482
rect 10498 22430 10500 22482
rect 10444 22148 10500 22430
rect 10444 22082 10500 22092
rect 10556 20132 10612 23772
rect 10668 23156 10724 25230
rect 10892 24948 10948 24958
rect 10668 23090 10724 23100
rect 10780 24612 10836 24622
rect 10780 24050 10836 24556
rect 10780 23998 10782 24050
rect 10834 23998 10836 24050
rect 10556 19012 10612 20076
rect 10556 18946 10612 18956
rect 10668 20018 10724 20030
rect 10668 19966 10670 20018
rect 10722 19966 10724 20018
rect 10668 18676 10724 19966
rect 10668 18610 10724 18620
rect 10332 18498 10388 18508
rect 9884 18450 9940 18462
rect 9884 18398 9886 18450
rect 9938 18398 9940 18450
rect 9884 15988 9940 18398
rect 10668 18450 10724 18462
rect 10668 18398 10670 18450
rect 10722 18398 10724 18450
rect 9996 18228 10052 18238
rect 9996 18226 10612 18228
rect 9996 18174 9998 18226
rect 10050 18174 10612 18226
rect 9996 18172 10612 18174
rect 9996 18162 10052 18172
rect 9996 16884 10052 16894
rect 9996 16790 10052 16828
rect 9884 15148 9940 15932
rect 10108 15876 10164 15886
rect 10108 15314 10164 15820
rect 10108 15262 10110 15314
rect 10162 15262 10164 15314
rect 10108 15250 10164 15262
rect 10556 15148 10612 18172
rect 10668 17890 10724 18398
rect 10668 17838 10670 17890
rect 10722 17838 10724 17890
rect 10668 17826 10724 17838
rect 10668 15876 10724 15886
rect 10668 15782 10724 15820
rect 10668 15316 10724 15326
rect 10668 15222 10724 15260
rect 9884 15092 10052 15148
rect 9884 14532 9940 14542
rect 9884 14438 9940 14476
rect 9996 14308 10052 15092
rect 9772 13682 9828 13692
rect 9884 14252 10052 14308
rect 10220 15092 10612 15148
rect 9884 13524 9940 14252
rect 9996 13748 10052 13758
rect 9996 13746 10164 13748
rect 9996 13694 9998 13746
rect 10050 13694 10164 13746
rect 9996 13692 10164 13694
rect 9996 13682 10052 13692
rect 9996 13524 10052 13534
rect 9884 13468 9996 13524
rect 9884 11508 9940 11518
rect 9660 10780 9828 10836
rect 9436 10724 9492 10734
rect 9324 10052 9380 10062
rect 9324 9156 9380 9996
rect 9324 9090 9380 9100
rect 9436 9042 9492 10668
rect 9660 10612 9716 10622
rect 9660 10518 9716 10556
rect 9772 10388 9828 10780
rect 9660 10332 9828 10388
rect 9436 8990 9438 9042
rect 9490 8990 9492 9042
rect 9436 8596 9492 8990
rect 9436 8530 9492 8540
rect 9548 9938 9604 9950
rect 9548 9886 9550 9938
rect 9602 9886 9604 9938
rect 9548 8372 9604 9886
rect 9436 8316 9604 8372
rect 9212 7746 9268 7756
rect 9324 8260 9380 8270
rect 8876 7644 9156 7700
rect 8764 7476 8820 7486
rect 8652 7474 8820 7476
rect 8652 7422 8766 7474
rect 8818 7422 8820 7474
rect 8652 7420 8820 7422
rect 8652 6804 8708 7420
rect 8764 7410 8820 7420
rect 8876 7028 8932 7644
rect 9100 7476 9156 7486
rect 9156 7420 9268 7476
rect 9100 7410 9156 7420
rect 8652 6738 8708 6748
rect 8764 6972 8932 7028
rect 8652 4228 8708 4238
rect 8652 4134 8708 4172
rect 8652 2772 8708 2782
rect 8652 2678 8708 2716
rect 8540 1922 8596 1932
rect 8764 1876 8820 6972
rect 8876 6802 8932 6814
rect 8876 6750 8878 6802
rect 8930 6750 8932 6802
rect 8876 6132 8932 6750
rect 9100 6692 9156 6702
rect 8876 6066 8932 6076
rect 8988 6690 9156 6692
rect 8988 6638 9102 6690
rect 9154 6638 9156 6690
rect 8988 6636 9156 6638
rect 8988 3108 9044 6636
rect 9100 6626 9156 6636
rect 9212 5906 9268 7420
rect 9212 5854 9214 5906
rect 9266 5854 9268 5906
rect 9100 5796 9156 5806
rect 9100 5702 9156 5740
rect 9100 5460 9156 5470
rect 9100 5010 9156 5404
rect 9100 4958 9102 5010
rect 9154 4958 9156 5010
rect 9100 4946 9156 4958
rect 9100 4676 9156 4686
rect 9100 4226 9156 4620
rect 9212 4564 9268 5854
rect 9324 4676 9380 8204
rect 9436 6916 9492 8316
rect 9436 6850 9492 6860
rect 9548 8146 9604 8158
rect 9548 8094 9550 8146
rect 9602 8094 9604 8146
rect 9548 7588 9604 8094
rect 9548 5460 9604 7532
rect 9660 5906 9716 10332
rect 9772 9828 9828 9838
rect 9772 9734 9828 9772
rect 9772 8372 9828 8382
rect 9772 8036 9828 8316
rect 9772 7970 9828 7980
rect 9772 7476 9828 7486
rect 9772 7382 9828 7420
rect 9660 5854 9662 5906
rect 9714 5854 9716 5906
rect 9660 5842 9716 5854
rect 9772 6580 9828 6590
rect 9772 5684 9828 6524
rect 9324 4610 9380 4620
rect 9436 5404 9548 5460
rect 9212 4338 9268 4508
rect 9212 4286 9214 4338
rect 9266 4286 9268 4338
rect 9212 4274 9268 4286
rect 9100 4174 9102 4226
rect 9154 4174 9156 4226
rect 9100 4162 9156 4174
rect 9436 4116 9492 5404
rect 9548 5394 9604 5404
rect 9660 5628 9828 5684
rect 9660 5572 9716 5628
rect 9548 5234 9604 5246
rect 9548 5182 9550 5234
rect 9602 5182 9604 5234
rect 9548 5124 9604 5182
rect 9548 5058 9604 5068
rect 9212 4060 9492 4116
rect 9548 4116 9604 4126
rect 8988 3042 9044 3052
rect 9100 3780 9156 3790
rect 8652 1820 8820 1876
rect 8316 1652 8372 1662
rect 8316 112 8372 1596
rect 8540 1652 8596 1662
rect 8540 112 8596 1596
rect 8652 1204 8708 1820
rect 9100 1764 9156 3724
rect 9212 2996 9268 4060
rect 9324 3442 9380 3454
rect 9324 3390 9326 3442
rect 9378 3390 9380 3442
rect 9324 3332 9380 3390
rect 9324 3266 9380 3276
rect 9212 2930 9268 2940
rect 9436 3220 9492 3230
rect 9212 2772 9268 2782
rect 9212 2210 9268 2716
rect 9436 2770 9492 3164
rect 9436 2718 9438 2770
rect 9490 2718 9492 2770
rect 9436 2706 9492 2718
rect 9548 2548 9604 4060
rect 9660 2660 9716 5516
rect 9772 4788 9828 4798
rect 9772 4338 9828 4732
rect 9772 4286 9774 4338
rect 9826 4286 9828 4338
rect 9772 4274 9828 4286
rect 9772 3780 9828 3790
rect 9884 3780 9940 11452
rect 9996 10612 10052 13468
rect 10108 12402 10164 13692
rect 10108 12350 10110 12402
rect 10162 12350 10164 12402
rect 10108 12338 10164 12350
rect 9996 10546 10052 10556
rect 10108 11506 10164 11518
rect 10108 11454 10110 11506
rect 10162 11454 10164 11506
rect 9996 9828 10052 9838
rect 9996 8596 10052 9772
rect 10108 9492 10164 11454
rect 10108 9426 10164 9436
rect 9996 8540 10164 8596
rect 9996 8372 10052 8382
rect 9996 8278 10052 8316
rect 10108 8148 10164 8540
rect 10220 8484 10276 15092
rect 10444 14756 10500 14766
rect 10444 13972 10500 14700
rect 10332 13746 10388 13758
rect 10332 13694 10334 13746
rect 10386 13694 10388 13746
rect 10332 13524 10388 13694
rect 10332 13458 10388 13468
rect 10332 12852 10388 12862
rect 10332 12758 10388 12796
rect 10444 11620 10500 13916
rect 10668 13636 10724 13646
rect 10556 11954 10612 11966
rect 10556 11902 10558 11954
rect 10610 11902 10612 11954
rect 10556 11732 10612 11902
rect 10556 11666 10612 11676
rect 10444 11554 10500 11564
rect 10444 11396 10500 11406
rect 10444 11302 10500 11340
rect 10444 10498 10500 10510
rect 10444 10446 10446 10498
rect 10498 10446 10500 10498
rect 10332 10388 10388 10398
rect 10332 10050 10388 10332
rect 10332 9998 10334 10050
rect 10386 9998 10388 10050
rect 10332 9986 10388 9998
rect 10444 9492 10500 10446
rect 10668 10164 10724 13580
rect 10780 13300 10836 23998
rect 10892 23042 10948 24892
rect 11004 23156 11060 23166
rect 11004 23062 11060 23100
rect 10892 22990 10894 23042
rect 10946 22990 10948 23042
rect 10892 22978 10948 22990
rect 11116 22820 11172 26124
rect 10892 22764 11172 22820
rect 10892 14868 10948 22764
rect 11228 20804 11284 20814
rect 11228 20710 11284 20748
rect 11228 19348 11284 19358
rect 11116 19236 11172 19246
rect 11116 19142 11172 19180
rect 10892 14802 10948 14812
rect 11004 18450 11060 18462
rect 11004 18398 11006 18450
rect 11058 18398 11060 18450
rect 11004 14644 11060 18398
rect 11228 18004 11284 19292
rect 11340 19236 11396 26348
rect 11452 19348 11508 27468
rect 11676 27188 11732 27198
rect 11564 26292 11620 26302
rect 11564 25508 11620 26236
rect 11564 25442 11620 25452
rect 11676 23378 11732 27132
rect 11900 27074 11956 27804
rect 11900 27022 11902 27074
rect 11954 27022 11956 27074
rect 11900 26292 11956 27022
rect 11900 26198 11956 26236
rect 12124 26404 12180 26414
rect 11900 25844 11956 25854
rect 11900 25396 11956 25788
rect 11676 23326 11678 23378
rect 11730 23326 11732 23378
rect 11676 23314 11732 23326
rect 11788 25394 11956 25396
rect 11788 25342 11902 25394
rect 11954 25342 11956 25394
rect 11788 25340 11956 25342
rect 11564 22596 11620 22606
rect 11564 20916 11620 22540
rect 11676 22148 11732 22158
rect 11676 22054 11732 22092
rect 11676 20916 11732 20926
rect 11564 20914 11732 20916
rect 11564 20862 11678 20914
rect 11730 20862 11732 20914
rect 11564 20860 11732 20862
rect 11676 20850 11732 20860
rect 11676 20244 11732 20254
rect 11676 20018 11732 20188
rect 11676 19966 11678 20018
rect 11730 19966 11732 20018
rect 11676 19954 11732 19966
rect 11564 19348 11620 19358
rect 11452 19346 11620 19348
rect 11452 19294 11566 19346
rect 11618 19294 11620 19346
rect 11452 19292 11620 19294
rect 11340 19180 11508 19236
rect 11228 17938 11284 17948
rect 11340 19012 11396 19022
rect 11340 17666 11396 18956
rect 11340 17614 11342 17666
rect 11394 17614 11396 17666
rect 11340 17602 11396 17614
rect 11452 17780 11508 19180
rect 11564 17892 11620 19292
rect 11564 17826 11620 17836
rect 11676 18340 11732 18350
rect 11340 17332 11396 17342
rect 11116 16660 11172 16670
rect 11116 16566 11172 16604
rect 11228 16212 11284 16222
rect 11228 16118 11284 16156
rect 11340 15988 11396 17276
rect 11004 14578 11060 14588
rect 11116 15932 11396 15988
rect 11116 15652 11172 15932
rect 10780 13234 10836 13244
rect 10892 14418 10948 14430
rect 10892 14366 10894 14418
rect 10946 14366 10948 14418
rect 10668 10098 10724 10108
rect 10780 13074 10836 13086
rect 10780 13022 10782 13074
rect 10834 13022 10836 13074
rect 10780 11844 10836 13022
rect 10892 12852 10948 14366
rect 10892 12786 10948 12796
rect 10892 12068 10948 12078
rect 10892 11974 10948 12012
rect 10444 9426 10500 9436
rect 10668 9826 10724 9838
rect 10668 9774 10670 9826
rect 10722 9774 10724 9826
rect 10668 9156 10724 9774
rect 10668 9090 10724 9100
rect 10220 8418 10276 8428
rect 10556 9042 10612 9054
rect 10556 8990 10558 9042
rect 10610 8990 10612 9042
rect 9996 8092 10164 8148
rect 9996 6580 10052 8092
rect 10556 8036 10612 8990
rect 10780 8372 10836 11788
rect 11004 11396 11060 11406
rect 11116 11396 11172 15596
rect 11340 14644 11396 14654
rect 11452 14644 11508 17724
rect 11564 17332 11620 17342
rect 11564 16994 11620 17276
rect 11564 16942 11566 16994
rect 11618 16942 11620 16994
rect 11564 16930 11620 16942
rect 11564 16212 11620 16222
rect 11564 16118 11620 16156
rect 11564 15988 11620 15998
rect 11564 15314 11620 15932
rect 11564 15262 11566 15314
rect 11618 15262 11620 15314
rect 11564 15250 11620 15262
rect 11340 14642 11508 14644
rect 11340 14590 11342 14642
rect 11394 14590 11508 14642
rect 11340 14588 11508 14590
rect 11340 14578 11396 14588
rect 11340 14420 11396 14430
rect 11228 13748 11284 13758
rect 11228 12516 11284 13692
rect 11340 13746 11396 14364
rect 11340 13694 11342 13746
rect 11394 13694 11396 13746
rect 11340 13682 11396 13694
rect 11228 12460 11396 12516
rect 11228 12292 11284 12302
rect 11228 12178 11284 12236
rect 11228 12126 11230 12178
rect 11282 12126 11284 12178
rect 11228 12114 11284 12126
rect 11004 11394 11172 11396
rect 11004 11342 11006 11394
rect 11058 11342 11172 11394
rect 11004 11340 11172 11342
rect 11004 11330 11060 11340
rect 11004 11060 11060 11070
rect 11004 10836 11060 11004
rect 11004 10610 11060 10780
rect 11004 10558 11006 10610
rect 11058 10558 11060 10610
rect 11004 10546 11060 10558
rect 10892 10500 10948 10510
rect 10892 10406 10948 10444
rect 11116 9940 11172 11340
rect 10780 8306 10836 8316
rect 10892 9884 11172 9940
rect 11228 11620 11284 11630
rect 10892 8148 10948 9884
rect 11004 9714 11060 9726
rect 11004 9662 11006 9714
rect 11058 9662 11060 9714
rect 11004 9044 11060 9662
rect 11004 8978 11060 8988
rect 11004 8818 11060 8830
rect 11004 8766 11006 8818
rect 11058 8766 11060 8818
rect 11004 8484 11060 8766
rect 11004 8418 11060 8428
rect 11116 8596 11172 8606
rect 11116 8482 11172 8540
rect 11116 8430 11118 8482
rect 11170 8430 11172 8482
rect 11116 8418 11172 8430
rect 10892 8092 11060 8148
rect 10556 7980 10948 8036
rect 10220 7700 10276 7710
rect 10108 6692 10164 6702
rect 10108 6598 10164 6636
rect 9996 6514 10052 6524
rect 10108 6020 10164 6030
rect 10220 6020 10276 7644
rect 10556 7588 10612 7598
rect 10556 7494 10612 7532
rect 10780 7140 10836 7150
rect 10108 6018 10276 6020
rect 10108 5966 10110 6018
rect 10162 5966 10276 6018
rect 10108 5964 10276 5966
rect 10332 6802 10388 6814
rect 10332 6750 10334 6802
rect 10386 6750 10388 6802
rect 10332 6020 10388 6750
rect 9772 3778 9940 3780
rect 9772 3726 9774 3778
rect 9826 3726 9940 3778
rect 9772 3724 9940 3726
rect 9996 5572 10052 5582
rect 9772 3714 9828 3724
rect 9884 2660 9940 2670
rect 9660 2658 9940 2660
rect 9660 2606 9886 2658
rect 9938 2606 9940 2658
rect 9660 2604 9940 2606
rect 9884 2594 9940 2604
rect 9212 2158 9214 2210
rect 9266 2158 9268 2210
rect 9212 2146 9268 2158
rect 9324 2492 9604 2548
rect 9100 1708 9268 1764
rect 8652 1138 8708 1148
rect 8764 1652 8820 1662
rect 8764 112 8820 1596
rect 8988 1428 9044 1438
rect 8988 112 9044 1372
rect 9212 112 9268 1708
rect 9324 1202 9380 2492
rect 9996 2436 10052 5516
rect 10108 4450 10164 5964
rect 10332 5954 10388 5964
rect 10556 5684 10612 5694
rect 10556 5590 10612 5628
rect 10668 5460 10724 5470
rect 10668 5346 10724 5404
rect 10668 5294 10670 5346
rect 10722 5294 10724 5346
rect 10668 5282 10724 5294
rect 10780 5124 10836 7084
rect 10892 6580 10948 7980
rect 11004 7812 11060 8092
rect 11004 7588 11060 7756
rect 11004 7522 11060 7532
rect 11004 7252 11060 7262
rect 11228 7252 11284 11564
rect 11340 10052 11396 12460
rect 11452 11618 11508 14588
rect 11452 11566 11454 11618
rect 11506 11566 11508 11618
rect 11452 11554 11508 11566
rect 11564 11954 11620 11966
rect 11564 11902 11566 11954
rect 11618 11902 11620 11954
rect 11564 10836 11620 11902
rect 11564 10770 11620 10780
rect 11564 10612 11620 10622
rect 11564 10518 11620 10556
rect 11340 9996 11508 10052
rect 11340 9826 11396 9838
rect 11340 9774 11342 9826
rect 11394 9774 11396 9826
rect 11340 8596 11396 9774
rect 11340 8530 11396 8540
rect 11060 7196 11284 7252
rect 11004 7158 11060 7196
rect 11340 6916 11396 6926
rect 11452 6916 11508 9996
rect 11564 8146 11620 8158
rect 11564 8094 11566 8146
rect 11618 8094 11620 8146
rect 11564 7924 11620 8094
rect 11564 7858 11620 7868
rect 11340 6914 11452 6916
rect 11340 6862 11342 6914
rect 11394 6862 11452 6914
rect 11340 6860 11452 6862
rect 11340 6850 11396 6860
rect 11452 6822 11508 6860
rect 11676 6692 11732 18284
rect 11788 15876 11844 25340
rect 11900 25330 11956 25340
rect 12124 24164 12180 26348
rect 12236 25506 12292 30158
rect 12236 25454 12238 25506
rect 12290 25454 12292 25506
rect 12236 25442 12292 25454
rect 12124 24098 12180 24108
rect 12236 25172 12292 25182
rect 11900 24052 11956 24062
rect 11900 19460 11956 23996
rect 12012 23716 12068 23726
rect 12012 23714 12180 23716
rect 12012 23662 12014 23714
rect 12066 23662 12180 23714
rect 12012 23660 12180 23662
rect 12012 23650 12068 23660
rect 12012 23044 12068 23054
rect 12012 22950 12068 22988
rect 11900 19394 11956 19404
rect 12012 22484 12068 22494
rect 11900 19236 11956 19246
rect 11900 19142 11956 19180
rect 11900 18564 11956 18574
rect 11900 17890 11956 18508
rect 12012 18452 12068 22428
rect 12124 20802 12180 23660
rect 12124 20750 12126 20802
rect 12178 20750 12180 20802
rect 12124 20738 12180 20750
rect 12012 18358 12068 18396
rect 12124 20580 12180 20590
rect 11900 17838 11902 17890
rect 11954 17838 11956 17890
rect 11900 16324 11956 17838
rect 11900 16258 11956 16268
rect 12012 16100 12068 16110
rect 11788 15810 11844 15820
rect 11900 15986 11956 15998
rect 11900 15934 11902 15986
rect 11954 15934 11956 15986
rect 11788 15428 11844 15438
rect 11788 10164 11844 15372
rect 11900 14980 11956 15934
rect 11900 14914 11956 14924
rect 11900 14308 11956 14318
rect 11900 13634 11956 14252
rect 11900 13582 11902 13634
rect 11954 13582 11956 13634
rect 11900 13570 11956 13582
rect 11900 13188 11956 13198
rect 12012 13188 12068 16044
rect 12124 15428 12180 20524
rect 12236 19012 12292 25116
rect 12348 22484 12404 35196
rect 12460 35028 12516 35066
rect 12460 34962 12516 34972
rect 12460 34804 12516 34814
rect 12460 30100 12516 34748
rect 12572 30436 12628 37324
rect 12684 36596 12740 36606
rect 12684 32452 12740 36540
rect 12908 34804 12964 34814
rect 12908 34710 12964 34748
rect 12796 33908 12852 33918
rect 12796 33814 12852 33852
rect 12796 33124 12852 33134
rect 12796 33122 13076 33124
rect 12796 33070 12798 33122
rect 12850 33070 13076 33122
rect 12796 33068 13076 33070
rect 12796 33058 12852 33068
rect 13020 32562 13076 33068
rect 13020 32510 13022 32562
rect 13074 32510 13076 32562
rect 13020 32498 13076 32510
rect 12908 32452 12964 32462
rect 12684 32450 12964 32452
rect 12684 32398 12910 32450
rect 12962 32398 12964 32450
rect 12684 32396 12964 32398
rect 12908 32386 12964 32396
rect 13132 32340 13188 40796
rect 13244 38836 13300 38846
rect 13244 38274 13300 38780
rect 13244 38222 13246 38274
rect 13298 38222 13300 38274
rect 13244 38210 13300 38222
rect 13356 36482 13412 44940
rect 13468 42084 13524 45164
rect 13804 44996 13860 45006
rect 13468 42018 13524 42028
rect 13580 44994 13860 44996
rect 13580 44942 13806 44994
rect 13858 44942 13860 44994
rect 13580 44940 13860 44942
rect 13468 40292 13524 40302
rect 13468 40198 13524 40236
rect 13356 36430 13358 36482
rect 13410 36430 13412 36482
rect 13356 35252 13412 36430
rect 13468 39172 13524 39182
rect 13468 36484 13524 39116
rect 13580 38388 13636 44940
rect 13804 44930 13860 44940
rect 14028 43428 14084 43438
rect 14140 43428 14196 50372
rect 14252 44324 14308 50876
rect 14588 50866 14644 50876
rect 14700 52836 14756 52846
rect 14364 50708 14420 50718
rect 14700 50708 14756 52780
rect 14812 52388 14868 59724
rect 14924 59220 14980 59230
rect 14924 57428 14980 59164
rect 15036 59106 15092 61404
rect 15484 61348 15540 63756
rect 15820 63698 15876 63710
rect 15820 63646 15822 63698
rect 15874 63646 15876 63698
rect 15708 63028 15764 63038
rect 15708 62934 15764 62972
rect 15820 62354 15876 63646
rect 15820 62302 15822 62354
rect 15874 62302 15876 62354
rect 15820 62290 15876 62302
rect 15932 63250 15988 63262
rect 15932 63198 15934 63250
rect 15986 63198 15988 63250
rect 15932 63140 15988 63198
rect 15708 61794 15764 61806
rect 15708 61742 15710 61794
rect 15762 61742 15764 61794
rect 15596 61572 15652 61582
rect 15596 61478 15652 61516
rect 15484 61292 15652 61348
rect 15372 60786 15428 60798
rect 15372 60734 15374 60786
rect 15426 60734 15428 60786
rect 15372 59220 15428 60734
rect 15596 60676 15652 61292
rect 15596 60610 15652 60620
rect 15372 59154 15428 59164
rect 15036 59054 15038 59106
rect 15090 59054 15092 59106
rect 15036 59042 15092 59054
rect 15260 58212 15316 58222
rect 15036 58210 15316 58212
rect 15036 58158 15262 58210
rect 15314 58158 15316 58210
rect 15036 58156 15316 58158
rect 15036 57650 15092 58156
rect 15260 58146 15316 58156
rect 15036 57598 15038 57650
rect 15090 57598 15092 57650
rect 15036 57586 15092 57598
rect 15372 57876 15428 57886
rect 15372 57650 15428 57820
rect 15372 57598 15374 57650
rect 15426 57598 15428 57650
rect 15372 57586 15428 57598
rect 15596 57428 15652 57438
rect 14924 57372 15092 57428
rect 14924 54516 14980 54526
rect 14924 54422 14980 54460
rect 14924 53844 14980 53854
rect 14924 52834 14980 53788
rect 14924 52782 14926 52834
rect 14978 52782 14980 52834
rect 14924 52770 14980 52782
rect 14924 52388 14980 52398
rect 14812 52386 14980 52388
rect 14812 52334 14926 52386
rect 14978 52334 14980 52386
rect 14812 52332 14980 52334
rect 14812 51380 14868 51390
rect 14812 51286 14868 51324
rect 14924 51044 14980 52332
rect 14924 50978 14980 50988
rect 15036 50820 15092 57372
rect 15596 57334 15652 57372
rect 15260 55076 15316 55086
rect 15260 54982 15316 55020
rect 14364 49252 14420 50652
rect 14588 50652 14756 50708
rect 14924 50764 15092 50820
rect 15148 54290 15204 54302
rect 15148 54238 15150 54290
rect 15202 54238 15204 54290
rect 14476 50036 14532 50046
rect 14476 49698 14532 49980
rect 14476 49646 14478 49698
rect 14530 49646 14532 49698
rect 14476 49634 14532 49646
rect 14364 49186 14420 49196
rect 14588 48804 14644 50652
rect 14812 50596 14868 50634
rect 14812 50530 14868 50540
rect 14924 50428 14980 50764
rect 14476 48748 14644 48804
rect 14700 50372 14980 50428
rect 15036 50596 15092 50606
rect 14364 48244 14420 48254
rect 14476 48244 14532 48748
rect 14364 48242 14532 48244
rect 14364 48190 14366 48242
rect 14418 48190 14532 48242
rect 14364 48188 14532 48190
rect 14588 48580 14644 48590
rect 14364 47796 14420 48188
rect 14364 47346 14420 47740
rect 14364 47294 14366 47346
rect 14418 47294 14420 47346
rect 14364 46676 14420 47294
rect 14476 46676 14532 46686
rect 14364 46674 14532 46676
rect 14364 46622 14478 46674
rect 14530 46622 14532 46674
rect 14364 46620 14532 46622
rect 14364 46564 14420 46620
rect 14476 46610 14532 46620
rect 14364 46498 14420 46508
rect 14588 46340 14644 48524
rect 14588 46274 14644 46284
rect 14252 44258 14308 44268
rect 14364 45220 14420 45230
rect 14364 44322 14420 45164
rect 14364 44270 14366 44322
rect 14418 44270 14420 44322
rect 14364 44100 14420 44270
rect 14364 44034 14420 44044
rect 14476 43540 14532 43550
rect 14476 43446 14532 43484
rect 14084 43372 14196 43428
rect 14028 43334 14084 43372
rect 13916 42754 13972 42766
rect 14476 42756 14532 42766
rect 13916 42702 13918 42754
rect 13970 42702 13972 42754
rect 13916 42532 13972 42702
rect 13916 42466 13972 42476
rect 14028 42754 14532 42756
rect 14028 42702 14478 42754
rect 14530 42702 14532 42754
rect 14028 42700 14532 42702
rect 14028 42308 14084 42700
rect 14476 42690 14532 42700
rect 14588 42756 14644 42766
rect 13804 42252 14084 42308
rect 13804 42194 13860 42252
rect 13804 42142 13806 42194
rect 13858 42142 13860 42194
rect 13804 42130 13860 42142
rect 14476 41972 14532 41982
rect 14476 41186 14532 41916
rect 14476 41134 14478 41186
rect 14530 41134 14532 41186
rect 13804 40516 13860 40526
rect 13804 39396 13860 40460
rect 14476 40516 14532 41134
rect 14588 40626 14644 42700
rect 14588 40574 14590 40626
rect 14642 40574 14644 40626
rect 14588 40562 14644 40574
rect 14476 40450 14532 40460
rect 14700 39956 14756 50372
rect 14812 49810 14868 49822
rect 14812 49758 14814 49810
rect 14866 49758 14868 49810
rect 14812 49700 14868 49758
rect 14812 49634 14868 49644
rect 15036 48580 15092 50540
rect 15036 48514 15092 48524
rect 15148 49924 15204 54238
rect 15596 53842 15652 53854
rect 15596 53790 15598 53842
rect 15650 53790 15652 53842
rect 15260 53730 15316 53742
rect 15260 53678 15262 53730
rect 15314 53678 15316 53730
rect 15260 52948 15316 53678
rect 15596 53508 15652 53790
rect 15596 53442 15652 53452
rect 15260 52882 15316 52892
rect 15372 52052 15428 52062
rect 15372 51958 15428 51996
rect 15260 50932 15316 50942
rect 15260 50482 15316 50876
rect 15260 50430 15262 50482
rect 15314 50430 15316 50482
rect 15260 50148 15316 50430
rect 15708 50428 15764 61742
rect 15932 61796 15988 63084
rect 15932 61730 15988 61740
rect 16044 62914 16100 62926
rect 16044 62862 16046 62914
rect 16098 62862 16100 62914
rect 15820 61572 15876 61582
rect 15820 60228 15876 61516
rect 16044 61570 16100 62862
rect 16268 62692 16324 62702
rect 16268 62354 16324 62636
rect 16268 62302 16270 62354
rect 16322 62302 16324 62354
rect 16268 62290 16324 62302
rect 16044 61518 16046 61570
rect 16098 61518 16100 61570
rect 16044 61506 16100 61518
rect 16156 62132 16212 62142
rect 15932 61348 15988 61358
rect 15932 61254 15988 61292
rect 15932 60676 15988 60686
rect 15932 60582 15988 60620
rect 15932 60228 15988 60238
rect 15820 60226 15988 60228
rect 15820 60174 15934 60226
rect 15986 60174 15988 60226
rect 15820 60172 15988 60174
rect 15932 60162 15988 60172
rect 16156 55468 16212 62076
rect 16268 58994 16324 59006
rect 16268 58942 16270 58994
rect 16322 58942 16324 58994
rect 16268 57650 16324 58942
rect 16268 57598 16270 57650
rect 16322 57598 16324 57650
rect 16268 57586 16324 57598
rect 16156 55412 16324 55468
rect 15820 54516 15876 54526
rect 15820 54514 16100 54516
rect 15820 54462 15822 54514
rect 15874 54462 16100 54514
rect 15820 54460 16100 54462
rect 15820 54450 15876 54460
rect 16044 53170 16100 54460
rect 16156 54514 16212 54526
rect 16156 54462 16158 54514
rect 16210 54462 16212 54514
rect 16156 53620 16212 54462
rect 16156 53554 16212 53564
rect 16044 53118 16046 53170
rect 16098 53118 16100 53170
rect 16044 53106 16100 53118
rect 15596 50372 15764 50428
rect 15820 51378 15876 51390
rect 15820 51326 15822 51378
rect 15874 51326 15876 51378
rect 15820 50484 15876 51326
rect 15820 50418 15876 50428
rect 15260 50082 15316 50092
rect 15484 50260 15540 50270
rect 15036 48356 15092 48366
rect 14924 48244 14980 48254
rect 14812 48020 14868 48030
rect 14812 47926 14868 47964
rect 14812 47684 14868 47694
rect 14924 47684 14980 48188
rect 14812 47682 14980 47684
rect 14812 47630 14814 47682
rect 14866 47630 14980 47682
rect 14812 47628 14980 47630
rect 14812 47618 14868 47628
rect 15036 47572 15092 48300
rect 14924 47516 15092 47572
rect 14924 47460 14980 47516
rect 14812 46452 14868 46462
rect 14812 44546 14868 46396
rect 14812 44494 14814 44546
rect 14866 44494 14868 44546
rect 14812 44482 14868 44494
rect 14812 43538 14868 43550
rect 14812 43486 14814 43538
rect 14866 43486 14868 43538
rect 14812 43092 14868 43486
rect 14812 43026 14868 43036
rect 14812 41298 14868 41310
rect 14812 41246 14814 41298
rect 14866 41246 14868 41298
rect 14812 40964 14868 41246
rect 14812 40898 14868 40908
rect 14588 39900 14756 39956
rect 13916 39620 13972 39630
rect 13916 39526 13972 39564
rect 13804 39340 13972 39396
rect 13580 38322 13636 38332
rect 13692 38722 13748 38734
rect 13692 38670 13694 38722
rect 13746 38670 13748 38722
rect 13692 37156 13748 38670
rect 13916 37940 13972 39340
rect 14028 38836 14084 38846
rect 14028 38742 14084 38780
rect 14476 38834 14532 38846
rect 14476 38782 14478 38834
rect 14530 38782 14532 38834
rect 14252 38388 14308 38398
rect 14252 38162 14308 38332
rect 14252 38110 14254 38162
rect 14306 38110 14308 38162
rect 14252 38098 14308 38110
rect 13916 37846 13972 37884
rect 14364 37940 14420 37950
rect 14252 37156 14308 37166
rect 13692 37154 14308 37156
rect 13692 37102 14254 37154
rect 14306 37102 14308 37154
rect 13692 37100 14308 37102
rect 13580 36484 13636 36494
rect 13468 36428 13580 36484
rect 13468 35700 13524 35710
rect 13580 35700 13636 36428
rect 14252 36148 14308 37100
rect 14364 36708 14420 37884
rect 14476 37268 14532 38782
rect 14476 37202 14532 37212
rect 14364 36652 14532 36708
rect 14364 36484 14420 36494
rect 14364 36390 14420 36428
rect 14252 36082 14308 36092
rect 13468 35698 13636 35700
rect 13468 35646 13470 35698
rect 13522 35646 13636 35698
rect 13468 35644 13636 35646
rect 13468 35634 13524 35644
rect 13356 35196 13524 35252
rect 13244 35028 13300 35038
rect 13244 34914 13300 34972
rect 13244 34862 13246 34914
rect 13298 34862 13300 34914
rect 13244 34850 13300 34862
rect 13468 34692 13524 35196
rect 13020 32284 13188 32340
rect 13244 34636 13524 34692
rect 13020 31220 13076 32284
rect 13132 31556 13188 31566
rect 13132 31462 13188 31500
rect 13244 31332 13300 34636
rect 12908 31164 13076 31220
rect 13132 31276 13300 31332
rect 13356 32788 13412 32798
rect 12796 30884 12852 30894
rect 12572 30380 12740 30436
rect 12460 26908 12516 30044
rect 12572 30210 12628 30222
rect 12572 30158 12574 30210
rect 12626 30158 12628 30210
rect 12572 27076 12628 30158
rect 12684 27860 12740 30380
rect 12796 30434 12852 30828
rect 12796 30382 12798 30434
rect 12850 30382 12852 30434
rect 12796 30370 12852 30382
rect 12908 29204 12964 31164
rect 13020 30994 13076 31006
rect 13020 30942 13022 30994
rect 13074 30942 13076 30994
rect 13020 29428 13076 30942
rect 13020 29362 13076 29372
rect 12908 29148 13076 29204
rect 12684 27794 12740 27804
rect 12908 28530 12964 28542
rect 12908 28478 12910 28530
rect 12962 28478 12964 28530
rect 12572 27010 12628 27020
rect 12684 26964 12740 26974
rect 12460 26852 12628 26908
rect 12348 22418 12404 22428
rect 12460 26292 12516 26302
rect 12348 22258 12404 22270
rect 12348 22206 12350 22258
rect 12402 22206 12404 22258
rect 12348 22036 12404 22206
rect 12348 21970 12404 21980
rect 12460 21476 12516 26236
rect 12572 25284 12628 26852
rect 12684 25508 12740 26908
rect 12908 25844 12964 28478
rect 13020 27524 13076 29148
rect 13132 28420 13188 31276
rect 13356 30882 13412 32732
rect 13356 30830 13358 30882
rect 13410 30830 13412 30882
rect 13356 30818 13412 30830
rect 13468 30210 13524 30222
rect 13468 30158 13470 30210
rect 13522 30158 13524 30210
rect 13468 29988 13524 30158
rect 13244 28644 13300 28654
rect 13244 28550 13300 28588
rect 13132 28364 13300 28420
rect 13020 27468 13188 27524
rect 13020 27300 13076 27310
rect 13020 27074 13076 27244
rect 13020 27022 13022 27074
rect 13074 27022 13076 27074
rect 13020 27010 13076 27022
rect 13132 26908 13188 27468
rect 12908 25778 12964 25788
rect 13020 26852 13188 26908
rect 12908 25620 12964 25630
rect 12908 25526 12964 25564
rect 12796 25508 12852 25518
rect 12684 25506 12852 25508
rect 12684 25454 12798 25506
rect 12850 25454 12852 25506
rect 12684 25452 12852 25454
rect 12572 25218 12628 25228
rect 12684 24500 12740 24510
rect 12460 21410 12516 21420
rect 12572 24164 12628 24174
rect 12460 20802 12516 20814
rect 12460 20750 12462 20802
rect 12514 20750 12516 20802
rect 12460 19796 12516 20750
rect 12460 19730 12516 19740
rect 12348 19572 12404 19582
rect 12572 19572 12628 24108
rect 12684 21140 12740 24444
rect 12796 23492 12852 25452
rect 13020 25060 13076 26852
rect 12908 25004 13076 25060
rect 12908 24052 12964 25004
rect 13020 24836 13076 24846
rect 13020 24742 13076 24780
rect 12908 23986 12964 23996
rect 13244 23492 13300 28364
rect 13468 25506 13524 29932
rect 13580 29428 13636 35644
rect 13916 36036 13972 36046
rect 13916 35474 13972 35980
rect 13916 35422 13918 35474
rect 13970 35422 13972 35474
rect 13916 35410 13972 35422
rect 13916 35140 13972 35150
rect 14476 35140 14532 36652
rect 13916 35046 13972 35084
rect 14252 35084 14532 35140
rect 13804 34916 13860 34926
rect 13804 34822 13860 34860
rect 14140 34132 14196 34142
rect 13692 33684 13748 33694
rect 13692 32786 13748 33628
rect 13692 32734 13694 32786
rect 13746 32734 13748 32786
rect 13692 32722 13748 32734
rect 14140 33346 14196 34076
rect 14140 33294 14142 33346
rect 14194 33294 14196 33346
rect 14140 32564 14196 33294
rect 13692 32508 14196 32564
rect 14252 32564 14308 35084
rect 13692 31444 13748 32508
rect 14252 32498 14308 32508
rect 14364 34914 14420 34926
rect 14364 34862 14366 34914
rect 14418 34862 14420 34914
rect 14028 32340 14084 32350
rect 14028 32246 14084 32284
rect 13804 32004 13860 32014
rect 14364 32004 14420 34862
rect 14588 32788 14644 39900
rect 14700 38724 14756 38762
rect 14924 38668 14980 47404
rect 15148 45108 15204 49868
rect 15372 49700 15428 49710
rect 15372 49606 15428 49644
rect 15260 48916 15316 48926
rect 15260 45332 15316 48860
rect 15260 45266 15316 45276
rect 15148 45052 15316 45108
rect 15036 44882 15092 44894
rect 15036 44830 15038 44882
rect 15090 44830 15092 44882
rect 15036 43540 15092 44830
rect 15036 43474 15092 43484
rect 15036 43316 15092 43326
rect 15036 43222 15092 43260
rect 15036 42980 15092 42990
rect 15148 42980 15204 42990
rect 15092 42978 15204 42980
rect 15092 42926 15150 42978
rect 15202 42926 15204 42978
rect 15092 42924 15204 42926
rect 15036 42914 15092 42924
rect 15148 42914 15204 42924
rect 15260 42754 15316 45052
rect 15484 44660 15540 50204
rect 15260 42702 15262 42754
rect 15314 42702 15316 42754
rect 15260 42690 15316 42702
rect 15372 44604 15540 44660
rect 15372 42532 15428 44604
rect 15148 42476 15428 42532
rect 15484 43988 15540 43998
rect 14700 38658 14756 38668
rect 14812 38612 14980 38668
rect 15036 41858 15092 41870
rect 15036 41806 15038 41858
rect 15090 41806 15092 41858
rect 14700 37266 14756 37278
rect 14700 37214 14702 37266
rect 14754 37214 14756 37266
rect 14700 36036 14756 37214
rect 14700 35970 14756 35980
rect 14812 36594 14868 38612
rect 15036 38052 15092 41806
rect 15036 37986 15092 37996
rect 15036 37268 15092 37278
rect 15036 37174 15092 37212
rect 14812 36542 14814 36594
rect 14866 36542 14868 36594
rect 14812 35028 14868 36542
rect 15036 36036 15092 36046
rect 15036 35922 15092 35980
rect 15036 35870 15038 35922
rect 15090 35870 15092 35922
rect 15036 35858 15092 35870
rect 14812 34962 14868 34972
rect 14924 34914 14980 34926
rect 14924 34862 14926 34914
rect 14978 34862 14980 34914
rect 14924 34244 14980 34862
rect 14980 34188 15092 34244
rect 14924 34178 14980 34188
rect 14700 34132 14756 34142
rect 14700 34038 14756 34076
rect 14700 33460 14756 33470
rect 14700 33458 14868 33460
rect 14700 33406 14702 33458
rect 14754 33406 14868 33458
rect 14700 33404 14868 33406
rect 14700 33394 14756 33404
rect 14588 32732 14756 32788
rect 13804 32002 14420 32004
rect 13804 31950 13806 32002
rect 13858 31950 14420 32002
rect 13804 31948 14420 31950
rect 13804 31938 13860 31948
rect 13692 31378 13748 31388
rect 14588 30772 14644 30782
rect 14476 30770 14644 30772
rect 14476 30718 14590 30770
rect 14642 30718 14644 30770
rect 14476 30716 14644 30718
rect 13804 30212 13860 30222
rect 13580 29362 13636 29372
rect 13692 30210 13860 30212
rect 13692 30158 13806 30210
rect 13858 30158 13860 30210
rect 13692 30156 13860 30158
rect 13468 25454 13470 25506
rect 13522 25454 13524 25506
rect 13468 25442 13524 25454
rect 13580 27748 13636 27758
rect 13692 27748 13748 30156
rect 13804 30146 13860 30156
rect 14252 30212 14308 30222
rect 14028 29428 14084 29438
rect 13804 28868 13860 28878
rect 13804 28642 13860 28812
rect 13916 28756 13972 28766
rect 13916 28662 13972 28700
rect 13804 28590 13806 28642
rect 13858 28590 13860 28642
rect 13804 28578 13860 28590
rect 13636 27692 13748 27748
rect 13916 28308 13972 28318
rect 13356 24610 13412 24622
rect 13356 24558 13358 24610
rect 13410 24558 13412 24610
rect 13356 24388 13412 24558
rect 13356 24322 13412 24332
rect 12796 23426 12852 23436
rect 13020 23436 13300 23492
rect 13020 22708 13076 23436
rect 13244 23268 13300 23278
rect 13020 22642 13076 22652
rect 13132 23042 13188 23054
rect 13132 22990 13134 23042
rect 13186 22990 13188 23042
rect 13132 22596 13188 22990
rect 13244 23042 13300 23212
rect 13244 22990 13246 23042
rect 13298 22990 13300 23042
rect 13244 22978 13300 22990
rect 13468 22932 13524 22942
rect 13132 22530 13188 22540
rect 13356 22930 13524 22932
rect 13356 22878 13470 22930
rect 13522 22878 13524 22930
rect 13356 22876 13524 22878
rect 12796 22484 12852 22494
rect 12796 22482 13076 22484
rect 12796 22430 12798 22482
rect 12850 22430 13076 22482
rect 12796 22428 13076 22430
rect 12796 22418 12852 22428
rect 13020 22372 13076 22428
rect 13020 22316 13300 22372
rect 13132 22148 13188 22158
rect 12796 21812 12852 21822
rect 12796 21474 12852 21756
rect 13132 21586 13188 22092
rect 13244 21924 13300 22316
rect 13244 21858 13300 21868
rect 13132 21534 13134 21586
rect 13186 21534 13188 21586
rect 13132 21522 13188 21534
rect 13356 21588 13412 22876
rect 13468 22866 13524 22876
rect 13468 22708 13524 22718
rect 13468 22148 13524 22652
rect 13468 22082 13524 22092
rect 13580 21924 13636 27692
rect 13916 27074 13972 28252
rect 13916 27022 13918 27074
rect 13970 27022 13972 27074
rect 13916 27010 13972 27022
rect 13916 26852 13972 26862
rect 13916 26402 13972 26796
rect 13916 26350 13918 26402
rect 13970 26350 13972 26402
rect 13916 26338 13972 26350
rect 14028 26292 14084 29372
rect 14140 27746 14196 27758
rect 14140 27694 14142 27746
rect 14194 27694 14196 27746
rect 14140 27412 14196 27694
rect 14140 26908 14196 27356
rect 14252 27300 14308 30156
rect 14364 29428 14420 29438
rect 14364 29334 14420 29372
rect 14252 27234 14308 27244
rect 14364 28868 14420 28878
rect 14140 26852 14308 26908
rect 14084 26236 14196 26292
rect 14028 26226 14084 26236
rect 14028 26066 14084 26078
rect 14028 26014 14030 26066
rect 14082 26014 14084 26066
rect 13916 25844 13972 25854
rect 13916 25508 13972 25788
rect 14028 25732 14084 26014
rect 14028 25666 14084 25676
rect 13804 25506 13972 25508
rect 13804 25454 13918 25506
rect 13970 25454 13972 25506
rect 13804 25452 13972 25454
rect 13580 21858 13636 21868
rect 13692 23042 13748 23054
rect 13692 22990 13694 23042
rect 13746 22990 13748 23042
rect 13580 21588 13636 21598
rect 13356 21586 13636 21588
rect 13356 21534 13582 21586
rect 13634 21534 13636 21586
rect 13356 21532 13636 21534
rect 13580 21522 13636 21532
rect 12796 21422 12798 21474
rect 12850 21422 12852 21474
rect 12796 21252 12852 21422
rect 12796 21186 12852 21196
rect 13468 21252 13524 21262
rect 12684 21074 12740 21084
rect 12348 19234 12404 19516
rect 12348 19182 12350 19234
rect 12402 19182 12404 19234
rect 12348 19170 12404 19182
rect 12460 19516 12628 19572
rect 12684 20914 12740 20926
rect 12684 20862 12686 20914
rect 12738 20862 12740 20914
rect 12236 18956 12404 19012
rect 12236 16100 12292 16110
rect 12236 16006 12292 16044
rect 12348 15876 12404 18956
rect 12460 18676 12516 19516
rect 12572 19348 12628 19358
rect 12572 19254 12628 19292
rect 12460 18620 12628 18676
rect 12124 15362 12180 15372
rect 12236 15820 12404 15876
rect 12460 18452 12516 18462
rect 12236 15148 12292 15820
rect 12460 15764 12516 18396
rect 11900 13186 12068 13188
rect 11900 13134 11902 13186
rect 11954 13134 12068 13186
rect 11900 13132 12068 13134
rect 12124 15092 12292 15148
rect 12348 15708 12516 15764
rect 11900 13122 11956 13132
rect 12124 13076 12180 15092
rect 12236 13636 12292 13646
rect 12236 13542 12292 13580
rect 12348 13524 12404 15708
rect 12572 15540 12628 18620
rect 12684 15652 12740 20862
rect 13132 20804 13188 20814
rect 13132 20710 13188 20748
rect 13132 20020 13188 20030
rect 13020 19964 13132 20020
rect 13020 19124 13076 19964
rect 13132 19926 13188 19964
rect 13244 19348 13300 19358
rect 13020 18564 13076 19068
rect 13020 18470 13076 18508
rect 13132 19234 13188 19246
rect 13132 19182 13134 19234
rect 13186 19182 13188 19234
rect 13020 17892 13076 17902
rect 13132 17892 13188 19182
rect 13020 17890 13188 17892
rect 13020 17838 13022 17890
rect 13074 17838 13188 17890
rect 13020 17836 13188 17838
rect 13020 17826 13076 17836
rect 12908 17108 12964 17118
rect 12908 17014 12964 17052
rect 12908 16212 12964 16222
rect 12908 16118 12964 16156
rect 12796 16098 12852 16110
rect 12796 16046 12798 16098
rect 12850 16046 12852 16098
rect 12796 15876 12852 16046
rect 12796 15810 12852 15820
rect 12684 15596 13076 15652
rect 12572 15484 12852 15540
rect 12460 15428 12516 15438
rect 12460 14980 12516 15372
rect 12460 14914 12516 14924
rect 12572 15316 12628 15326
rect 12460 14756 12516 14766
rect 12460 14662 12516 14700
rect 12348 13458 12404 13468
rect 12460 14196 12516 14206
rect 12460 13300 12516 14140
rect 12012 13020 12180 13076
rect 12348 13244 12516 13300
rect 12012 12740 12068 13020
rect 11900 12628 11956 12638
rect 11900 12292 11956 12572
rect 11900 12226 11956 12236
rect 11900 11954 11956 11966
rect 11900 11902 11902 11954
rect 11954 11902 11956 11954
rect 11900 10948 11956 11902
rect 12012 11956 12068 12684
rect 12124 12180 12180 12190
rect 12124 12086 12180 12124
rect 12012 11890 12068 11900
rect 11900 10882 11956 10892
rect 12012 11396 12068 11406
rect 12348 11396 12404 13244
rect 12572 13188 12628 15260
rect 11900 10498 11956 10510
rect 11900 10446 11902 10498
rect 11954 10446 11956 10498
rect 11900 10388 11956 10446
rect 11900 10322 11956 10332
rect 11788 10108 11956 10164
rect 11788 9828 11844 9838
rect 11900 9828 11956 10108
rect 12012 10050 12068 11340
rect 12012 9998 12014 10050
rect 12066 9998 12068 10050
rect 12012 9986 12068 9998
rect 12124 11340 12404 11396
rect 12460 13132 12628 13188
rect 12684 14532 12740 14542
rect 12124 9828 12180 11340
rect 12348 11060 12404 11070
rect 11900 9772 12068 9828
rect 11788 9734 11844 9772
rect 11900 9604 11956 9614
rect 11900 8258 11956 9548
rect 11900 8206 11902 8258
rect 11954 8206 11956 8258
rect 11900 8194 11956 8206
rect 10892 6486 10948 6524
rect 11340 6636 11732 6692
rect 10892 5682 10948 5694
rect 11228 5684 11284 5694
rect 10892 5630 10894 5682
rect 10946 5630 10948 5682
rect 10892 5460 10948 5630
rect 10892 5394 10948 5404
rect 11004 5682 11284 5684
rect 11004 5630 11230 5682
rect 11282 5630 11284 5682
rect 11004 5628 11284 5630
rect 10108 4398 10110 4450
rect 10162 4398 10164 4450
rect 10108 4386 10164 4398
rect 10444 5068 10836 5124
rect 10108 2996 10164 3006
rect 10108 2772 10164 2940
rect 10108 2770 10276 2772
rect 10108 2718 10110 2770
rect 10162 2718 10276 2770
rect 10108 2716 10276 2718
rect 10108 2706 10164 2716
rect 9884 2380 10052 2436
rect 9548 2098 9604 2110
rect 9548 2046 9550 2098
rect 9602 2046 9604 2098
rect 9548 1764 9604 2046
rect 9548 1698 9604 1708
rect 9324 1150 9326 1202
rect 9378 1150 9380 1202
rect 9324 1138 9380 1150
rect 9660 1652 9716 1662
rect 9436 980 9492 990
rect 9436 112 9492 924
rect 9548 978 9604 990
rect 9548 926 9550 978
rect 9602 926 9604 978
rect 9548 420 9604 926
rect 9548 354 9604 364
rect 9660 112 9716 1596
rect 9884 112 9940 2380
rect 10220 2100 10276 2716
rect 10220 2034 10276 2044
rect 10444 2098 10500 5068
rect 10556 4340 10612 4350
rect 10556 4246 10612 4284
rect 10892 4228 10948 4238
rect 11004 4228 11060 5628
rect 11228 5618 11284 5628
rect 11228 5124 11284 5134
rect 11228 5030 11284 5068
rect 10892 4226 11060 4228
rect 10892 4174 10894 4226
rect 10946 4174 11060 4226
rect 10892 4172 11060 4174
rect 10892 4162 10948 4172
rect 11228 4116 11284 4126
rect 11228 4022 11284 4060
rect 10668 4004 10724 4014
rect 10556 2770 10612 2782
rect 10556 2718 10558 2770
rect 10610 2718 10612 2770
rect 10556 2436 10612 2718
rect 10556 2370 10612 2380
rect 10444 2046 10446 2098
rect 10498 2046 10500 2098
rect 10444 1988 10500 2046
rect 10444 1922 10500 1932
rect 10108 1876 10164 1914
rect 10108 1810 10164 1820
rect 10108 1652 10164 1662
rect 10108 112 10164 1596
rect 10332 1652 10388 1662
rect 10220 1202 10276 1214
rect 10220 1150 10222 1202
rect 10274 1150 10276 1202
rect 10220 1092 10276 1150
rect 10220 1026 10276 1036
rect 10332 112 10388 1596
rect 10668 1090 10724 3948
rect 10892 3780 10948 3790
rect 10892 3686 10948 3724
rect 11228 3556 11284 3566
rect 10892 3332 10948 3342
rect 10892 2882 10948 3276
rect 11228 2884 11284 3500
rect 11340 2996 11396 6636
rect 12012 5906 12068 9772
rect 12124 9762 12180 9772
rect 12236 10948 12292 10958
rect 12124 9044 12180 9054
rect 12124 8950 12180 8988
rect 12124 8372 12180 8382
rect 12124 7698 12180 8316
rect 12124 7646 12126 7698
rect 12178 7646 12180 7698
rect 12124 7634 12180 7646
rect 12236 7476 12292 10892
rect 12348 8258 12404 11004
rect 12460 10388 12516 13132
rect 12572 12852 12628 12862
rect 12572 12758 12628 12796
rect 12460 10164 12516 10332
rect 12460 10098 12516 10108
rect 12572 11170 12628 11182
rect 12572 11118 12574 11170
rect 12626 11118 12628 11170
rect 12572 9826 12628 11118
rect 12684 10500 12740 14476
rect 12796 12740 12852 15484
rect 12908 15204 12964 15242
rect 12908 15138 12964 15148
rect 12908 14980 12964 14990
rect 12908 14418 12964 14924
rect 12908 14366 12910 14418
rect 12962 14366 12964 14418
rect 12908 12852 12964 14366
rect 13020 13636 13076 15596
rect 13020 13570 13076 13580
rect 13020 13300 13076 13310
rect 13020 13186 13076 13244
rect 13020 13134 13022 13186
rect 13074 13134 13076 13186
rect 13020 13076 13076 13134
rect 13020 13010 13076 13020
rect 12908 12796 13188 12852
rect 12796 12684 13076 12740
rect 12796 12292 12852 12302
rect 12796 10948 12852 12236
rect 12796 10882 12852 10892
rect 12908 11954 12964 11966
rect 12908 11902 12910 11954
rect 12962 11902 12964 11954
rect 12908 10612 12964 11902
rect 12908 10546 12964 10556
rect 13020 10610 13076 12684
rect 13020 10558 13022 10610
rect 13074 10558 13076 10610
rect 13020 10546 13076 10558
rect 12796 10500 12852 10510
rect 12684 10498 12852 10500
rect 12684 10446 12798 10498
rect 12850 10446 12852 10498
rect 12684 10444 12852 10446
rect 12796 10434 12852 10444
rect 13020 9828 13076 9838
rect 12572 9774 12574 9826
rect 12626 9774 12628 9826
rect 12572 9762 12628 9774
rect 12908 9826 13076 9828
rect 12908 9774 13022 9826
rect 13074 9774 13076 9826
rect 12908 9772 13076 9774
rect 12572 9156 12628 9166
rect 12572 8370 12628 9100
rect 12572 8318 12574 8370
rect 12626 8318 12628 8370
rect 12572 8306 12628 8318
rect 12796 8818 12852 8830
rect 12796 8766 12798 8818
rect 12850 8766 12852 8818
rect 12348 8206 12350 8258
rect 12402 8206 12404 8258
rect 12348 8194 12404 8206
rect 12796 8260 12852 8766
rect 12796 8194 12852 8204
rect 12908 8036 12964 9772
rect 13020 9762 13076 9772
rect 13132 9604 13188 12796
rect 13020 9548 13188 9604
rect 13020 8932 13076 9548
rect 13020 8866 13076 8876
rect 13132 8820 13188 8830
rect 13132 8726 13188 8764
rect 13020 8372 13076 8382
rect 13020 8278 13076 8316
rect 12908 7970 12964 7980
rect 13244 7924 13300 19292
rect 13468 19012 13524 21196
rect 13692 21028 13748 22990
rect 13804 21812 13860 25452
rect 13916 25442 13972 25452
rect 14140 24836 14196 26236
rect 14252 25060 14308 26852
rect 14252 24994 14308 25004
rect 14140 23940 14196 24780
rect 14140 23874 14196 23884
rect 14364 23380 14420 28812
rect 14476 27858 14532 30716
rect 14588 30706 14644 30716
rect 14700 28980 14756 32732
rect 14812 31892 14868 33404
rect 14812 31826 14868 31836
rect 14924 32564 14980 32574
rect 14924 31890 14980 32508
rect 14924 31838 14926 31890
rect 14978 31838 14980 31890
rect 14812 30212 14868 30222
rect 14812 30118 14868 30156
rect 14812 29316 14868 29326
rect 14924 29316 14980 31838
rect 15036 30324 15092 34188
rect 15148 33124 15204 42476
rect 15372 42082 15428 42094
rect 15372 42030 15374 42082
rect 15426 42030 15428 42082
rect 15372 41972 15428 42030
rect 15372 41906 15428 41916
rect 15260 38836 15316 38846
rect 15260 37268 15316 38780
rect 15372 38834 15428 38846
rect 15372 38782 15374 38834
rect 15426 38782 15428 38834
rect 15372 38276 15428 38782
rect 15484 38500 15540 43932
rect 15484 38434 15540 38444
rect 15484 38276 15540 38286
rect 15372 38274 15540 38276
rect 15372 38222 15486 38274
rect 15538 38222 15540 38274
rect 15372 38220 15540 38222
rect 15484 38210 15540 38220
rect 15260 37212 15428 37268
rect 15260 37044 15316 37054
rect 15260 36950 15316 36988
rect 15260 33908 15316 33918
rect 15260 33814 15316 33852
rect 15148 33058 15204 33068
rect 15148 32788 15204 32798
rect 15148 32674 15204 32732
rect 15148 32622 15150 32674
rect 15202 32622 15204 32674
rect 15148 32452 15204 32622
rect 15148 32386 15204 32396
rect 15372 31892 15428 37212
rect 15596 33236 15652 50372
rect 15820 49810 15876 49822
rect 15820 49758 15822 49810
rect 15874 49758 15876 49810
rect 15820 48468 15876 49758
rect 16156 49812 16212 49822
rect 16156 49718 16212 49756
rect 16268 49700 16324 55412
rect 16380 54516 16436 74396
rect 16492 58884 16548 76526
rect 16828 76244 16884 77198
rect 17052 77810 17108 77822
rect 17052 77758 17054 77810
rect 17106 77758 17108 77810
rect 16940 76466 16996 76478
rect 16940 76414 16942 76466
rect 16994 76414 16996 76466
rect 16940 76356 16996 76414
rect 17052 76356 17108 77758
rect 16940 76300 17108 76356
rect 16828 76188 16996 76244
rect 16828 75124 16884 75134
rect 16716 74788 16772 74798
rect 16716 74694 16772 74732
rect 16716 74340 16772 74350
rect 16716 74246 16772 74284
rect 16604 74116 16660 74126
rect 16604 74004 16660 74060
rect 16828 74004 16884 75068
rect 16604 73948 16884 74004
rect 16604 73892 16660 73948
rect 16604 73836 16884 73892
rect 16716 73332 16772 73342
rect 16716 71762 16772 73276
rect 16716 71710 16718 71762
rect 16770 71710 16772 71762
rect 16716 67732 16772 71710
rect 16828 73330 16884 73836
rect 16828 73278 16830 73330
rect 16882 73278 16884 73330
rect 16828 71764 16884 73278
rect 16828 70532 16884 71708
rect 16940 71428 16996 76188
rect 17052 75570 17108 75582
rect 17052 75518 17054 75570
rect 17106 75518 17108 75570
rect 17052 75124 17108 75518
rect 17052 75058 17108 75068
rect 17052 74900 17108 74910
rect 17052 74806 17108 74844
rect 17052 74676 17108 74686
rect 17052 74338 17108 74620
rect 17052 74286 17054 74338
rect 17106 74286 17108 74338
rect 17052 74274 17108 74286
rect 16940 71362 16996 71372
rect 17052 74116 17108 74126
rect 16828 70466 16884 70476
rect 16940 69972 16996 69982
rect 16828 69970 16996 69972
rect 16828 69918 16942 69970
rect 16994 69918 16996 69970
rect 16828 69916 16996 69918
rect 16828 68626 16884 69916
rect 16940 69906 16996 69916
rect 16940 69412 16996 69422
rect 16940 69318 16996 69356
rect 16828 68574 16830 68626
rect 16882 68574 16884 68626
rect 16828 68562 16884 68574
rect 16828 68068 16884 68078
rect 16828 67954 16884 68012
rect 16828 67902 16830 67954
rect 16882 67902 16884 67954
rect 16828 67890 16884 67902
rect 16716 67666 16772 67676
rect 17052 67172 17108 74060
rect 16828 67116 17108 67172
rect 17164 67228 17220 85372
rect 17276 84532 17332 89292
rect 17500 89010 17556 89516
rect 17500 88958 17502 89010
rect 17554 88958 17556 89010
rect 17500 88946 17556 88958
rect 17388 88900 17444 88910
rect 17388 88806 17444 88844
rect 17500 88788 17556 88798
rect 17500 87444 17556 88732
rect 17388 86884 17444 86894
rect 17388 85316 17444 86828
rect 17388 85222 17444 85260
rect 17276 84466 17332 84476
rect 17276 84308 17332 84318
rect 17276 84306 17444 84308
rect 17276 84254 17278 84306
rect 17330 84254 17444 84306
rect 17276 84252 17444 84254
rect 17276 84242 17332 84252
rect 17276 80946 17332 80958
rect 17276 80894 17278 80946
rect 17330 80894 17332 80946
rect 17276 79602 17332 80894
rect 17276 79550 17278 79602
rect 17330 79550 17332 79602
rect 17276 79538 17332 79550
rect 17276 79044 17332 79054
rect 17276 76466 17332 78988
rect 17388 78596 17444 84252
rect 17500 83972 17556 87388
rect 17500 83906 17556 83916
rect 17500 83524 17556 83534
rect 17612 83524 17668 89628
rect 17500 83522 17668 83524
rect 17500 83470 17502 83522
rect 17554 83470 17668 83522
rect 17500 83468 17668 83470
rect 17724 84308 17780 90188
rect 17836 85988 17892 85998
rect 17836 85708 17892 85932
rect 17948 85876 18004 91196
rect 18284 91140 18340 93100
rect 18060 91084 18340 91140
rect 18060 89348 18116 91084
rect 18060 89282 18116 89292
rect 18172 90356 18228 90366
rect 18172 89234 18228 90300
rect 18172 89182 18174 89234
rect 18226 89182 18228 89234
rect 18172 89170 18228 89182
rect 18284 89906 18340 89918
rect 18284 89854 18286 89906
rect 18338 89854 18340 89906
rect 18284 88788 18340 89854
rect 18284 88722 18340 88732
rect 18396 88340 18452 93212
rect 18508 92820 18564 96012
rect 18620 96002 18676 96012
rect 18508 92754 18564 92764
rect 18620 93714 18676 93726
rect 18620 93662 18622 93714
rect 18674 93662 18676 93714
rect 18508 92596 18564 92606
rect 18508 90748 18564 92540
rect 18620 92146 18676 93662
rect 18732 92932 18788 96796
rect 18956 96180 19012 96190
rect 18956 96086 19012 96124
rect 18956 95508 19012 95518
rect 18844 95058 18900 95070
rect 18844 95006 18846 95058
rect 18898 95006 18900 95058
rect 18844 94500 18900 95006
rect 18844 94434 18900 94444
rect 18732 92876 18900 92932
rect 18732 92708 18788 92718
rect 18732 92614 18788 92652
rect 18620 92094 18622 92146
rect 18674 92094 18676 92146
rect 18620 91588 18676 92094
rect 18620 91522 18676 91532
rect 18732 91362 18788 91374
rect 18732 91310 18734 91362
rect 18786 91310 18788 91362
rect 18732 91140 18788 91310
rect 18732 91074 18788 91084
rect 18844 91364 18900 92876
rect 18508 90692 18676 90748
rect 18508 88788 18564 88798
rect 18508 88694 18564 88732
rect 18396 88246 18452 88284
rect 18060 88114 18116 88126
rect 18060 88062 18062 88114
rect 18114 88062 18116 88114
rect 18060 87668 18116 88062
rect 18116 87612 18340 87668
rect 18060 87602 18116 87612
rect 18284 87442 18340 87612
rect 18284 87390 18286 87442
rect 18338 87390 18340 87442
rect 18284 87378 18340 87390
rect 18172 85876 18228 85886
rect 17948 85874 18228 85876
rect 17948 85822 18174 85874
rect 18226 85822 18228 85874
rect 17948 85820 18228 85822
rect 17836 85652 18004 85708
rect 17724 83634 17780 84252
rect 17724 83582 17726 83634
rect 17778 83582 17780 83634
rect 17500 79044 17556 83468
rect 17724 83412 17780 83582
rect 17612 83356 17780 83412
rect 17836 84084 17892 84094
rect 17612 79156 17668 83356
rect 17724 82964 17780 82974
rect 17836 82964 17892 84028
rect 17724 82962 17892 82964
rect 17724 82910 17726 82962
rect 17778 82910 17892 82962
rect 17724 82908 17892 82910
rect 17724 82898 17780 82908
rect 17948 82348 18004 85652
rect 18060 84308 18116 84318
rect 18060 84214 18116 84252
rect 17612 79090 17668 79100
rect 17724 82292 18004 82348
rect 18060 82852 18116 82862
rect 17500 78818 17556 78988
rect 17724 79042 17780 82292
rect 17836 79604 17892 79614
rect 17836 79510 17892 79548
rect 17724 78990 17726 79042
rect 17778 78990 17780 79042
rect 17500 78766 17502 78818
rect 17554 78766 17556 78818
rect 17500 78754 17556 78766
rect 17612 78820 17668 78830
rect 17388 78540 17556 78596
rect 17388 77364 17444 77374
rect 17388 77270 17444 77308
rect 17276 76414 17278 76466
rect 17330 76414 17332 76466
rect 17276 76356 17332 76414
rect 17276 76290 17332 76300
rect 17500 76244 17556 78540
rect 17612 78258 17668 78764
rect 17612 78206 17614 78258
rect 17666 78206 17668 78258
rect 17612 78194 17668 78206
rect 17388 76242 17556 76244
rect 17388 76190 17502 76242
rect 17554 76190 17556 76242
rect 17388 76188 17556 76190
rect 17388 75572 17444 76188
rect 17500 76178 17556 76188
rect 17612 77364 17668 77374
rect 17388 75506 17444 75516
rect 17500 75908 17556 75918
rect 17500 74564 17556 75852
rect 17388 74508 17556 74564
rect 17612 74898 17668 77308
rect 17724 76580 17780 78990
rect 17724 76514 17780 76524
rect 17948 76468 18004 76478
rect 17612 74846 17614 74898
rect 17666 74846 17668 74898
rect 17388 74116 17444 74508
rect 17612 74452 17668 74846
rect 17836 75124 17892 75134
rect 17724 74676 17780 74686
rect 17724 74582 17780 74620
rect 17388 74050 17444 74060
rect 17500 74396 17668 74452
rect 17276 73106 17332 73118
rect 17276 73054 17278 73106
rect 17330 73054 17332 73106
rect 17276 70084 17332 73054
rect 17388 72772 17444 72782
rect 17388 72678 17444 72716
rect 17332 70028 17444 70084
rect 17276 70018 17332 70028
rect 17276 69524 17332 69534
rect 17276 69430 17332 69468
rect 17276 68964 17332 68974
rect 17276 68626 17332 68908
rect 17276 68574 17278 68626
rect 17330 68574 17332 68626
rect 17276 68562 17332 68574
rect 17164 67162 17220 67172
rect 17276 67842 17332 67854
rect 17276 67790 17278 67842
rect 17330 67790 17332 67842
rect 16828 63812 16884 67116
rect 17164 67058 17220 67070
rect 17164 67006 17166 67058
rect 17218 67006 17220 67058
rect 17164 66948 17220 67006
rect 17164 66882 17220 66892
rect 16828 63140 16884 63756
rect 16828 63074 16884 63084
rect 16940 65604 16996 65614
rect 16940 63138 16996 65548
rect 17276 65492 17332 67790
rect 17388 66724 17444 70028
rect 17388 66658 17444 66668
rect 17388 65492 17444 65502
rect 17276 65490 17444 65492
rect 17276 65438 17390 65490
rect 17442 65438 17444 65490
rect 17276 65436 17444 65438
rect 17388 65426 17444 65436
rect 17500 65268 17556 74396
rect 17724 74116 17780 74126
rect 17612 74004 17668 74014
rect 17612 73910 17668 73948
rect 17724 72770 17780 74060
rect 17724 72718 17726 72770
rect 17778 72718 17780 72770
rect 17724 72706 17780 72718
rect 17612 72212 17668 72222
rect 17612 71762 17668 72156
rect 17612 71710 17614 71762
rect 17666 71710 17668 71762
rect 17612 68852 17668 71710
rect 17724 70196 17780 70206
rect 17724 70102 17780 70140
rect 17612 68786 17668 68796
rect 17836 68180 17892 75068
rect 17724 68124 17892 68180
rect 17612 67842 17668 67854
rect 17612 67790 17614 67842
rect 17666 67790 17668 67842
rect 17612 67508 17668 67790
rect 17612 67442 17668 67452
rect 16940 63086 16942 63138
rect 16994 63086 16996 63138
rect 16940 63074 16996 63086
rect 17164 65212 17556 65268
rect 16828 62692 16884 62702
rect 16828 61570 16884 62636
rect 16828 61518 16830 61570
rect 16882 61518 16884 61570
rect 16828 61506 16884 61518
rect 16940 62132 16996 62142
rect 16716 61348 16772 61358
rect 16716 61254 16772 61292
rect 16604 60228 16660 60238
rect 16604 60004 16660 60172
rect 16940 60114 16996 62076
rect 17164 61684 17220 65212
rect 17388 63924 17444 63934
rect 17724 63924 17780 68124
rect 17836 67956 17892 67966
rect 17836 67862 17892 67900
rect 17836 66834 17892 66846
rect 17836 66782 17838 66834
rect 17890 66782 17892 66834
rect 17836 66276 17892 66782
rect 17836 66210 17892 66220
rect 17388 63810 17444 63868
rect 17388 63758 17390 63810
rect 17442 63758 17444 63810
rect 17388 63746 17444 63758
rect 17612 63868 17780 63924
rect 17388 63588 17444 63598
rect 17276 62356 17332 62394
rect 17276 62290 17332 62300
rect 17388 62188 17444 63532
rect 17500 63364 17556 63374
rect 17500 63270 17556 63308
rect 17276 62132 17444 62188
rect 17500 63140 17556 63150
rect 17276 61908 17332 62132
rect 17276 61842 17332 61852
rect 17164 61618 17220 61628
rect 17052 61572 17108 61582
rect 17052 61478 17108 61516
rect 17164 61346 17220 61358
rect 17164 61294 17166 61346
rect 17218 61294 17220 61346
rect 17164 61012 17220 61294
rect 17164 60946 17220 60956
rect 17388 61236 17444 61246
rect 17052 60564 17108 60574
rect 17052 60562 17332 60564
rect 17052 60510 17054 60562
rect 17106 60510 17332 60562
rect 17052 60508 17332 60510
rect 17052 60498 17108 60508
rect 16940 60062 16942 60114
rect 16994 60062 16996 60114
rect 16940 60050 16996 60062
rect 16604 59910 16660 59948
rect 17276 60002 17332 60508
rect 17276 59950 17278 60002
rect 17330 59950 17332 60002
rect 17276 59938 17332 59950
rect 16828 59220 16884 59230
rect 16828 59126 16884 59164
rect 16492 58818 16548 58828
rect 16716 59108 16772 59118
rect 16716 58658 16772 59052
rect 17388 59106 17444 61180
rect 17500 60116 17556 63084
rect 17612 62188 17668 63868
rect 17724 63700 17780 63710
rect 17724 63606 17780 63644
rect 17948 62188 18004 76412
rect 18060 75908 18116 82796
rect 18172 82292 18228 85820
rect 18508 84868 18564 84878
rect 18396 84866 18564 84868
rect 18396 84814 18510 84866
rect 18562 84814 18564 84866
rect 18396 84812 18564 84814
rect 18396 83522 18452 84812
rect 18508 84802 18564 84812
rect 18620 84868 18676 90692
rect 18732 90692 18788 90702
rect 18732 89794 18788 90636
rect 18844 90580 18900 91308
rect 18844 90486 18900 90524
rect 18732 89742 18734 89794
rect 18786 89742 18788 89794
rect 18732 89730 18788 89742
rect 18732 89012 18788 89022
rect 18732 85708 18788 88956
rect 18844 87220 18900 87230
rect 18844 87126 18900 87164
rect 18844 86772 18900 86782
rect 18956 86772 19012 95452
rect 18844 86770 19012 86772
rect 18844 86718 18846 86770
rect 18898 86718 19012 86770
rect 18844 86716 19012 86718
rect 18844 86706 18900 86716
rect 18956 86660 19012 86716
rect 18956 86594 19012 86604
rect 19068 86324 19124 97358
rect 19292 94500 19348 98140
rect 19516 97468 19572 99148
rect 19404 97412 19572 97468
rect 19404 97410 19460 97412
rect 19404 97358 19406 97410
rect 19458 97358 19460 97410
rect 19404 97346 19460 97358
rect 19516 97076 19572 97086
rect 19516 96850 19572 97020
rect 19516 96798 19518 96850
rect 19570 96798 19572 96850
rect 19516 96786 19572 96798
rect 19516 95956 19572 95966
rect 19516 95862 19572 95900
rect 19628 94724 19684 103964
rect 19628 94658 19684 94668
rect 19740 94612 19796 104636
rect 19852 98868 19908 106428
rect 19964 104020 20020 109452
rect 20076 109170 20132 109182
rect 20076 109118 20078 109170
rect 20130 109118 20132 109170
rect 20076 107604 20132 109118
rect 20076 107538 20132 107548
rect 20188 105924 20244 111806
rect 20300 110402 20356 112476
rect 20412 111076 20468 113036
rect 20524 112420 20580 114380
rect 20636 112644 20692 114800
rect 20636 112578 20692 112588
rect 20748 112756 20804 112766
rect 20636 112420 20692 112430
rect 20524 112418 20692 112420
rect 20524 112366 20638 112418
rect 20690 112366 20692 112418
rect 20524 112364 20692 112366
rect 20636 112354 20692 112364
rect 20748 111746 20804 112700
rect 20748 111694 20750 111746
rect 20802 111694 20804 111746
rect 20748 111682 20804 111694
rect 20412 111010 20468 111020
rect 20524 111636 20580 111646
rect 20300 110350 20302 110402
rect 20354 110350 20356 110402
rect 20300 110338 20356 110350
rect 20076 105868 20244 105924
rect 20076 105140 20132 105868
rect 20076 105074 20132 105084
rect 20524 104130 20580 111580
rect 20636 111524 20692 111534
rect 20636 110850 20692 111468
rect 20860 111188 20916 114800
rect 20860 111122 20916 111132
rect 20972 112306 21028 112318
rect 20972 112254 20974 112306
rect 21026 112254 21028 112306
rect 20860 110964 20916 110974
rect 20636 110798 20638 110850
rect 20690 110798 20692 110850
rect 20636 110786 20692 110798
rect 20748 110962 20916 110964
rect 20748 110910 20862 110962
rect 20914 110910 20916 110962
rect 20748 110908 20916 110910
rect 20636 110290 20692 110302
rect 20636 110238 20638 110290
rect 20690 110238 20692 110290
rect 20636 109284 20692 110238
rect 20636 109218 20692 109228
rect 20524 104078 20526 104130
rect 20578 104078 20580 104130
rect 20524 104066 20580 104078
rect 19964 103964 20132 104020
rect 19964 103796 20020 103806
rect 19964 103702 20020 103740
rect 19852 98802 19908 98812
rect 19964 99204 20020 99214
rect 19964 98530 20020 99148
rect 19964 98478 19966 98530
rect 20018 98478 20020 98530
rect 19964 98466 20020 98478
rect 19852 98196 19908 98206
rect 19852 98102 19908 98140
rect 19852 96626 19908 96638
rect 19852 96574 19854 96626
rect 19906 96574 19908 96626
rect 19852 95284 19908 96574
rect 19964 96292 20020 96302
rect 20076 96292 20132 103964
rect 20020 96236 20132 96292
rect 20300 98868 20356 98878
rect 19964 96198 20020 96236
rect 19852 95218 19908 95228
rect 19964 95058 20020 95070
rect 19964 95006 19966 95058
rect 20018 95006 20020 95058
rect 19740 94556 19908 94612
rect 19292 94444 19684 94500
rect 19292 94276 19348 94286
rect 19292 94182 19348 94220
rect 19180 93492 19236 93502
rect 19180 93398 19236 93436
rect 19516 93492 19572 93502
rect 19516 93398 19572 93436
rect 19404 92708 19460 92718
rect 19292 92484 19348 92494
rect 19180 91922 19236 91934
rect 19180 91870 19182 91922
rect 19234 91870 19236 91922
rect 19180 90916 19236 91870
rect 19292 91700 19348 92428
rect 19292 91634 19348 91644
rect 19180 90850 19236 90860
rect 19404 89794 19460 92652
rect 19516 91924 19572 91934
rect 19516 91830 19572 91868
rect 19516 91700 19572 91710
rect 19516 89906 19572 91644
rect 19516 89854 19518 89906
rect 19570 89854 19572 89906
rect 19516 89842 19572 89854
rect 19404 89742 19406 89794
rect 19458 89742 19460 89794
rect 19404 89730 19460 89742
rect 19628 88228 19684 94444
rect 19740 94386 19796 94398
rect 19740 94334 19742 94386
rect 19794 94334 19796 94386
rect 19740 93156 19796 94334
rect 19740 93042 19796 93100
rect 19740 92990 19742 93042
rect 19794 92990 19796 93042
rect 19740 92978 19796 92990
rect 19852 92596 19908 94556
rect 19964 94500 20020 95006
rect 19964 94434 20020 94444
rect 20076 94724 20132 94734
rect 19852 92530 19908 92540
rect 19740 91364 19796 91374
rect 19740 91270 19796 91308
rect 20076 91028 20132 94668
rect 20188 94500 20244 94538
rect 20188 94434 20244 94444
rect 20188 94276 20244 94286
rect 20188 92930 20244 94220
rect 20188 92878 20190 92930
rect 20242 92878 20244 92930
rect 20188 92866 20244 92878
rect 19404 88172 19684 88228
rect 19852 90972 20132 91028
rect 20188 91476 20244 91486
rect 19292 88004 19348 88014
rect 19292 86658 19348 87948
rect 19292 86606 19294 86658
rect 19346 86606 19348 86658
rect 19292 86594 19348 86606
rect 19068 86268 19348 86324
rect 19180 85988 19236 85998
rect 19068 85762 19124 85774
rect 19068 85710 19070 85762
rect 19122 85710 19124 85762
rect 18732 85652 19012 85708
rect 18620 84802 18676 84812
rect 18732 84084 18788 84094
rect 18396 83470 18398 83522
rect 18450 83470 18452 83522
rect 18396 83458 18452 83470
rect 18508 84082 18788 84084
rect 18508 84030 18734 84082
rect 18786 84030 18788 84082
rect 18508 84028 18788 84030
rect 18508 83300 18564 84028
rect 18732 84018 18788 84028
rect 18284 83244 18564 83300
rect 18732 83522 18788 83534
rect 18732 83470 18734 83522
rect 18786 83470 18788 83522
rect 18284 82738 18340 83244
rect 18284 82686 18286 82738
rect 18338 82686 18340 82738
rect 18284 82674 18340 82686
rect 18508 82516 18564 82526
rect 18508 82422 18564 82460
rect 18172 82226 18228 82236
rect 18396 81396 18452 81406
rect 18396 80386 18452 81340
rect 18396 80334 18398 80386
rect 18450 80334 18452 80386
rect 18396 80322 18452 80334
rect 18620 79604 18676 79614
rect 18508 79602 18676 79604
rect 18508 79550 18622 79602
rect 18674 79550 18676 79602
rect 18508 79548 18676 79550
rect 18172 78820 18228 78830
rect 18172 78726 18228 78764
rect 18508 77252 18564 79548
rect 18620 79538 18676 79548
rect 18732 79604 18788 83470
rect 18844 80836 18900 80846
rect 18844 80610 18900 80780
rect 18844 80558 18846 80610
rect 18898 80558 18900 80610
rect 18844 80546 18900 80558
rect 18732 78820 18788 79548
rect 18396 77196 18564 77252
rect 18620 78818 18788 78820
rect 18620 78766 18734 78818
rect 18786 78766 18788 78818
rect 18620 78764 18788 78766
rect 18172 77028 18228 77038
rect 18172 76466 18228 76972
rect 18172 76414 18174 76466
rect 18226 76414 18228 76466
rect 18172 76402 18228 76414
rect 18396 76468 18452 77196
rect 18508 77028 18564 77038
rect 18508 76934 18564 76972
rect 18396 76402 18452 76412
rect 18620 76468 18676 78764
rect 18732 78754 18788 78764
rect 18732 78260 18788 78270
rect 18732 77812 18788 78204
rect 18732 77718 18788 77756
rect 18620 76466 18788 76468
rect 18620 76414 18622 76466
rect 18674 76414 18788 76466
rect 18620 76412 18788 76414
rect 18620 76402 18676 76412
rect 18060 75842 18116 75852
rect 18620 75684 18676 75694
rect 18396 75682 18676 75684
rect 18396 75630 18622 75682
rect 18674 75630 18676 75682
rect 18396 75628 18676 75630
rect 18396 74898 18452 75628
rect 18620 75618 18676 75628
rect 18732 75124 18788 76412
rect 18732 75058 18788 75068
rect 18844 76356 18900 76366
rect 18396 74846 18398 74898
rect 18450 74846 18452 74898
rect 18396 74834 18452 74846
rect 18844 74898 18900 76300
rect 18844 74846 18846 74898
rect 18898 74846 18900 74898
rect 18844 74834 18900 74846
rect 18396 74228 18452 74238
rect 18060 74114 18116 74126
rect 18060 74062 18062 74114
rect 18114 74062 18116 74114
rect 18060 73556 18116 74062
rect 18396 74114 18452 74172
rect 18396 74062 18398 74114
rect 18450 74062 18452 74114
rect 18396 74050 18452 74062
rect 18620 74226 18676 74238
rect 18620 74174 18622 74226
rect 18674 74174 18676 74226
rect 18620 74116 18676 74174
rect 18620 74050 18676 74060
rect 18060 73490 18116 73500
rect 18172 74004 18228 74014
rect 18172 70308 18228 73948
rect 18396 73556 18452 73566
rect 18396 73462 18452 73500
rect 18844 72660 18900 72670
rect 18956 72660 19012 85652
rect 19068 84532 19124 85710
rect 19068 84466 19124 84476
rect 19068 84306 19124 84318
rect 19068 84254 19070 84306
rect 19122 84254 19124 84306
rect 19068 84196 19124 84254
rect 19068 84130 19124 84140
rect 19180 79044 19236 85932
rect 19292 84420 19348 86268
rect 19404 85988 19460 88172
rect 19628 88004 19684 88014
rect 19628 87910 19684 87948
rect 19628 87108 19684 87118
rect 19628 86658 19684 87052
rect 19852 87108 19908 90972
rect 20076 90804 20132 90814
rect 19852 87042 19908 87052
rect 19964 87218 20020 87230
rect 19964 87166 19966 87218
rect 20018 87166 20020 87218
rect 19852 86772 19908 86782
rect 19852 86678 19908 86716
rect 19628 86606 19630 86658
rect 19682 86606 19684 86658
rect 19628 86594 19684 86606
rect 19964 86436 20020 87166
rect 19404 85922 19460 85932
rect 19852 86380 20020 86436
rect 19628 85874 19684 85886
rect 19628 85822 19630 85874
rect 19682 85822 19684 85874
rect 19404 85764 19460 85802
rect 19404 85698 19460 85708
rect 19628 85316 19684 85822
rect 19852 85708 19908 86380
rect 19964 86100 20020 86110
rect 20076 86100 20132 90748
rect 20188 89794 20244 91420
rect 20188 89742 20190 89794
rect 20242 89742 20244 89794
rect 20188 89730 20244 89742
rect 19964 86098 20132 86100
rect 19964 86046 19966 86098
rect 20018 86046 20132 86098
rect 19964 86044 20132 86046
rect 20188 87108 20244 87118
rect 19964 86034 20020 86044
rect 19852 85652 20020 85708
rect 19628 85250 19684 85260
rect 19740 85092 19796 85102
rect 19740 84998 19796 85036
rect 19964 85092 20020 85652
rect 19964 85026 20020 85036
rect 20188 85090 20244 87052
rect 20188 85038 20190 85090
rect 20242 85038 20244 85090
rect 20188 85026 20244 85038
rect 19404 84978 19460 84990
rect 19404 84926 19406 84978
rect 19458 84926 19460 84978
rect 19404 84756 19460 84926
rect 19404 84690 19460 84700
rect 19852 84868 19908 84878
rect 19292 84354 19348 84364
rect 19628 84644 19684 84654
rect 19292 84194 19348 84206
rect 19292 84142 19294 84194
rect 19346 84142 19348 84194
rect 19292 84084 19348 84142
rect 19628 84194 19684 84588
rect 19628 84142 19630 84194
rect 19682 84142 19684 84194
rect 19628 84130 19684 84142
rect 19740 84420 19796 84430
rect 19292 84018 19348 84028
rect 19740 83522 19796 84364
rect 19740 83470 19742 83522
rect 19794 83470 19796 83522
rect 19516 83300 19572 83310
rect 19516 82068 19572 83244
rect 19516 82012 19684 82068
rect 19404 81956 19460 81966
rect 19404 81862 19460 81900
rect 18620 72658 19012 72660
rect 18620 72606 18846 72658
rect 18898 72606 19012 72658
rect 18620 72604 19012 72606
rect 19068 78988 19236 79044
rect 19292 81284 19348 81294
rect 18396 72548 18452 72558
rect 18284 72546 18452 72548
rect 18284 72494 18398 72546
rect 18450 72494 18452 72546
rect 18284 72492 18452 72494
rect 18284 71764 18340 72492
rect 18396 72482 18452 72492
rect 18284 71670 18340 71708
rect 18060 70252 18228 70308
rect 18060 68068 18116 70252
rect 18172 70084 18228 70094
rect 18172 69990 18228 70028
rect 18508 69186 18564 69198
rect 18508 69134 18510 69186
rect 18562 69134 18564 69186
rect 18284 68964 18340 68974
rect 18060 68002 18116 68012
rect 18172 68852 18228 68862
rect 18172 67508 18228 68796
rect 18284 67620 18340 68908
rect 18396 68626 18452 68638
rect 18396 68574 18398 68626
rect 18450 68574 18452 68626
rect 18396 68292 18452 68574
rect 18396 68226 18452 68236
rect 18396 67844 18452 67854
rect 18508 67844 18564 69134
rect 18396 67842 18564 67844
rect 18396 67790 18398 67842
rect 18450 67790 18564 67842
rect 18396 67788 18564 67790
rect 18396 67778 18452 67788
rect 18284 67564 18564 67620
rect 18172 67442 18228 67452
rect 18284 67172 18340 67182
rect 18172 67060 18228 67070
rect 18172 66386 18228 67004
rect 18172 66334 18174 66386
rect 18226 66334 18228 66386
rect 18172 66322 18228 66334
rect 18172 65604 18228 65614
rect 18172 63922 18228 65548
rect 18172 63870 18174 63922
rect 18226 63870 18228 63922
rect 18172 63858 18228 63870
rect 18284 65602 18340 67116
rect 18508 66500 18564 67564
rect 18508 66434 18564 66444
rect 18508 66276 18564 66286
rect 18508 66182 18564 66220
rect 18284 65550 18286 65602
rect 18338 65550 18340 65602
rect 18284 63700 18340 65550
rect 17612 62132 17780 62188
rect 17724 61908 17780 62132
rect 17724 61842 17780 61852
rect 17836 62132 18004 62188
rect 18060 63644 18340 63700
rect 18508 66052 18564 66062
rect 18060 62466 18116 63644
rect 18060 62414 18062 62466
rect 18114 62414 18116 62466
rect 17612 61796 17668 61806
rect 17612 61702 17668 61740
rect 17724 61458 17780 61470
rect 17724 61406 17726 61458
rect 17778 61406 17780 61458
rect 17612 61124 17668 61134
rect 17612 60786 17668 61068
rect 17724 61012 17780 61406
rect 17836 61124 17892 62132
rect 17948 61908 18004 61918
rect 17948 61236 18004 61852
rect 18060 61348 18116 62414
rect 18396 63364 18452 63374
rect 18396 62242 18452 63308
rect 18396 62190 18398 62242
rect 18450 62190 18452 62242
rect 18396 62178 18452 62190
rect 18172 61684 18228 61694
rect 18172 61590 18228 61628
rect 18060 61292 18228 61348
rect 18172 61236 18228 61292
rect 17948 61180 18116 61236
rect 18172 61180 18340 61236
rect 17836 61068 18004 61124
rect 17724 60946 17780 60956
rect 17612 60734 17614 60786
rect 17666 60734 17668 60786
rect 17612 60722 17668 60734
rect 17836 60900 17892 60910
rect 17500 60050 17556 60060
rect 17724 60340 17780 60350
rect 17388 59054 17390 59106
rect 17442 59054 17444 59106
rect 17388 59042 17444 59054
rect 16716 58606 16718 58658
rect 16770 58606 16772 58658
rect 16716 58594 16772 58606
rect 17052 58660 17108 58670
rect 17052 58566 17108 58604
rect 16716 57650 16772 57662
rect 16716 57598 16718 57650
rect 16770 57598 16772 57650
rect 16716 57204 16772 57598
rect 16716 57138 16772 57148
rect 17724 57650 17780 60284
rect 17836 60002 17892 60844
rect 17948 60340 18004 61068
rect 17948 60274 18004 60284
rect 17836 59950 17838 60002
rect 17890 59950 17892 60002
rect 17836 59938 17892 59950
rect 17948 60114 18004 60126
rect 17948 60062 17950 60114
rect 18002 60062 18004 60114
rect 17948 58660 18004 60062
rect 17948 58594 18004 58604
rect 17724 57598 17726 57650
rect 17778 57598 17780 57650
rect 17724 55468 17780 57598
rect 17500 55412 17780 55468
rect 16380 50260 16436 54460
rect 17164 54516 17220 54526
rect 17164 54422 17220 54460
rect 17164 53732 17220 53742
rect 16492 53396 16548 53406
rect 16492 52946 16548 53340
rect 16492 52894 16494 52946
rect 16546 52894 16548 52946
rect 16492 52882 16548 52894
rect 16828 52724 16884 52734
rect 16828 52630 16884 52668
rect 16828 52500 16884 52510
rect 16828 52162 16884 52444
rect 17052 52276 17108 52286
rect 17052 52182 17108 52220
rect 16828 52110 16830 52162
rect 16882 52110 16884 52162
rect 16828 52098 16884 52110
rect 16940 51154 16996 51166
rect 16940 51102 16942 51154
rect 16994 51102 16996 51154
rect 16380 50194 16436 50204
rect 16828 50370 16884 50382
rect 16828 50318 16830 50370
rect 16882 50318 16884 50370
rect 16828 49810 16884 50318
rect 16828 49758 16830 49810
rect 16882 49758 16884 49810
rect 16828 49746 16884 49758
rect 16156 49588 16212 49598
rect 15932 48468 15988 48478
rect 15820 48466 15988 48468
rect 15820 48414 15934 48466
rect 15986 48414 15988 48466
rect 15820 48412 15988 48414
rect 15932 48402 15988 48412
rect 15932 47460 15988 47470
rect 15932 47366 15988 47404
rect 16044 46450 16100 46462
rect 16044 46398 16046 46450
rect 16098 46398 16100 46450
rect 16044 46116 16100 46398
rect 16044 46050 16100 46060
rect 15932 44100 15988 44110
rect 15708 44098 15988 44100
rect 15708 44046 15934 44098
rect 15986 44046 15988 44098
rect 15708 44044 15988 44046
rect 15708 43538 15764 44044
rect 15932 44034 15988 44044
rect 15708 43486 15710 43538
rect 15762 43486 15764 43538
rect 15708 43474 15764 43486
rect 16044 43538 16100 43550
rect 16044 43486 16046 43538
rect 16098 43486 16100 43538
rect 16044 43204 16100 43486
rect 16044 43138 16100 43148
rect 16156 42868 16212 49532
rect 15820 42812 16212 42868
rect 15708 42756 15764 42766
rect 15708 42662 15764 42700
rect 15820 41524 15876 42812
rect 16156 42644 16212 42654
rect 15820 40404 15876 41468
rect 15820 40338 15876 40348
rect 15932 42642 16212 42644
rect 15932 42590 16158 42642
rect 16210 42590 16212 42642
rect 15932 42588 16212 42590
rect 15932 40292 15988 42588
rect 16156 42578 16212 42588
rect 16268 41860 16324 49644
rect 16380 49588 16436 49598
rect 16380 49494 16436 49532
rect 16604 48580 16660 48590
rect 16604 48354 16660 48524
rect 16604 48302 16606 48354
rect 16658 48302 16660 48354
rect 16604 47908 16660 48302
rect 16940 48356 16996 51102
rect 16940 48290 16996 48300
rect 16604 47842 16660 47852
rect 16828 48244 16884 48254
rect 16604 47348 16660 47358
rect 16380 46564 16436 46574
rect 16380 46470 16436 46508
rect 16604 46450 16660 47292
rect 16604 46398 16606 46450
rect 16658 46398 16660 46450
rect 16268 41794 16324 41804
rect 16380 46004 16436 46014
rect 16380 41636 16436 45948
rect 16604 46004 16660 46398
rect 16604 45938 16660 45948
rect 16716 47346 16772 47358
rect 16716 47294 16718 47346
rect 16770 47294 16772 47346
rect 16604 45556 16660 45566
rect 16604 42980 16660 45500
rect 16604 42914 16660 42924
rect 16492 42082 16548 42094
rect 16492 42030 16494 42082
rect 16546 42030 16548 42082
rect 16492 41972 16548 42030
rect 16492 41906 16548 41916
rect 16380 41580 16660 41636
rect 16044 40964 16100 40974
rect 16044 40962 16548 40964
rect 16044 40910 16046 40962
rect 16098 40910 16548 40962
rect 16044 40908 16548 40910
rect 16044 40898 16100 40908
rect 16268 40516 16324 40526
rect 15932 40226 15988 40236
rect 16156 40290 16212 40302
rect 16156 40238 16158 40290
rect 16210 40238 16212 40290
rect 15708 38836 15764 38846
rect 15708 38742 15764 38780
rect 16044 38500 16100 38510
rect 15932 37266 15988 37278
rect 15932 37214 15934 37266
rect 15986 37214 15988 37266
rect 15932 36708 15988 37214
rect 16044 36932 16100 38444
rect 16156 37380 16212 40238
rect 16268 38668 16324 40460
rect 16492 40402 16548 40908
rect 16492 40350 16494 40402
rect 16546 40350 16548 40402
rect 16492 40338 16548 40350
rect 16604 38668 16660 41580
rect 16716 40516 16772 47294
rect 16828 46116 16884 48188
rect 16940 48132 16996 48142
rect 17164 48132 17220 53676
rect 17276 51156 17332 51166
rect 17276 51062 17332 51100
rect 17500 50428 17556 55412
rect 17948 51604 18004 51614
rect 17948 50818 18004 51548
rect 17948 50766 17950 50818
rect 18002 50766 18004 50818
rect 17948 50708 18004 50766
rect 17948 50642 18004 50652
rect 17948 50484 18004 50494
rect 17500 50372 17668 50428
rect 17388 49810 17444 49822
rect 17388 49758 17390 49810
rect 17442 49758 17444 49810
rect 17388 48916 17444 49758
rect 17388 48850 17444 48860
rect 16940 48130 17220 48132
rect 16940 48078 16942 48130
rect 16994 48078 17220 48130
rect 16940 48076 17220 48078
rect 16940 46452 16996 48076
rect 17500 47572 17556 47582
rect 17052 47460 17108 47470
rect 17052 47366 17108 47404
rect 17500 47458 17556 47516
rect 17500 47406 17502 47458
rect 17554 47406 17556 47458
rect 17500 47394 17556 47406
rect 16940 46396 17108 46452
rect 16828 46060 16996 46116
rect 16828 44322 16884 44334
rect 16828 44270 16830 44322
rect 16882 44270 16884 44322
rect 16828 41972 16884 44270
rect 16828 41906 16884 41916
rect 16940 41858 16996 46060
rect 16940 41806 16942 41858
rect 16994 41806 16996 41858
rect 16940 41794 16996 41806
rect 17052 40964 17108 46396
rect 17276 46340 17332 46350
rect 17276 44434 17332 46284
rect 17276 44382 17278 44434
rect 17330 44382 17332 44434
rect 17276 44370 17332 44382
rect 17388 45106 17444 45118
rect 17388 45054 17390 45106
rect 17442 45054 17444 45106
rect 17164 43540 17220 43550
rect 17164 43446 17220 43484
rect 17388 43316 17444 45054
rect 17612 43652 17668 50372
rect 17836 49140 17892 49150
rect 17724 47570 17780 47582
rect 17724 47518 17726 47570
rect 17778 47518 17780 47570
rect 17724 43764 17780 47518
rect 17836 46340 17892 49084
rect 17948 48580 18004 50428
rect 17948 48514 18004 48524
rect 17836 46284 18004 46340
rect 17836 46116 17892 46126
rect 17836 46022 17892 46060
rect 17836 44996 17892 45006
rect 17948 44996 18004 46284
rect 18060 45108 18116 61180
rect 18172 60676 18228 60686
rect 18172 60582 18228 60620
rect 18284 59892 18340 61180
rect 18508 60788 18564 65996
rect 18620 63476 18676 72604
rect 18844 72594 18900 72604
rect 18844 71538 18900 71550
rect 18844 71486 18846 71538
rect 18898 71486 18900 71538
rect 18732 69860 18788 69870
rect 18732 66052 18788 69804
rect 18844 69524 18900 71486
rect 18844 69458 18900 69468
rect 18956 70866 19012 70878
rect 18956 70814 18958 70866
rect 19010 70814 19012 70866
rect 18956 70532 19012 70814
rect 18956 68964 19012 70476
rect 18956 68898 19012 68908
rect 19068 68740 19124 78988
rect 18844 68684 19124 68740
rect 19180 78036 19236 78046
rect 19292 78036 19348 81228
rect 19180 78034 19348 78036
rect 19180 77982 19182 78034
rect 19234 77982 19348 78034
rect 19180 77980 19348 77982
rect 19180 70196 19236 77980
rect 19628 77924 19684 82012
rect 19628 77858 19684 77868
rect 19740 78818 19796 83470
rect 19740 78766 19742 78818
rect 19794 78766 19796 78818
rect 19404 76804 19460 76814
rect 19292 74114 19348 74126
rect 19292 74062 19294 74114
rect 19346 74062 19348 74114
rect 19292 71988 19348 74062
rect 19404 73948 19460 76748
rect 19516 76468 19572 76478
rect 19740 76468 19796 78766
rect 19572 76412 19796 76468
rect 19516 76374 19572 76412
rect 19740 75124 19796 75134
rect 19740 74898 19796 75068
rect 19740 74846 19742 74898
rect 19794 74846 19796 74898
rect 19740 74834 19796 74846
rect 19740 74116 19796 74154
rect 19740 74050 19796 74060
rect 19404 73892 19796 73948
rect 19292 71922 19348 71932
rect 19180 69410 19236 70140
rect 19628 71876 19684 71886
rect 19292 69972 19348 69982
rect 19292 69970 19460 69972
rect 19292 69918 19294 69970
rect 19346 69918 19460 69970
rect 19292 69916 19460 69918
rect 19292 69906 19348 69916
rect 19180 69358 19182 69410
rect 19234 69358 19236 69410
rect 18844 68180 18900 68684
rect 18844 68114 18900 68124
rect 18956 68514 19012 68526
rect 18956 68462 18958 68514
rect 19010 68462 19012 68514
rect 18844 67842 18900 67854
rect 18844 67790 18846 67842
rect 18898 67790 18900 67842
rect 18844 67732 18900 67790
rect 18844 67666 18900 67676
rect 18956 67172 19012 68462
rect 19068 68516 19124 68526
rect 19068 68422 19124 68460
rect 19180 68292 19236 69358
rect 19292 69188 19348 69198
rect 19292 68626 19348 69132
rect 19292 68574 19294 68626
rect 19346 68574 19348 68626
rect 19292 68562 19348 68574
rect 19180 68236 19348 68292
rect 18732 65986 18788 65996
rect 18844 67116 19012 67172
rect 19180 68068 19236 68078
rect 18844 67060 18900 67116
rect 18732 65266 18788 65278
rect 18732 65214 18734 65266
rect 18786 65214 18788 65266
rect 18732 65156 18788 65214
rect 18732 65090 18788 65100
rect 18844 64932 18900 67004
rect 19068 66946 19124 66958
rect 19068 66894 19070 66946
rect 19122 66894 19124 66946
rect 18956 66500 19012 66510
rect 18956 66274 19012 66444
rect 18956 66222 18958 66274
rect 19010 66222 19012 66274
rect 18956 66210 19012 66222
rect 19068 66052 19124 66894
rect 19180 66498 19236 68012
rect 19292 67172 19348 68236
rect 19404 67844 19460 69916
rect 19516 69524 19572 69534
rect 19516 69430 19572 69468
rect 19628 68852 19684 71820
rect 19740 70082 19796 73892
rect 19852 70532 19908 84812
rect 20076 84756 20132 84766
rect 20076 82348 20132 84700
rect 20076 82292 20244 82348
rect 19964 82068 20020 82078
rect 19964 80836 20020 82012
rect 19964 80770 20020 80780
rect 19964 80162 20020 80174
rect 19964 80110 19966 80162
rect 20018 80110 20020 80162
rect 19964 79604 20020 80110
rect 19964 79538 20020 79548
rect 20076 79268 20132 79278
rect 19964 77252 20020 77262
rect 19964 77158 20020 77196
rect 20076 75906 20132 79212
rect 20188 78932 20244 82292
rect 20300 80612 20356 98812
rect 20748 97468 20804 110908
rect 20860 110898 20916 110908
rect 20972 110740 21028 112254
rect 21084 111972 21140 114800
rect 21308 113652 21364 114800
rect 21308 113596 21476 113652
rect 21308 113426 21364 113438
rect 21308 113374 21310 113426
rect 21362 113374 21364 113426
rect 21084 111906 21140 111916
rect 21196 113316 21252 113326
rect 21196 111970 21252 113260
rect 21308 113092 21364 113374
rect 21420 113204 21476 113596
rect 21532 113540 21588 114800
rect 21532 113474 21588 113484
rect 21756 113428 21812 114800
rect 21756 113362 21812 113372
rect 21868 114100 21924 114110
rect 21420 113148 21588 113204
rect 21308 113036 21476 113092
rect 21308 112868 21364 112878
rect 21308 112418 21364 112812
rect 21308 112366 21310 112418
rect 21362 112366 21364 112418
rect 21308 112354 21364 112366
rect 21196 111918 21198 111970
rect 21250 111918 21252 111970
rect 21196 111906 21252 111918
rect 20860 110684 21028 110740
rect 21084 111076 21140 111086
rect 20860 108836 20916 110684
rect 20860 108770 20916 108780
rect 20972 110290 21028 110302
rect 20972 110238 20974 110290
rect 21026 110238 21028 110290
rect 20860 104132 20916 104142
rect 20860 104038 20916 104076
rect 20972 100324 21028 110238
rect 21084 100996 21140 111020
rect 21308 110964 21364 110974
rect 21308 110870 21364 110908
rect 21084 100930 21140 100940
rect 21196 110178 21252 110190
rect 21196 110126 21198 110178
rect 21250 110126 21252 110178
rect 20972 100258 21028 100268
rect 21196 98868 21252 110126
rect 21420 105476 21476 113036
rect 21532 112084 21588 113148
rect 21756 113202 21812 113214
rect 21756 113150 21758 113202
rect 21810 113150 21812 113202
rect 21756 112756 21812 113150
rect 21868 112756 21924 114044
rect 21980 112980 22036 114800
rect 21980 112914 22036 112924
rect 22204 112756 22260 114800
rect 22428 114100 22484 114800
rect 22428 114034 22484 114044
rect 22316 113876 22372 113886
rect 22316 113538 22372 113820
rect 22652 113876 22708 114800
rect 22876 114548 22932 114800
rect 22876 114482 22932 114492
rect 22988 114660 23044 114670
rect 22652 113810 22708 113820
rect 22316 113486 22318 113538
rect 22370 113486 22372 113538
rect 22316 113474 22372 113486
rect 22988 113538 23044 114604
rect 22988 113486 22990 113538
rect 23042 113486 23044 113538
rect 22988 113474 23044 113486
rect 23100 113540 23156 114800
rect 23324 114436 23380 114800
rect 23324 114370 23380 114380
rect 23100 113484 23492 113540
rect 21868 112700 22036 112756
rect 21532 112018 21588 112028
rect 21644 112306 21700 112318
rect 21644 112254 21646 112306
rect 21698 112254 21700 112306
rect 21532 111860 21588 111870
rect 21532 111766 21588 111804
rect 21644 110964 21700 112254
rect 21756 111076 21812 112700
rect 21980 112418 22036 112700
rect 22204 112690 22260 112700
rect 22540 113314 22596 113326
rect 22540 113262 22542 113314
rect 22594 113262 22596 113314
rect 21980 112366 21982 112418
rect 22034 112366 22036 112418
rect 21980 112354 22036 112366
rect 22316 112308 22372 112318
rect 22316 112306 22484 112308
rect 22316 112254 22318 112306
rect 22370 112254 22484 112306
rect 22316 112252 22484 112254
rect 22316 112242 22372 112252
rect 21868 111972 21924 111982
rect 21868 111878 21924 111916
rect 22204 111860 22260 111870
rect 22204 111766 22260 111804
rect 22204 111524 22260 111534
rect 21756 111010 21812 111020
rect 21980 111188 22036 111198
rect 21532 110908 21700 110964
rect 21980 110962 22036 111132
rect 21980 110910 21982 110962
rect 22034 110910 22036 110962
rect 21532 110292 21588 110908
rect 21980 110898 22036 110910
rect 22092 110852 22148 110862
rect 21644 110740 21700 110750
rect 21644 110738 21812 110740
rect 21644 110686 21646 110738
rect 21698 110686 21812 110738
rect 21644 110684 21812 110686
rect 21644 110674 21700 110684
rect 21644 110516 21700 110526
rect 21644 110402 21700 110460
rect 21644 110350 21646 110402
rect 21698 110350 21700 110402
rect 21644 110338 21700 110350
rect 21532 110226 21588 110236
rect 21756 106260 21812 110684
rect 21980 110404 22036 110414
rect 22092 110404 22148 110796
rect 21980 110402 22148 110404
rect 21980 110350 21982 110402
rect 22034 110350 22148 110402
rect 21980 110348 22148 110350
rect 21980 110338 22036 110348
rect 22204 110292 22260 111468
rect 22316 110964 22372 110974
rect 22316 110850 22372 110908
rect 22316 110798 22318 110850
rect 22370 110798 22372 110850
rect 22316 110786 22372 110798
rect 22092 110236 22260 110292
rect 22092 109228 22148 110236
rect 22316 110178 22372 110190
rect 22316 110126 22318 110178
rect 22370 110126 22372 110178
rect 22316 110068 22372 110126
rect 22316 110002 22372 110012
rect 21756 106194 21812 106204
rect 21980 109172 22148 109228
rect 22204 109956 22260 109966
rect 21420 105410 21476 105420
rect 21868 105474 21924 105486
rect 21868 105422 21870 105474
rect 21922 105422 21924 105474
rect 21868 104356 21924 105422
rect 21868 104290 21924 104300
rect 21196 98802 21252 98812
rect 21980 97858 22036 109172
rect 22092 105700 22148 105710
rect 22204 105700 22260 109900
rect 22428 107380 22484 112252
rect 22540 111972 22596 113262
rect 22876 113316 22932 113326
rect 23212 113316 23268 113326
rect 22652 112306 22708 112318
rect 22652 112254 22654 112306
rect 22706 112254 22708 112306
rect 22652 112196 22708 112254
rect 22652 112130 22708 112140
rect 22764 112084 22820 112094
rect 22540 111916 22708 111972
rect 22428 107314 22484 107324
rect 22540 111746 22596 111758
rect 22540 111694 22542 111746
rect 22594 111694 22596 111746
rect 22092 105698 22260 105700
rect 22092 105646 22094 105698
rect 22146 105646 22260 105698
rect 22092 105644 22260 105646
rect 22092 105634 22148 105644
rect 22540 103348 22596 111694
rect 22652 110628 22708 111916
rect 22764 110962 22820 112028
rect 22876 111970 22932 113260
rect 23100 113314 23268 113316
rect 23100 113262 23214 113314
rect 23266 113262 23268 113314
rect 23100 113260 23268 113262
rect 22876 111918 22878 111970
rect 22930 111918 22932 111970
rect 22876 111906 22932 111918
rect 22988 112306 23044 112318
rect 22988 112254 22990 112306
rect 23042 112254 23044 112306
rect 22988 111188 23044 112254
rect 22764 110910 22766 110962
rect 22818 110910 22820 110962
rect 22764 110898 22820 110910
rect 22876 111132 23044 111188
rect 22652 110562 22708 110572
rect 22652 110404 22708 110414
rect 22652 110310 22708 110348
rect 22428 103292 22596 103348
rect 22652 106148 22708 106158
rect 21980 97806 21982 97858
rect 22034 97806 22036 97858
rect 21980 97794 22036 97806
rect 22204 99762 22260 99774
rect 22204 99710 22206 99762
rect 22258 99710 22260 99762
rect 20412 97412 20804 97468
rect 21756 97634 21812 97646
rect 21756 97582 21758 97634
rect 21810 97582 21812 97634
rect 20412 90804 20468 97412
rect 21756 96740 21812 97582
rect 22204 97468 22260 99710
rect 20748 96628 20804 96638
rect 20748 96626 21364 96628
rect 20748 96574 20750 96626
rect 20802 96574 21364 96626
rect 20748 96572 21364 96574
rect 20748 96562 20804 96572
rect 20972 95956 21028 95966
rect 20636 95170 20692 95182
rect 20636 95118 20638 95170
rect 20690 95118 20692 95170
rect 20412 90738 20468 90748
rect 20524 94948 20580 94958
rect 20524 94498 20580 94892
rect 20524 94446 20526 94498
rect 20578 94446 20580 94498
rect 20524 92930 20580 94446
rect 20524 92878 20526 92930
rect 20578 92878 20580 92930
rect 20524 90580 20580 92878
rect 20412 90524 20580 90580
rect 20636 92034 20692 95118
rect 20748 94612 20804 94622
rect 20748 94610 20916 94612
rect 20748 94558 20750 94610
rect 20802 94558 20916 94610
rect 20748 94556 20916 94558
rect 20748 94546 20804 94556
rect 20636 91982 20638 92034
rect 20690 91982 20692 92034
rect 20636 90580 20692 91982
rect 20412 85708 20468 90524
rect 20524 89570 20580 89582
rect 20524 89518 20526 89570
rect 20578 89518 20580 89570
rect 20524 87556 20580 89518
rect 20636 89460 20692 90524
rect 20748 93042 20804 93054
rect 20748 92990 20750 93042
rect 20802 92990 20804 93042
rect 20748 90468 20804 92990
rect 20860 93044 20916 94556
rect 20860 92978 20916 92988
rect 20860 92820 20916 92830
rect 20860 90804 20916 92764
rect 20860 90738 20916 90748
rect 20972 91364 21028 95900
rect 21084 95842 21140 95854
rect 21084 95790 21086 95842
rect 21138 95790 21140 95842
rect 21084 95284 21140 95790
rect 21084 95282 21252 95284
rect 21084 95230 21086 95282
rect 21138 95230 21252 95282
rect 21084 95228 21252 95230
rect 21084 95218 21140 95228
rect 21084 93940 21140 93950
rect 21084 92820 21140 93884
rect 21196 93042 21252 95228
rect 21196 92990 21198 93042
rect 21250 92990 21252 93042
rect 21196 92978 21252 92990
rect 21308 94498 21364 96572
rect 21756 95956 21812 96684
rect 21980 97412 22260 97468
rect 21868 96628 21924 96638
rect 21868 96534 21924 96572
rect 21756 95862 21812 95900
rect 21308 94446 21310 94498
rect 21362 94446 21364 94498
rect 21084 92764 21252 92820
rect 21084 92148 21140 92158
rect 21084 92054 21140 92092
rect 21196 91924 21252 92764
rect 21308 92148 21364 94446
rect 21308 92082 21364 92092
rect 21420 95282 21476 95294
rect 21420 95230 21422 95282
rect 21474 95230 21476 95282
rect 21420 92146 21476 95230
rect 21644 95058 21700 95070
rect 21644 95006 21646 95058
rect 21698 95006 21700 95058
rect 21644 92932 21700 95006
rect 21644 92866 21700 92876
rect 21868 94498 21924 94510
rect 21868 94446 21870 94498
rect 21922 94446 21924 94498
rect 21868 92930 21924 94446
rect 21868 92878 21870 92930
rect 21922 92878 21924 92930
rect 21644 92708 21700 92718
rect 21420 92094 21422 92146
rect 21474 92094 21476 92146
rect 21196 91868 21364 91924
rect 21084 91364 21140 91374
rect 20972 91362 21140 91364
rect 20972 91310 21086 91362
rect 21138 91310 21140 91362
rect 20972 91308 21140 91310
rect 20972 90692 21028 91308
rect 21084 91298 21140 91308
rect 20972 90626 21028 90636
rect 21196 90692 21252 90702
rect 21196 90468 21252 90636
rect 20748 90412 21252 90468
rect 20636 89394 20692 89404
rect 20524 87490 20580 87500
rect 20636 89236 20692 89246
rect 20524 87220 20580 87230
rect 20524 86658 20580 87164
rect 20524 86606 20526 86658
rect 20578 86606 20580 86658
rect 20524 86594 20580 86606
rect 20412 85652 20580 85708
rect 20412 85316 20468 85326
rect 20412 85222 20468 85260
rect 20524 83636 20580 85652
rect 20636 84418 20692 89180
rect 21196 88228 21252 88238
rect 21196 88134 21252 88172
rect 21308 88004 21364 91868
rect 21420 90244 21476 92094
rect 21532 92372 21588 92382
rect 21532 91474 21588 92316
rect 21644 92034 21700 92652
rect 21868 92260 21924 92878
rect 21868 92194 21924 92204
rect 21644 91982 21646 92034
rect 21698 91982 21700 92034
rect 21644 91970 21700 91982
rect 21756 92148 21812 92158
rect 21532 91422 21534 91474
rect 21586 91422 21588 91474
rect 21532 90916 21588 91422
rect 21756 91252 21812 92092
rect 21980 91700 22036 97412
rect 22204 96852 22260 96862
rect 22204 96292 22260 96796
rect 22316 96850 22372 96862
rect 22316 96798 22318 96850
rect 22370 96798 22372 96850
rect 22316 96740 22372 96798
rect 22316 96674 22372 96684
rect 22204 96290 22372 96292
rect 22204 96238 22206 96290
rect 22258 96238 22372 96290
rect 22204 96236 22372 96238
rect 22204 96226 22260 96236
rect 22204 95282 22260 95294
rect 22204 95230 22206 95282
rect 22258 95230 22260 95282
rect 22092 94500 22148 94510
rect 22092 92146 22148 94444
rect 22204 94276 22260 95230
rect 22204 94210 22260 94220
rect 22316 94108 22372 96236
rect 22428 94276 22484 103292
rect 22540 99876 22596 99886
rect 22652 99876 22708 106092
rect 22876 104916 22932 111132
rect 22988 110964 23044 110974
rect 22988 110850 23044 110908
rect 22988 110798 22990 110850
rect 23042 110798 23044 110850
rect 22988 110786 23044 110798
rect 22876 104850 22932 104860
rect 22988 109394 23044 109406
rect 22988 109342 22990 109394
rect 23042 109342 23044 109394
rect 22540 99874 22708 99876
rect 22540 99822 22542 99874
rect 22594 99822 22708 99874
rect 22540 99820 22708 99822
rect 22540 99810 22596 99820
rect 22988 97748 23044 109342
rect 23100 106372 23156 113260
rect 23212 113250 23268 113260
rect 23436 113092 23492 113484
rect 23548 113204 23604 114800
rect 23772 114324 23828 114800
rect 23996 114772 24052 114800
rect 23996 114706 24052 114716
rect 23772 114258 23828 114268
rect 24220 114212 24276 114800
rect 24220 114146 24276 114156
rect 24444 113988 24500 114800
rect 24668 114660 24724 114800
rect 24668 114594 24724 114604
rect 24444 113922 24500 113932
rect 24464 113708 24728 113718
rect 24520 113652 24568 113708
rect 24624 113652 24672 113708
rect 24464 113642 24728 113652
rect 24556 113540 24612 113550
rect 24556 113446 24612 113484
rect 23884 113428 23940 113438
rect 23548 113138 23604 113148
rect 23660 113426 23940 113428
rect 23660 113374 23886 113426
rect 23938 113374 23940 113426
rect 23660 113372 23940 113374
rect 23436 113026 23492 113036
rect 23324 112980 23380 112990
rect 23324 112418 23380 112924
rect 23324 112366 23326 112418
rect 23378 112366 23380 112418
rect 23324 112354 23380 112366
rect 23548 112530 23604 112542
rect 23548 112478 23550 112530
rect 23602 112478 23604 112530
rect 23324 111748 23380 111758
rect 23212 111746 23380 111748
rect 23212 111694 23326 111746
rect 23378 111694 23380 111746
rect 23212 111692 23380 111694
rect 23212 111412 23268 111692
rect 23324 111682 23380 111692
rect 23212 111346 23268 111356
rect 23324 111300 23380 111310
rect 23324 110962 23380 111244
rect 23324 110910 23326 110962
rect 23378 110910 23380 110962
rect 23324 110898 23380 110910
rect 23324 110628 23380 110638
rect 23212 109396 23268 109406
rect 23212 109282 23268 109340
rect 23212 109230 23214 109282
rect 23266 109230 23268 109282
rect 23212 109218 23268 109230
rect 23100 106306 23156 106316
rect 23324 105868 23380 110572
rect 23548 110404 23604 112478
rect 23660 112420 23716 113372
rect 23884 113362 23940 113372
rect 24668 113428 24724 113438
rect 24220 113314 24276 113326
rect 24220 113262 24222 113314
rect 24274 113262 24276 113314
rect 23804 112924 24068 112934
rect 23860 112868 23908 112924
rect 23964 112868 24012 112924
rect 23804 112858 24068 112868
rect 23660 112354 23716 112364
rect 23996 112756 24052 112766
rect 23996 112418 24052 112700
rect 24220 112756 24276 113262
rect 24220 112690 24276 112700
rect 24332 112868 24388 112878
rect 24220 112532 24276 112542
rect 23996 112366 23998 112418
rect 24050 112366 24052 112418
rect 23996 112354 24052 112366
rect 24108 112530 24276 112532
rect 24108 112478 24222 112530
rect 24274 112478 24276 112530
rect 24108 112476 24276 112478
rect 23660 111858 23716 111870
rect 23660 111806 23662 111858
rect 23714 111806 23716 111858
rect 23660 111636 23716 111806
rect 23660 111570 23716 111580
rect 23996 111524 24052 111534
rect 24108 111524 24164 112476
rect 24220 112466 24276 112476
rect 24052 111468 24164 111524
rect 24220 112308 24276 112318
rect 23996 111458 24052 111468
rect 23804 111356 24068 111366
rect 23860 111300 23908 111356
rect 23964 111300 24012 111356
rect 23804 111290 24068 111300
rect 23884 111188 23940 111198
rect 23660 111076 23716 111086
rect 23660 110850 23716 111020
rect 23660 110798 23662 110850
rect 23714 110798 23716 110850
rect 23660 110786 23716 110798
rect 23548 110338 23604 110348
rect 23884 110402 23940 111132
rect 23996 110964 24052 110974
rect 23996 110870 24052 110908
rect 23884 110350 23886 110402
rect 23938 110350 23940 110402
rect 23884 110338 23940 110350
rect 23548 110178 23604 110190
rect 23548 110126 23550 110178
rect 23602 110126 23604 110178
rect 23548 109172 23604 110126
rect 23804 109788 24068 109798
rect 23860 109732 23908 109788
rect 23964 109732 24012 109788
rect 23804 109722 24068 109732
rect 23548 109170 23716 109172
rect 23548 109118 23550 109170
rect 23602 109118 23716 109170
rect 23548 109116 23716 109118
rect 23548 108836 23604 109116
rect 23492 108780 23604 108836
rect 23492 108734 23548 108780
rect 23436 108722 23548 108734
rect 23436 108670 23438 108722
rect 23490 108670 23548 108722
rect 23436 108668 23548 108670
rect 23436 108658 23492 108668
rect 23660 108388 23716 109116
rect 23660 108322 23716 108332
rect 23804 108220 24068 108230
rect 23860 108164 23908 108220
rect 23964 108164 24012 108220
rect 23804 108154 24068 108164
rect 23804 106652 24068 106662
rect 23860 106596 23908 106652
rect 23964 106596 24012 106652
rect 23804 106586 24068 106596
rect 23324 105812 23492 105868
rect 22988 97682 23044 97692
rect 23436 97468 23492 105812
rect 24220 105812 24276 112252
rect 24332 110850 24388 112812
rect 24668 112418 24724 113372
rect 24780 113316 24836 113326
rect 24780 113222 24836 113260
rect 24892 112532 24948 114800
rect 25116 113092 25172 114800
rect 25116 113026 25172 113036
rect 25228 113202 25284 113214
rect 25228 113150 25230 113202
rect 25282 113150 25284 113202
rect 24892 112466 24948 112476
rect 24668 112366 24670 112418
rect 24722 112366 24724 112418
rect 24668 112354 24724 112366
rect 24892 112308 24948 112318
rect 24464 112140 24728 112150
rect 24520 112084 24568 112140
rect 24624 112084 24672 112140
rect 24464 112074 24728 112084
rect 24892 111970 24948 112252
rect 24892 111918 24894 111970
rect 24946 111918 24948 111970
rect 24892 111906 24948 111918
rect 25004 112306 25060 112318
rect 25004 112254 25006 112306
rect 25058 112254 25060 112306
rect 24332 110798 24334 110850
rect 24386 110798 24388 110850
rect 24332 110786 24388 110798
rect 24556 111746 24612 111758
rect 24556 111694 24558 111746
rect 24610 111694 24612 111746
rect 24556 110740 24612 111694
rect 24668 111748 24724 111758
rect 24668 110962 24724 111692
rect 25004 111636 25060 112254
rect 24668 110910 24670 110962
rect 24722 110910 24724 110962
rect 24668 110898 24724 110910
rect 24780 111580 25060 111636
rect 25116 111972 25172 111982
rect 24780 110852 24836 111580
rect 24780 110786 24836 110796
rect 24892 111412 24948 111422
rect 24556 110674 24612 110684
rect 24464 110572 24728 110582
rect 24520 110516 24568 110572
rect 24624 110516 24672 110572
rect 24464 110506 24728 110516
rect 24892 110402 24948 111356
rect 25004 111188 25060 111198
rect 25004 110850 25060 111132
rect 25116 111076 25172 111916
rect 25116 111010 25172 111020
rect 25228 111746 25284 113150
rect 25340 112644 25396 114800
rect 25452 114100 25508 114110
rect 25452 113538 25508 114044
rect 25452 113486 25454 113538
rect 25506 113486 25508 113538
rect 25452 113474 25508 113486
rect 25564 112756 25620 114800
rect 25564 112690 25620 112700
rect 25676 113876 25732 113886
rect 25340 112578 25396 112588
rect 25564 112420 25620 112430
rect 25676 112420 25732 113820
rect 25788 113652 25844 114800
rect 25788 113586 25844 113596
rect 26012 113540 26068 114800
rect 28476 114772 28532 114782
rect 26012 113474 26068 113484
rect 26124 114548 26180 114558
rect 26124 113538 26180 114492
rect 26124 113486 26126 113538
rect 26178 113486 26180 113538
rect 26124 113474 26180 113486
rect 26796 114436 26852 114446
rect 26796 113538 26852 114380
rect 28364 114324 28420 114334
rect 26796 113486 26798 113538
rect 26850 113486 26852 113538
rect 26796 113474 26852 113486
rect 27692 113988 27748 113998
rect 27692 113538 27748 113932
rect 27692 113486 27694 113538
rect 27746 113486 27748 113538
rect 27692 113474 27748 113486
rect 28364 113538 28420 114268
rect 28364 113486 28366 113538
rect 28418 113486 28420 113538
rect 28364 113474 28420 113486
rect 25788 113316 25844 113326
rect 25788 113314 25956 113316
rect 25788 113262 25790 113314
rect 25842 113262 25956 113314
rect 25788 113260 25956 113262
rect 25788 113250 25844 113260
rect 25564 112418 25732 112420
rect 25564 112366 25566 112418
rect 25618 112366 25732 112418
rect 25564 112364 25732 112366
rect 25788 112530 25844 112542
rect 25788 112478 25790 112530
rect 25842 112478 25844 112530
rect 25564 112354 25620 112364
rect 25340 112306 25396 112318
rect 25340 112254 25342 112306
rect 25394 112254 25396 112306
rect 25340 112084 25396 112254
rect 25340 112018 25396 112028
rect 25564 111860 25620 111870
rect 25564 111766 25620 111804
rect 25228 111694 25230 111746
rect 25282 111694 25284 111746
rect 25004 110798 25006 110850
rect 25058 110798 25060 110850
rect 25004 110786 25060 110798
rect 25228 110516 25284 111694
rect 25676 111300 25732 111310
rect 25564 111076 25620 111086
rect 25340 110738 25396 110750
rect 25340 110686 25342 110738
rect 25394 110686 25396 110738
rect 25340 110628 25396 110686
rect 25340 110562 25396 110572
rect 24892 110350 24894 110402
rect 24946 110350 24948 110402
rect 24892 110338 24948 110350
rect 25116 110460 25284 110516
rect 24668 110180 24724 110190
rect 24668 110086 24724 110124
rect 24464 109004 24728 109014
rect 24520 108948 24568 109004
rect 24624 108948 24672 109004
rect 24464 108938 24728 108948
rect 25116 108500 25172 110460
rect 25564 110402 25620 111020
rect 25676 110850 25732 111244
rect 25676 110798 25678 110850
rect 25730 110798 25732 110850
rect 25676 110786 25732 110798
rect 25564 110350 25566 110402
rect 25618 110350 25620 110402
rect 25564 110338 25620 110350
rect 25228 110292 25284 110302
rect 25228 110198 25284 110236
rect 25340 110068 25396 110078
rect 25228 109170 25284 109182
rect 25228 109118 25230 109170
rect 25282 109118 25284 109170
rect 25228 109060 25284 109118
rect 25228 108994 25284 109004
rect 25116 108406 25172 108444
rect 25116 107940 25172 107950
rect 24464 107436 24728 107446
rect 24520 107380 24568 107436
rect 24624 107380 24672 107436
rect 24464 107370 24728 107380
rect 25116 107266 25172 107884
rect 25116 107214 25118 107266
rect 25170 107214 25172 107266
rect 25116 106932 25172 107214
rect 25116 106866 25172 106876
rect 24464 105868 24728 105878
rect 24520 105812 24568 105868
rect 24624 105812 24672 105868
rect 24464 105802 24728 105812
rect 24220 105746 24276 105756
rect 23804 105084 24068 105094
rect 23860 105028 23908 105084
rect 23964 105028 24012 105084
rect 23804 105018 24068 105028
rect 24464 104300 24728 104310
rect 24520 104244 24568 104300
rect 24624 104244 24672 104300
rect 24464 104234 24728 104244
rect 23804 103516 24068 103526
rect 23860 103460 23908 103516
rect 23964 103460 24012 103516
rect 23804 103450 24068 103460
rect 24464 102732 24728 102742
rect 24520 102676 24568 102732
rect 24624 102676 24672 102732
rect 24464 102666 24728 102676
rect 23804 101948 24068 101958
rect 23860 101892 23908 101948
rect 23964 101892 24012 101948
rect 23804 101882 24068 101892
rect 24464 101164 24728 101174
rect 24520 101108 24568 101164
rect 24624 101108 24672 101164
rect 24464 101098 24728 101108
rect 23804 100380 24068 100390
rect 23860 100324 23908 100380
rect 23964 100324 24012 100380
rect 23804 100314 24068 100324
rect 24464 99596 24728 99606
rect 24520 99540 24568 99596
rect 24624 99540 24672 99596
rect 24464 99530 24728 99540
rect 23804 98812 24068 98822
rect 23860 98756 23908 98812
rect 23964 98756 24012 98812
rect 23804 98746 24068 98756
rect 24464 98028 24728 98038
rect 24520 97972 24568 98028
rect 24624 97972 24672 98028
rect 24464 97962 24728 97972
rect 22988 97412 23492 97468
rect 22876 95282 22932 95294
rect 22876 95230 22878 95282
rect 22930 95230 22932 95282
rect 22764 94500 22820 94510
rect 22428 94210 22484 94220
rect 22652 94498 22820 94500
rect 22652 94446 22766 94498
rect 22818 94446 22820 94498
rect 22652 94444 22820 94446
rect 22092 92094 22094 92146
rect 22146 92094 22148 92146
rect 22092 92082 22148 92094
rect 22204 94052 22372 94108
rect 21980 91634 22036 91644
rect 21532 90850 21588 90860
rect 21644 91196 21812 91252
rect 21532 90692 21588 90702
rect 21532 90466 21588 90636
rect 21532 90414 21534 90466
rect 21586 90414 21588 90466
rect 21532 90402 21588 90414
rect 21420 90188 21588 90244
rect 21420 89010 21476 89022
rect 21420 88958 21422 89010
rect 21474 88958 21476 89010
rect 21420 88228 21476 88958
rect 21420 88162 21476 88172
rect 21308 87948 21476 88004
rect 21308 87332 21364 87342
rect 20748 87220 20804 87230
rect 20748 87126 20804 87164
rect 20860 86658 20916 86670
rect 20860 86606 20862 86658
rect 20914 86606 20916 86658
rect 20860 86436 20916 86606
rect 20860 86370 20916 86380
rect 20860 86212 20916 86222
rect 20748 85764 20804 85802
rect 20748 85698 20804 85708
rect 20636 84366 20638 84418
rect 20690 84366 20692 84418
rect 20636 84354 20692 84366
rect 20860 83636 20916 86156
rect 21308 85764 21364 87276
rect 20972 85092 21028 85102
rect 20972 84306 21028 85036
rect 20972 84254 20974 84306
rect 21026 84254 21028 84306
rect 20972 84242 21028 84254
rect 21084 85090 21140 85102
rect 21084 85038 21086 85090
rect 21138 85038 21140 85090
rect 21084 84308 21140 85038
rect 21084 84242 21140 84252
rect 21196 84980 21252 84990
rect 20524 83580 20692 83636
rect 20412 83522 20468 83534
rect 20412 83470 20414 83522
rect 20466 83470 20468 83522
rect 20412 81956 20468 83470
rect 20412 81890 20468 81900
rect 20524 82180 20580 82190
rect 20300 80546 20356 80556
rect 20412 80500 20468 80510
rect 20524 80500 20580 82124
rect 20412 80498 20580 80500
rect 20412 80446 20414 80498
rect 20466 80446 20580 80498
rect 20412 80444 20580 80446
rect 20412 80434 20468 80444
rect 20300 78932 20356 78942
rect 20244 78930 20356 78932
rect 20244 78878 20302 78930
rect 20354 78878 20356 78930
rect 20244 78876 20356 78878
rect 20188 78838 20244 78876
rect 20300 78866 20356 78876
rect 20524 78820 20580 80444
rect 20636 79714 20692 83580
rect 20748 83634 20916 83636
rect 20748 83582 20862 83634
rect 20914 83582 20916 83634
rect 20748 83580 20916 83582
rect 20748 79828 20804 83580
rect 20860 83570 20916 83580
rect 21196 82180 21252 84924
rect 21196 82114 21252 82124
rect 21196 81956 21252 81966
rect 21084 81732 21140 81742
rect 20972 81730 21140 81732
rect 20972 81678 21086 81730
rect 21138 81678 21140 81730
rect 20972 81676 21140 81678
rect 20860 81284 20916 81294
rect 20860 81190 20916 81228
rect 20860 80388 20916 80398
rect 20972 80388 21028 81676
rect 21084 81666 21140 81676
rect 21196 81172 21252 81900
rect 21196 81058 21252 81116
rect 21196 81006 21198 81058
rect 21250 81006 21252 81058
rect 21196 80994 21252 81006
rect 21308 81060 21364 85708
rect 21420 85708 21476 87948
rect 21532 85876 21588 90188
rect 21532 85810 21588 85820
rect 21420 85652 21588 85708
rect 21420 85090 21476 85102
rect 21420 85038 21422 85090
rect 21474 85038 21476 85090
rect 21420 84980 21476 85038
rect 21420 84914 21476 84924
rect 21308 80994 21364 81004
rect 21420 84756 21476 84766
rect 21420 84306 21476 84700
rect 21420 84254 21422 84306
rect 21474 84254 21476 84306
rect 21420 80836 21476 84254
rect 21532 81284 21588 85652
rect 21644 84756 21700 91196
rect 22092 91140 22148 91150
rect 21868 90916 21924 90926
rect 21756 90804 21812 90814
rect 21756 88450 21812 90748
rect 21756 88398 21758 88450
rect 21810 88398 21812 88450
rect 21756 87332 21812 88398
rect 21756 87266 21812 87276
rect 21868 87330 21924 90860
rect 22092 90466 22148 91084
rect 22204 90916 22260 94052
rect 22204 90850 22260 90860
rect 22316 92932 22372 92942
rect 22652 92932 22708 94444
rect 22764 94434 22820 94444
rect 22764 94276 22820 94286
rect 22764 93826 22820 94220
rect 22764 93774 22766 93826
rect 22818 93774 22820 93826
rect 22764 93762 22820 93774
rect 22764 92932 22820 92942
rect 22652 92930 22820 92932
rect 22652 92878 22766 92930
rect 22818 92878 22820 92930
rect 22652 92876 22820 92878
rect 22316 90690 22372 92876
rect 22652 92148 22708 92158
rect 22652 92054 22708 92092
rect 22764 91364 22820 92876
rect 22876 92146 22932 95230
rect 22876 92094 22878 92146
rect 22930 92094 22932 92146
rect 22876 92082 22932 92094
rect 22764 91308 22932 91364
rect 22764 91140 22820 91150
rect 22764 91046 22820 91084
rect 22316 90638 22318 90690
rect 22370 90638 22372 90690
rect 22316 90626 22372 90638
rect 22092 90414 22094 90466
rect 22146 90414 22148 90466
rect 22092 90402 22148 90414
rect 22204 90580 22260 90590
rect 21980 89012 22036 89022
rect 21980 88898 22036 88956
rect 21980 88846 21982 88898
rect 22034 88846 22036 88898
rect 21980 88834 22036 88846
rect 21868 87278 21870 87330
rect 21922 87278 21924 87330
rect 21868 86884 21924 87278
rect 21868 86818 21924 86828
rect 21868 86658 21924 86670
rect 21868 86606 21870 86658
rect 21922 86606 21924 86658
rect 21868 86212 21924 86606
rect 21868 86146 21924 86156
rect 21644 84690 21700 84700
rect 21868 85650 21924 85662
rect 21868 85598 21870 85650
rect 21922 85598 21924 85650
rect 21644 84532 21700 84542
rect 21644 84194 21700 84476
rect 21644 84142 21646 84194
rect 21698 84142 21700 84194
rect 21644 84130 21700 84142
rect 21644 81732 21700 81742
rect 21644 81730 21812 81732
rect 21644 81678 21646 81730
rect 21698 81678 21812 81730
rect 21644 81676 21812 81678
rect 21644 81666 21700 81676
rect 21532 81228 21700 81284
rect 21308 80780 21476 80836
rect 21532 81060 21588 81070
rect 20860 80386 21028 80388
rect 20860 80334 20862 80386
rect 20914 80334 21028 80386
rect 20860 80332 21028 80334
rect 21196 80386 21252 80398
rect 21196 80334 21198 80386
rect 21250 80334 21252 80386
rect 20860 80322 20916 80332
rect 20748 79772 20916 79828
rect 20636 79662 20638 79714
rect 20690 79662 20692 79714
rect 20636 79650 20692 79662
rect 20412 78764 20524 78820
rect 20300 78596 20356 78606
rect 20188 77700 20244 77710
rect 20188 77474 20244 77644
rect 20188 77422 20190 77474
rect 20242 77422 20244 77474
rect 20188 77410 20244 77422
rect 20076 75854 20078 75906
rect 20130 75854 20132 75906
rect 20076 75842 20132 75854
rect 20188 75460 20244 75470
rect 20188 74116 20244 75404
rect 20076 72548 20132 72558
rect 20076 72454 20132 72492
rect 19964 71988 20020 71998
rect 19964 71894 20020 71932
rect 19852 70466 19908 70476
rect 20188 70196 20244 74060
rect 20300 73948 20356 78540
rect 20412 77364 20468 78764
rect 20524 78754 20580 78764
rect 20748 79604 20804 79614
rect 20748 78818 20804 79548
rect 20748 78766 20750 78818
rect 20802 78766 20804 78818
rect 20748 78754 20804 78766
rect 20860 78148 20916 79772
rect 20972 79604 21028 79614
rect 20972 79510 21028 79548
rect 21084 78818 21140 78830
rect 21084 78766 21086 78818
rect 21138 78766 21140 78818
rect 21084 78596 21140 78766
rect 21084 78530 21140 78540
rect 20412 77298 20468 77308
rect 20524 78092 20916 78148
rect 20524 76356 20580 78092
rect 21196 78036 21252 80334
rect 21308 79604 21364 80780
rect 21420 80612 21476 80622
rect 21420 80518 21476 80556
rect 21420 79604 21476 79614
rect 21308 79602 21476 79604
rect 21308 79550 21422 79602
rect 21474 79550 21476 79602
rect 21308 79548 21476 79550
rect 20860 77980 21252 78036
rect 21308 78930 21364 78942
rect 21308 78878 21310 78930
rect 21362 78878 21364 78930
rect 20748 77810 20804 77822
rect 20748 77758 20750 77810
rect 20802 77758 20804 77810
rect 20748 77588 20804 77758
rect 20748 77522 20804 77532
rect 20748 77364 20804 77374
rect 20636 77252 20692 77262
rect 20636 77158 20692 77196
rect 20748 76468 20804 77308
rect 20524 76290 20580 76300
rect 20636 76412 20804 76468
rect 20412 75796 20468 75806
rect 20636 75796 20692 76412
rect 20748 76244 20804 76254
rect 20748 76150 20804 76188
rect 20748 75796 20804 75806
rect 20636 75794 20804 75796
rect 20636 75742 20750 75794
rect 20802 75742 20804 75794
rect 20636 75740 20804 75742
rect 20412 75702 20468 75740
rect 20524 75012 20580 75022
rect 20300 73892 20468 73948
rect 20188 70130 20244 70140
rect 19740 70030 19742 70082
rect 19794 70030 19796 70082
rect 19740 70018 19796 70030
rect 20076 69972 20132 69982
rect 20076 69878 20132 69916
rect 19404 67778 19460 67788
rect 19516 68796 19684 68852
rect 19404 67172 19460 67182
rect 19348 67170 19460 67172
rect 19348 67118 19406 67170
rect 19458 67118 19460 67170
rect 19348 67116 19460 67118
rect 19292 67078 19348 67116
rect 19404 67106 19460 67116
rect 19516 66948 19572 68796
rect 19964 68740 20020 68750
rect 19964 68646 20020 68684
rect 19628 68626 19684 68638
rect 19628 68574 19630 68626
rect 19682 68574 19684 68626
rect 19628 67284 19684 68574
rect 19740 68626 19796 68638
rect 19740 68574 19742 68626
rect 19794 68574 19796 68626
rect 19740 67396 19796 68574
rect 20076 68628 20132 68638
rect 20076 68534 20132 68572
rect 20188 68292 20244 68302
rect 19964 67842 20020 67854
rect 19964 67790 19966 67842
rect 20018 67790 20020 67842
rect 19964 67508 20020 67790
rect 19964 67442 20020 67452
rect 19740 67330 19796 67340
rect 19628 67218 19684 67228
rect 19180 66446 19182 66498
rect 19234 66446 19236 66498
rect 19180 66434 19236 66446
rect 19404 66892 19572 66948
rect 19068 65986 19124 65996
rect 18844 64876 19012 64932
rect 18844 64706 18900 64718
rect 18844 64654 18846 64706
rect 18898 64654 18900 64706
rect 18732 63812 18788 63822
rect 18732 63718 18788 63756
rect 18620 63420 18788 63476
rect 18620 62914 18676 62926
rect 18620 62862 18622 62914
rect 18674 62862 18676 62914
rect 18620 61570 18676 62862
rect 18620 61518 18622 61570
rect 18674 61518 18676 61570
rect 18620 61506 18676 61518
rect 18508 60722 18564 60732
rect 18732 61460 18788 63420
rect 18732 60676 18788 61404
rect 18732 60610 18788 60620
rect 18284 59826 18340 59836
rect 18508 60002 18564 60014
rect 18508 59950 18510 60002
rect 18562 59950 18564 60002
rect 18508 59442 18564 59950
rect 18732 60004 18788 60014
rect 18732 59556 18788 59948
rect 18732 59490 18788 59500
rect 18508 59390 18510 59442
rect 18562 59390 18564 59442
rect 18508 59378 18564 59390
rect 18844 55468 18900 64654
rect 18956 63252 19012 64876
rect 19068 64820 19124 64830
rect 19068 64726 19124 64764
rect 19180 63700 19236 63710
rect 19068 63252 19124 63262
rect 18956 63250 19124 63252
rect 18956 63198 19070 63250
rect 19122 63198 19124 63250
rect 18956 63196 19124 63198
rect 18956 62244 19012 62254
rect 18956 61570 19012 62188
rect 19068 62132 19124 63196
rect 19068 61796 19124 62076
rect 19068 61730 19124 61740
rect 19180 61794 19236 63644
rect 19180 61742 19182 61794
rect 19234 61742 19236 61794
rect 19180 61730 19236 61742
rect 18956 61518 18958 61570
rect 19010 61518 19012 61570
rect 18956 61506 19012 61518
rect 19068 61124 19124 61134
rect 18956 60004 19012 60014
rect 18956 59910 19012 59948
rect 18732 55412 18900 55468
rect 18956 59332 19012 59342
rect 18956 57762 19012 59276
rect 19068 58434 19124 61068
rect 19292 60788 19348 60798
rect 19292 60694 19348 60732
rect 19292 60228 19348 60238
rect 19068 58382 19070 58434
rect 19122 58382 19124 58434
rect 19068 58370 19124 58382
rect 19180 59556 19236 59566
rect 18956 57710 18958 57762
rect 19010 57710 19012 57762
rect 18956 57090 19012 57710
rect 18956 57038 18958 57090
rect 19010 57038 19012 57090
rect 18956 56194 19012 57038
rect 18956 56142 18958 56194
rect 19010 56142 19012 56194
rect 18956 55522 19012 56142
rect 18956 55470 18958 55522
rect 19010 55470 19012 55522
rect 18956 55458 19012 55470
rect 18732 54852 18788 55412
rect 18732 54786 18788 54796
rect 18172 54180 18228 54190
rect 18172 50428 18228 54124
rect 18396 50484 18452 50522
rect 18172 50372 18340 50428
rect 18396 50418 18452 50428
rect 18172 48018 18228 48030
rect 18172 47966 18174 48018
rect 18226 47966 18228 48018
rect 18172 47570 18228 47966
rect 18172 47518 18174 47570
rect 18226 47518 18228 47570
rect 18172 47506 18228 47518
rect 18060 45042 18116 45052
rect 18172 45666 18228 45678
rect 18172 45614 18174 45666
rect 18226 45614 18228 45666
rect 17836 44994 18004 44996
rect 17836 44942 17838 44994
rect 17890 44942 18004 44994
rect 17836 44940 18004 44942
rect 17836 44930 17892 44940
rect 17724 43708 17892 43764
rect 17612 43586 17668 43596
rect 17724 43538 17780 43550
rect 17724 43486 17726 43538
rect 17778 43486 17780 43538
rect 17724 43316 17780 43486
rect 17836 43428 17892 43708
rect 17836 43362 17892 43372
rect 17388 43260 17780 43316
rect 17612 41972 17668 43260
rect 17948 43204 18004 44940
rect 18172 43988 18228 45614
rect 18172 43922 18228 43932
rect 18284 43428 18340 50372
rect 18396 50148 18452 50158
rect 18396 49810 18452 50092
rect 18396 49758 18398 49810
rect 18450 49758 18452 49810
rect 18396 49746 18452 49758
rect 18956 48244 19012 48254
rect 18956 48130 19012 48188
rect 18956 48078 18958 48130
rect 19010 48078 19012 48130
rect 18956 48066 19012 48078
rect 18620 48018 18676 48030
rect 18620 47966 18622 48018
rect 18674 47966 18676 48018
rect 18620 46900 18676 47966
rect 18620 46834 18676 46844
rect 18732 47460 18788 47470
rect 17612 41906 17668 41916
rect 17724 43148 18004 43204
rect 18172 43426 18340 43428
rect 18172 43374 18286 43426
rect 18338 43374 18340 43426
rect 18172 43372 18340 43374
rect 17052 40898 17108 40908
rect 16716 40450 16772 40460
rect 17164 40516 17220 40526
rect 16940 40404 16996 40414
rect 16996 40348 17108 40404
rect 16940 40310 16996 40348
rect 16268 38612 16436 38668
rect 16156 37314 16212 37324
rect 16268 38388 16324 38398
rect 16268 37266 16324 38332
rect 16268 37214 16270 37266
rect 16322 37214 16324 37266
rect 16268 37202 16324 37214
rect 16044 36876 16212 36932
rect 16044 36708 16100 36718
rect 15932 36706 16100 36708
rect 15932 36654 16046 36706
rect 16098 36654 16100 36706
rect 15932 36652 16100 36654
rect 16044 36642 16100 36652
rect 16044 35586 16100 35598
rect 16044 35534 16046 35586
rect 16098 35534 16100 35586
rect 15708 35474 15764 35486
rect 15708 35422 15710 35474
rect 15762 35422 15764 35474
rect 15708 33460 15764 35422
rect 15932 35476 15988 35486
rect 15932 35382 15988 35420
rect 16044 35364 16100 35534
rect 16044 35298 16100 35308
rect 15932 35140 15988 35150
rect 15932 34914 15988 35084
rect 15932 34862 15934 34914
rect 15986 34862 15988 34914
rect 15932 34850 15988 34862
rect 15708 33394 15764 33404
rect 15260 31836 15428 31892
rect 15484 33180 15652 33236
rect 15148 31220 15204 31230
rect 15148 31126 15204 31164
rect 15036 30258 15092 30268
rect 14812 29314 14980 29316
rect 14812 29262 14814 29314
rect 14866 29262 14980 29314
rect 14812 29260 14980 29262
rect 14812 29250 14868 29260
rect 14700 28924 14868 28980
rect 14476 27806 14478 27858
rect 14530 27806 14532 27858
rect 14476 27794 14532 27806
rect 14588 28642 14644 28654
rect 14588 28590 14590 28642
rect 14642 28590 14644 28642
rect 14588 26908 14644 28590
rect 14700 28644 14756 28654
rect 14700 27186 14756 28588
rect 14700 27134 14702 27186
rect 14754 27134 14756 27186
rect 14700 27122 14756 27134
rect 14700 26964 14756 26974
rect 14588 26852 14756 26908
rect 14476 26292 14532 26302
rect 14476 26198 14532 26236
rect 14588 24948 14644 24958
rect 14700 24948 14756 26852
rect 14588 24946 14756 24948
rect 14588 24894 14590 24946
rect 14642 24894 14756 24946
rect 14588 24892 14756 24894
rect 14588 24882 14644 24892
rect 14476 24724 14532 24734
rect 14476 23938 14532 24668
rect 14812 24276 14868 28924
rect 14924 28868 14980 28878
rect 14924 27858 14980 28812
rect 14924 27806 14926 27858
rect 14978 27806 14980 27858
rect 14924 27794 14980 27806
rect 15036 28642 15092 28654
rect 15036 28590 15038 28642
rect 15090 28590 15092 28642
rect 15036 27636 15092 28590
rect 14924 27580 15092 27636
rect 15148 27634 15204 27646
rect 15148 27582 15150 27634
rect 15202 27582 15204 27634
rect 14924 25844 14980 27580
rect 15148 27412 15204 27582
rect 15260 27636 15316 31836
rect 15372 31668 15428 31678
rect 15372 31574 15428 31612
rect 15484 31444 15540 33180
rect 15820 33124 15876 33134
rect 15596 33122 15876 33124
rect 15596 33070 15822 33122
rect 15874 33070 15876 33122
rect 15596 33068 15876 33070
rect 15596 32562 15652 33068
rect 15820 33058 15876 33068
rect 15932 32564 15988 32574
rect 15596 32510 15598 32562
rect 15650 32510 15652 32562
rect 15596 32498 15652 32510
rect 15820 32562 15988 32564
rect 15820 32510 15934 32562
rect 15986 32510 15988 32562
rect 15820 32508 15988 32510
rect 15260 27570 15316 27580
rect 15372 31388 15540 31444
rect 15596 32340 15652 32350
rect 15036 27356 15204 27412
rect 15036 26964 15092 27356
rect 15148 27188 15204 27198
rect 15148 27094 15204 27132
rect 15260 27076 15316 27086
rect 15260 26982 15316 27020
rect 15036 26908 15204 26964
rect 15036 26068 15092 26078
rect 15036 25974 15092 26012
rect 14924 25778 14980 25788
rect 14476 23886 14478 23938
rect 14530 23886 14532 23938
rect 14476 23874 14532 23886
rect 14700 24220 14868 24276
rect 14924 25508 14980 25518
rect 14924 25284 14980 25452
rect 14364 23314 14420 23324
rect 14028 23266 14084 23278
rect 14028 23214 14030 23266
rect 14082 23214 14084 23266
rect 13916 23156 13972 23166
rect 13916 22930 13972 23100
rect 13916 22878 13918 22930
rect 13970 22878 13972 22930
rect 13916 22820 13972 22878
rect 13916 22754 13972 22764
rect 14028 22708 14084 23214
rect 14588 23156 14644 23194
rect 14588 23090 14644 23100
rect 14364 23044 14420 23054
rect 14364 22950 14420 22988
rect 14028 22652 14196 22708
rect 14140 22372 14196 22652
rect 14364 22372 14420 22382
rect 14140 22370 14420 22372
rect 14140 22318 14366 22370
rect 14418 22318 14420 22370
rect 14140 22316 14420 22318
rect 14364 22306 14420 22316
rect 13916 22148 13972 22158
rect 14364 22148 14420 22158
rect 13916 22146 14308 22148
rect 13916 22094 13918 22146
rect 13970 22094 14308 22146
rect 13916 22092 14308 22094
rect 13916 22082 13972 22092
rect 13804 21746 13860 21756
rect 14140 21588 14196 21598
rect 13804 21362 13860 21374
rect 13804 21310 13806 21362
rect 13858 21310 13860 21362
rect 13804 21252 13860 21310
rect 13804 21186 13860 21196
rect 13916 21140 13972 21150
rect 13692 20972 13860 21028
rect 13692 19908 13748 19918
rect 13692 19814 13748 19852
rect 13580 19460 13636 19470
rect 13580 19236 13636 19404
rect 13580 19142 13636 19180
rect 13468 18956 13636 19012
rect 13468 18340 13524 18350
rect 13468 18246 13524 18284
rect 13468 16098 13524 16110
rect 13468 16046 13470 16098
rect 13522 16046 13524 16098
rect 13468 14756 13524 16046
rect 13580 14980 13636 18956
rect 13804 17890 13860 20972
rect 13916 20804 13972 21084
rect 14140 21140 14196 21532
rect 14252 21586 14308 22092
rect 14252 21534 14254 21586
rect 14306 21534 14308 21586
rect 14252 21522 14308 21534
rect 14364 21588 14420 22092
rect 14700 21812 14756 24220
rect 14812 24052 14868 24062
rect 14812 23958 14868 23996
rect 14924 23492 14980 25228
rect 15148 23548 15204 26908
rect 14924 23426 14980 23436
rect 15036 23492 15204 23548
rect 15260 26292 15316 26302
rect 15260 23492 15316 26236
rect 15372 24052 15428 31388
rect 15484 30994 15540 31006
rect 15484 30942 15486 30994
rect 15538 30942 15540 30994
rect 15484 25620 15540 30942
rect 15596 27636 15652 32284
rect 15708 31556 15764 31566
rect 15708 30882 15764 31500
rect 15708 30830 15710 30882
rect 15762 30830 15764 30882
rect 15708 30818 15764 30830
rect 15820 29316 15876 32508
rect 15932 32498 15988 32508
rect 16156 32450 16212 36876
rect 16380 36484 16436 38612
rect 16156 32398 16158 32450
rect 16210 32398 16212 32450
rect 16156 32386 16212 32398
rect 16268 36428 16436 36484
rect 16492 38612 16660 38668
rect 16716 38834 16772 38846
rect 16716 38782 16718 38834
rect 16770 38782 16772 38834
rect 16268 32228 16324 36428
rect 16380 35700 16436 35710
rect 16380 35606 16436 35644
rect 16492 34132 16548 38612
rect 16716 37268 16772 38782
rect 16604 35586 16660 35598
rect 16604 35534 16606 35586
rect 16658 35534 16660 35586
rect 16604 34804 16660 35534
rect 16716 35028 16772 37212
rect 16828 36258 16884 36270
rect 16828 36206 16830 36258
rect 16882 36206 16884 36258
rect 16828 35700 16884 36206
rect 16940 36036 16996 36046
rect 16940 35922 16996 35980
rect 16940 35870 16942 35922
rect 16994 35870 16996 35922
rect 16940 35858 16996 35870
rect 17052 35812 17108 40348
rect 17164 40290 17220 40460
rect 17164 40238 17166 40290
rect 17218 40238 17220 40290
rect 17164 40226 17220 40238
rect 17388 40292 17444 40302
rect 17276 37268 17332 37278
rect 17276 37174 17332 37212
rect 17052 35746 17108 35756
rect 17276 36036 17332 36046
rect 16828 35476 16884 35644
rect 17164 35700 17220 35738
rect 17164 35634 17220 35644
rect 17164 35476 17220 35486
rect 16828 35410 16884 35420
rect 17052 35474 17220 35476
rect 17052 35422 17166 35474
rect 17218 35422 17220 35474
rect 17052 35420 17220 35422
rect 16716 34972 16884 35028
rect 16828 34916 16884 34972
rect 16828 34860 16996 34916
rect 16604 34738 16660 34748
rect 16716 34802 16772 34814
rect 16716 34750 16718 34802
rect 16770 34750 16772 34802
rect 16716 34468 16772 34750
rect 16828 34692 16884 34702
rect 16828 34598 16884 34636
rect 16716 34402 16772 34412
rect 16828 34244 16884 34254
rect 16828 34150 16884 34188
rect 16492 34066 16548 34076
rect 16380 33906 16436 33918
rect 16380 33854 16382 33906
rect 16434 33854 16436 33906
rect 16380 32564 16436 33854
rect 16716 33234 16772 33246
rect 16716 33182 16718 33234
rect 16770 33182 16772 33234
rect 16716 33124 16772 33182
rect 16828 33236 16884 33246
rect 16828 33142 16884 33180
rect 16716 33058 16772 33068
rect 16940 32900 16996 34860
rect 17052 33346 17108 35420
rect 17164 35410 17220 35420
rect 17276 35308 17332 35980
rect 17164 35252 17332 35308
rect 17388 35252 17444 40236
rect 17500 39956 17556 39966
rect 17500 38724 17556 39900
rect 17500 36820 17556 38668
rect 17500 36754 17556 36764
rect 17724 35924 17780 43148
rect 17836 42642 17892 42654
rect 17836 42590 17838 42642
rect 17890 42590 17892 42642
rect 17836 41972 17892 42590
rect 17836 41906 17892 41916
rect 18060 41748 18116 41758
rect 17836 41746 18116 41748
rect 17836 41694 18062 41746
rect 18114 41694 18116 41746
rect 17836 41692 18116 41694
rect 17836 40402 17892 41692
rect 18060 41682 18116 41692
rect 18172 41524 18228 43372
rect 18284 43362 18340 43372
rect 18508 44098 18564 44110
rect 18508 44046 18510 44098
rect 18562 44046 18564 44098
rect 18284 42756 18340 42766
rect 18508 42756 18564 44046
rect 18284 42754 18564 42756
rect 18284 42702 18286 42754
rect 18338 42702 18564 42754
rect 18284 42700 18564 42702
rect 18284 42690 18340 42700
rect 17836 40350 17838 40402
rect 17890 40350 17892 40402
rect 17836 40338 17892 40350
rect 17948 41468 18228 41524
rect 17836 38052 17892 38062
rect 17836 37044 17892 37996
rect 17948 37268 18004 41468
rect 18508 41186 18564 42700
rect 18508 41134 18510 41186
rect 18562 41134 18564 41186
rect 18508 41122 18564 41134
rect 18620 43428 18676 43438
rect 18620 42754 18676 43372
rect 18620 42702 18622 42754
rect 18674 42702 18676 42754
rect 18060 41074 18116 41086
rect 18060 41022 18062 41074
rect 18114 41022 18116 41074
rect 18060 37604 18116 41022
rect 18172 40404 18228 40414
rect 18172 40310 18228 40348
rect 18620 40292 18676 42702
rect 18732 41972 18788 47404
rect 18844 46002 18900 46014
rect 18844 45950 18846 46002
rect 18898 45950 18900 46002
rect 18844 44212 18900 45950
rect 18956 45890 19012 45902
rect 18956 45838 18958 45890
rect 19010 45838 19012 45890
rect 18956 45330 19012 45838
rect 18956 45278 18958 45330
rect 19010 45278 19012 45330
rect 18956 45266 19012 45278
rect 18844 44156 19124 44212
rect 18844 43988 18900 43998
rect 18844 42978 18900 43932
rect 18844 42926 18846 42978
rect 18898 42926 18900 42978
rect 18844 42914 18900 42926
rect 18732 41906 18788 41916
rect 18956 41858 19012 41870
rect 18956 41806 18958 41858
rect 19010 41806 19012 41858
rect 18844 41186 18900 41198
rect 18844 41134 18846 41186
rect 18898 41134 18900 41186
rect 18844 40852 18900 41134
rect 18844 40786 18900 40796
rect 18956 40516 19012 41806
rect 19068 41410 19124 44156
rect 19068 41358 19070 41410
rect 19122 41358 19124 41410
rect 19068 41346 19124 41358
rect 19180 40740 19236 59500
rect 19292 53844 19348 60172
rect 19404 60004 19460 66892
rect 19964 66500 20020 66510
rect 19852 66274 19908 66286
rect 19852 66222 19854 66274
rect 19906 66222 19908 66274
rect 19852 65714 19908 66222
rect 19852 65662 19854 65714
rect 19906 65662 19908 65714
rect 19852 65650 19908 65662
rect 19628 64706 19684 64718
rect 19628 64654 19630 64706
rect 19682 64654 19684 64706
rect 19628 64036 19684 64654
rect 19516 63138 19572 63150
rect 19516 63086 19518 63138
rect 19570 63086 19572 63138
rect 19516 62580 19572 63086
rect 19628 62916 19684 63980
rect 19852 63700 19908 63710
rect 19628 62850 19684 62860
rect 19740 63698 19908 63700
rect 19740 63646 19854 63698
rect 19906 63646 19908 63698
rect 19740 63644 19908 63646
rect 19628 62580 19684 62590
rect 19516 62578 19684 62580
rect 19516 62526 19630 62578
rect 19682 62526 19684 62578
rect 19516 62524 19684 62526
rect 19628 62514 19684 62524
rect 19740 61570 19796 63644
rect 19852 63634 19908 63644
rect 19964 63138 20020 66444
rect 20188 66274 20244 68236
rect 20412 67956 20468 73892
rect 20524 73220 20580 74956
rect 20636 74114 20692 74126
rect 20636 74062 20638 74114
rect 20690 74062 20692 74114
rect 20636 73444 20692 74062
rect 20636 73378 20692 73388
rect 20636 73220 20692 73230
rect 20524 73218 20692 73220
rect 20524 73166 20638 73218
rect 20690 73166 20692 73218
rect 20524 73164 20692 73166
rect 20636 73154 20692 73164
rect 20412 67890 20468 67900
rect 20524 72436 20580 72446
rect 20748 72436 20804 75740
rect 20860 72772 20916 77980
rect 21196 77588 21252 77598
rect 21196 77362 21252 77532
rect 21196 77310 21198 77362
rect 21250 77310 21252 77362
rect 21196 77298 21252 77310
rect 20972 77140 21028 77150
rect 21308 77140 21364 78878
rect 21420 77364 21476 79548
rect 21420 77298 21476 77308
rect 20972 77138 21364 77140
rect 20972 77086 20974 77138
rect 21026 77086 21364 77138
rect 20972 77084 21364 77086
rect 20972 77074 21028 77084
rect 21532 77028 21588 81004
rect 21644 79604 21700 81228
rect 21756 80500 21812 81676
rect 21868 80724 21924 85598
rect 21980 85652 22036 85662
rect 21980 81284 22036 85596
rect 22092 84308 22148 84318
rect 22092 83746 22148 84252
rect 22092 83694 22094 83746
rect 22146 83694 22148 83746
rect 22092 83682 22148 83694
rect 22036 81228 22148 81284
rect 21980 81218 22036 81228
rect 21868 80658 21924 80668
rect 21868 80500 21924 80510
rect 21756 80498 21924 80500
rect 21756 80446 21870 80498
rect 21922 80446 21924 80498
rect 21756 80444 21924 80446
rect 21868 80434 21924 80444
rect 21980 80500 22036 80510
rect 21980 80276 22036 80444
rect 21868 80220 22036 80276
rect 21644 79548 21812 79604
rect 21644 79378 21700 79390
rect 21644 79326 21646 79378
rect 21698 79326 21700 79378
rect 21644 77362 21700 79326
rect 21644 77310 21646 77362
rect 21698 77310 21700 77362
rect 21644 77298 21700 77310
rect 21196 76972 21588 77028
rect 21084 76244 21140 76254
rect 21084 75682 21140 76188
rect 21084 75630 21086 75682
rect 21138 75630 21140 75682
rect 21084 75618 21140 75630
rect 21084 74116 21140 74126
rect 20972 73108 21028 73118
rect 20972 73014 21028 73052
rect 20860 72716 21028 72772
rect 20860 72548 20916 72558
rect 20860 72454 20916 72492
rect 20524 72434 20804 72436
rect 20524 72382 20526 72434
rect 20578 72382 20804 72434
rect 20524 72380 20804 72382
rect 20412 67730 20468 67742
rect 20412 67678 20414 67730
rect 20466 67678 20468 67730
rect 20412 67060 20468 67678
rect 20412 66994 20468 67004
rect 20188 66222 20190 66274
rect 20242 66222 20244 66274
rect 20188 66210 20244 66222
rect 20524 66052 20580 72380
rect 20860 71652 20916 71662
rect 20636 70084 20692 70094
rect 20636 68738 20692 70028
rect 20636 68686 20638 68738
rect 20690 68686 20692 68738
rect 20636 68404 20692 68686
rect 20636 68338 20692 68348
rect 20748 69186 20804 69198
rect 20748 69134 20750 69186
rect 20802 69134 20804 69186
rect 20748 68068 20804 69134
rect 20748 68002 20804 68012
rect 20188 65996 20580 66052
rect 20636 67956 20692 67966
rect 20076 64818 20132 64830
rect 20076 64766 20078 64818
rect 20130 64766 20132 64818
rect 20076 63588 20132 64766
rect 20076 63522 20132 63532
rect 20076 63364 20132 63374
rect 20188 63364 20244 65996
rect 20636 65940 20692 67900
rect 20748 67844 20804 67854
rect 20748 67750 20804 67788
rect 20076 63362 20244 63364
rect 20076 63310 20078 63362
rect 20130 63310 20244 63362
rect 20076 63308 20244 63310
rect 20300 65884 20692 65940
rect 20748 67172 20804 67182
rect 20076 63298 20132 63308
rect 20300 63252 20356 65884
rect 20636 65268 20692 65278
rect 19964 63086 19966 63138
rect 20018 63086 20020 63138
rect 19740 61518 19742 61570
rect 19794 61518 19796 61570
rect 19740 61506 19796 61518
rect 19852 62916 19908 62926
rect 19404 59948 19572 60004
rect 19404 58548 19460 58558
rect 19404 58454 19460 58492
rect 19292 53778 19348 53788
rect 19516 57316 19572 59948
rect 19292 52052 19348 52062
rect 19292 44322 19348 51996
rect 19516 50036 19572 57260
rect 19404 49026 19460 49038
rect 19404 48974 19406 49026
rect 19458 48974 19460 49026
rect 19404 47796 19460 48974
rect 19404 47730 19460 47740
rect 19516 44548 19572 49980
rect 19740 49140 19796 49150
rect 19740 49046 19796 49084
rect 19740 47458 19796 47470
rect 19740 47406 19742 47458
rect 19794 47406 19796 47458
rect 19740 47348 19796 47406
rect 19740 47282 19796 47292
rect 19516 44482 19572 44492
rect 19740 45780 19796 45790
rect 19852 45780 19908 62860
rect 19964 62692 20020 63086
rect 19964 59332 20020 62636
rect 20188 63196 20356 63252
rect 20412 65266 20692 65268
rect 20412 65214 20638 65266
rect 20690 65214 20692 65266
rect 20412 65212 20692 65214
rect 20188 62244 20244 63196
rect 20412 63140 20468 65212
rect 20636 65202 20692 65212
rect 20748 63812 20804 67116
rect 20748 63746 20804 63756
rect 20188 62178 20244 62188
rect 20300 63084 20468 63140
rect 20748 63138 20804 63150
rect 20748 63086 20750 63138
rect 20802 63086 20804 63138
rect 20076 60004 20132 60014
rect 20076 60002 20244 60004
rect 20076 59950 20078 60002
rect 20130 59950 20244 60002
rect 20076 59948 20244 59950
rect 20076 59938 20132 59948
rect 20188 59556 20244 59948
rect 20188 59490 20244 59500
rect 19964 59266 20020 59276
rect 20300 53956 20356 63084
rect 20636 62242 20692 62254
rect 20636 62190 20638 62242
rect 20690 62190 20692 62242
rect 20636 62020 20692 62190
rect 20524 61964 20636 62020
rect 20524 61684 20580 61964
rect 20636 61954 20692 61964
rect 20524 61618 20580 61628
rect 20636 61796 20692 61806
rect 20412 61570 20468 61582
rect 20412 61518 20414 61570
rect 20466 61518 20468 61570
rect 20412 60900 20468 61518
rect 20412 60834 20468 60844
rect 20636 60898 20692 61740
rect 20636 60846 20638 60898
rect 20690 60846 20692 60898
rect 20636 60834 20692 60846
rect 20300 53890 20356 53900
rect 20412 60676 20468 60686
rect 20300 51940 20356 51950
rect 20188 49028 20244 49038
rect 20188 47012 20244 48972
rect 20188 46946 20244 46956
rect 20076 46002 20132 46014
rect 20076 45950 20078 46002
rect 20130 45950 20132 46002
rect 20076 45892 20132 45950
rect 20076 45826 20132 45836
rect 19740 45778 19908 45780
rect 19740 45726 19742 45778
rect 19794 45726 19908 45778
rect 19740 45724 19908 45726
rect 19740 45220 19796 45724
rect 19292 44270 19294 44322
rect 19346 44270 19348 44322
rect 19292 44258 19348 44270
rect 19404 44212 19460 44222
rect 19404 44118 19460 44156
rect 19740 44100 19796 45164
rect 19852 44548 19908 44558
rect 19852 44454 19908 44492
rect 19740 44034 19796 44044
rect 19404 43314 19460 43326
rect 19404 43262 19406 43314
rect 19458 43262 19460 43314
rect 19404 42754 19460 43262
rect 19852 42756 19908 42766
rect 19404 42702 19406 42754
rect 19458 42702 19460 42754
rect 19292 41860 19348 41870
rect 19292 41766 19348 41804
rect 19404 41300 19460 42702
rect 19740 42754 19908 42756
rect 19740 42702 19854 42754
rect 19906 42702 19908 42754
rect 19740 42700 19908 42702
rect 19740 42084 19796 42700
rect 19852 42690 19908 42700
rect 20188 42756 20244 42766
rect 19628 41970 19684 41982
rect 19628 41918 19630 41970
rect 19682 41918 19684 41970
rect 19628 41860 19684 41918
rect 19628 41794 19684 41804
rect 19516 41300 19572 41310
rect 19404 41298 19572 41300
rect 19404 41246 19518 41298
rect 19570 41246 19572 41298
rect 19404 41244 19572 41246
rect 19516 41234 19572 41244
rect 19180 40684 19348 40740
rect 18956 40450 19012 40460
rect 18620 40226 18676 40236
rect 19180 40402 19236 40414
rect 19180 40350 19182 40402
rect 19234 40350 19236 40402
rect 19180 38668 19236 40350
rect 18508 38612 19236 38668
rect 18060 37538 18116 37548
rect 18396 38276 18452 38286
rect 18396 37940 18452 38220
rect 17948 37202 18004 37212
rect 18060 37268 18116 37278
rect 18060 37266 18340 37268
rect 18060 37214 18062 37266
rect 18114 37214 18340 37266
rect 18060 37212 18340 37214
rect 18060 37202 18116 37212
rect 17836 36988 18228 37044
rect 18060 36820 18116 36830
rect 17948 36708 18004 36718
rect 17948 36614 18004 36652
rect 17724 35858 17780 35868
rect 17612 35812 17668 35822
rect 17164 34914 17220 35252
rect 17388 35186 17444 35196
rect 17500 35476 17556 35486
rect 17500 35028 17556 35420
rect 17388 35026 17556 35028
rect 17388 34974 17502 35026
rect 17554 34974 17556 35026
rect 17388 34972 17556 34974
rect 17164 34862 17166 34914
rect 17218 34862 17220 34914
rect 17164 34850 17220 34862
rect 17276 34916 17332 34926
rect 17276 34822 17332 34860
rect 17052 33294 17054 33346
rect 17106 33294 17108 33346
rect 17052 33282 17108 33294
rect 17164 34132 17220 34142
rect 16716 32844 16996 32900
rect 16380 32498 16436 32508
rect 16604 32564 16660 32574
rect 16604 32470 16660 32508
rect 16044 32172 16324 32228
rect 16044 31890 16100 32172
rect 16044 31838 16046 31890
rect 16098 31838 16100 31890
rect 15932 31668 15988 31678
rect 15932 30772 15988 31612
rect 16044 31332 16100 31838
rect 16156 31780 16212 31790
rect 16156 31686 16212 31724
rect 16044 31266 16100 31276
rect 16156 31444 16212 31454
rect 16044 30884 16100 30894
rect 16044 30790 16100 30828
rect 15932 30706 15988 30716
rect 16156 30548 16212 31388
rect 16604 30994 16660 31006
rect 16604 30942 16606 30994
rect 16658 30942 16660 30994
rect 15932 30492 16212 30548
rect 16380 30772 16436 30782
rect 15932 30322 15988 30492
rect 16268 30436 16324 30446
rect 16268 30342 16324 30380
rect 15932 30270 15934 30322
rect 15986 30270 15988 30322
rect 15932 30258 15988 30270
rect 16044 30324 16100 30334
rect 16044 30230 16100 30268
rect 15708 29260 15876 29316
rect 15708 28868 15764 29260
rect 15932 29204 15988 29214
rect 15708 28802 15764 28812
rect 15820 29202 15988 29204
rect 15820 29150 15934 29202
rect 15986 29150 15988 29202
rect 15820 29148 15988 29150
rect 15820 27858 15876 29148
rect 15932 29138 15988 29148
rect 15820 27806 15822 27858
rect 15874 27806 15876 27858
rect 15820 27794 15876 27806
rect 15932 28642 15988 28654
rect 15932 28590 15934 28642
rect 15986 28590 15988 28642
rect 15596 27580 15876 27636
rect 15708 27074 15764 27086
rect 15708 27022 15710 27074
rect 15762 27022 15764 27074
rect 15708 26964 15764 27022
rect 15708 26898 15764 26908
rect 15820 26292 15876 27580
rect 15820 26226 15876 26236
rect 15820 26068 15876 26078
rect 15596 25844 15652 25854
rect 15596 25730 15652 25788
rect 15596 25678 15598 25730
rect 15650 25678 15652 25730
rect 15596 25666 15652 25678
rect 15484 25554 15540 25564
rect 15708 25508 15764 25518
rect 15708 25414 15764 25452
rect 15820 25506 15876 26012
rect 15820 25454 15822 25506
rect 15874 25454 15876 25506
rect 15820 25172 15876 25454
rect 15932 25284 15988 28590
rect 16156 28420 16212 28430
rect 16156 27858 16212 28364
rect 16156 27806 16158 27858
rect 16210 27806 16212 27858
rect 16156 27794 16212 27806
rect 16156 27636 16212 27646
rect 16156 27186 16212 27580
rect 16156 27134 16158 27186
rect 16210 27134 16212 27186
rect 16156 26852 16212 27134
rect 16156 26786 16212 26796
rect 16268 27076 16324 27086
rect 16156 26516 16212 26526
rect 16268 26516 16324 27020
rect 16156 26514 16324 26516
rect 16156 26462 16158 26514
rect 16210 26462 16324 26514
rect 16156 26460 16324 26462
rect 16156 26450 16212 26460
rect 16380 26292 16436 30716
rect 16604 30436 16660 30942
rect 16604 30370 16660 30380
rect 16716 26740 16772 32844
rect 17164 32788 17220 34076
rect 17276 34132 17332 34142
rect 17388 34132 17444 34972
rect 17500 34962 17556 34972
rect 17612 34916 17668 35756
rect 17836 35812 17892 35822
rect 17724 35700 17780 35710
rect 17836 35700 17892 35756
rect 17724 35698 17892 35700
rect 17724 35646 17726 35698
rect 17778 35646 17892 35698
rect 17724 35644 17892 35646
rect 17724 35140 17780 35644
rect 18060 35586 18116 36764
rect 18060 35534 18062 35586
rect 18114 35534 18116 35586
rect 18060 35522 18116 35534
rect 17724 35074 17780 35084
rect 17948 35364 18004 35374
rect 17836 35028 17892 35038
rect 17836 34934 17892 34972
rect 17612 34860 17780 34916
rect 17612 34132 17668 34142
rect 17276 34130 17556 34132
rect 17276 34078 17278 34130
rect 17330 34078 17556 34130
rect 17276 34076 17556 34078
rect 17276 34066 17332 34076
rect 17500 33684 17556 34076
rect 17612 34038 17668 34076
rect 17724 33796 17780 34860
rect 17836 34132 17892 34142
rect 17948 34132 18004 35308
rect 18060 34914 18116 34926
rect 18060 34862 18062 34914
rect 18114 34862 18116 34914
rect 18060 34804 18116 34862
rect 18060 34738 18116 34748
rect 18172 34802 18228 36988
rect 18284 36372 18340 37212
rect 18396 37154 18452 37884
rect 18396 37102 18398 37154
rect 18450 37102 18452 37154
rect 18396 37090 18452 37102
rect 18396 36372 18452 36382
rect 18284 36370 18452 36372
rect 18284 36318 18398 36370
rect 18450 36318 18452 36370
rect 18284 36316 18452 36318
rect 18172 34750 18174 34802
rect 18226 34750 18228 34802
rect 18172 34738 18228 34750
rect 18284 36036 18340 36046
rect 18172 34132 18228 34142
rect 17948 34076 18116 34132
rect 17836 34018 17892 34076
rect 17836 33966 17838 34018
rect 17890 33966 17892 34018
rect 17836 33954 17892 33966
rect 18060 33908 18116 34076
rect 17948 33852 18116 33908
rect 17724 33740 17892 33796
rect 16940 32732 17220 32788
rect 17388 33628 17780 33684
rect 16828 29540 16884 29550
rect 16828 29446 16884 29484
rect 16940 29428 16996 32732
rect 17276 32564 17332 32574
rect 17276 32470 17332 32508
rect 17388 31890 17444 33628
rect 17724 33570 17780 33628
rect 17724 33518 17726 33570
rect 17778 33518 17780 33570
rect 17500 33346 17556 33358
rect 17500 33294 17502 33346
rect 17554 33294 17556 33346
rect 17500 33236 17556 33294
rect 17724 33348 17780 33518
rect 17724 33282 17780 33292
rect 17500 32900 17556 33180
rect 17500 32834 17556 32844
rect 17612 33234 17668 33246
rect 17612 33182 17614 33234
rect 17666 33182 17668 33234
rect 17388 31838 17390 31890
rect 17442 31838 17444 31890
rect 17388 31826 17444 31838
rect 17052 31780 17108 31818
rect 17108 31724 17332 31780
rect 17052 31714 17108 31724
rect 17052 31556 17108 31566
rect 17052 31462 17108 31500
rect 17164 31108 17220 31118
rect 17164 31014 17220 31052
rect 17052 30996 17108 31006
rect 17052 30324 17108 30940
rect 17276 30994 17332 31724
rect 17612 31778 17668 33182
rect 17612 31726 17614 31778
rect 17666 31726 17668 31778
rect 17612 31714 17668 31726
rect 17724 33124 17780 33134
rect 17724 31220 17780 33068
rect 17276 30942 17278 30994
rect 17330 30942 17332 30994
rect 17276 30930 17332 30942
rect 17388 31164 17780 31220
rect 17052 29428 17108 30268
rect 17276 30212 17332 30222
rect 17276 30118 17332 30156
rect 17276 29988 17332 29998
rect 17164 29428 17220 29438
rect 17052 29426 17220 29428
rect 17052 29374 17166 29426
rect 17218 29374 17220 29426
rect 17052 29372 17220 29374
rect 16940 29362 16996 29372
rect 17164 29362 17220 29372
rect 17164 27860 17220 27870
rect 17052 27858 17220 27860
rect 17052 27806 17166 27858
rect 17218 27806 17220 27858
rect 17052 27804 17220 27806
rect 17052 27300 17108 27804
rect 17164 27794 17220 27804
rect 16940 27188 16996 27198
rect 16940 27094 16996 27132
rect 16828 27076 16884 27086
rect 16828 26982 16884 27020
rect 16716 26674 16772 26684
rect 16380 26226 16436 26236
rect 17052 26180 17108 27244
rect 17164 26292 17220 26302
rect 17164 26198 17220 26236
rect 16828 26124 17108 26180
rect 16604 26068 16660 26078
rect 16604 25974 16660 26012
rect 16716 26066 16772 26078
rect 16716 26014 16718 26066
rect 16770 26014 16772 26066
rect 16716 25844 16772 26014
rect 16828 26066 16884 26124
rect 16828 26014 16830 26066
rect 16882 26014 16884 26066
rect 16828 26002 16884 26014
rect 16716 25788 16996 25844
rect 15932 25218 15988 25228
rect 16044 25618 16100 25630
rect 16044 25566 16046 25618
rect 16098 25566 16100 25618
rect 15372 23986 15428 23996
rect 15484 25116 15876 25172
rect 15484 23604 15540 25116
rect 16044 25060 16100 25566
rect 16268 25508 16324 25518
rect 16716 25508 16772 25518
rect 16268 25506 16772 25508
rect 16268 25454 16270 25506
rect 16322 25454 16718 25506
rect 16770 25454 16772 25506
rect 16268 25452 16772 25454
rect 16268 25442 16324 25452
rect 16716 25442 16772 25452
rect 16940 25506 16996 25788
rect 17276 25730 17332 29932
rect 17388 29652 17444 31164
rect 17388 29586 17444 29596
rect 17500 30996 17556 31006
rect 17388 29428 17444 29438
rect 17388 27972 17444 29372
rect 17500 28866 17556 30940
rect 17724 30882 17780 31164
rect 17724 30830 17726 30882
rect 17778 30830 17780 30882
rect 17724 30818 17780 30830
rect 17836 30660 17892 33740
rect 17948 32004 18004 33852
rect 18060 33684 18116 33694
rect 18060 33346 18116 33628
rect 18060 33294 18062 33346
rect 18114 33294 18116 33346
rect 18060 33236 18116 33294
rect 18060 33170 18116 33180
rect 18172 32788 18228 34076
rect 18284 34018 18340 35980
rect 18396 35812 18452 36316
rect 18396 35746 18452 35756
rect 18284 33966 18286 34018
rect 18338 33966 18340 34018
rect 18284 33684 18340 33966
rect 18284 33618 18340 33628
rect 18396 35588 18452 35598
rect 18284 33460 18340 33470
rect 18284 33366 18340 33404
rect 18172 32732 18340 32788
rect 18172 32564 18228 32574
rect 18172 32470 18228 32508
rect 18060 32004 18116 32014
rect 17948 32002 18116 32004
rect 17948 31950 18062 32002
rect 18114 31950 18116 32002
rect 17948 31948 18116 31950
rect 18060 31938 18116 31948
rect 18284 32002 18340 32732
rect 18284 31950 18286 32002
rect 18338 31950 18340 32002
rect 18284 31938 18340 31950
rect 17724 30604 17892 30660
rect 17948 31780 18004 31790
rect 17612 29988 17668 29998
rect 17612 29894 17668 29932
rect 17612 29428 17668 29438
rect 17612 29334 17668 29372
rect 17500 28814 17502 28866
rect 17554 28814 17556 28866
rect 17500 28802 17556 28814
rect 17388 26908 17444 27916
rect 17612 28756 17668 28766
rect 17612 27074 17668 28700
rect 17612 27022 17614 27074
rect 17666 27022 17668 27074
rect 17612 27010 17668 27022
rect 17724 26908 17780 30604
rect 17836 30436 17892 30446
rect 17836 30342 17892 30380
rect 17836 30212 17892 30222
rect 17836 30118 17892 30156
rect 17836 29316 17892 29326
rect 17948 29316 18004 31724
rect 18172 31668 18228 31678
rect 18396 31668 18452 35532
rect 18508 33572 18564 38612
rect 19292 38388 19348 40684
rect 19404 40292 19460 40302
rect 19404 38500 19460 40236
rect 19740 38668 19796 42028
rect 19964 41746 20020 41758
rect 19964 41694 19966 41746
rect 20018 41694 20020 41746
rect 19964 40404 20020 41694
rect 19964 40338 20020 40348
rect 20188 41186 20244 42700
rect 20188 41134 20190 41186
rect 20242 41134 20244 41186
rect 19740 38612 20020 38668
rect 19404 38444 19796 38500
rect 19292 38332 19460 38388
rect 18620 38276 18676 38286
rect 18620 38274 19348 38276
rect 18620 38222 18622 38274
rect 18674 38222 19348 38274
rect 18620 38220 19348 38222
rect 18620 38210 18676 38220
rect 18732 38050 18788 38062
rect 18732 37998 18734 38050
rect 18786 37998 18788 38050
rect 18620 37826 18676 37838
rect 18620 37774 18622 37826
rect 18674 37774 18676 37826
rect 18620 35028 18676 37774
rect 18732 37828 18788 37998
rect 19180 37938 19236 37950
rect 19180 37886 19182 37938
rect 19234 37886 19236 37938
rect 19068 37828 19124 37838
rect 18732 37826 19124 37828
rect 18732 37774 19070 37826
rect 19122 37774 19124 37826
rect 18732 37772 19124 37774
rect 18732 35364 18788 37772
rect 19068 37762 19124 37772
rect 19180 36596 19236 37886
rect 18732 35298 18788 35308
rect 19068 36258 19124 36270
rect 19068 36206 19070 36258
rect 19122 36206 19124 36258
rect 18620 34962 18676 34972
rect 18732 35140 18788 35150
rect 18732 34802 18788 35084
rect 19068 34916 19124 36206
rect 19180 35700 19236 36540
rect 19292 36036 19348 38220
rect 19404 37828 19460 38332
rect 19404 37762 19460 37772
rect 19516 38050 19572 38062
rect 19516 37998 19518 38050
rect 19570 37998 19572 38050
rect 19404 36260 19460 36270
rect 19404 36166 19460 36204
rect 19292 35922 19348 35980
rect 19292 35870 19294 35922
rect 19346 35870 19348 35922
rect 19292 35858 19348 35870
rect 19236 35644 19348 35700
rect 19180 35606 19236 35644
rect 19068 34850 19124 34860
rect 19180 35026 19236 35038
rect 19180 34974 19182 35026
rect 19234 34974 19236 35026
rect 18732 34750 18734 34802
rect 18786 34750 18788 34802
rect 18732 33796 18788 34750
rect 18956 34692 19012 34702
rect 19180 34692 19236 34974
rect 18844 34132 18900 34142
rect 18844 34038 18900 34076
rect 18732 33730 18788 33740
rect 18508 33516 18900 33572
rect 18508 33348 18564 33358
rect 18564 33292 18676 33348
rect 18508 33254 18564 33292
rect 18620 32564 18676 33292
rect 18732 33234 18788 33246
rect 18732 33182 18734 33234
rect 18786 33182 18788 33234
rect 18732 33124 18788 33182
rect 18732 33058 18788 33068
rect 18732 32564 18788 32574
rect 18620 32562 18788 32564
rect 18620 32510 18734 32562
rect 18786 32510 18788 32562
rect 18620 32508 18788 32510
rect 18732 32498 18788 32508
rect 18844 32564 18900 33516
rect 18956 33346 19012 34636
rect 19068 34636 19236 34692
rect 19068 34580 19124 34636
rect 19292 34580 19348 35644
rect 19068 34514 19124 34524
rect 19180 34524 19348 34580
rect 19404 35028 19460 35038
rect 19068 33572 19124 33610
rect 19068 33506 19124 33516
rect 18956 33294 18958 33346
rect 19010 33294 19012 33346
rect 18956 33012 19012 33294
rect 19180 33124 19236 34524
rect 19292 33572 19348 33582
rect 19292 33458 19348 33516
rect 19292 33406 19294 33458
rect 19346 33406 19348 33458
rect 19292 33394 19348 33406
rect 19180 33058 19236 33068
rect 18956 32946 19012 32956
rect 19292 32788 19348 32798
rect 19404 32788 19460 34972
rect 19516 33572 19572 37998
rect 19740 37156 19796 38444
rect 19852 38052 19908 38062
rect 19852 37958 19908 37996
rect 19628 37042 19684 37054
rect 19628 36990 19630 37042
rect 19682 36990 19684 37042
rect 19628 36596 19684 36990
rect 19628 36502 19684 36540
rect 19740 36372 19796 37100
rect 19964 36820 20020 38612
rect 20188 38388 20244 41134
rect 20188 38322 20244 38332
rect 20300 38276 20356 51884
rect 20412 44436 20468 60620
rect 20636 60228 20692 60238
rect 20748 60228 20804 63086
rect 20636 60226 20804 60228
rect 20636 60174 20638 60226
rect 20690 60174 20804 60226
rect 20636 60172 20804 60174
rect 20636 60162 20692 60172
rect 20636 59332 20692 59342
rect 20636 58658 20692 59276
rect 20636 58606 20638 58658
rect 20690 58606 20692 58658
rect 20636 58594 20692 58606
rect 20860 58548 20916 71596
rect 20972 68852 21028 72716
rect 21084 71764 21140 74060
rect 21084 71670 21140 71708
rect 21196 71652 21252 76972
rect 21532 76804 21588 76814
rect 21420 76468 21476 76478
rect 21308 76356 21364 76366
rect 21308 73948 21364 76300
rect 21420 74116 21476 76412
rect 21532 75682 21588 76748
rect 21756 76020 21812 79548
rect 21868 77922 21924 80220
rect 22092 79828 22148 81228
rect 22204 80836 22260 90524
rect 22652 90356 22708 90366
rect 22652 90262 22708 90300
rect 22876 89236 22932 91308
rect 22876 89170 22932 89180
rect 22988 89012 23044 97412
rect 23804 97244 24068 97254
rect 23860 97188 23908 97244
rect 23964 97188 24012 97244
rect 23804 97178 24068 97188
rect 24464 96460 24728 96470
rect 24520 96404 24568 96460
rect 24624 96404 24672 96460
rect 24464 96394 24728 96404
rect 23324 95842 23380 95854
rect 23324 95790 23326 95842
rect 23378 95790 23380 95842
rect 23324 95060 23380 95790
rect 23804 95676 24068 95686
rect 23860 95620 23908 95676
rect 23964 95620 24012 95676
rect 23804 95610 24068 95620
rect 23324 94994 23380 95004
rect 23772 95282 23828 95294
rect 23772 95230 23774 95282
rect 23826 95230 23828 95282
rect 23772 94836 23828 95230
rect 24892 95060 24948 95070
rect 24464 94892 24728 94902
rect 24520 94836 24568 94892
rect 24624 94836 24672 94892
rect 24464 94826 24728 94836
rect 23660 94724 23716 94734
rect 23660 94630 23716 94668
rect 23324 94612 23380 94622
rect 23324 94518 23380 94556
rect 23772 94276 23828 94780
rect 23660 94220 23828 94276
rect 23660 92148 23716 94220
rect 23804 94108 24068 94118
rect 23860 94052 23908 94108
rect 23964 94052 24012 94108
rect 23804 94042 24068 94052
rect 24464 93324 24728 93334
rect 24520 93268 24568 93324
rect 24624 93268 24672 93324
rect 24464 93258 24728 93268
rect 24668 93044 24724 93054
rect 24668 92950 24724 92988
rect 24892 92930 24948 95004
rect 24892 92878 24894 92930
rect 24946 92878 24948 92930
rect 24892 92866 24948 92878
rect 23804 92540 24068 92550
rect 23860 92484 23908 92540
rect 23964 92484 24012 92540
rect 23804 92474 24068 92484
rect 23660 92146 24276 92148
rect 23660 92094 23662 92146
rect 23714 92094 24276 92146
rect 23660 92092 24276 92094
rect 23660 92082 23716 92092
rect 23804 90972 24068 90982
rect 23860 90916 23908 90972
rect 23964 90916 24012 90972
rect 23804 90906 24068 90916
rect 23804 89404 24068 89414
rect 23860 89348 23908 89404
rect 23964 89348 24012 89404
rect 23804 89338 24068 89348
rect 22428 88956 23044 89012
rect 22316 87668 22372 87678
rect 22316 87554 22372 87612
rect 22316 87502 22318 87554
rect 22370 87502 22372 87554
rect 22316 85986 22372 87502
rect 22316 85934 22318 85986
rect 22370 85934 22372 85986
rect 22316 85922 22372 85934
rect 22428 82628 22484 88956
rect 23100 88788 23156 88798
rect 22764 88786 23156 88788
rect 22764 88734 23102 88786
rect 23154 88734 23156 88786
rect 22764 88732 23156 88734
rect 22652 86660 22708 86670
rect 22540 86434 22596 86446
rect 22540 86382 22542 86434
rect 22594 86382 22596 86434
rect 22540 86212 22596 86382
rect 22540 86146 22596 86156
rect 22540 85876 22596 85886
rect 22540 85092 22596 85820
rect 22540 84998 22596 85036
rect 22428 82562 22484 82572
rect 22652 84306 22708 86604
rect 22764 86658 22820 88732
rect 23100 88722 23156 88732
rect 22876 88004 22932 88014
rect 22876 88002 23044 88004
rect 22876 87950 22878 88002
rect 22930 87950 23044 88002
rect 22876 87948 23044 87950
rect 22876 87938 22932 87948
rect 22876 87444 22932 87454
rect 22876 87350 22932 87388
rect 22764 86606 22766 86658
rect 22818 86606 22820 86658
rect 22764 85876 22820 86606
rect 22876 86882 22932 86894
rect 22876 86830 22878 86882
rect 22930 86830 22932 86882
rect 22876 86100 22932 86830
rect 22988 86660 23044 87948
rect 23804 87836 24068 87846
rect 23860 87780 23908 87836
rect 23964 87780 24012 87836
rect 23804 87770 24068 87780
rect 23884 87556 23940 87566
rect 23212 87444 23268 87454
rect 23212 87330 23268 87388
rect 23212 87278 23214 87330
rect 23266 87278 23268 87330
rect 23212 87266 23268 87278
rect 23884 87330 23940 87500
rect 23884 87278 23886 87330
rect 23938 87278 23940 87330
rect 23884 87266 23940 87278
rect 23548 87218 23604 87230
rect 23548 87166 23550 87218
rect 23602 87166 23604 87218
rect 23548 86996 23604 87166
rect 23548 86930 23604 86940
rect 23436 86772 23492 86782
rect 23436 86678 23492 86716
rect 22988 86658 23156 86660
rect 22988 86606 22990 86658
rect 23042 86606 23156 86658
rect 22988 86604 23156 86606
rect 22988 86594 23044 86604
rect 22876 86034 22932 86044
rect 22988 85988 23044 85998
rect 22764 85316 22820 85820
rect 22876 85876 22932 85886
rect 22988 85876 23044 85932
rect 22876 85874 23044 85876
rect 22876 85822 22878 85874
rect 22930 85822 23044 85874
rect 22876 85820 23044 85822
rect 23100 85874 23156 86604
rect 23548 86658 23604 86670
rect 23548 86606 23550 86658
rect 23602 86606 23604 86658
rect 23436 86434 23492 86446
rect 23436 86382 23438 86434
rect 23490 86382 23492 86434
rect 23324 86100 23380 86110
rect 23324 86006 23380 86044
rect 23436 85988 23492 86382
rect 23548 86100 23604 86606
rect 23996 86546 24052 86558
rect 23996 86494 23998 86546
rect 24050 86494 24052 86546
rect 23884 86436 23940 86446
rect 23548 86034 23604 86044
rect 23660 86434 23940 86436
rect 23660 86382 23886 86434
rect 23938 86382 23940 86434
rect 23660 86380 23940 86382
rect 23436 85922 23492 85932
rect 23100 85822 23102 85874
rect 23154 85822 23156 85874
rect 22876 85810 22932 85820
rect 23100 85810 23156 85822
rect 23548 85876 23604 85886
rect 23660 85876 23716 86380
rect 23884 86370 23940 86380
rect 23996 86436 24052 86494
rect 23996 86370 24052 86380
rect 23804 86268 24068 86278
rect 23860 86212 23908 86268
rect 23964 86212 24012 86268
rect 23804 86202 24068 86212
rect 23772 85876 23828 85886
rect 23660 85874 23828 85876
rect 23660 85822 23774 85874
rect 23826 85822 23828 85874
rect 23660 85820 23828 85822
rect 23548 85782 23604 85820
rect 23772 85810 23828 85820
rect 24108 85764 24164 85802
rect 24108 85698 24164 85708
rect 23884 85652 23940 85662
rect 23884 85558 23940 85596
rect 23100 85316 23156 85326
rect 22764 85260 23044 85316
rect 22988 85202 23044 85260
rect 23100 85222 23156 85260
rect 23548 85316 23604 85326
rect 23548 85222 23604 85260
rect 22988 85150 22990 85202
rect 23042 85150 23044 85202
rect 22988 85138 23044 85150
rect 23884 85204 23940 85214
rect 23884 85110 23940 85148
rect 22652 84254 22654 84306
rect 22706 84254 22708 84306
rect 22540 82514 22596 82526
rect 22540 82462 22542 82514
rect 22594 82462 22596 82514
rect 22540 82068 22596 82462
rect 22540 82002 22596 82012
rect 22652 81284 22708 84254
rect 23436 85092 23492 85102
rect 23324 83522 23380 83534
rect 23324 83470 23326 83522
rect 23378 83470 23380 83522
rect 22876 82628 22932 82638
rect 22876 82534 22932 82572
rect 22540 81228 22708 81284
rect 22764 82068 22820 82078
rect 23324 82068 23380 83470
rect 22764 82066 23380 82068
rect 22764 82014 22766 82066
rect 22818 82014 23380 82066
rect 22764 82012 23380 82014
rect 22428 80948 22484 80958
rect 22428 80854 22484 80892
rect 22204 80770 22260 80780
rect 22092 79762 22148 79772
rect 22204 80164 22260 80174
rect 22092 79492 22148 79502
rect 21980 79490 22148 79492
rect 21980 79438 22094 79490
rect 22146 79438 22148 79490
rect 21980 79436 22148 79438
rect 21980 78818 22036 79436
rect 22092 79426 22148 79436
rect 21980 78766 21982 78818
rect 22034 78766 22036 78818
rect 21980 78754 22036 78766
rect 22092 78932 22148 78942
rect 21868 77870 21870 77922
rect 21922 77870 21924 77922
rect 21868 77858 21924 77870
rect 22092 77476 22148 78876
rect 22092 77410 22148 77420
rect 21868 76356 21924 76366
rect 21868 76262 21924 76300
rect 21532 75630 21534 75682
rect 21586 75630 21588 75682
rect 21532 75618 21588 75630
rect 21644 75964 21812 76020
rect 21420 74050 21476 74060
rect 21644 73948 21700 75964
rect 21756 75796 21812 75806
rect 21756 75702 21812 75740
rect 21756 74226 21812 74238
rect 21756 74174 21758 74226
rect 21810 74174 21812 74226
rect 21756 73948 21812 74174
rect 22204 73948 22260 80108
rect 22428 79828 22484 79838
rect 22316 79604 22372 79614
rect 22316 79510 22372 79548
rect 22316 78820 22372 78830
rect 22316 78726 22372 78764
rect 22428 78034 22484 79772
rect 22428 77982 22430 78034
rect 22482 77982 22484 78034
rect 22428 77970 22484 77982
rect 22316 76468 22372 76478
rect 22316 76374 22372 76412
rect 22428 75682 22484 75694
rect 22428 75630 22430 75682
rect 22482 75630 22484 75682
rect 22428 74340 22484 75630
rect 22428 74274 22484 74284
rect 21308 73892 21476 73948
rect 21644 73892 21812 73948
rect 21308 72660 21364 72670
rect 21308 72546 21364 72604
rect 21308 72494 21310 72546
rect 21362 72494 21364 72546
rect 21308 72482 21364 72494
rect 21420 72324 21476 73892
rect 21532 73108 21588 73118
rect 21532 72770 21588 73052
rect 21532 72718 21534 72770
rect 21586 72718 21588 72770
rect 21532 72706 21588 72718
rect 21196 71586 21252 71596
rect 21308 72268 21476 72324
rect 21196 71428 21252 71438
rect 21084 70978 21140 70990
rect 21084 70926 21086 70978
rect 21138 70926 21140 70978
rect 21084 69412 21140 70926
rect 21084 69346 21140 69356
rect 21196 70194 21252 71372
rect 21308 71092 21364 72268
rect 21420 71652 21476 71662
rect 21420 71558 21476 71596
rect 21532 71092 21588 71102
rect 21308 71090 21588 71092
rect 21308 71038 21534 71090
rect 21586 71038 21588 71090
rect 21308 71036 21588 71038
rect 21196 70142 21198 70194
rect 21250 70142 21252 70194
rect 20972 68786 21028 68796
rect 21084 68964 21140 68974
rect 21084 68626 21140 68908
rect 21084 68574 21086 68626
rect 21138 68574 21140 68626
rect 21084 68562 21140 68574
rect 21196 68404 21252 70142
rect 21308 69186 21364 69198
rect 21308 69134 21310 69186
rect 21362 69134 21364 69186
rect 21308 68964 21364 69134
rect 21308 68898 21364 68908
rect 21420 68628 21476 68638
rect 21084 68348 21252 68404
rect 21308 68626 21476 68628
rect 21308 68574 21422 68626
rect 21474 68574 21476 68626
rect 21308 68572 21476 68574
rect 20972 68292 21028 68302
rect 20972 66724 21028 68236
rect 21084 67172 21140 68348
rect 21308 67956 21364 68572
rect 21420 68562 21476 68572
rect 21420 68404 21476 68414
rect 21420 68066 21476 68348
rect 21420 68014 21422 68066
rect 21474 68014 21476 68066
rect 21420 68002 21476 68014
rect 21308 67890 21364 67900
rect 21196 67842 21252 67854
rect 21196 67790 21198 67842
rect 21250 67790 21252 67842
rect 21196 67620 21252 67790
rect 21196 67554 21252 67564
rect 21084 67078 21140 67116
rect 21196 67284 21252 67294
rect 20972 66668 21140 66724
rect 20972 66500 21028 66510
rect 20972 65378 21028 66444
rect 20972 65326 20974 65378
rect 21026 65326 21028 65378
rect 20972 65314 21028 65326
rect 20972 64036 21028 64046
rect 20972 63942 21028 63980
rect 20972 63812 21028 63822
rect 20972 61124 21028 63756
rect 21084 63138 21140 66668
rect 21196 66274 21252 67228
rect 21420 66948 21476 66958
rect 21532 66948 21588 71036
rect 21644 69972 21700 69982
rect 21644 68514 21700 69916
rect 21756 69970 21812 73892
rect 21756 69918 21758 69970
rect 21810 69918 21812 69970
rect 21756 69860 21812 69918
rect 21756 69794 21812 69804
rect 21980 73892 22260 73948
rect 21644 68462 21646 68514
rect 21698 68462 21700 68514
rect 21644 68450 21700 68462
rect 21756 68852 21812 68862
rect 21196 66222 21198 66274
rect 21250 66222 21252 66274
rect 21196 64708 21252 66222
rect 21308 66946 21588 66948
rect 21308 66894 21422 66946
rect 21474 66894 21588 66946
rect 21308 66892 21588 66894
rect 21308 65156 21364 66892
rect 21420 66882 21476 66892
rect 21756 66836 21812 68796
rect 21868 68068 21924 68078
rect 21868 67954 21924 68012
rect 21868 67902 21870 67954
rect 21922 67902 21924 67954
rect 21868 67890 21924 67902
rect 21308 65090 21364 65100
rect 21532 66780 21812 66836
rect 21868 67508 21924 67518
rect 21196 64652 21476 64708
rect 21308 64484 21364 64494
rect 21084 63086 21086 63138
rect 21138 63086 21140 63138
rect 21084 62580 21140 63086
rect 21084 62514 21140 62524
rect 21196 64482 21364 64484
rect 21196 64430 21310 64482
rect 21362 64430 21364 64482
rect 21196 64428 21364 64430
rect 21084 62356 21140 62366
rect 21196 62356 21252 64428
rect 21308 64418 21364 64428
rect 21308 63810 21364 63822
rect 21308 63758 21310 63810
rect 21362 63758 21364 63810
rect 21308 63476 21364 63758
rect 21308 63410 21364 63420
rect 21420 63140 21476 64652
rect 21420 63074 21476 63084
rect 21084 62354 21252 62356
rect 21084 62302 21086 62354
rect 21138 62302 21252 62354
rect 21084 62300 21252 62302
rect 21420 62692 21476 62702
rect 21084 62290 21140 62300
rect 20972 61058 21028 61068
rect 21196 62132 21252 62142
rect 21196 61570 21252 62076
rect 21196 61518 21198 61570
rect 21250 61518 21252 61570
rect 20972 60788 21028 60798
rect 20972 60694 21028 60732
rect 20860 58482 20916 58492
rect 21196 57204 21252 61518
rect 21420 60786 21476 62636
rect 21532 62354 21588 66780
rect 21868 66724 21924 67452
rect 21756 66668 21924 66724
rect 21756 62804 21812 66668
rect 21644 62748 21812 62804
rect 21644 62468 21700 62748
rect 21644 62402 21700 62412
rect 21756 62580 21812 62590
rect 21532 62302 21534 62354
rect 21586 62302 21588 62354
rect 21532 62290 21588 62302
rect 21644 62244 21700 62282
rect 21644 62178 21700 62188
rect 21756 62132 21812 62524
rect 21980 62188 22036 73892
rect 22540 72772 22596 81228
rect 22652 80836 22708 80846
rect 22652 80386 22708 80780
rect 22764 80500 22820 82012
rect 23212 81844 23268 81854
rect 23212 81750 23268 81788
rect 22764 80434 22820 80444
rect 22876 80724 22932 80734
rect 22652 80334 22654 80386
rect 22706 80334 22708 80386
rect 22652 79602 22708 80334
rect 22652 79550 22654 79602
rect 22706 79550 22708 79602
rect 22652 79538 22708 79550
rect 22876 78932 22932 80668
rect 23436 80612 23492 85036
rect 23804 84700 24068 84710
rect 23860 84644 23908 84700
rect 23964 84644 24012 84700
rect 23804 84634 24068 84644
rect 23660 84308 23716 84318
rect 22876 78866 22932 78876
rect 23324 80556 23492 80612
rect 23548 84306 23716 84308
rect 23548 84254 23662 84306
rect 23714 84254 23716 84306
rect 23548 84252 23716 84254
rect 23324 78820 23380 80556
rect 23548 80388 23604 84252
rect 23660 84242 23716 84252
rect 23660 84084 23716 84094
rect 23660 83746 23716 84028
rect 23660 83694 23662 83746
rect 23714 83694 23716 83746
rect 23660 83682 23716 83694
rect 23804 83132 24068 83142
rect 23860 83076 23908 83132
rect 23964 83076 24012 83132
rect 23804 83066 24068 83076
rect 23804 81564 24068 81574
rect 23860 81508 23908 81564
rect 23964 81508 24012 81564
rect 23804 81498 24068 81508
rect 23548 79604 23604 80332
rect 23804 79996 24068 80006
rect 23860 79940 23908 79996
rect 23964 79940 24012 79996
rect 23804 79930 24068 79940
rect 23772 79604 23828 79614
rect 23548 79548 23772 79604
rect 23772 79510 23828 79548
rect 22988 78818 23380 78820
rect 22988 78766 23326 78818
rect 23378 78766 23380 78818
rect 22988 78764 23380 78766
rect 22988 75682 23044 78764
rect 23324 78754 23380 78764
rect 23804 78428 24068 78438
rect 23860 78372 23908 78428
rect 23964 78372 24012 78428
rect 23804 78362 24068 78372
rect 23804 76860 24068 76870
rect 23860 76804 23908 76860
rect 23964 76804 24012 76860
rect 23804 76794 24068 76804
rect 23772 75684 23828 75694
rect 22988 75630 22990 75682
rect 23042 75630 23044 75682
rect 22988 75460 23044 75630
rect 22988 75394 23044 75404
rect 23660 75682 23828 75684
rect 23660 75630 23774 75682
rect 23826 75630 23828 75682
rect 23660 75628 23828 75630
rect 22876 74898 22932 74910
rect 22876 74846 22878 74898
rect 22930 74846 22932 74898
rect 22092 72716 22596 72772
rect 22652 73332 22708 73342
rect 22092 72324 22148 72716
rect 22204 72548 22260 72558
rect 22204 72546 22484 72548
rect 22204 72494 22206 72546
rect 22258 72494 22484 72546
rect 22204 72492 22484 72494
rect 22204 72482 22260 72492
rect 22092 72268 22260 72324
rect 22204 66612 22260 72268
rect 22428 71988 22484 72492
rect 22652 72546 22708 73276
rect 22652 72494 22654 72546
rect 22706 72494 22708 72546
rect 22652 72482 22708 72494
rect 22652 71988 22708 71998
rect 22428 71986 22708 71988
rect 22428 71934 22654 71986
rect 22706 71934 22708 71986
rect 22428 71932 22708 71934
rect 22652 71922 22708 71932
rect 22764 70756 22820 70766
rect 22316 70754 22820 70756
rect 22316 70702 22766 70754
rect 22818 70702 22820 70754
rect 22316 70700 22820 70702
rect 22316 68626 22372 70700
rect 22764 70690 22820 70700
rect 22876 70196 22932 74846
rect 23324 74676 23380 74686
rect 22988 74340 23044 74350
rect 22988 74246 23044 74284
rect 23324 73218 23380 74620
rect 23324 73166 23326 73218
rect 23378 73166 23380 73218
rect 23324 73154 23380 73166
rect 23436 74116 23492 74126
rect 22988 73106 23044 73118
rect 22988 73054 22990 73106
rect 23042 73054 23044 73106
rect 22988 71876 23044 73054
rect 22988 71810 23044 71820
rect 23212 71764 23268 71774
rect 23212 71762 23380 71764
rect 23212 71710 23214 71762
rect 23266 71710 23380 71762
rect 23212 71708 23380 71710
rect 23212 71698 23268 71708
rect 22764 70140 22932 70196
rect 22428 69860 22484 69870
rect 22428 69634 22484 69804
rect 22428 69582 22430 69634
rect 22482 69582 22484 69634
rect 22428 69570 22484 69582
rect 22316 68574 22318 68626
rect 22370 68574 22372 68626
rect 22316 68562 22372 68574
rect 22652 68404 22708 68414
rect 22428 68292 22484 68302
rect 22428 67842 22484 68236
rect 22428 67790 22430 67842
rect 22482 67790 22484 67842
rect 22428 67778 22484 67790
rect 22652 67396 22708 68348
rect 22652 67170 22708 67340
rect 22652 67118 22654 67170
rect 22706 67118 22708 67170
rect 22652 67106 22708 67118
rect 22204 66556 22708 66612
rect 22540 63700 22596 63710
rect 22316 63698 22596 63700
rect 22316 63646 22542 63698
rect 22594 63646 22596 63698
rect 22316 63644 22596 63646
rect 22092 63140 22148 63150
rect 22148 63084 22260 63140
rect 22092 63046 22148 63084
rect 21980 62132 22148 62188
rect 21756 62076 21924 62132
rect 21420 60734 21422 60786
rect 21474 60734 21476 60786
rect 21420 60722 21476 60734
rect 21644 62020 21700 62030
rect 21644 60674 21700 61964
rect 21644 60622 21646 60674
rect 21698 60622 21700 60674
rect 21644 60610 21700 60622
rect 21756 60788 21812 60798
rect 21084 57148 21196 57204
rect 20972 55858 21028 55870
rect 20972 55806 20974 55858
rect 21026 55806 21028 55858
rect 20972 51828 21028 55806
rect 20972 51762 21028 51772
rect 20860 45668 20916 45678
rect 20412 44370 20468 44380
rect 20524 44548 20580 44558
rect 20524 42084 20580 44492
rect 20636 43428 20692 43438
rect 20636 43426 20804 43428
rect 20636 43374 20638 43426
rect 20690 43374 20804 43426
rect 20636 43372 20804 43374
rect 20636 43362 20692 43372
rect 20412 42028 20580 42084
rect 20412 41412 20468 42028
rect 20636 41972 20692 41982
rect 20412 41346 20468 41356
rect 20524 41916 20636 41972
rect 20524 38388 20580 41916
rect 20636 41878 20692 41916
rect 20636 40740 20692 40750
rect 20748 40740 20804 43372
rect 20860 42980 20916 45612
rect 20972 44098 21028 44110
rect 20972 44046 20974 44098
rect 21026 44046 21028 44098
rect 20972 43538 21028 44046
rect 20972 43486 20974 43538
rect 21026 43486 21028 43538
rect 20972 43474 21028 43486
rect 20860 42924 21028 42980
rect 20692 40684 20804 40740
rect 20860 42754 20916 42766
rect 20860 42702 20862 42754
rect 20914 42702 20916 42754
rect 20860 41636 20916 42702
rect 20972 41972 21028 42924
rect 20972 41878 21028 41916
rect 21084 41748 21140 57148
rect 21196 57138 21252 57148
rect 21644 59556 21700 59566
rect 21756 59556 21812 60732
rect 21868 60676 21924 62076
rect 22092 61348 22148 62132
rect 21868 60610 21924 60620
rect 21980 61292 22148 61348
rect 21868 60114 21924 60126
rect 21868 60062 21870 60114
rect 21922 60062 21924 60114
rect 21868 60004 21924 60062
rect 21868 59938 21924 59948
rect 21700 59500 21812 59556
rect 21308 56084 21364 56094
rect 21308 55970 21364 56028
rect 21308 55918 21310 55970
rect 21362 55918 21364 55970
rect 21308 55906 21364 55918
rect 21420 53732 21476 53742
rect 21420 53638 21476 53676
rect 21308 45668 21364 45678
rect 21308 45574 21364 45612
rect 21532 44098 21588 44110
rect 21532 44046 21534 44098
rect 21586 44046 21588 44098
rect 21420 43538 21476 43550
rect 21420 43486 21422 43538
rect 21474 43486 21476 43538
rect 21420 42196 21476 43486
rect 21532 43540 21588 44046
rect 21532 43474 21588 43484
rect 21644 43426 21700 59500
rect 21980 55468 22036 61292
rect 22204 60788 22260 63084
rect 22316 62354 22372 63644
rect 22540 63634 22596 63644
rect 22316 62302 22318 62354
rect 22370 62302 22372 62354
rect 22316 62290 22372 62302
rect 22652 62354 22708 66556
rect 22652 62302 22654 62354
rect 22706 62302 22708 62354
rect 22652 62290 22708 62302
rect 22764 61236 22820 70140
rect 22876 69970 22932 69982
rect 22876 69918 22878 69970
rect 22930 69918 22932 69970
rect 22876 69748 22932 69918
rect 22876 69692 23268 69748
rect 22876 69412 22932 69422
rect 22876 69318 22932 69356
rect 23100 68740 23156 68750
rect 23212 68740 23268 69692
rect 23156 68684 23268 68740
rect 22876 68626 22932 68638
rect 22876 68574 22878 68626
rect 22930 68574 22932 68626
rect 22876 67732 22932 68574
rect 22876 67666 22932 67676
rect 23100 67170 23156 68684
rect 23100 67118 23102 67170
rect 23154 67118 23156 67170
rect 23100 67106 23156 67118
rect 23212 68516 23268 68526
rect 23212 67170 23268 68460
rect 23212 67118 23214 67170
rect 23266 67118 23268 67170
rect 23212 67106 23268 67118
rect 23324 62188 23380 71708
rect 23436 71650 23492 74060
rect 23436 71598 23438 71650
rect 23490 71598 23492 71650
rect 23436 71586 23492 71598
rect 23660 72546 23716 75628
rect 23772 75618 23828 75628
rect 23804 75292 24068 75302
rect 23860 75236 23908 75292
rect 23964 75236 24012 75292
rect 23804 75226 24068 75236
rect 23804 73724 24068 73734
rect 23860 73668 23908 73724
rect 23964 73668 24012 73724
rect 23804 73658 24068 73668
rect 23660 72494 23662 72546
rect 23714 72494 23716 72546
rect 23436 69186 23492 69198
rect 23436 69134 23438 69186
rect 23490 69134 23492 69186
rect 23436 68516 23492 69134
rect 23436 68450 23492 68460
rect 23660 68626 23716 72494
rect 23804 72156 24068 72166
rect 23860 72100 23908 72156
rect 23964 72100 24012 72156
rect 23804 72090 24068 72100
rect 23804 70588 24068 70598
rect 23860 70532 23908 70588
rect 23964 70532 24012 70588
rect 23804 70522 24068 70532
rect 23772 69412 23828 69422
rect 24220 69412 24276 92092
rect 24464 91756 24728 91766
rect 24520 91700 24568 91756
rect 24624 91700 24672 91756
rect 24464 91690 24728 91700
rect 24464 90188 24728 90198
rect 24520 90132 24568 90188
rect 24624 90132 24672 90188
rect 24464 90122 24728 90132
rect 24332 89012 24388 89022
rect 24332 85316 24388 88956
rect 24892 88788 24948 88798
rect 24464 88620 24728 88630
rect 24520 88564 24568 88620
rect 24624 88564 24672 88620
rect 24464 88554 24728 88564
rect 24464 87052 24728 87062
rect 24520 86996 24568 87052
rect 24624 86996 24672 87052
rect 24464 86986 24728 86996
rect 24444 85764 24500 85802
rect 24444 85698 24500 85708
rect 24464 85484 24728 85494
rect 24520 85428 24568 85484
rect 24624 85428 24672 85484
rect 24464 85418 24728 85428
rect 24332 85250 24388 85260
rect 24464 83916 24728 83926
rect 24520 83860 24568 83916
rect 24624 83860 24672 83916
rect 24464 83850 24728 83860
rect 24464 82348 24728 82358
rect 24520 82292 24568 82348
rect 24624 82292 24672 82348
rect 24464 82282 24728 82292
rect 24464 80780 24728 80790
rect 24520 80724 24568 80780
rect 24624 80724 24672 80780
rect 24464 80714 24728 80724
rect 24464 79212 24728 79222
rect 24520 79156 24568 79212
rect 24624 79156 24672 79212
rect 24464 79146 24728 79156
rect 24464 77644 24728 77654
rect 24520 77588 24568 77644
rect 24624 77588 24672 77644
rect 24464 77578 24728 77588
rect 24464 76076 24728 76086
rect 24520 76020 24568 76076
rect 24624 76020 24672 76076
rect 24464 76010 24728 76020
rect 24464 74508 24728 74518
rect 24520 74452 24568 74508
rect 24624 74452 24672 74508
rect 24464 74442 24728 74452
rect 24464 72940 24728 72950
rect 24520 72884 24568 72940
rect 24624 72884 24672 72940
rect 24464 72874 24728 72884
rect 24464 71372 24728 71382
rect 24520 71316 24568 71372
rect 24624 71316 24672 71372
rect 24464 71306 24728 71316
rect 24464 69804 24728 69814
rect 24520 69748 24568 69804
rect 24624 69748 24672 69804
rect 24464 69738 24728 69748
rect 23772 69410 24276 69412
rect 23772 69358 23774 69410
rect 23826 69358 24276 69410
rect 23772 69356 24276 69358
rect 23772 69346 23828 69356
rect 23772 69188 23828 69198
rect 23772 69186 24836 69188
rect 23772 69134 23774 69186
rect 23826 69134 24836 69186
rect 23772 69132 24836 69134
rect 23772 69122 23828 69132
rect 23804 69020 24068 69030
rect 23860 68964 23908 69020
rect 23964 68964 24012 69020
rect 23804 68954 24068 68964
rect 24220 68964 24276 68974
rect 23660 68574 23662 68626
rect 23714 68574 23716 68626
rect 23436 67842 23492 67854
rect 23436 67790 23438 67842
rect 23490 67790 23492 67842
rect 23436 67284 23492 67790
rect 23660 67508 23716 68574
rect 24220 68626 24276 68908
rect 24332 68852 24388 68862
rect 24332 68738 24388 68796
rect 24332 68686 24334 68738
rect 24386 68686 24388 68738
rect 24332 68674 24388 68686
rect 24220 68574 24222 68626
rect 24274 68574 24276 68626
rect 24220 68562 24276 68574
rect 24668 68628 24724 68638
rect 24668 68534 24724 68572
rect 24780 68626 24836 69132
rect 24780 68574 24782 68626
rect 24834 68574 24836 68626
rect 24780 68562 24836 68574
rect 24444 68514 24500 68526
rect 24444 68462 24446 68514
rect 24498 68462 24500 68514
rect 24444 68404 24500 68462
rect 24444 68338 24500 68348
rect 24464 68236 24728 68246
rect 24520 68180 24568 68236
rect 24624 68180 24672 68236
rect 24464 68170 24728 68180
rect 23660 67442 23716 67452
rect 23804 67452 24068 67462
rect 23860 67396 23908 67452
rect 23964 67396 24012 67452
rect 23804 67386 24068 67396
rect 23436 67218 23492 67228
rect 24464 66668 24728 66678
rect 24520 66612 24568 66668
rect 24624 66612 24672 66668
rect 24464 66602 24728 66612
rect 23804 65884 24068 65894
rect 23860 65828 23908 65884
rect 23964 65828 24012 65884
rect 23804 65818 24068 65828
rect 24464 65100 24728 65110
rect 24520 65044 24568 65100
rect 24624 65044 24672 65100
rect 24464 65034 24728 65044
rect 23804 64316 24068 64326
rect 23860 64260 23908 64316
rect 23964 64260 24012 64316
rect 23804 64250 24068 64260
rect 24464 63532 24728 63542
rect 24520 63476 24568 63532
rect 24624 63476 24672 63532
rect 24464 63466 24728 63476
rect 23804 62748 24068 62758
rect 23860 62692 23908 62748
rect 23964 62692 24012 62748
rect 23804 62682 24068 62692
rect 23772 62356 23828 62366
rect 23772 62262 23828 62300
rect 22764 61170 22820 61180
rect 22988 62132 23380 62188
rect 22204 60722 22260 60732
rect 22428 60900 22484 60910
rect 22092 60674 22148 60686
rect 22092 60622 22094 60674
rect 22146 60622 22148 60674
rect 22092 59332 22148 60622
rect 22204 59892 22260 59902
rect 22204 59798 22260 59836
rect 22092 59266 22148 59276
rect 21980 55412 22260 55468
rect 21756 53842 21812 53854
rect 21756 53790 21758 53842
rect 21810 53790 21812 53842
rect 21756 53732 21812 53790
rect 21756 53666 21812 53676
rect 21644 43374 21646 43426
rect 21698 43374 21700 43426
rect 21644 43362 21700 43374
rect 21868 44884 21924 44894
rect 20636 40514 20692 40684
rect 20636 40462 20638 40514
rect 20690 40462 20692 40514
rect 20636 38668 20692 40462
rect 20860 40292 20916 41580
rect 20972 41692 21140 41748
rect 21196 42140 21476 42196
rect 21532 42530 21588 42542
rect 21532 42478 21534 42530
rect 21586 42478 21588 42530
rect 20972 40628 21028 41692
rect 21084 41188 21140 41198
rect 21084 41094 21140 41132
rect 20972 40572 21140 40628
rect 20972 40404 21028 40414
rect 20972 40310 21028 40348
rect 20860 40226 20916 40236
rect 20860 39060 20916 39070
rect 20860 38834 20916 39004
rect 20860 38782 20862 38834
rect 20914 38782 20916 38834
rect 20636 38612 20804 38668
rect 20524 38332 20692 38388
rect 20300 38220 20580 38276
rect 20076 38164 20132 38174
rect 20076 38162 20356 38164
rect 20076 38110 20078 38162
rect 20130 38110 20356 38162
rect 20076 38108 20356 38110
rect 20076 38098 20132 38108
rect 20076 37938 20132 37950
rect 20076 37886 20078 37938
rect 20130 37886 20132 37938
rect 20076 36932 20132 37886
rect 20076 36876 20244 36932
rect 19964 36764 20132 36820
rect 19628 36316 19796 36372
rect 19964 36594 20020 36606
rect 19964 36542 19966 36594
rect 20018 36542 20020 36594
rect 19628 33908 19684 36316
rect 19964 36148 20020 36542
rect 19964 36082 20020 36092
rect 19740 35588 19796 35598
rect 19740 35494 19796 35532
rect 19852 35474 19908 35486
rect 19852 35422 19854 35474
rect 19906 35422 19908 35474
rect 19852 34356 19908 35422
rect 19852 34290 19908 34300
rect 19964 35474 20020 35486
rect 19964 35422 19966 35474
rect 20018 35422 20020 35474
rect 19628 33842 19684 33852
rect 19852 34130 19908 34142
rect 19852 34078 19854 34130
rect 19906 34078 19908 34130
rect 19740 33684 19796 33694
rect 19852 33684 19908 34078
rect 19796 33628 19908 33684
rect 19740 33618 19796 33628
rect 19516 33516 19684 33572
rect 19628 33458 19684 33516
rect 19964 33460 20020 35422
rect 19628 33406 19630 33458
rect 19682 33406 19684 33458
rect 19628 33394 19684 33406
rect 19740 33404 20020 33460
rect 19516 33348 19572 33358
rect 19516 33254 19572 33292
rect 19740 33124 19796 33404
rect 20076 33348 20132 36764
rect 20188 35364 20244 36876
rect 20188 35298 20244 35308
rect 19964 33292 20132 33348
rect 20188 35140 20244 35150
rect 19852 33236 19908 33246
rect 19852 33142 19908 33180
rect 19292 32786 19460 32788
rect 19292 32734 19294 32786
rect 19346 32734 19460 32786
rect 19292 32732 19460 32734
rect 19516 33068 19796 33124
rect 19292 32722 19348 32732
rect 18956 32564 19012 32574
rect 18844 32562 19012 32564
rect 18844 32510 18958 32562
rect 19010 32510 19012 32562
rect 18844 32508 19012 32510
rect 18172 31666 18452 31668
rect 18172 31614 18174 31666
rect 18226 31614 18452 31666
rect 18172 31612 18452 31614
rect 18172 31602 18228 31612
rect 18620 31554 18676 31566
rect 18620 31502 18622 31554
rect 18674 31502 18676 31554
rect 18172 31444 18228 31454
rect 18060 30994 18116 31006
rect 18060 30942 18062 30994
rect 18114 30942 18116 30994
rect 18060 30212 18116 30942
rect 18060 30146 18116 30156
rect 18172 29988 18228 31388
rect 18508 31220 18564 31230
rect 18508 31126 18564 31164
rect 18620 31108 18676 31502
rect 18620 31042 18676 31052
rect 18732 31554 18788 31566
rect 18732 31502 18734 31554
rect 18786 31502 18788 31554
rect 18396 30100 18452 30110
rect 18396 30006 18452 30044
rect 17836 29314 18004 29316
rect 17836 29262 17838 29314
rect 17890 29262 18004 29314
rect 17836 29260 18004 29262
rect 18060 29932 18228 29988
rect 18284 29988 18340 29998
rect 17836 29250 17892 29260
rect 17388 26852 17556 26908
rect 17724 26852 17892 26908
rect 17276 25678 17278 25730
rect 17330 25678 17332 25730
rect 17276 25666 17332 25678
rect 16940 25454 16942 25506
rect 16994 25454 16996 25506
rect 16940 25442 16996 25454
rect 17164 25506 17220 25518
rect 17164 25454 17166 25506
rect 17218 25454 17220 25506
rect 16380 25284 16436 25294
rect 15596 25004 16100 25060
rect 16268 25172 16324 25182
rect 15596 24946 15652 25004
rect 15596 24894 15598 24946
rect 15650 24894 15652 24946
rect 15596 24882 15652 24894
rect 16156 24948 16212 24958
rect 16044 23714 16100 23726
rect 16044 23662 16046 23714
rect 16098 23662 16100 23714
rect 16044 23604 16100 23662
rect 15372 23548 16100 23604
rect 15372 23492 15652 23548
rect 14812 23156 14868 23166
rect 14868 23100 14980 23156
rect 14812 23090 14868 23100
rect 14924 23042 14980 23100
rect 14924 22990 14926 23042
rect 14978 22990 14980 23042
rect 14924 22978 14980 22990
rect 15036 23044 15092 23492
rect 15260 23426 15316 23436
rect 15596 23380 15652 23492
rect 15372 23324 15652 23380
rect 16044 23380 16100 23390
rect 16156 23380 16212 24892
rect 16044 23378 16212 23380
rect 16044 23326 16046 23378
rect 16098 23326 16212 23378
rect 16044 23324 16212 23326
rect 15260 23156 15316 23166
rect 15372 23156 15428 23324
rect 16044 23314 16100 23324
rect 15260 23154 15428 23156
rect 15260 23102 15262 23154
rect 15314 23102 15428 23154
rect 15260 23100 15428 23102
rect 15484 23156 15540 23166
rect 15260 23090 15316 23100
rect 15484 23062 15540 23100
rect 15036 22978 15092 22988
rect 15596 23044 15652 23054
rect 15596 23042 15764 23044
rect 15596 22990 15598 23042
rect 15650 22990 15764 23042
rect 15596 22988 15764 22990
rect 15596 22978 15652 22988
rect 14812 22930 14868 22942
rect 14812 22878 14814 22930
rect 14866 22878 14868 22930
rect 14812 22820 14868 22878
rect 15596 22820 15652 22830
rect 14812 22764 15092 22820
rect 14924 22596 14980 22606
rect 14924 22502 14980 22540
rect 14812 22370 14868 22382
rect 14812 22318 14814 22370
rect 14866 22318 14868 22370
rect 14812 22148 14868 22318
rect 14812 22082 14868 22092
rect 15036 22370 15092 22764
rect 15036 22318 15038 22370
rect 15090 22318 15092 22370
rect 14364 21522 14420 21532
rect 14588 21756 14756 21812
rect 14812 21924 14868 21934
rect 14140 21074 14196 21084
rect 13916 20710 13972 20748
rect 14476 20468 14532 20478
rect 14476 19236 14532 20412
rect 14588 19460 14644 21756
rect 14700 21588 14756 21598
rect 14700 20802 14756 21532
rect 14812 21586 14868 21868
rect 14812 21534 14814 21586
rect 14866 21534 14868 21586
rect 14812 21522 14868 21534
rect 14700 20750 14702 20802
rect 14754 20750 14756 20802
rect 14700 20738 14756 20750
rect 14812 21028 14868 21038
rect 14812 20242 14868 20972
rect 14812 20190 14814 20242
rect 14866 20190 14868 20242
rect 14812 20178 14868 20190
rect 15036 19460 15092 22318
rect 15596 22370 15652 22764
rect 15708 22596 15764 22988
rect 16268 22708 16324 25116
rect 15708 22530 15764 22540
rect 15820 22652 16324 22708
rect 15596 22318 15598 22370
rect 15650 22318 15652 22370
rect 15596 22306 15652 22318
rect 15372 22260 15428 22270
rect 15372 20804 15428 22204
rect 15820 21924 15876 22652
rect 16156 22484 16212 22494
rect 16044 22482 16212 22484
rect 16044 22430 16158 22482
rect 16210 22430 16212 22482
rect 16044 22428 16212 22430
rect 15708 21868 15876 21924
rect 15932 22370 15988 22382
rect 15932 22318 15934 22370
rect 15986 22318 15988 22370
rect 15708 20916 15764 21868
rect 15820 21700 15876 21710
rect 15820 21586 15876 21644
rect 15820 21534 15822 21586
rect 15874 21534 15876 21586
rect 15820 21522 15876 21534
rect 15708 20850 15764 20860
rect 15260 20748 15428 20804
rect 15932 20802 15988 22318
rect 16044 20916 16100 22428
rect 16156 22418 16212 22428
rect 16044 20850 16100 20860
rect 16156 22258 16212 22270
rect 16156 22206 16158 22258
rect 16210 22206 16212 22258
rect 16156 20914 16212 22206
rect 16380 22260 16436 25228
rect 17164 24948 17220 25454
rect 17388 25508 17444 25518
rect 17388 25414 17444 25452
rect 17164 24882 17220 24892
rect 17276 24724 17332 24734
rect 17276 24630 17332 24668
rect 16716 24612 16772 24622
rect 16716 24518 16772 24556
rect 17500 23940 17556 26852
rect 17724 26292 17780 26302
rect 17724 25730 17780 26236
rect 17724 25678 17726 25730
rect 17778 25678 17780 25730
rect 17724 25666 17780 25678
rect 16940 23884 17556 23940
rect 17724 24724 17780 24734
rect 16828 23154 16884 23166
rect 16828 23102 16830 23154
rect 16882 23102 16884 23154
rect 16716 23044 16772 23054
rect 16380 22194 16436 22204
rect 16604 23042 16772 23044
rect 16604 22990 16718 23042
rect 16770 22990 16772 23042
rect 16604 22988 16772 22990
rect 16604 21812 16660 22988
rect 16716 22978 16772 22988
rect 16828 22260 16884 23102
rect 16940 22594 16996 23884
rect 17164 23716 17220 23726
rect 16940 22542 16942 22594
rect 16994 22542 16996 22594
rect 16940 22484 16996 22542
rect 16940 22418 16996 22428
rect 17052 23156 17108 23166
rect 16828 22194 16884 22204
rect 17052 22258 17108 23100
rect 17052 22206 17054 22258
rect 17106 22206 17108 22258
rect 17052 22194 17108 22206
rect 16156 20862 16158 20914
rect 16210 20862 16212 20914
rect 16156 20850 16212 20862
rect 16268 21756 16660 21812
rect 16716 22146 16772 22158
rect 16716 22094 16718 22146
rect 16770 22094 16772 22146
rect 15932 20750 15934 20802
rect 15986 20750 15988 20802
rect 15260 20020 15316 20748
rect 15708 20692 15764 20702
rect 15260 19954 15316 19964
rect 15372 20578 15428 20590
rect 15372 20526 15374 20578
rect 15426 20526 15428 20578
rect 15148 19460 15204 19470
rect 14588 19404 14756 19460
rect 15036 19458 15204 19460
rect 15036 19406 15150 19458
rect 15202 19406 15204 19458
rect 15036 19404 15204 19406
rect 14588 19236 14644 19246
rect 14476 19234 14644 19236
rect 14476 19182 14590 19234
rect 14642 19182 14644 19234
rect 14476 19180 14644 19182
rect 14588 19170 14644 19180
rect 13804 17838 13806 17890
rect 13858 17838 13860 17890
rect 13804 17826 13860 17838
rect 13916 18788 13972 18798
rect 13692 17778 13748 17790
rect 13692 17726 13694 17778
rect 13746 17726 13748 17778
rect 13692 15148 13748 17726
rect 13916 17778 13972 18732
rect 14588 18788 14644 18798
rect 13916 17726 13918 17778
rect 13970 17726 13972 17778
rect 13916 17714 13972 17726
rect 14476 18564 14532 18574
rect 14476 17666 14532 18508
rect 14588 18450 14644 18732
rect 14588 18398 14590 18450
rect 14642 18398 14644 18450
rect 14588 18386 14644 18398
rect 14476 17614 14478 17666
rect 14530 17614 14532 17666
rect 14476 17602 14532 17614
rect 14700 17668 14756 19404
rect 15148 19394 15204 19404
rect 15260 19122 15316 19134
rect 15260 19070 15262 19122
rect 15314 19070 15316 19122
rect 15148 19012 15204 19022
rect 15148 18564 15204 18956
rect 15260 18788 15316 19070
rect 15260 18722 15316 18732
rect 15260 18564 15316 18574
rect 15204 18562 15316 18564
rect 15204 18510 15262 18562
rect 15314 18510 15316 18562
rect 15204 18508 15316 18510
rect 15148 18470 15204 18508
rect 15260 18498 15316 18508
rect 15372 18564 15428 20526
rect 15596 20580 15652 20590
rect 15596 20486 15652 20524
rect 15596 20018 15652 20030
rect 15596 19966 15598 20018
rect 15650 19966 15652 20018
rect 15372 18498 15428 18508
rect 15484 19908 15540 19918
rect 14588 16884 14644 16894
rect 14700 16884 14756 17612
rect 14924 17780 14980 17790
rect 14924 17108 14980 17724
rect 14924 17042 14980 17052
rect 15036 17220 15092 17230
rect 14588 16882 14756 16884
rect 14588 16830 14590 16882
rect 14642 16830 14756 16882
rect 14588 16828 14756 16830
rect 14588 16818 14644 16828
rect 14140 16770 14196 16782
rect 14140 16718 14142 16770
rect 14194 16718 14196 16770
rect 14028 16100 14084 16110
rect 13916 16044 14028 16100
rect 13916 15316 13972 16044
rect 14028 16006 14084 16044
rect 13916 15250 13972 15260
rect 14028 15428 14084 15438
rect 14028 15202 14084 15372
rect 14028 15150 14030 15202
rect 14082 15150 14084 15202
rect 13692 15092 13860 15148
rect 14028 15138 14084 15150
rect 14140 15204 14196 16718
rect 13580 14924 13748 14980
rect 13468 14690 13524 14700
rect 13356 14530 13412 14542
rect 13356 14478 13358 14530
rect 13410 14478 13412 14530
rect 13356 13188 13412 14478
rect 13580 14532 13636 14542
rect 13356 13122 13412 13132
rect 13468 13746 13524 13758
rect 13468 13694 13470 13746
rect 13522 13694 13524 13746
rect 13468 13412 13524 13694
rect 13468 12852 13524 13356
rect 13468 12786 13524 12796
rect 13468 11396 13524 11406
rect 13580 11396 13636 14476
rect 13468 11394 13636 11396
rect 13468 11342 13470 11394
rect 13522 11342 13636 11394
rect 13468 11340 13636 11342
rect 13692 14530 13748 14924
rect 13692 14478 13694 14530
rect 13746 14478 13748 14530
rect 13692 11396 13748 14478
rect 13804 13524 13860 15092
rect 14028 14868 14084 14878
rect 13916 14756 13972 14766
rect 13916 14662 13972 14700
rect 13916 13972 13972 13982
rect 13916 13634 13972 13916
rect 13916 13582 13918 13634
rect 13970 13582 13972 13634
rect 13916 13570 13972 13582
rect 13804 13458 13860 13468
rect 13804 13300 13860 13310
rect 13804 11788 13860 13244
rect 13916 12964 13972 12974
rect 14028 12964 14084 14812
rect 14140 13412 14196 15148
rect 14364 16660 14420 16670
rect 14140 13356 14308 13412
rect 14140 13188 14196 13198
rect 14140 13094 14196 13132
rect 14028 12908 14196 12964
rect 13916 12068 13972 12908
rect 14028 12068 14084 12078
rect 13916 12012 14028 12068
rect 14028 11974 14084 12012
rect 13804 11732 14084 11788
rect 13916 11508 13972 11518
rect 13916 11414 13972 11452
rect 13692 11340 13860 11396
rect 13468 11330 13524 11340
rect 13468 10612 13524 10622
rect 13132 7868 13300 7924
rect 13356 8260 13412 8270
rect 13132 7588 13188 7868
rect 12012 5854 12014 5906
rect 12066 5854 12068 5906
rect 12012 5842 12068 5854
rect 12124 7420 12292 7476
rect 13020 7532 13188 7588
rect 11564 5684 11620 5694
rect 11900 5684 11956 5694
rect 11564 5682 11732 5684
rect 11564 5630 11566 5682
rect 11618 5630 11732 5682
rect 11564 5628 11732 5630
rect 11564 5618 11620 5628
rect 11564 5122 11620 5134
rect 11564 5070 11566 5122
rect 11618 5070 11620 5122
rect 11564 4676 11620 5070
rect 11564 4610 11620 4620
rect 11564 4340 11620 4350
rect 11564 4246 11620 4284
rect 11452 3559 11508 3594
rect 11452 3556 11454 3559
rect 11506 3556 11508 3559
rect 11452 3490 11508 3500
rect 11340 2930 11396 2940
rect 11676 2884 11732 5628
rect 11900 4226 11956 5628
rect 12124 5122 12180 7420
rect 12236 7252 12292 7262
rect 12236 5794 12292 7196
rect 12460 6692 12516 6702
rect 12460 6598 12516 6636
rect 12236 5742 12238 5794
rect 12290 5742 12292 5794
rect 12236 5730 12292 5742
rect 12908 6578 12964 6590
rect 12908 6526 12910 6578
rect 12962 6526 12964 6578
rect 12908 6468 12964 6526
rect 12236 5236 12292 5246
rect 12236 5142 12292 5180
rect 12124 5070 12126 5122
rect 12178 5070 12180 5122
rect 12124 5058 12180 5070
rect 12684 5122 12740 5134
rect 12684 5070 12686 5122
rect 12738 5070 12740 5122
rect 12236 4340 12292 4350
rect 12236 4246 12292 4284
rect 11900 4174 11902 4226
rect 11954 4174 11956 4226
rect 11900 4162 11956 4174
rect 12684 3780 12740 5070
rect 12908 5124 12964 6412
rect 12908 5058 12964 5068
rect 12684 3714 12740 3724
rect 10892 2830 10894 2882
rect 10946 2830 10948 2882
rect 10892 2818 10948 2830
rect 11116 2882 11284 2884
rect 11116 2830 11230 2882
rect 11282 2830 11284 2882
rect 11116 2828 11284 2830
rect 10668 1038 10670 1090
rect 10722 1038 10724 1090
rect 10668 1026 10724 1038
rect 11004 980 11060 990
rect 10780 644 10836 654
rect 10556 532 10612 542
rect 10556 112 10612 476
rect 10780 112 10836 588
rect 11004 112 11060 924
rect 11116 308 11172 2828
rect 11228 2818 11284 2828
rect 11452 2828 11732 2884
rect 11788 3556 11844 3566
rect 11452 1876 11508 2828
rect 11676 2660 11732 2670
rect 11564 2548 11620 2558
rect 11564 2454 11620 2492
rect 11676 2210 11732 2604
rect 11788 2548 11844 3500
rect 12348 3554 12404 3566
rect 12348 3502 12350 3554
rect 12402 3502 12404 3554
rect 12348 3388 12404 3502
rect 11788 2482 11844 2492
rect 11900 3332 12404 3388
rect 12908 3554 12964 3566
rect 12908 3502 12910 3554
rect 12962 3502 12964 3554
rect 11676 2158 11678 2210
rect 11730 2158 11732 2210
rect 11676 2146 11732 2158
rect 11788 2212 11844 2222
rect 11452 1820 11620 1876
rect 11116 242 11172 252
rect 11228 1652 11284 1662
rect 11228 112 11284 1596
rect 11452 1652 11508 1662
rect 11452 112 11508 1596
rect 11564 1316 11620 1820
rect 11564 1250 11620 1260
rect 11676 1540 11732 1550
rect 11676 112 11732 1484
rect 11788 1426 11844 2156
rect 11900 1876 11956 3332
rect 12012 2772 12068 2782
rect 12012 2770 12404 2772
rect 12012 2718 12014 2770
rect 12066 2718 12404 2770
rect 12012 2716 12404 2718
rect 12012 2706 12068 2716
rect 12348 2660 12404 2716
rect 12796 2660 12852 2670
rect 12348 2658 12852 2660
rect 12348 2606 12798 2658
rect 12850 2606 12852 2658
rect 12348 2604 12852 2606
rect 12796 2594 12852 2604
rect 12236 2546 12292 2558
rect 12236 2494 12238 2546
rect 12290 2494 12292 2546
rect 11900 1820 12068 1876
rect 11788 1374 11790 1426
rect 11842 1374 11844 1426
rect 11788 1362 11844 1374
rect 11900 1652 11956 1662
rect 11900 112 11956 1596
rect 12012 1428 12068 1820
rect 12012 1362 12068 1372
rect 12124 1652 12180 1662
rect 12124 112 12180 1596
rect 12236 644 12292 2494
rect 12908 2212 12964 3502
rect 13020 2770 13076 7532
rect 13356 7476 13412 8204
rect 13244 7364 13300 7374
rect 13244 7270 13300 7308
rect 13356 7140 13412 7420
rect 13132 7084 13412 7140
rect 13132 5124 13188 7084
rect 13356 6690 13412 6702
rect 13356 6638 13358 6690
rect 13410 6638 13412 6690
rect 13244 5682 13300 5694
rect 13244 5630 13246 5682
rect 13298 5630 13300 5682
rect 13244 5348 13300 5630
rect 13244 5282 13300 5292
rect 13244 5124 13300 5134
rect 13132 5122 13300 5124
rect 13132 5070 13246 5122
rect 13298 5070 13300 5122
rect 13132 5068 13300 5070
rect 13244 5058 13300 5068
rect 13356 5124 13412 6638
rect 13468 5906 13524 10556
rect 13580 9940 13636 11340
rect 13580 9874 13636 9884
rect 13692 10610 13748 10622
rect 13692 10558 13694 10610
rect 13746 10558 13748 10610
rect 13692 9492 13748 10558
rect 13692 9426 13748 9436
rect 13580 9156 13636 9166
rect 13580 9062 13636 9100
rect 13580 8258 13636 8270
rect 13580 8206 13582 8258
rect 13634 8206 13636 8258
rect 13580 8036 13636 8206
rect 13580 7588 13636 7980
rect 13804 7924 13860 11340
rect 13916 10948 13972 10958
rect 13916 9604 13972 10892
rect 14028 9828 14084 11732
rect 14140 10948 14196 12908
rect 14140 10882 14196 10892
rect 14140 10500 14196 10510
rect 14252 10500 14308 13356
rect 14364 10612 14420 16604
rect 14924 16098 14980 16110
rect 14924 16046 14926 16098
rect 14978 16046 14980 16098
rect 14476 15652 14532 15662
rect 14476 15426 14532 15596
rect 14476 15374 14478 15426
rect 14530 15374 14532 15426
rect 14476 12290 14532 15374
rect 14588 14530 14644 14542
rect 14588 14478 14590 14530
rect 14642 14478 14644 14530
rect 14588 14084 14644 14478
rect 14812 14420 14868 14430
rect 14924 14420 14980 16046
rect 15036 15202 15092 17164
rect 15036 15150 15038 15202
rect 15090 15150 15092 15202
rect 15036 15138 15092 15150
rect 15484 15204 15540 19852
rect 15596 19796 15652 19966
rect 15596 19012 15652 19740
rect 15708 19346 15764 20636
rect 15932 19572 15988 20750
rect 16044 20692 16100 20702
rect 16044 20578 16100 20636
rect 16044 20526 16046 20578
rect 16098 20526 16100 20578
rect 16044 20514 16100 20526
rect 16044 19908 16100 19918
rect 16044 19814 16100 19852
rect 15932 19516 16100 19572
rect 15708 19294 15710 19346
rect 15762 19294 15764 19346
rect 15708 19282 15764 19294
rect 15932 19348 15988 19358
rect 15932 19254 15988 19292
rect 15596 18946 15652 18956
rect 15596 18340 15652 18378
rect 15596 18274 15652 18284
rect 15484 15138 15540 15148
rect 15596 18116 15652 18126
rect 15596 15148 15652 18060
rect 16044 17890 16100 19516
rect 16268 19458 16324 21756
rect 16716 21700 16772 22094
rect 17164 21812 17220 23660
rect 17724 23604 17780 24668
rect 17724 23538 17780 23548
rect 17276 23154 17332 23166
rect 17276 23102 17278 23154
rect 17330 23102 17332 23154
rect 17276 22820 17332 23102
rect 17500 23156 17556 23166
rect 17500 23062 17556 23100
rect 17612 22930 17668 22942
rect 17612 22878 17614 22930
rect 17666 22878 17668 22930
rect 17276 22764 17556 22820
rect 16268 19406 16270 19458
rect 16322 19406 16324 19458
rect 16268 19394 16324 19406
rect 16380 21644 16772 21700
rect 16828 21756 17220 21812
rect 17276 22260 17332 22270
rect 16828 21698 16884 21756
rect 16828 21646 16830 21698
rect 16882 21646 16884 21698
rect 16380 21362 16436 21644
rect 16828 21634 16884 21646
rect 17164 21588 17220 21598
rect 16940 21586 17220 21588
rect 16940 21534 17166 21586
rect 17218 21534 17220 21586
rect 16940 21532 17220 21534
rect 16492 21476 16548 21486
rect 16492 21474 16772 21476
rect 16492 21422 16494 21474
rect 16546 21422 16772 21474
rect 16492 21420 16772 21422
rect 16492 21410 16548 21420
rect 16380 21310 16382 21362
rect 16434 21310 16436 21362
rect 16156 19346 16212 19358
rect 16156 19294 16158 19346
rect 16210 19294 16212 19346
rect 16156 19012 16212 19294
rect 16380 19012 16436 21310
rect 16604 21252 16660 21262
rect 16156 18956 16436 19012
rect 16492 21028 16548 21038
rect 16044 17838 16046 17890
rect 16098 17838 16100 17890
rect 16044 17826 16100 17838
rect 16156 18228 16212 18238
rect 15932 15316 15988 15326
rect 15932 15148 15988 15260
rect 15372 15090 15428 15102
rect 15596 15092 15876 15148
rect 15932 15092 16100 15148
rect 15372 15038 15374 15090
rect 15426 15038 15428 15090
rect 15372 14756 15428 15038
rect 15372 14690 15428 14700
rect 14868 14364 14980 14420
rect 15036 14530 15092 14542
rect 15036 14478 15038 14530
rect 15090 14478 15092 14530
rect 15036 14420 15092 14478
rect 14812 14354 14868 14364
rect 15036 14354 15092 14364
rect 14588 14018 14644 14028
rect 15036 14084 15092 14094
rect 15036 13970 15092 14028
rect 15036 13918 15038 13970
rect 15090 13918 15092 13970
rect 15036 13906 15092 13918
rect 14700 13748 14756 13758
rect 14476 12238 14478 12290
rect 14530 12238 14532 12290
rect 14476 12226 14532 12238
rect 14588 13636 14644 13646
rect 14364 10546 14420 10556
rect 14140 10498 14308 10500
rect 14140 10446 14142 10498
rect 14194 10446 14308 10498
rect 14140 10444 14308 10446
rect 14140 10434 14196 10444
rect 14252 10388 14308 10444
rect 14252 10322 14308 10332
rect 14588 10164 14644 13580
rect 14700 11060 14756 13692
rect 15708 12516 15764 12526
rect 15708 11396 15764 12460
rect 15708 11330 15764 11340
rect 14700 10994 14756 11004
rect 15036 11170 15092 11182
rect 15036 11118 15038 11170
rect 15090 11118 15092 11170
rect 14028 9734 14084 9772
rect 14140 10108 14644 10164
rect 14924 10836 14980 10846
rect 13916 9548 14084 9604
rect 13916 9044 13972 9054
rect 13916 8950 13972 8988
rect 13804 7858 13860 7868
rect 13580 7522 13636 7532
rect 13692 7476 13748 7486
rect 13580 7250 13636 7262
rect 13580 7198 13582 7250
rect 13634 7198 13636 7250
rect 13580 7028 13636 7198
rect 13580 6962 13636 6972
rect 13692 6690 13748 7420
rect 13916 7252 13972 7262
rect 13916 7158 13972 7196
rect 13916 6916 13972 6926
rect 14028 6916 14084 9548
rect 13916 6914 14084 6916
rect 13916 6862 13918 6914
rect 13970 6862 14084 6914
rect 13916 6860 14084 6862
rect 13916 6850 13972 6860
rect 13692 6638 13694 6690
rect 13746 6638 13748 6690
rect 13692 6626 13748 6638
rect 13468 5854 13470 5906
rect 13522 5854 13524 5906
rect 13468 5842 13524 5854
rect 13580 6580 13636 6590
rect 13580 6356 13636 6524
rect 13356 5058 13412 5068
rect 13468 5460 13524 5470
rect 13356 4340 13412 4350
rect 13356 4246 13412 4284
rect 13020 2718 13022 2770
rect 13074 2718 13076 2770
rect 13020 2706 13076 2718
rect 13132 4114 13188 4126
rect 13132 4062 13134 4114
rect 13186 4062 13188 4114
rect 12908 2146 12964 2156
rect 12796 2100 12852 2110
rect 12796 2006 12852 2044
rect 12348 1988 12404 1998
rect 12348 1894 12404 1932
rect 12236 578 12292 588
rect 12348 1652 12404 1662
rect 12348 112 12404 1596
rect 12572 1652 12628 1662
rect 12572 112 12628 1596
rect 12796 1652 12852 1662
rect 12684 1202 12740 1214
rect 12684 1150 12686 1202
rect 12738 1150 12740 1202
rect 12684 1092 12740 1150
rect 12684 1026 12740 1036
rect 12796 112 12852 1596
rect 13020 1652 13076 1662
rect 13020 112 13076 1596
rect 13132 1204 13188 4062
rect 13356 3444 13412 3454
rect 13244 2996 13300 3006
rect 13244 1988 13300 2940
rect 13356 2436 13412 3388
rect 13468 2548 13524 5404
rect 13580 5348 13636 6300
rect 14140 5906 14196 10108
rect 14924 10050 14980 10780
rect 14924 9998 14926 10050
rect 14978 9998 14980 10050
rect 14924 9986 14980 9998
rect 14588 9938 14644 9950
rect 14588 9886 14590 9938
rect 14642 9886 14644 9938
rect 14588 9268 14644 9886
rect 14588 9202 14644 9212
rect 14700 9492 14756 9502
rect 14476 9156 14532 9166
rect 14364 9044 14420 9054
rect 14364 8950 14420 8988
rect 14476 7588 14532 9100
rect 14588 8932 14644 8942
rect 14588 8838 14644 8876
rect 14588 8260 14644 8270
rect 14588 8166 14644 8204
rect 14588 7588 14644 7598
rect 14476 7586 14644 7588
rect 14476 7534 14590 7586
rect 14642 7534 14644 7586
rect 14476 7532 14644 7534
rect 14140 5854 14142 5906
rect 14194 5854 14196 5906
rect 14140 5842 14196 5854
rect 14252 7250 14308 7262
rect 14252 7198 14254 7250
rect 14306 7198 14308 7250
rect 14252 5908 14308 7198
rect 14364 6692 14420 6702
rect 14364 6598 14420 6636
rect 14476 6468 14532 7532
rect 14588 7522 14644 7532
rect 14476 6402 14532 6412
rect 14700 6356 14756 9436
rect 15036 7474 15092 11118
rect 15708 11172 15764 11182
rect 15708 10498 15764 11116
rect 15708 10446 15710 10498
rect 15762 10446 15764 10498
rect 15708 10434 15764 10446
rect 15260 10388 15316 10398
rect 15148 10386 15316 10388
rect 15148 10334 15262 10386
rect 15314 10334 15316 10386
rect 15148 10332 15316 10334
rect 15148 9042 15204 10332
rect 15260 10322 15316 10332
rect 15708 10164 15764 10174
rect 15260 9938 15316 9950
rect 15260 9886 15262 9938
rect 15314 9886 15316 9938
rect 15260 9716 15316 9886
rect 15484 9828 15540 9838
rect 15260 9650 15316 9660
rect 15372 9826 15540 9828
rect 15372 9774 15486 9826
rect 15538 9774 15540 9826
rect 15372 9772 15540 9774
rect 15148 8990 15150 9042
rect 15202 8990 15204 9042
rect 15148 8978 15204 8990
rect 15036 7422 15038 7474
rect 15090 7422 15092 7474
rect 15036 7410 15092 7422
rect 15148 8370 15204 8382
rect 15148 8318 15150 8370
rect 15202 8318 15204 8370
rect 15148 6804 15204 8318
rect 15372 7700 15428 9772
rect 15484 9762 15540 9772
rect 15596 9042 15652 9054
rect 15596 8990 15598 9042
rect 15650 8990 15652 9042
rect 15484 8820 15540 8830
rect 15484 8370 15540 8764
rect 15484 8318 15486 8370
rect 15538 8318 15540 8370
rect 15484 8306 15540 8318
rect 15596 8148 15652 8990
rect 15148 6738 15204 6748
rect 15260 7644 15428 7700
rect 15484 8092 15652 8148
rect 14924 6690 14980 6702
rect 14924 6638 14926 6690
rect 14978 6638 14980 6690
rect 14700 6290 14756 6300
rect 14812 6468 14868 6478
rect 14812 6018 14868 6412
rect 14812 5966 14814 6018
rect 14866 5966 14868 6018
rect 14812 5954 14868 5966
rect 14252 5852 14420 5908
rect 13916 5684 13972 5694
rect 13916 5682 14196 5684
rect 13916 5630 13918 5682
rect 13970 5630 14196 5682
rect 13916 5628 14196 5630
rect 13916 5618 13972 5628
rect 13580 5282 13636 5292
rect 14028 5348 14084 5358
rect 13916 5124 13972 5134
rect 13580 4564 13636 4574
rect 13580 3778 13636 4508
rect 13580 3726 13582 3778
rect 13634 3726 13636 3778
rect 13580 3714 13636 3726
rect 13692 3556 13748 3566
rect 13692 3462 13748 3500
rect 13692 2996 13748 3006
rect 13692 2882 13748 2940
rect 13692 2830 13694 2882
rect 13746 2830 13748 2882
rect 13692 2818 13748 2830
rect 13468 2492 13748 2548
rect 13356 2380 13524 2436
rect 13244 1922 13300 1932
rect 13132 1138 13188 1148
rect 13244 1652 13300 1662
rect 13132 978 13188 990
rect 13132 926 13134 978
rect 13186 926 13188 978
rect 13132 308 13188 926
rect 13132 242 13188 252
rect 13244 112 13300 1596
rect 13468 112 13524 2380
rect 13692 112 13748 2492
rect 13916 2210 13972 5068
rect 14028 4338 14084 5292
rect 14028 4286 14030 4338
rect 14082 4286 14084 4338
rect 14028 2996 14084 4286
rect 14028 2930 14084 2940
rect 14140 2772 14196 5628
rect 14252 5124 14308 5134
rect 14252 5030 14308 5068
rect 14140 2706 14196 2716
rect 14252 3554 14308 3566
rect 14252 3502 14254 3554
rect 14306 3502 14308 3554
rect 13916 2158 13918 2210
rect 13970 2158 13972 2210
rect 13916 2146 13972 2158
rect 14028 2660 14084 2670
rect 13916 1316 13972 1326
rect 13916 112 13972 1260
rect 14028 308 14084 2604
rect 14028 242 14084 252
rect 14140 2548 14196 2558
rect 14140 112 14196 2492
rect 14252 1426 14308 3502
rect 14364 2212 14420 5852
rect 14700 5684 14756 5694
rect 14476 4114 14532 4126
rect 14476 4062 14478 4114
rect 14530 4062 14532 4114
rect 14476 4004 14532 4062
rect 14476 3938 14532 3948
rect 14588 3556 14644 3566
rect 14588 3462 14644 3500
rect 14700 2660 14756 5628
rect 14924 5572 14980 6638
rect 15260 6132 15316 7644
rect 15372 7476 15428 7486
rect 15372 7382 15428 7420
rect 14924 5506 14980 5516
rect 15148 6076 15316 6132
rect 15036 5234 15092 5246
rect 15036 5182 15038 5234
rect 15090 5182 15092 5234
rect 15036 3108 15092 5182
rect 15148 4900 15204 6076
rect 15148 4834 15204 4844
rect 15260 5906 15316 5918
rect 15260 5854 15262 5906
rect 15314 5854 15316 5906
rect 15148 3554 15204 3566
rect 15148 3502 15150 3554
rect 15202 3502 15204 3554
rect 15148 3444 15204 3502
rect 15148 3378 15204 3388
rect 14700 2594 14756 2604
rect 14924 3052 15092 3108
rect 14364 2156 14532 2212
rect 14364 1988 14420 1998
rect 14364 1894 14420 1932
rect 14476 1764 14532 2156
rect 14252 1374 14254 1426
rect 14306 1374 14308 1426
rect 14252 1362 14308 1374
rect 14364 1708 14532 1764
rect 14700 2098 14756 2110
rect 14700 2046 14702 2098
rect 14754 2046 14756 2098
rect 14364 112 14420 1708
rect 14700 1652 14756 2046
rect 14700 1586 14756 1596
rect 14812 1204 14868 1214
rect 14812 1110 14868 1148
rect 14812 980 14868 990
rect 14924 980 14980 3052
rect 15260 2994 15316 5854
rect 15484 5572 15540 8092
rect 15596 7924 15652 7934
rect 15596 7362 15652 7868
rect 15596 7310 15598 7362
rect 15650 7310 15652 7362
rect 15596 7298 15652 7310
rect 15596 5908 15652 5918
rect 15596 5814 15652 5852
rect 15708 5796 15764 10108
rect 15820 8370 15876 15092
rect 15820 8318 15822 8370
rect 15874 8318 15876 8370
rect 15820 8306 15876 8318
rect 15932 14530 15988 14542
rect 15932 14478 15934 14530
rect 15986 14478 15988 14530
rect 15932 8148 15988 14478
rect 16044 13412 16100 15092
rect 16044 13346 16100 13356
rect 16044 10386 16100 10398
rect 16044 10334 16046 10386
rect 16098 10334 16100 10386
rect 16044 10276 16100 10334
rect 16044 10210 16100 10220
rect 16156 9380 16212 18172
rect 16268 15204 16324 15242
rect 16268 15138 16324 15148
rect 15820 8092 15988 8148
rect 16044 9324 16212 9380
rect 16380 12180 16436 12190
rect 15820 6356 15876 8092
rect 15932 6690 15988 6702
rect 15932 6638 15934 6690
rect 15986 6638 15988 6690
rect 15932 6580 15988 6638
rect 15932 6514 15988 6524
rect 15820 6300 15988 6356
rect 15820 5796 15876 5806
rect 15708 5794 15876 5796
rect 15708 5742 15822 5794
rect 15874 5742 15876 5794
rect 15708 5740 15876 5742
rect 15820 5730 15876 5740
rect 15932 5572 15988 6300
rect 15484 5506 15540 5516
rect 15708 5516 15988 5572
rect 15372 5348 15428 5358
rect 15372 5254 15428 5292
rect 15708 5348 15764 5516
rect 15260 2942 15262 2994
rect 15314 2942 15316 2994
rect 15260 2930 15316 2942
rect 15372 5124 15428 5134
rect 15036 2884 15092 2894
rect 15036 2210 15092 2828
rect 15036 2158 15038 2210
rect 15090 2158 15092 2210
rect 15036 2146 15092 2158
rect 15260 2324 15316 2334
rect 14868 924 14980 980
rect 15036 980 15092 990
rect 14812 914 14868 924
rect 15036 886 15092 924
rect 14588 756 14644 766
rect 14588 112 14644 700
rect 15036 756 15092 766
rect 14812 420 14868 430
rect 14812 112 14868 364
rect 15036 112 15092 700
rect 15260 112 15316 2268
rect 15372 2210 15428 5068
rect 15596 4564 15652 4574
rect 15596 4470 15652 4508
rect 15372 2158 15374 2210
rect 15426 2158 15428 2210
rect 15372 2146 15428 2158
rect 15484 3666 15540 3678
rect 15484 3614 15486 3666
rect 15538 3614 15540 3666
rect 15372 1764 15428 1774
rect 15372 868 15428 1708
rect 15484 1202 15540 3614
rect 15708 3388 15764 5292
rect 15932 5236 15988 5246
rect 15820 5122 15876 5134
rect 15820 5070 15822 5122
rect 15874 5070 15876 5122
rect 15820 3778 15876 5070
rect 15820 3726 15822 3778
rect 15874 3726 15876 3778
rect 15820 3714 15876 3726
rect 15484 1150 15486 1202
rect 15538 1150 15540 1202
rect 15484 1138 15540 1150
rect 15596 3332 15764 3388
rect 15372 812 15540 868
rect 15484 112 15540 812
rect 15596 532 15652 3332
rect 15708 2772 15764 2782
rect 15708 2678 15764 2716
rect 15932 2660 15988 5180
rect 16044 3554 16100 9324
rect 16156 8258 16212 8270
rect 16156 8206 16158 8258
rect 16210 8206 16212 8258
rect 16156 6692 16212 8206
rect 16268 8036 16324 8046
rect 16268 7474 16324 7980
rect 16268 7422 16270 7474
rect 16322 7422 16324 7474
rect 16268 7410 16324 7422
rect 16156 6626 16212 6636
rect 16268 5794 16324 5806
rect 16268 5742 16270 5794
rect 16322 5742 16324 5794
rect 16156 5234 16212 5246
rect 16156 5182 16158 5234
rect 16210 5182 16212 5234
rect 16156 4004 16212 5182
rect 16268 4564 16324 5742
rect 16268 4498 16324 4508
rect 16268 4340 16324 4350
rect 16380 4340 16436 12124
rect 16492 5124 16548 20972
rect 16604 16324 16660 21196
rect 16716 20188 16772 21420
rect 16828 21028 16884 21038
rect 16940 21028 16996 21532
rect 17164 21522 17220 21532
rect 16828 21026 16996 21028
rect 16828 20974 16830 21026
rect 16882 20974 16996 21026
rect 16828 20972 16996 20974
rect 16828 20962 16884 20972
rect 17052 20804 17108 20814
rect 16716 20132 16884 20188
rect 16828 18676 16884 20132
rect 16940 19796 16996 19806
rect 16940 19234 16996 19740
rect 16940 19182 16942 19234
rect 16994 19182 16996 19234
rect 16940 19170 16996 19182
rect 17052 18900 17108 20748
rect 17164 20132 17220 20142
rect 17276 20132 17332 22204
rect 17164 20130 17332 20132
rect 17164 20078 17166 20130
rect 17218 20078 17332 20130
rect 17164 20076 17332 20078
rect 17388 21812 17444 21822
rect 17164 19348 17220 20076
rect 17164 19282 17220 19292
rect 17388 19458 17444 21756
rect 17388 19406 17390 19458
rect 17442 19406 17444 19458
rect 17388 19236 17444 19406
rect 17388 19170 17444 19180
rect 17052 18844 17444 18900
rect 17276 18676 17332 18686
rect 16828 18674 17332 18676
rect 16828 18622 16830 18674
rect 16882 18622 17278 18674
rect 17330 18622 17332 18674
rect 16828 18620 17332 18622
rect 16828 18610 16884 18620
rect 17276 18610 17332 18620
rect 16940 18452 16996 18462
rect 16716 17892 16772 17902
rect 16716 17666 16772 17836
rect 16940 17890 16996 18396
rect 17388 18340 17444 18844
rect 17500 18562 17556 22764
rect 17612 22596 17668 22878
rect 17612 22530 17668 22540
rect 17612 22260 17668 22270
rect 17612 22166 17668 22204
rect 17724 21588 17780 21598
rect 17836 21588 17892 26852
rect 17948 26852 18004 26862
rect 17948 26758 18004 26796
rect 18060 26628 18116 29932
rect 18284 29426 18340 29932
rect 18284 29374 18286 29426
rect 18338 29374 18340 29426
rect 18284 29362 18340 29374
rect 18732 29540 18788 31502
rect 18844 31444 18900 32508
rect 18956 32498 19012 32508
rect 19404 32562 19460 32574
rect 19404 32510 19406 32562
rect 19458 32510 19460 32562
rect 19068 31892 19124 31902
rect 19068 31798 19124 31836
rect 19292 31780 19348 31790
rect 19292 31686 19348 31724
rect 19404 31556 19460 32510
rect 19516 32338 19572 33068
rect 19852 32564 19908 32574
rect 19516 32286 19518 32338
rect 19570 32286 19572 32338
rect 19516 32274 19572 32286
rect 19740 32452 19796 32462
rect 19404 31490 19460 31500
rect 19516 31778 19572 31790
rect 19516 31726 19518 31778
rect 19570 31726 19572 31778
rect 18844 31378 18900 31388
rect 19516 31108 19572 31726
rect 19628 31668 19684 31678
rect 19628 31574 19684 31612
rect 19740 31444 19796 32396
rect 19404 31052 19572 31108
rect 19628 31388 19796 31444
rect 19292 30882 19348 30894
rect 19292 30830 19294 30882
rect 19346 30830 19348 30882
rect 18844 30772 18900 30782
rect 18844 30678 18900 30716
rect 18844 30548 18900 30558
rect 18844 30434 18900 30492
rect 18844 30382 18846 30434
rect 18898 30382 18900 30434
rect 18844 30370 18900 30382
rect 18620 28868 18676 28878
rect 18620 28774 18676 28812
rect 18396 28644 18452 28654
rect 18396 27858 18452 28588
rect 18396 27806 18398 27858
rect 18450 27806 18452 27858
rect 18396 26908 18452 27806
rect 18508 28532 18564 28542
rect 18508 27186 18564 28476
rect 18732 27972 18788 29484
rect 19068 30100 19124 30110
rect 18844 29428 18900 29438
rect 18844 29334 18900 29372
rect 19068 28532 19124 30044
rect 19068 28438 19124 28476
rect 19180 28084 19236 28094
rect 18732 27916 18900 27972
rect 18732 27748 18788 27758
rect 18732 27654 18788 27692
rect 18732 27524 18788 27534
rect 18620 27300 18676 27310
rect 18620 27206 18676 27244
rect 18508 27134 18510 27186
rect 18562 27134 18564 27186
rect 18508 27122 18564 27134
rect 18732 26964 18788 27468
rect 18844 27076 18900 27916
rect 19180 27298 19236 28028
rect 19292 27636 19348 30830
rect 19292 27570 19348 27580
rect 19404 27412 19460 31052
rect 19516 30882 19572 30894
rect 19516 30830 19518 30882
rect 19570 30830 19572 30882
rect 19516 29988 19572 30830
rect 19628 30100 19684 31388
rect 19628 30034 19684 30044
rect 19740 30994 19796 31006
rect 19740 30942 19742 30994
rect 19794 30942 19796 30994
rect 19516 29428 19572 29932
rect 19516 28532 19572 29372
rect 19628 28756 19684 28766
rect 19740 28756 19796 30942
rect 19852 29426 19908 32508
rect 19964 30212 20020 33292
rect 20076 33124 20132 33134
rect 20076 33030 20132 33068
rect 20076 30996 20132 31006
rect 20076 30902 20132 30940
rect 20076 30770 20132 30782
rect 20076 30718 20078 30770
rect 20130 30718 20132 30770
rect 20076 30548 20132 30718
rect 20076 30482 20132 30492
rect 19964 30156 20132 30212
rect 19852 29374 19854 29426
rect 19906 29374 19908 29426
rect 19852 28868 19908 29374
rect 19852 28802 19908 28812
rect 19964 29988 20020 29998
rect 19628 28754 19796 28756
rect 19628 28702 19630 28754
rect 19682 28702 19796 28754
rect 19628 28700 19796 28702
rect 19628 28690 19684 28700
rect 19964 28642 20020 29932
rect 19964 28590 19966 28642
rect 20018 28590 20020 28642
rect 19740 28532 19796 28542
rect 19516 28530 19796 28532
rect 19516 28478 19742 28530
rect 19794 28478 19796 28530
rect 19516 28476 19796 28478
rect 19516 28084 19572 28476
rect 19740 28466 19796 28476
rect 19964 28308 20020 28590
rect 20076 28644 20132 30156
rect 20076 28578 20132 28588
rect 19516 28018 19572 28028
rect 19740 28252 20020 28308
rect 20076 28420 20132 28430
rect 19180 27246 19182 27298
rect 19234 27246 19236 27298
rect 19180 27234 19236 27246
rect 19292 27356 19460 27412
rect 19292 27300 19348 27356
rect 19292 27188 19348 27244
rect 19628 27188 19684 27198
rect 19292 27186 19684 27188
rect 19292 27134 19294 27186
rect 19346 27134 19630 27186
rect 19682 27134 19684 27186
rect 19292 27132 19684 27134
rect 19292 27122 19348 27132
rect 19628 27122 19684 27132
rect 19740 27186 19796 28252
rect 19964 28084 20020 28094
rect 19964 27990 20020 28028
rect 19740 27134 19742 27186
rect 19794 27134 19796 27186
rect 19740 27122 19796 27134
rect 19852 27748 19908 27758
rect 18844 27010 18900 27020
rect 19180 27076 19236 27086
rect 18620 26908 18788 26964
rect 18396 26852 18564 26908
rect 18060 26572 18228 26628
rect 18060 26068 18116 26078
rect 17948 25732 18004 25742
rect 17948 25638 18004 25676
rect 18060 25618 18116 26012
rect 18060 25566 18062 25618
rect 18114 25566 18116 25618
rect 18060 25554 18116 25566
rect 17724 21586 17836 21588
rect 17724 21534 17726 21586
rect 17778 21534 17836 21586
rect 17724 21532 17836 21534
rect 17724 21522 17780 21532
rect 17836 21522 17892 21532
rect 17948 24612 18004 24622
rect 17836 21362 17892 21374
rect 17836 21310 17838 21362
rect 17890 21310 17892 21362
rect 17500 18510 17502 18562
rect 17554 18510 17556 18562
rect 17500 18498 17556 18510
rect 17612 20916 17668 20926
rect 17612 20130 17668 20860
rect 17612 20078 17614 20130
rect 17666 20078 17668 20130
rect 17500 18340 17556 18350
rect 17388 18338 17556 18340
rect 17388 18286 17502 18338
rect 17554 18286 17556 18338
rect 17388 18284 17556 18286
rect 17500 18274 17556 18284
rect 17612 18004 17668 20078
rect 17724 19906 17780 19918
rect 17724 19854 17726 19906
rect 17778 19854 17780 19906
rect 17724 19460 17780 19854
rect 17724 19394 17780 19404
rect 16940 17838 16942 17890
rect 16994 17838 16996 17890
rect 16940 17826 16996 17838
rect 17052 17948 17668 18004
rect 17724 19236 17780 19246
rect 17052 17778 17108 17948
rect 17724 17892 17780 19180
rect 17836 18228 17892 21310
rect 17948 19908 18004 24556
rect 18060 24388 18116 24398
rect 18060 23044 18116 24332
rect 18172 23716 18228 26572
rect 18172 23650 18228 23660
rect 18284 26404 18340 26414
rect 18060 22978 18116 22988
rect 18060 22596 18116 22606
rect 18284 22596 18340 26348
rect 18508 25396 18564 26852
rect 18620 26850 18676 26908
rect 18620 26798 18622 26850
rect 18674 26798 18676 26850
rect 18620 26786 18676 26798
rect 19068 26852 19124 26862
rect 18732 26516 18788 26526
rect 18620 25396 18676 25406
rect 18508 25340 18620 25396
rect 18060 22594 18340 22596
rect 18060 22542 18062 22594
rect 18114 22542 18340 22594
rect 18060 22540 18340 22542
rect 18396 23940 18452 23950
rect 18396 23156 18452 23884
rect 18060 22530 18116 22540
rect 18060 22372 18116 22382
rect 18060 20914 18116 22316
rect 18396 22260 18452 23100
rect 18396 21812 18452 22204
rect 18396 21756 18564 21812
rect 18060 20862 18062 20914
rect 18114 20862 18116 20914
rect 18060 20850 18116 20862
rect 18172 21588 18228 21598
rect 17948 19842 18004 19852
rect 18060 20580 18116 20590
rect 17948 19124 18004 19134
rect 17948 18450 18004 19068
rect 18060 18562 18116 20524
rect 18060 18510 18062 18562
rect 18114 18510 18116 18562
rect 18060 18498 18116 18510
rect 17948 18398 17950 18450
rect 18002 18398 18004 18450
rect 17948 18386 18004 18398
rect 17836 18162 17892 18172
rect 17052 17726 17054 17778
rect 17106 17726 17108 17778
rect 17052 17714 17108 17726
rect 17612 17836 17780 17892
rect 16716 17614 16718 17666
rect 16770 17614 16772 17666
rect 16716 17602 16772 17614
rect 16716 16324 16772 16334
rect 16604 16322 16772 16324
rect 16604 16270 16718 16322
rect 16770 16270 16772 16322
rect 16604 16268 16772 16270
rect 16716 16258 16772 16268
rect 17388 16210 17444 16222
rect 17388 16158 17390 16210
rect 17442 16158 17444 16210
rect 17052 16098 17108 16110
rect 17052 16046 17054 16098
rect 17106 16046 17108 16098
rect 17052 15652 17108 16046
rect 17052 15586 17108 15596
rect 17388 15540 17444 16158
rect 17388 15474 17444 15484
rect 17500 15092 17556 15102
rect 17388 15090 17556 15092
rect 17388 15038 17502 15090
rect 17554 15038 17556 15090
rect 17388 15036 17556 15038
rect 17164 14532 17220 14542
rect 17388 14532 17444 15036
rect 17500 15026 17556 15036
rect 17164 14530 17444 14532
rect 17164 14478 17166 14530
rect 17218 14478 17444 14530
rect 17164 14476 17444 14478
rect 17500 14532 17556 14542
rect 17164 14466 17220 14476
rect 17500 14438 17556 14476
rect 16716 14420 16772 14430
rect 16716 14418 16884 14420
rect 16716 14366 16718 14418
rect 16770 14366 16884 14418
rect 16716 14364 16884 14366
rect 16716 14354 16772 14364
rect 16604 13748 16660 13758
rect 16828 13748 16884 14364
rect 16604 13746 16772 13748
rect 16604 13694 16606 13746
rect 16658 13694 16772 13746
rect 16604 13692 16772 13694
rect 16604 13682 16660 13692
rect 16604 13524 16660 13534
rect 16604 9042 16660 13468
rect 16716 13412 16772 13692
rect 16828 13682 16884 13692
rect 16940 13636 16996 13646
rect 16940 13542 16996 13580
rect 17276 13636 17332 13646
rect 16716 12180 16772 13356
rect 17052 13074 17108 13086
rect 17052 13022 17054 13074
rect 17106 13022 17108 13074
rect 16716 12086 16772 12124
rect 16828 12628 16884 12638
rect 16716 10052 16772 10062
rect 16716 9958 16772 9996
rect 16604 8990 16606 9042
rect 16658 8990 16660 9042
rect 16604 6580 16660 8990
rect 16828 9044 16884 12572
rect 17052 12404 17108 13022
rect 17052 12338 17108 12348
rect 17164 11954 17220 11966
rect 17164 11902 17166 11954
rect 17218 11902 17220 11954
rect 17164 11732 17220 11902
rect 17164 11666 17220 11676
rect 16828 8978 16884 8988
rect 16940 10610 16996 10622
rect 16940 10558 16942 10610
rect 16994 10558 16996 10610
rect 16940 9828 16996 10558
rect 17276 10498 17332 13580
rect 17388 12962 17444 12974
rect 17388 12910 17390 12962
rect 17442 12910 17444 12962
rect 17388 11620 17444 12910
rect 17612 11844 17668 17836
rect 18060 16882 18116 16894
rect 18060 16830 18062 16882
rect 18114 16830 18116 16882
rect 17948 16660 18004 16670
rect 17724 16100 17780 16110
rect 17724 16098 17892 16100
rect 17724 16046 17726 16098
rect 17778 16046 17892 16098
rect 17724 16044 17892 16046
rect 17724 16034 17780 16044
rect 17724 15652 17780 15662
rect 17724 14754 17780 15596
rect 17724 14702 17726 14754
rect 17778 14702 17780 14754
rect 17724 14690 17780 14702
rect 17724 13748 17780 13758
rect 17724 13074 17780 13692
rect 17836 13524 17892 16044
rect 17836 13458 17892 13468
rect 17948 15428 18004 16604
rect 17724 13022 17726 13074
rect 17778 13022 17780 13074
rect 17724 13010 17780 13022
rect 17612 11778 17668 11788
rect 17724 12740 17780 12750
rect 17388 11554 17444 11564
rect 17276 10446 17278 10498
rect 17330 10446 17332 10498
rect 17276 10434 17332 10446
rect 17388 10386 17444 10398
rect 17388 10334 17390 10386
rect 17442 10334 17444 10386
rect 16828 8036 16884 8046
rect 16828 7942 16884 7980
rect 16940 7812 16996 9772
rect 16940 7746 16996 7756
rect 17052 9826 17108 9838
rect 17052 9774 17054 9826
rect 17106 9774 17108 9826
rect 16716 7474 16772 7486
rect 16716 7422 16718 7474
rect 16770 7422 16772 7474
rect 16716 6692 16772 7422
rect 16940 6692 16996 6702
rect 16716 6690 16996 6692
rect 16716 6638 16942 6690
rect 16994 6638 16996 6690
rect 16716 6636 16996 6638
rect 16604 6514 16660 6524
rect 16828 5906 16884 6636
rect 16940 6626 16996 6636
rect 16828 5854 16830 5906
rect 16882 5854 16884 5906
rect 16828 5572 16884 5854
rect 16828 5506 16884 5516
rect 16940 6356 16996 6366
rect 16492 5058 16548 5068
rect 16324 4284 16436 4340
rect 16268 4246 16324 4284
rect 16604 4226 16660 4238
rect 16604 4174 16606 4226
rect 16658 4174 16660 4226
rect 16156 3948 16324 4004
rect 16044 3502 16046 3554
rect 16098 3502 16100 3554
rect 16044 3490 16100 3502
rect 16268 3388 16324 3948
rect 16156 3332 16324 3388
rect 16604 3388 16660 4174
rect 16940 3780 16996 6300
rect 17052 5012 17108 9774
rect 17276 9156 17332 9166
rect 17276 9062 17332 9100
rect 17388 8932 17444 10334
rect 17388 8484 17444 8876
rect 17388 8418 17444 8428
rect 17724 8036 17780 12684
rect 17948 11732 18004 15372
rect 18060 15988 18116 16830
rect 18060 15316 18116 15932
rect 18060 15222 18116 15260
rect 18172 15764 18228 21532
rect 18396 21588 18452 21598
rect 18396 21494 18452 21532
rect 18508 21364 18564 21756
rect 18396 21308 18564 21364
rect 18396 20802 18452 21308
rect 18396 20750 18398 20802
rect 18450 20750 18452 20802
rect 18396 20738 18452 20750
rect 18396 20018 18452 20030
rect 18396 19966 18398 20018
rect 18450 19966 18452 20018
rect 18396 19908 18452 19966
rect 18396 19842 18452 19852
rect 18620 19908 18676 25340
rect 18620 19842 18676 19852
rect 18284 19460 18340 19470
rect 18284 18674 18340 19404
rect 18508 19460 18564 19470
rect 18508 19366 18564 19404
rect 18284 18622 18286 18674
rect 18338 18622 18340 18674
rect 18284 18610 18340 18622
rect 18508 18004 18564 18014
rect 18284 17778 18340 17790
rect 18284 17726 18286 17778
rect 18338 17726 18340 17778
rect 18284 17444 18340 17726
rect 18284 17378 18340 17388
rect 18508 16884 18564 17948
rect 18620 17780 18676 17790
rect 18620 17686 18676 17724
rect 18508 16770 18564 16828
rect 18508 16718 18510 16770
rect 18562 16718 18564 16770
rect 18508 16706 18564 16718
rect 18172 15148 18228 15708
rect 18620 15204 18676 15214
rect 18732 15204 18788 26460
rect 18956 25284 19012 25294
rect 18844 23044 18900 23054
rect 18844 22148 18900 22988
rect 18844 22082 18900 22092
rect 18844 19794 18900 19806
rect 18844 19742 18846 19794
rect 18898 19742 18900 19794
rect 18844 16772 18900 19742
rect 18956 19348 19012 25228
rect 19068 21586 19124 26796
rect 19180 26850 19236 27020
rect 19180 26798 19182 26850
rect 19234 26798 19236 26850
rect 19180 26786 19236 26798
rect 19516 26964 19572 26974
rect 19852 26908 19908 27692
rect 20076 27300 20132 28364
rect 20076 27234 20132 27244
rect 19516 25284 19572 26908
rect 19516 25218 19572 25228
rect 19740 26852 19908 26908
rect 19404 23938 19460 23950
rect 19404 23886 19406 23938
rect 19458 23886 19460 23938
rect 19404 23268 19460 23886
rect 19628 23938 19684 23950
rect 19628 23886 19630 23938
rect 19682 23886 19684 23938
rect 19068 21534 19070 21586
rect 19122 21534 19124 21586
rect 19068 19572 19124 21534
rect 19180 22146 19236 22158
rect 19180 22094 19182 22146
rect 19234 22094 19236 22146
rect 19180 21588 19236 22094
rect 19180 21522 19236 21532
rect 19292 21252 19348 21262
rect 19180 20690 19236 20702
rect 19180 20638 19182 20690
rect 19234 20638 19236 20690
rect 19180 19908 19236 20638
rect 19180 19842 19236 19852
rect 19068 19506 19124 19516
rect 18956 19292 19124 19348
rect 18956 17892 19012 17902
rect 18956 17778 19012 17836
rect 18956 17726 18958 17778
rect 19010 17726 19012 17778
rect 18956 17714 19012 17726
rect 18844 16706 18900 16716
rect 18620 15202 18788 15204
rect 18620 15150 18622 15202
rect 18674 15150 18788 15202
rect 18620 15148 18788 15150
rect 18172 15092 18564 15148
rect 18620 15138 18676 15148
rect 18172 14530 18228 14542
rect 18172 14478 18174 14530
rect 18226 14478 18228 14530
rect 18172 13970 18228 14478
rect 18172 13918 18174 13970
rect 18226 13918 18228 13970
rect 18172 13906 18228 13918
rect 18396 14532 18452 14542
rect 18284 13860 18340 13870
rect 18172 12962 18228 12974
rect 18172 12910 18174 12962
rect 18226 12910 18228 12962
rect 18172 12404 18228 12910
rect 18284 12852 18340 13804
rect 18284 12786 18340 12796
rect 18284 12404 18340 12414
rect 18172 12402 18340 12404
rect 18172 12350 18286 12402
rect 18338 12350 18340 12402
rect 18172 12348 18340 12350
rect 18284 12338 18340 12348
rect 17948 11666 18004 11676
rect 18172 11508 18228 11518
rect 18396 11508 18452 14476
rect 18508 14196 18564 15092
rect 18732 14868 18788 15148
rect 18732 14802 18788 14812
rect 18956 15876 19012 15886
rect 19068 15876 19124 19292
rect 19012 15820 19124 15876
rect 19180 18900 19236 18910
rect 18732 14532 18788 14542
rect 18732 14438 18788 14476
rect 18508 14140 18900 14196
rect 18732 13524 18788 13534
rect 18732 13186 18788 13468
rect 18732 13134 18734 13186
rect 18786 13134 18788 13186
rect 18732 13122 18788 13134
rect 18620 12964 18676 12974
rect 18732 12964 18788 12974
rect 18620 12962 18732 12964
rect 18620 12910 18622 12962
rect 18674 12910 18732 12962
rect 18620 12908 18732 12910
rect 18620 12898 18676 12908
rect 18172 11506 18452 11508
rect 18172 11454 18174 11506
rect 18226 11454 18452 11506
rect 18172 11452 18452 11454
rect 18620 12068 18676 12078
rect 18172 11442 18228 11452
rect 18508 11394 18564 11406
rect 18508 11342 18510 11394
rect 18562 11342 18564 11394
rect 18508 10834 18564 11342
rect 18508 10782 18510 10834
rect 18562 10782 18564 10834
rect 18508 10770 18564 10782
rect 18508 10388 18564 10398
rect 18396 9940 18452 9950
rect 18060 9828 18116 9838
rect 18060 9734 18116 9772
rect 17948 8372 18004 8382
rect 17612 7474 17668 7486
rect 17612 7422 17614 7474
rect 17666 7422 17668 7474
rect 17500 7140 17556 7150
rect 17500 5234 17556 7084
rect 17612 6580 17668 7422
rect 17724 6692 17780 7980
rect 17836 8316 17948 8372
rect 17836 7252 17892 8316
rect 17948 8278 18004 8316
rect 18396 8258 18452 9884
rect 18508 9938 18564 10332
rect 18508 9886 18510 9938
rect 18562 9886 18564 9938
rect 18508 9874 18564 9886
rect 18508 8932 18564 8942
rect 18620 8932 18676 12012
rect 18508 8930 18676 8932
rect 18508 8878 18510 8930
rect 18562 8878 18676 8930
rect 18508 8876 18676 8878
rect 18508 8866 18564 8876
rect 18396 8206 18398 8258
rect 18450 8206 18452 8258
rect 18396 8148 18452 8206
rect 18396 7586 18452 8092
rect 18396 7534 18398 7586
rect 18450 7534 18452 7586
rect 18396 7522 18452 7534
rect 18508 8708 18564 8718
rect 17836 7186 17892 7196
rect 18060 6804 18116 6814
rect 17724 6636 17892 6692
rect 17668 6524 17780 6580
rect 17612 6514 17668 6524
rect 17724 5908 17780 6524
rect 17836 6356 17892 6636
rect 18060 6690 18116 6748
rect 18060 6638 18062 6690
rect 18114 6638 18116 6690
rect 18060 6626 18116 6638
rect 18284 6580 18340 6590
rect 17836 6300 18116 6356
rect 17836 5908 17892 5918
rect 17724 5906 17892 5908
rect 17724 5854 17838 5906
rect 17890 5854 17892 5906
rect 17724 5852 17892 5854
rect 17836 5842 17892 5852
rect 17500 5182 17502 5234
rect 17554 5182 17556 5234
rect 17052 4946 17108 4956
rect 17164 5010 17220 5022
rect 17164 4958 17166 5010
rect 17218 4958 17220 5010
rect 17164 4564 17220 4958
rect 17164 4498 17220 4508
rect 17052 3780 17108 3790
rect 16940 3778 17108 3780
rect 16940 3726 17054 3778
rect 17106 3726 17108 3778
rect 16940 3724 17108 3726
rect 17052 3714 17108 3724
rect 16828 3556 16884 3566
rect 16828 3462 16884 3500
rect 16604 3332 16772 3388
rect 16044 2660 16100 2670
rect 15932 2658 16100 2660
rect 15932 2606 16046 2658
rect 16098 2606 16100 2658
rect 15932 2604 16100 2606
rect 16044 2594 16100 2604
rect 15708 2212 15764 2222
rect 15708 2118 15764 2156
rect 16044 2100 16100 2110
rect 16044 2006 16100 2044
rect 16156 1764 16212 3332
rect 16716 3108 16772 3332
rect 16604 2996 16660 3006
rect 16604 2882 16660 2940
rect 16604 2830 16606 2882
rect 16658 2830 16660 2882
rect 16604 2818 16660 2830
rect 16716 2884 16772 3052
rect 16716 2818 16772 2828
rect 17052 2884 17108 2894
rect 17052 2658 17108 2828
rect 17052 2606 17054 2658
rect 17106 2606 17108 2658
rect 17052 2594 17108 2606
rect 16940 2548 16996 2558
rect 16828 2100 16884 2110
rect 15932 1708 16212 1764
rect 16716 2098 16884 2100
rect 16716 2046 16830 2098
rect 16882 2046 16884 2098
rect 16716 2044 16884 2046
rect 15708 978 15764 990
rect 15708 926 15710 978
rect 15762 926 15764 978
rect 15708 868 15764 926
rect 15708 802 15764 812
rect 15596 466 15652 476
rect 15708 644 15764 654
rect 15708 112 15764 588
rect 15932 112 15988 1708
rect 16604 980 16660 990
rect 16380 978 16660 980
rect 16380 926 16606 978
rect 16658 926 16660 978
rect 16380 924 16660 926
rect 16156 868 16212 878
rect 16156 112 16212 812
rect 16380 112 16436 924
rect 16604 914 16660 924
rect 16716 756 16772 2044
rect 16828 2034 16884 2044
rect 16940 1316 16996 2492
rect 17500 2212 17556 5182
rect 17836 5460 17892 5470
rect 17724 5124 17780 5134
rect 17724 3666 17780 5068
rect 17836 4562 17892 5404
rect 17836 4510 17838 4562
rect 17890 4510 17892 4562
rect 17836 4498 17892 4510
rect 17724 3614 17726 3666
rect 17778 3614 17780 3666
rect 17724 3602 17780 3614
rect 17500 2146 17556 2156
rect 17612 2996 17668 3006
rect 17164 2100 17220 2110
rect 17164 2006 17220 2044
rect 17612 1986 17668 2940
rect 17612 1934 17614 1986
rect 17666 1934 17668 1986
rect 17612 1922 17668 1934
rect 16604 700 16772 756
rect 16828 1260 16996 1316
rect 17836 1876 17892 1886
rect 17836 1314 17892 1820
rect 17836 1262 17838 1314
rect 17890 1262 17892 1314
rect 16604 112 16660 700
rect 16828 112 16884 1260
rect 17836 1250 17892 1262
rect 17500 1092 17556 1102
rect 18060 1092 18116 6300
rect 18284 5124 18340 6524
rect 18284 5058 18340 5068
rect 18396 5682 18452 5694
rect 18396 5630 18398 5682
rect 18450 5630 18452 5682
rect 18284 4340 18340 4350
rect 18284 4246 18340 4284
rect 18396 3668 18452 5630
rect 18396 3602 18452 3612
rect 18172 3554 18228 3566
rect 18172 3502 18174 3554
rect 18226 3502 18228 3554
rect 18172 2994 18228 3502
rect 18508 3554 18564 8652
rect 18732 7700 18788 12908
rect 18844 11396 18900 14140
rect 18956 12964 19012 15820
rect 18956 12898 19012 12908
rect 19068 14868 19124 14878
rect 18956 11396 19012 11406
rect 18844 11394 19012 11396
rect 18844 11342 18958 11394
rect 19010 11342 19012 11394
rect 18844 11340 19012 11342
rect 18844 9156 18900 9166
rect 18844 9062 18900 9100
rect 18956 8708 19012 11340
rect 18956 8642 19012 8652
rect 19068 8372 19124 14812
rect 19180 13188 19236 18844
rect 19180 13122 19236 13132
rect 19180 11620 19236 11630
rect 19180 11526 19236 11564
rect 19068 8306 19124 8316
rect 19180 9492 19236 9502
rect 19180 9044 19236 9436
rect 19180 8258 19236 8988
rect 19180 8206 19182 8258
rect 19234 8206 19236 8258
rect 19180 8194 19236 8206
rect 18732 7634 18788 7644
rect 18844 7476 18900 7486
rect 18844 7362 18900 7420
rect 18844 7310 18846 7362
rect 18898 7310 18900 7362
rect 18844 7298 18900 7310
rect 18956 7364 19012 7374
rect 18620 6692 18676 6702
rect 18620 6690 18788 6692
rect 18620 6638 18622 6690
rect 18674 6638 18788 6690
rect 18620 6636 18788 6638
rect 18620 6626 18676 6636
rect 18620 5906 18676 5918
rect 18620 5854 18622 5906
rect 18674 5854 18676 5906
rect 18620 4676 18676 5854
rect 18732 5346 18788 6636
rect 18956 6356 19012 7308
rect 19068 6802 19124 6814
rect 19068 6750 19070 6802
rect 19122 6750 19124 6802
rect 19068 6692 19124 6750
rect 19068 6626 19124 6636
rect 19180 6690 19236 6702
rect 19180 6638 19182 6690
rect 19234 6638 19236 6690
rect 19180 6580 19236 6638
rect 19180 6514 19236 6524
rect 19292 6468 19348 21196
rect 19404 18228 19460 23212
rect 19516 23714 19572 23726
rect 19516 23662 19518 23714
rect 19570 23662 19572 23714
rect 19516 21924 19572 23662
rect 19516 21858 19572 21868
rect 19628 21140 19684 23886
rect 19628 21074 19684 21084
rect 19740 22258 19796 26852
rect 20188 24388 20244 35084
rect 20300 35138 20356 38108
rect 20524 36372 20580 38220
rect 20524 36306 20580 36316
rect 20300 35086 20302 35138
rect 20354 35086 20356 35138
rect 20300 32564 20356 35086
rect 20300 32498 20356 32508
rect 20524 35364 20580 35374
rect 20524 32562 20580 35308
rect 20524 32510 20526 32562
rect 20578 32510 20580 32562
rect 20524 32498 20580 32510
rect 20636 32340 20692 38332
rect 20748 35924 20804 38612
rect 20860 37938 20916 38782
rect 21084 38164 21140 40572
rect 21084 38098 21140 38108
rect 20860 37886 20862 37938
rect 20914 37886 20916 37938
rect 20860 37492 20916 37886
rect 20860 37436 21140 37492
rect 20748 35858 20804 35868
rect 20860 37266 20916 37278
rect 20860 37214 20862 37266
rect 20914 37214 20916 37266
rect 20860 36482 20916 37214
rect 20860 36430 20862 36482
rect 20914 36430 20916 36482
rect 20748 35476 20804 35486
rect 20748 35026 20804 35420
rect 20860 35252 20916 36430
rect 20860 35186 20916 35196
rect 20972 35812 21028 35822
rect 20748 34974 20750 35026
rect 20802 34974 20804 35026
rect 20748 33458 20804 34974
rect 20972 34242 21028 35756
rect 21084 34692 21140 37436
rect 21196 35140 21252 42140
rect 21308 41972 21364 41982
rect 21308 40740 21364 41916
rect 21420 41970 21476 41982
rect 21420 41918 21422 41970
rect 21474 41918 21476 41970
rect 21420 41524 21476 41918
rect 21532 41972 21588 42478
rect 21532 41906 21588 41916
rect 21644 41860 21700 41870
rect 21644 41766 21700 41804
rect 21420 41458 21476 41468
rect 21756 41748 21812 41758
rect 21756 41410 21812 41692
rect 21756 41358 21758 41410
rect 21810 41358 21812 41410
rect 21756 41346 21812 41358
rect 21308 40674 21364 40684
rect 21532 40852 21588 40862
rect 21532 40402 21588 40796
rect 21532 40350 21534 40402
rect 21586 40350 21588 40402
rect 21532 40338 21588 40350
rect 21644 40516 21700 40526
rect 21308 40292 21364 40302
rect 21308 38388 21364 40236
rect 21644 40290 21700 40460
rect 21644 40238 21646 40290
rect 21698 40238 21700 40290
rect 21644 40226 21700 40238
rect 21420 38724 21476 38762
rect 21868 38724 21924 44828
rect 22204 44548 22260 55412
rect 22204 44482 22260 44492
rect 22316 45890 22372 45902
rect 22316 45838 22318 45890
rect 22370 45838 22372 45890
rect 22092 43540 22148 43550
rect 22092 43446 22148 43484
rect 22316 42420 22372 45838
rect 21476 38668 21924 38724
rect 21980 42364 22372 42420
rect 21420 38658 21476 38668
rect 21308 38332 21588 38388
rect 21308 38162 21364 38174
rect 21308 38110 21310 38162
rect 21362 38110 21364 38162
rect 21308 37940 21364 38110
rect 21308 37874 21364 37884
rect 21308 37492 21364 37502
rect 21308 36820 21364 37436
rect 21420 37044 21476 37054
rect 21420 36950 21476 36988
rect 21308 36764 21476 36820
rect 21308 36594 21364 36606
rect 21308 36542 21310 36594
rect 21362 36542 21364 36594
rect 21308 36372 21364 36542
rect 21308 36306 21364 36316
rect 21420 35924 21476 36764
rect 21196 35074 21252 35084
rect 21308 35868 21476 35924
rect 21196 34916 21252 34926
rect 21308 34916 21364 35868
rect 21420 35700 21476 35710
rect 21532 35700 21588 38332
rect 21980 37940 22036 42364
rect 22092 41972 22148 41982
rect 22092 41858 22148 41916
rect 22092 41806 22094 41858
rect 22146 41806 22148 41858
rect 22092 40516 22148 41806
rect 22428 40964 22484 60844
rect 22652 60786 22708 60798
rect 22652 60734 22654 60786
rect 22706 60734 22708 60786
rect 22652 60676 22708 60734
rect 22652 60610 22708 60620
rect 22988 55468 23044 62132
rect 24464 61964 24728 61974
rect 24520 61908 24568 61964
rect 24624 61908 24672 61964
rect 24464 61898 24728 61908
rect 23804 61180 24068 61190
rect 23860 61124 23908 61180
rect 23964 61124 24012 61180
rect 23804 61114 24068 61124
rect 23660 60788 23716 60798
rect 23660 60694 23716 60732
rect 24464 60396 24728 60406
rect 24520 60340 24568 60396
rect 24624 60340 24672 60396
rect 24464 60330 24728 60340
rect 23804 59612 24068 59622
rect 23860 59556 23908 59612
rect 23964 59556 24012 59612
rect 23804 59546 24068 59556
rect 24464 58828 24728 58838
rect 24520 58772 24568 58828
rect 24624 58772 24672 58828
rect 24464 58762 24728 58772
rect 23804 58044 24068 58054
rect 23860 57988 23908 58044
rect 23964 57988 24012 58044
rect 23804 57978 24068 57988
rect 22540 55412 23044 55468
rect 23436 57876 23492 57886
rect 22540 45892 22596 55412
rect 22652 47460 22708 47470
rect 22652 46114 22708 47404
rect 23212 46452 23268 46462
rect 23212 46358 23268 46396
rect 22652 46062 22654 46114
rect 22706 46062 22708 46114
rect 22652 46050 22708 46062
rect 22764 46228 22820 46238
rect 22652 45892 22708 45902
rect 22540 45836 22652 45892
rect 22428 40898 22484 40908
rect 22540 44548 22596 44558
rect 22092 40450 22148 40460
rect 22204 40740 22260 40750
rect 22540 40740 22596 44492
rect 22652 44546 22708 45836
rect 22652 44494 22654 44546
rect 22706 44494 22708 44546
rect 22652 44482 22708 44494
rect 22652 43538 22708 43550
rect 22652 43486 22654 43538
rect 22706 43486 22708 43538
rect 22652 42084 22708 43486
rect 22764 42866 22820 46172
rect 23212 45220 23268 45230
rect 23100 44212 23156 44222
rect 23100 44118 23156 44156
rect 22764 42814 22766 42866
rect 22818 42814 22820 42866
rect 22764 42802 22820 42814
rect 23212 42756 23268 45164
rect 23212 42754 23380 42756
rect 23212 42702 23214 42754
rect 23266 42702 23380 42754
rect 23212 42700 23380 42702
rect 23212 42690 23268 42700
rect 22652 41970 22708 42028
rect 22652 41918 22654 41970
rect 22706 41918 22708 41970
rect 22652 41906 22708 41918
rect 22876 41412 22932 41422
rect 22876 41318 22932 41356
rect 23324 41186 23380 42700
rect 23324 41134 23326 41186
rect 23378 41134 23380 41186
rect 23324 41122 23380 41134
rect 22204 40402 22260 40684
rect 22204 40350 22206 40402
rect 22258 40350 22260 40402
rect 22204 40338 22260 40350
rect 22428 40684 22596 40740
rect 22988 40852 23044 40862
rect 21980 37874 22036 37884
rect 22204 38388 22260 38398
rect 21756 35700 21812 35710
rect 21532 35698 21812 35700
rect 21532 35646 21758 35698
rect 21810 35646 21812 35698
rect 21532 35644 21812 35646
rect 21420 35606 21476 35644
rect 21532 34916 21588 34926
rect 21308 34914 21588 34916
rect 21308 34862 21534 34914
rect 21586 34862 21588 34914
rect 21308 34860 21588 34862
rect 21196 34822 21252 34860
rect 21084 34636 21364 34692
rect 20972 34190 20974 34242
rect 21026 34190 21028 34242
rect 20972 34178 21028 34190
rect 21196 34356 21252 34366
rect 20748 33406 20750 33458
rect 20802 33406 20804 33458
rect 20748 33394 20804 33406
rect 21084 33684 21140 33694
rect 21084 33346 21140 33628
rect 21084 33294 21086 33346
rect 21138 33294 21140 33346
rect 21084 33282 21140 33294
rect 20412 32284 20692 32340
rect 20748 32900 20804 32910
rect 20300 30436 20356 30446
rect 20300 30210 20356 30380
rect 20300 30158 20302 30210
rect 20354 30158 20356 30210
rect 20300 30146 20356 30158
rect 20300 28868 20356 28878
rect 20300 27412 20356 28812
rect 20300 27346 20356 27356
rect 20300 26292 20356 26302
rect 20300 25396 20356 26236
rect 20300 25302 20356 25340
rect 20076 24332 20244 24388
rect 19740 22206 19742 22258
rect 19794 22206 19796 22258
rect 19516 20916 19572 20926
rect 19516 20822 19572 20860
rect 19740 19124 19796 22206
rect 19852 24050 19908 24062
rect 19852 23998 19854 24050
rect 19906 23998 19908 24050
rect 19852 21812 19908 23998
rect 20076 23492 20132 24332
rect 20412 24276 20468 32284
rect 20524 31668 20580 31678
rect 20524 28308 20580 31612
rect 20636 30772 20692 30782
rect 20636 29652 20692 30716
rect 20748 30434 20804 32844
rect 21084 32676 21140 32686
rect 21084 32582 21140 32620
rect 20972 32564 21028 32574
rect 20972 32470 21028 32508
rect 21196 32562 21252 34300
rect 21196 32510 21198 32562
rect 21250 32510 21252 32562
rect 21196 32498 21252 32510
rect 20748 30382 20750 30434
rect 20802 30382 20804 30434
rect 20748 30370 20804 30382
rect 20860 31892 20916 31902
rect 20860 30210 20916 31836
rect 21308 31556 21364 34636
rect 21420 34244 21476 34254
rect 21420 34130 21476 34188
rect 21420 34078 21422 34130
rect 21474 34078 21476 34130
rect 21420 34066 21476 34078
rect 21532 33346 21588 34860
rect 21532 33294 21534 33346
rect 21586 33294 21588 33346
rect 21532 33282 21588 33294
rect 21644 34132 21700 35644
rect 21756 35634 21812 35644
rect 21980 35476 22036 35486
rect 21980 35382 22036 35420
rect 21756 35140 21812 35150
rect 21756 35138 21924 35140
rect 21756 35086 21758 35138
rect 21810 35086 21924 35138
rect 21756 35084 21924 35086
rect 21756 35074 21812 35084
rect 21868 35028 21924 35084
rect 21868 34962 21924 34972
rect 22092 34580 22148 34590
rect 21756 34132 21812 34142
rect 21644 34130 21812 34132
rect 21644 34078 21758 34130
rect 21810 34078 21812 34130
rect 21644 34076 21812 34078
rect 21644 33348 21700 34076
rect 21756 34066 21812 34076
rect 21980 34132 22036 34142
rect 21868 34020 21924 34030
rect 21756 33572 21812 33582
rect 21868 33572 21924 33964
rect 21980 34018 22036 34076
rect 21980 33966 21982 34018
rect 22034 33966 22036 34018
rect 21980 33954 22036 33966
rect 21756 33570 21924 33572
rect 21756 33518 21758 33570
rect 21810 33518 21924 33570
rect 21756 33516 21924 33518
rect 21756 33506 21812 33516
rect 21644 33292 21812 33348
rect 21644 33012 21700 33022
rect 21532 31778 21588 31790
rect 21532 31726 21534 31778
rect 21586 31726 21588 31778
rect 21532 31556 21588 31726
rect 21196 31500 21588 31556
rect 20860 30158 20862 30210
rect 20914 30158 20916 30210
rect 20860 30146 20916 30158
rect 20972 30996 21028 31006
rect 20972 30210 21028 30940
rect 20972 30158 20974 30210
rect 21026 30158 21028 30210
rect 20748 29652 20804 29662
rect 20636 29650 20804 29652
rect 20636 29598 20750 29650
rect 20802 29598 20804 29650
rect 20636 29596 20804 29598
rect 20748 29586 20804 29596
rect 20636 29428 20692 29438
rect 20636 29334 20692 29372
rect 20972 29314 21028 30158
rect 20972 29262 20974 29314
rect 21026 29262 21028 29314
rect 20972 29250 21028 29262
rect 21196 29092 21252 31500
rect 21644 31444 21700 32956
rect 21308 31388 21700 31444
rect 21308 30322 21364 31388
rect 21308 30270 21310 30322
rect 21362 30270 21364 30322
rect 21308 30258 21364 30270
rect 21420 30322 21476 30334
rect 21420 30270 21422 30322
rect 21474 30270 21476 30322
rect 21420 30212 21476 30270
rect 21420 30146 21476 30156
rect 21644 30210 21700 30222
rect 21644 30158 21646 30210
rect 21698 30158 21700 30210
rect 21308 29540 21364 29550
rect 21308 29426 21364 29484
rect 21308 29374 21310 29426
rect 21362 29374 21364 29426
rect 21308 29362 21364 29374
rect 21644 29428 21700 30158
rect 21644 29362 21700 29372
rect 21532 29316 21588 29326
rect 21532 29222 21588 29260
rect 21420 29202 21476 29214
rect 21420 29150 21422 29202
rect 21474 29150 21476 29202
rect 20972 29036 21252 29092
rect 21308 29092 21364 29102
rect 20860 28532 20916 28542
rect 20860 28438 20916 28476
rect 20524 28252 20916 28308
rect 20636 28084 20692 28094
rect 20636 27858 20692 28028
rect 20860 27970 20916 28252
rect 20860 27918 20862 27970
rect 20914 27918 20916 27970
rect 20860 27906 20916 27918
rect 20636 27806 20638 27858
rect 20690 27806 20692 27858
rect 20636 27794 20692 27806
rect 20748 27634 20804 27646
rect 20748 27582 20750 27634
rect 20802 27582 20804 27634
rect 20524 27412 20580 27422
rect 20524 24724 20580 27356
rect 20748 26852 20804 27582
rect 20972 26908 21028 29036
rect 21308 28866 21364 29036
rect 21308 28814 21310 28866
rect 21362 28814 21364 28866
rect 21308 28802 21364 28814
rect 21084 27860 21140 27870
rect 21084 27766 21140 27804
rect 21308 27860 21364 27870
rect 21420 27860 21476 29150
rect 21756 29092 21812 33292
rect 21868 32562 21924 32574
rect 21868 32510 21870 32562
rect 21922 32510 21924 32562
rect 21868 32452 21924 32510
rect 21868 32386 21924 32396
rect 22092 32002 22148 34524
rect 22204 32116 22260 38332
rect 22428 38052 22484 40684
rect 22764 40402 22820 40414
rect 22764 40350 22766 40402
rect 22818 40350 22820 40402
rect 22540 38612 22596 38622
rect 22540 38610 22708 38612
rect 22540 38558 22542 38610
rect 22594 38558 22708 38610
rect 22540 38556 22708 38558
rect 22540 38546 22596 38556
rect 22428 37986 22484 37996
rect 22428 37828 22484 37838
rect 22316 37826 22484 37828
rect 22316 37774 22430 37826
rect 22482 37774 22484 37826
rect 22316 37772 22484 37774
rect 22316 34244 22372 37772
rect 22428 37762 22484 37772
rect 22540 37044 22596 37054
rect 22428 37042 22596 37044
rect 22428 36990 22542 37042
rect 22594 36990 22596 37042
rect 22428 36988 22596 36990
rect 22428 35700 22484 36988
rect 22540 36978 22596 36988
rect 22428 34914 22484 35644
rect 22428 34862 22430 34914
rect 22482 34862 22484 34914
rect 22428 34850 22484 34862
rect 22540 36258 22596 36270
rect 22540 36206 22542 36258
rect 22594 36206 22596 36258
rect 22540 35698 22596 36206
rect 22540 35646 22542 35698
rect 22594 35646 22596 35698
rect 22540 34916 22596 35646
rect 22540 34850 22596 34860
rect 22316 33346 22372 34188
rect 22652 34130 22708 38556
rect 22764 37492 22820 40350
rect 22764 37426 22820 37436
rect 22988 35698 23044 40796
rect 22988 35646 22990 35698
rect 23042 35646 23044 35698
rect 22652 34078 22654 34130
rect 22706 34078 22708 34130
rect 22652 33684 22708 34078
rect 22652 33618 22708 33628
rect 22764 34914 22820 34926
rect 22764 34862 22766 34914
rect 22818 34862 22820 34914
rect 22764 33908 22820 34862
rect 22988 34132 23044 35646
rect 22316 33294 22318 33346
rect 22370 33294 22372 33346
rect 22316 33282 22372 33294
rect 22764 33346 22820 33852
rect 22764 33294 22766 33346
rect 22818 33294 22820 33346
rect 22764 33282 22820 33294
rect 22876 34130 23044 34132
rect 22876 34078 22990 34130
rect 23042 34078 23044 34130
rect 22876 34076 23044 34078
rect 22316 32340 22372 32350
rect 22316 32246 22372 32284
rect 22204 32060 22372 32116
rect 22092 31950 22094 32002
rect 22146 31950 22148 32002
rect 22092 31938 22148 31950
rect 21868 30548 21924 30558
rect 21868 29426 21924 30492
rect 21868 29374 21870 29426
rect 21922 29374 21924 29426
rect 21868 29362 21924 29374
rect 22204 29428 22260 29438
rect 22204 29334 22260 29372
rect 21308 27858 21476 27860
rect 21308 27806 21310 27858
rect 21362 27806 21476 27858
rect 21308 27804 21476 27806
rect 21532 29036 21812 29092
rect 22092 29202 22148 29214
rect 22092 29150 22094 29202
rect 22146 29150 22148 29202
rect 21308 27794 21364 27804
rect 21084 27300 21140 27310
rect 21084 27206 21140 27244
rect 21196 26962 21252 26974
rect 21196 26910 21198 26962
rect 21250 26910 21252 26962
rect 20972 26852 21140 26908
rect 20748 26786 20804 26796
rect 20748 26516 20804 26526
rect 20636 26460 20748 26516
rect 20636 24948 20692 26460
rect 20748 26422 20804 26460
rect 20748 26180 20804 26190
rect 20748 25730 20804 26124
rect 20748 25678 20750 25730
rect 20802 25678 20804 25730
rect 20748 25666 20804 25678
rect 20636 24892 20804 24948
rect 20636 24724 20692 24734
rect 20524 24722 20692 24724
rect 20524 24670 20638 24722
rect 20690 24670 20692 24722
rect 20524 24668 20692 24670
rect 20636 24658 20692 24668
rect 20748 24612 20804 24892
rect 20860 24836 20916 24846
rect 20860 24742 20916 24780
rect 20972 24612 21028 24622
rect 20748 24610 21028 24612
rect 20748 24558 20974 24610
rect 21026 24558 21028 24610
rect 20748 24556 21028 24558
rect 20972 24546 21028 24556
rect 20076 23426 20132 23436
rect 20188 24220 20468 24276
rect 19964 22930 20020 22942
rect 19964 22878 19966 22930
rect 20018 22878 20020 22930
rect 19964 22372 20020 22878
rect 20076 22372 20132 22382
rect 19964 22370 20132 22372
rect 19964 22318 20078 22370
rect 20130 22318 20132 22370
rect 19964 22316 20132 22318
rect 20076 22306 20132 22316
rect 19852 21756 20020 21812
rect 19852 21588 19908 21598
rect 19852 21364 19908 21532
rect 19852 21298 19908 21308
rect 19852 21140 19908 21150
rect 19852 19908 19908 21084
rect 19964 20356 20020 21756
rect 20020 20300 20132 20356
rect 19964 20290 20020 20300
rect 19964 19908 20020 19918
rect 19852 19906 20020 19908
rect 19852 19854 19966 19906
rect 20018 19854 20020 19906
rect 19852 19852 20020 19854
rect 19964 19842 20020 19852
rect 19852 19572 19908 19582
rect 19852 19458 19908 19516
rect 19852 19406 19854 19458
rect 19906 19406 19908 19458
rect 19852 19394 19908 19406
rect 19964 19460 20020 19470
rect 19964 19366 20020 19404
rect 20076 19346 20132 20300
rect 20076 19294 20078 19346
rect 20130 19294 20132 19346
rect 20076 19282 20132 19294
rect 19740 19068 19908 19124
rect 19404 18172 19796 18228
rect 19404 17668 19460 17678
rect 19404 17666 19684 17668
rect 19404 17614 19406 17666
rect 19458 17614 19684 17666
rect 19404 17612 19684 17614
rect 19404 17602 19460 17612
rect 19628 17108 19684 17612
rect 19740 17666 19796 18172
rect 19740 17614 19742 17666
rect 19794 17614 19796 17666
rect 19740 17602 19796 17614
rect 19852 17556 19908 19068
rect 20188 17892 20244 24220
rect 20300 24050 20356 24062
rect 20300 23998 20302 24050
rect 20354 23998 20356 24050
rect 20300 23716 20356 23998
rect 21084 24052 21140 26852
rect 21196 25844 21252 26910
rect 21308 26964 21364 27002
rect 21308 26898 21364 26908
rect 21196 25788 21476 25844
rect 21420 24946 21476 25788
rect 21420 24894 21422 24946
rect 21474 24894 21476 24946
rect 21420 24882 21476 24894
rect 21084 23996 21476 24052
rect 20412 23828 20468 23838
rect 20412 23734 20468 23772
rect 21196 23828 21252 23838
rect 21196 23826 21364 23828
rect 21196 23774 21198 23826
rect 21250 23774 21364 23826
rect 21196 23772 21364 23774
rect 21196 23762 21252 23772
rect 20300 23650 20356 23660
rect 20524 23716 20580 23726
rect 20524 23714 20692 23716
rect 20524 23662 20526 23714
rect 20578 23662 20692 23714
rect 20524 23660 20692 23662
rect 20524 23650 20580 23660
rect 20524 23492 20580 23502
rect 20524 22820 20580 23436
rect 20524 22370 20580 22764
rect 20524 22318 20526 22370
rect 20578 22318 20580 22370
rect 20524 22306 20580 22318
rect 20524 22148 20580 22158
rect 20244 17836 20468 17892
rect 20188 17826 20244 17836
rect 19964 17780 20020 17790
rect 19964 17686 20020 17724
rect 19852 17500 20020 17556
rect 19740 17108 19796 17118
rect 19628 17106 19796 17108
rect 19628 17054 19742 17106
rect 19794 17054 19796 17106
rect 19628 17052 19796 17054
rect 19740 17042 19796 17052
rect 19852 16324 19908 16334
rect 19852 16230 19908 16268
rect 19404 15988 19460 15998
rect 19404 15894 19460 15932
rect 19964 15148 20020 17500
rect 20188 17108 20244 17118
rect 19740 15092 19796 15102
rect 19404 15090 19796 15092
rect 19404 15038 19742 15090
rect 19794 15038 19796 15090
rect 19404 15036 19796 15038
rect 19404 12962 19460 15036
rect 19740 15026 19796 15036
rect 19852 15092 20020 15148
rect 20076 16884 20132 16894
rect 19740 14530 19796 14542
rect 19740 14478 19742 14530
rect 19794 14478 19796 14530
rect 19740 14308 19796 14478
rect 19740 13300 19796 14252
rect 19740 13234 19796 13244
rect 19404 12910 19406 12962
rect 19458 12910 19460 12962
rect 19404 12898 19460 12910
rect 19404 11508 19460 11518
rect 19404 7476 19460 11452
rect 19740 11394 19796 11406
rect 19740 11342 19742 11394
rect 19794 11342 19796 11394
rect 19740 10050 19796 11342
rect 19740 9998 19742 10050
rect 19794 9998 19796 10050
rect 19740 9986 19796 9998
rect 19852 9044 19908 15092
rect 19964 12964 20020 12974
rect 19964 12870 20020 12908
rect 20076 9044 20132 16828
rect 20188 12068 20244 17052
rect 20412 15148 20468 17836
rect 20524 17444 20580 22092
rect 20636 21028 20692 23660
rect 20748 22930 20804 22942
rect 20748 22878 20750 22930
rect 20802 22878 20804 22930
rect 20748 22708 20804 22878
rect 20748 22652 21252 22708
rect 20748 22482 20804 22494
rect 20748 22430 20750 22482
rect 20802 22430 20804 22482
rect 20748 21252 20804 22430
rect 21196 22482 21252 22652
rect 21196 22430 21198 22482
rect 21250 22430 21252 22482
rect 21196 22418 21252 22430
rect 21308 22260 21364 23772
rect 20972 22204 21364 22260
rect 20972 21698 21028 22204
rect 21420 22148 21476 23996
rect 20972 21646 20974 21698
rect 21026 21646 21028 21698
rect 20972 21634 21028 21646
rect 21084 22092 21476 22148
rect 20748 21186 20804 21196
rect 20860 21586 20916 21598
rect 20860 21534 20862 21586
rect 20914 21534 20916 21586
rect 20748 21028 20804 21038
rect 20636 21026 20804 21028
rect 20636 20974 20750 21026
rect 20802 20974 20804 21026
rect 20636 20972 20804 20974
rect 20636 20356 20692 20366
rect 20636 20242 20692 20300
rect 20636 20190 20638 20242
rect 20690 20190 20692 20242
rect 20636 20178 20692 20190
rect 20748 20130 20804 20972
rect 20748 20078 20750 20130
rect 20802 20078 20804 20130
rect 20748 20066 20804 20078
rect 20860 20020 20916 21534
rect 20860 19954 20916 19964
rect 21084 17780 21140 22092
rect 21196 21924 21252 21934
rect 21196 20914 21252 21868
rect 21420 21476 21476 21486
rect 21420 21382 21476 21420
rect 21196 20862 21198 20914
rect 21250 20862 21252 20914
rect 21196 20850 21252 20862
rect 21308 21140 21364 21150
rect 21308 20802 21364 21084
rect 21532 21028 21588 29036
rect 22092 28756 22148 29150
rect 21644 28700 22148 28756
rect 21644 27858 21700 28700
rect 22316 28308 22372 32060
rect 22540 29314 22596 29326
rect 22540 29262 22542 29314
rect 22594 29262 22596 29314
rect 22092 28252 22372 28308
rect 22428 28418 22484 28430
rect 22428 28366 22430 28418
rect 22482 28366 22484 28418
rect 21868 28084 21924 28094
rect 21868 27990 21924 28028
rect 21980 27972 22036 27982
rect 21980 27878 22036 27916
rect 21644 27806 21646 27858
rect 21698 27806 21700 27858
rect 21644 27794 21700 27806
rect 21644 26962 21700 26974
rect 21644 26910 21646 26962
rect 21698 26910 21700 26962
rect 21644 26516 21700 26910
rect 21756 26964 21812 27002
rect 22092 26908 22148 28252
rect 22428 27972 22484 28366
rect 22540 28084 22596 29262
rect 22540 28018 22596 28028
rect 22428 27906 22484 27916
rect 21756 26898 21812 26908
rect 21644 26450 21700 26460
rect 21980 26852 22148 26908
rect 22204 26964 22260 26974
rect 22876 26908 22932 34076
rect 22988 34066 23044 34076
rect 23100 40404 23156 40414
rect 21868 26066 21924 26078
rect 21868 26014 21870 26066
rect 21922 26014 21924 26066
rect 21868 25956 21924 26014
rect 21868 25890 21924 25900
rect 21868 25508 21924 25518
rect 21868 25414 21924 25452
rect 21644 24836 21700 24846
rect 21644 24742 21700 24780
rect 21868 24610 21924 24622
rect 21868 24558 21870 24610
rect 21922 24558 21924 24610
rect 21644 24276 21700 24286
rect 21644 24050 21700 24220
rect 21644 23998 21646 24050
rect 21698 23998 21700 24050
rect 21644 23986 21700 23998
rect 21756 23828 21812 23838
rect 21308 20750 21310 20802
rect 21362 20750 21364 20802
rect 21308 20738 21364 20750
rect 21420 20972 21588 21028
rect 21644 23604 21700 23614
rect 21420 19908 21476 20972
rect 21532 20804 21588 20814
rect 21532 20710 21588 20748
rect 21644 20580 21700 23548
rect 21756 20802 21812 23772
rect 21868 23380 21924 24558
rect 21868 23314 21924 23324
rect 21868 23044 21924 23054
rect 21868 22950 21924 22988
rect 21980 22370 22036 26852
rect 22204 25732 22260 26908
rect 22428 26852 22932 26908
rect 22988 32340 23044 32350
rect 22316 26292 22372 26302
rect 22316 26198 22372 26236
rect 22316 25732 22372 25742
rect 22204 25730 22372 25732
rect 22204 25678 22318 25730
rect 22370 25678 22372 25730
rect 22204 25676 22372 25678
rect 22316 25666 22372 25676
rect 22092 25508 22148 25518
rect 22092 24722 22148 25452
rect 22204 25282 22260 25294
rect 22204 25230 22206 25282
rect 22258 25230 22260 25282
rect 22204 24946 22260 25230
rect 22204 24894 22206 24946
rect 22258 24894 22260 24946
rect 22204 24882 22260 24894
rect 22092 24670 22094 24722
rect 22146 24670 22148 24722
rect 22092 24658 22148 24670
rect 22428 23380 22484 26852
rect 22540 25508 22596 25518
rect 22540 25414 22596 25452
rect 22764 25506 22820 25518
rect 22764 25454 22766 25506
rect 22818 25454 22820 25506
rect 22764 25284 22820 25454
rect 22764 25218 22820 25228
rect 22988 24276 23044 32284
rect 21980 22318 21982 22370
rect 22034 22318 22036 22370
rect 21980 22306 22036 22318
rect 22316 23324 22484 23380
rect 22540 24220 23044 24276
rect 21756 20750 21758 20802
rect 21810 20750 21812 20802
rect 21756 20738 21812 20750
rect 22092 22036 22148 22046
rect 21644 20524 21812 20580
rect 20972 17724 21140 17780
rect 21196 19852 21476 19908
rect 20636 17668 20692 17678
rect 20636 17666 20916 17668
rect 20636 17614 20638 17666
rect 20690 17614 20916 17666
rect 20636 17612 20916 17614
rect 20636 17602 20692 17612
rect 20524 17388 20804 17444
rect 20636 16772 20692 16782
rect 20412 15092 20580 15148
rect 20412 14644 20468 14654
rect 20188 12002 20244 12012
rect 20300 13636 20356 13646
rect 19628 8988 19908 9044
rect 19964 8988 20132 9044
rect 20188 9716 20244 9726
rect 20300 9716 20356 13580
rect 20412 13524 20468 14588
rect 20412 13458 20468 13468
rect 20188 9714 20356 9716
rect 20188 9662 20190 9714
rect 20242 9662 20356 9714
rect 20188 9660 20356 9662
rect 20412 12964 20468 12974
rect 20412 11394 20468 12908
rect 20412 11342 20414 11394
rect 20466 11342 20468 11394
rect 19516 8372 19572 8382
rect 19516 8278 19572 8316
rect 19404 7410 19460 7420
rect 19628 6692 19684 8988
rect 19740 8820 19796 8830
rect 19740 8818 19908 8820
rect 19740 8766 19742 8818
rect 19794 8766 19908 8818
rect 19740 8764 19908 8766
rect 19740 8754 19796 8764
rect 19740 8260 19796 8270
rect 19740 6916 19796 8204
rect 19740 6850 19796 6860
rect 19628 6626 19684 6636
rect 19740 6690 19796 6702
rect 19740 6638 19742 6690
rect 19794 6638 19796 6690
rect 19292 6412 19684 6468
rect 18956 6300 19460 6356
rect 18844 5908 18900 5918
rect 18844 5684 18900 5852
rect 19404 5794 19460 6300
rect 19628 5906 19684 6412
rect 19628 5854 19630 5906
rect 19682 5854 19684 5906
rect 19628 5842 19684 5854
rect 19404 5742 19406 5794
rect 19458 5742 19460 5794
rect 19404 5730 19460 5742
rect 18844 5618 18900 5628
rect 19068 5684 19124 5694
rect 18732 5294 18734 5346
rect 18786 5294 18788 5346
rect 18732 5282 18788 5294
rect 18956 4900 19012 4910
rect 18620 4620 18788 4676
rect 18508 3502 18510 3554
rect 18562 3502 18564 3554
rect 18508 3490 18564 3502
rect 18620 4114 18676 4126
rect 18620 4062 18622 4114
rect 18674 4062 18676 4114
rect 18172 2942 18174 2994
rect 18226 2942 18228 2994
rect 18172 2930 18228 2942
rect 18620 2996 18676 4062
rect 18732 3778 18788 4620
rect 18956 4226 19012 4844
rect 18956 4174 18958 4226
rect 19010 4174 19012 4226
rect 18956 4162 19012 4174
rect 18732 3726 18734 3778
rect 18786 3726 18788 3778
rect 18732 3714 18788 3726
rect 18844 4004 18900 4014
rect 18620 2930 18676 2940
rect 18620 2772 18676 2782
rect 18620 2678 18676 2716
rect 18284 2660 18340 2670
rect 18172 2212 18228 2222
rect 18172 2118 18228 2156
rect 18172 1092 18228 1102
rect 18060 1090 18228 1092
rect 18060 1038 18174 1090
rect 18226 1038 18228 1090
rect 18060 1036 18228 1038
rect 16940 980 16996 990
rect 16940 886 16996 924
rect 17276 980 17332 990
rect 17052 532 17108 542
rect 17052 112 17108 476
rect 17276 112 17332 924
rect 17500 112 17556 1036
rect 18172 1026 18228 1036
rect 18284 868 18340 2604
rect 18620 2324 18676 2334
rect 18172 812 18340 868
rect 18396 868 18452 878
rect 17948 644 18004 654
rect 17724 196 17780 206
rect 17724 112 17780 140
rect 17948 112 18004 588
rect 18172 112 18228 812
rect 18396 112 18452 812
rect 18620 112 18676 2268
rect 18844 112 18900 3948
rect 18956 2660 19012 2670
rect 19068 2660 19124 5628
rect 19404 5572 19460 5582
rect 19404 5234 19460 5516
rect 19740 5460 19796 6638
rect 19740 5394 19796 5404
rect 19404 5182 19406 5234
rect 19458 5182 19460 5234
rect 19404 5170 19460 5182
rect 19852 5236 19908 8764
rect 19964 8260 20020 8988
rect 20076 8820 20132 8830
rect 20076 8726 20132 8764
rect 19964 8194 20020 8204
rect 20076 7812 20132 7822
rect 19964 7588 20020 7598
rect 20076 7588 20132 7756
rect 19964 7586 20132 7588
rect 19964 7534 19966 7586
rect 20018 7534 20132 7586
rect 19964 7532 20132 7534
rect 19964 7522 20020 7532
rect 20076 7140 20132 7150
rect 19964 6916 20020 6926
rect 19964 5908 20020 6860
rect 20076 6802 20132 7084
rect 20076 6750 20078 6802
rect 20130 6750 20132 6802
rect 20076 6738 20132 6750
rect 20188 6580 20244 9660
rect 20412 7588 20468 11342
rect 20524 10612 20580 15092
rect 20524 7588 20580 10556
rect 20636 10388 20692 16716
rect 20748 14418 20804 17388
rect 20860 16324 20916 17612
rect 20972 16548 21028 17724
rect 21196 17668 21252 19852
rect 20972 16482 21028 16492
rect 21084 17666 21252 17668
rect 21084 17614 21198 17666
rect 21250 17614 21252 17666
rect 21084 17612 21252 17614
rect 20972 16324 21028 16334
rect 20860 16322 21028 16324
rect 20860 16270 20974 16322
rect 21026 16270 21028 16322
rect 20860 16268 21028 16270
rect 20972 16258 21028 16268
rect 21084 15148 21140 17612
rect 21196 17602 21252 17612
rect 21644 17108 21700 17118
rect 21196 16548 21252 16558
rect 21196 16100 21252 16492
rect 21196 15426 21252 16044
rect 21196 15374 21198 15426
rect 21250 15374 21252 15426
rect 21196 15362 21252 15374
rect 21532 15874 21588 15886
rect 21532 15822 21534 15874
rect 21586 15822 21588 15874
rect 21084 15092 21252 15148
rect 21084 14532 21140 14542
rect 20748 14366 20750 14418
rect 20802 14366 20804 14418
rect 20748 13636 20804 14366
rect 20748 13542 20804 13580
rect 20860 14530 21140 14532
rect 20860 14478 21086 14530
rect 21138 14478 21140 14530
rect 20860 14476 21140 14478
rect 20748 13300 20804 13310
rect 20748 12962 20804 13244
rect 20748 12910 20750 12962
rect 20802 12910 20804 12962
rect 20748 12898 20804 12910
rect 20748 12404 20804 12414
rect 20860 12404 20916 14476
rect 21084 14466 21140 14476
rect 21196 14532 21252 15092
rect 21532 14756 21588 15822
rect 21644 15202 21700 17052
rect 21644 15150 21646 15202
rect 21698 15150 21700 15202
rect 21644 15138 21700 15150
rect 21756 14868 21812 20524
rect 21980 20578 22036 20590
rect 21980 20526 21982 20578
rect 22034 20526 22036 20578
rect 21980 19460 22036 20526
rect 21980 19394 22036 19404
rect 21980 17668 22036 17678
rect 21532 14690 21588 14700
rect 21644 14812 21812 14868
rect 21868 17666 22036 17668
rect 21868 17614 21982 17666
rect 22034 17614 22036 17666
rect 21868 17612 22036 17614
rect 21196 14466 21252 14476
rect 21532 14530 21588 14542
rect 21532 14478 21534 14530
rect 21586 14478 21588 14530
rect 21532 14420 21588 14478
rect 21196 13748 21252 13758
rect 21196 13746 21476 13748
rect 21196 13694 21198 13746
rect 21250 13694 21476 13746
rect 21196 13692 21476 13694
rect 21196 13682 21252 13692
rect 21308 13524 21364 13534
rect 20748 12402 20916 12404
rect 20748 12350 20750 12402
rect 20802 12350 20916 12402
rect 20748 12348 20916 12350
rect 21196 13300 21252 13310
rect 20748 12338 20804 12348
rect 21196 11394 21252 13244
rect 21196 11342 21198 11394
rect 21250 11342 21252 11394
rect 21196 11284 21252 11342
rect 21196 11218 21252 11228
rect 21196 10612 21252 10622
rect 20748 10500 20804 10510
rect 20748 10406 20804 10444
rect 20636 10322 20692 10332
rect 21196 10050 21252 10556
rect 21196 9998 21198 10050
rect 21250 9998 21252 10050
rect 21196 9986 21252 9998
rect 21308 9940 21364 13468
rect 21420 13186 21476 13692
rect 21420 13134 21422 13186
rect 21474 13134 21476 13186
rect 21420 13122 21476 13134
rect 21532 13746 21588 14364
rect 21532 13694 21534 13746
rect 21586 13694 21588 13746
rect 21308 9884 21476 9940
rect 20636 9826 20692 9838
rect 20636 9774 20638 9826
rect 20690 9774 20692 9826
rect 20636 8484 20692 9774
rect 21084 9814 21140 9826
rect 21084 9762 21086 9814
rect 21138 9762 21140 9814
rect 21084 9716 21140 9762
rect 21084 9650 21140 9660
rect 21308 9716 21364 9726
rect 20860 9044 20916 9054
rect 20860 8950 20916 8988
rect 21196 8930 21252 8942
rect 21196 8878 21198 8930
rect 21250 8878 21252 8930
rect 21196 8596 21252 8878
rect 21196 8530 21252 8540
rect 20748 8484 20804 8494
rect 20636 8482 20804 8484
rect 20636 8430 20750 8482
rect 20802 8430 20804 8482
rect 20636 8428 20804 8430
rect 20748 8418 20804 8428
rect 21084 8148 21140 8158
rect 20748 7812 20804 7822
rect 20636 7588 20692 7598
rect 20524 7586 20692 7588
rect 20524 7534 20638 7586
rect 20690 7534 20692 7586
rect 20524 7532 20692 7534
rect 20188 6514 20244 6524
rect 20300 7028 20356 7038
rect 20412 7028 20468 7532
rect 20356 6972 20468 7028
rect 20524 7364 20580 7374
rect 19964 5842 20020 5852
rect 19852 5180 20132 5236
rect 19740 5124 19796 5134
rect 19516 5122 19796 5124
rect 19516 5070 19742 5122
rect 19794 5070 19796 5122
rect 19516 5068 19796 5070
rect 19292 4340 19348 4350
rect 19292 4246 19348 4284
rect 18956 2658 19124 2660
rect 18956 2606 18958 2658
rect 19010 2606 19124 2658
rect 18956 2604 19124 2606
rect 19180 3554 19236 3566
rect 19180 3502 19182 3554
rect 19234 3502 19236 3554
rect 18956 2594 19012 2604
rect 19180 2212 19236 3502
rect 19404 3444 19460 3454
rect 19292 2548 19348 2558
rect 19292 2454 19348 2492
rect 19292 2212 19348 2222
rect 19180 2210 19348 2212
rect 19180 2158 19294 2210
rect 19346 2158 19348 2210
rect 19180 2156 19348 2158
rect 19292 2146 19348 2156
rect 19404 1988 19460 3388
rect 19068 1932 19460 1988
rect 19068 112 19124 1932
rect 19516 1876 19572 5068
rect 19740 5058 19796 5068
rect 19852 5012 19908 5022
rect 19628 4452 19684 4462
rect 19628 4338 19684 4396
rect 19628 4286 19630 4338
rect 19682 4286 19684 4338
rect 19628 4274 19684 4286
rect 19852 3388 19908 4956
rect 19964 4900 20020 4910
rect 19964 4226 20020 4844
rect 20076 4676 20132 5180
rect 20300 5124 20356 6972
rect 20524 6804 20580 7308
rect 20636 7140 20692 7532
rect 20636 7074 20692 7084
rect 20412 6580 20468 6590
rect 20412 5572 20468 6524
rect 20412 5506 20468 5516
rect 20076 4610 20132 4620
rect 20188 5122 20356 5124
rect 20188 5070 20302 5122
rect 20354 5070 20356 5122
rect 20188 5068 20356 5070
rect 20188 4452 20244 5068
rect 20300 5058 20356 5068
rect 20412 5234 20468 5246
rect 20412 5182 20414 5234
rect 20466 5182 20468 5234
rect 19964 4174 19966 4226
rect 20018 4174 20020 4226
rect 19964 4162 20020 4174
rect 20076 4396 20244 4452
rect 20300 4676 20356 4686
rect 19964 3556 20020 3566
rect 20076 3556 20132 4396
rect 19964 3554 20132 3556
rect 19964 3502 19966 3554
rect 20018 3502 20132 3554
rect 19964 3500 20132 3502
rect 19964 3490 20020 3500
rect 19740 3332 19908 3388
rect 19628 2996 19684 3006
rect 19628 2770 19684 2940
rect 19628 2718 19630 2770
rect 19682 2718 19684 2770
rect 19628 2706 19684 2718
rect 19516 1820 19684 1876
rect 19404 1428 19460 1438
rect 19628 1428 19684 1820
rect 19404 1426 19684 1428
rect 19404 1374 19406 1426
rect 19458 1374 19684 1426
rect 19404 1372 19684 1374
rect 19404 1362 19460 1372
rect 19292 1316 19348 1326
rect 19740 1316 19796 3332
rect 19852 2548 19908 2558
rect 19852 1986 19908 2492
rect 19852 1934 19854 1986
rect 19906 1934 19908 1986
rect 19852 1764 19908 1934
rect 20188 2436 20244 2446
rect 19852 1698 19908 1708
rect 19964 1876 20020 1886
rect 19292 112 19348 1260
rect 19516 1260 19796 1316
rect 19964 1316 20020 1820
rect 20188 1426 20244 2380
rect 20188 1374 20190 1426
rect 20242 1374 20244 1426
rect 20188 1362 20244 1374
rect 19516 112 19572 1260
rect 19964 1250 20020 1260
rect 20300 756 20356 4620
rect 20412 4340 20468 5182
rect 20412 4274 20468 4284
rect 20524 4116 20580 6748
rect 20748 6690 20804 7756
rect 20972 7476 21028 7486
rect 20748 6638 20750 6690
rect 20802 6638 20804 6690
rect 20748 6626 20804 6638
rect 20860 7474 21028 7476
rect 20860 7422 20974 7474
rect 21026 7422 21028 7474
rect 20860 7420 21028 7422
rect 20748 6132 20804 6142
rect 20860 6132 20916 7420
rect 20972 7410 21028 7420
rect 21084 7252 21140 8092
rect 20748 6130 20916 6132
rect 20748 6078 20750 6130
rect 20802 6078 20916 6130
rect 20748 6076 20916 6078
rect 20972 7196 21140 7252
rect 20748 6066 20804 6076
rect 20412 4060 20580 4116
rect 20748 5572 20804 5582
rect 20412 2210 20468 4060
rect 20412 2158 20414 2210
rect 20466 2158 20468 2210
rect 20412 2146 20468 2158
rect 20524 3668 20580 3678
rect 20524 1764 20580 3612
rect 20748 3554 20804 5516
rect 20748 3502 20750 3554
rect 20802 3502 20804 3554
rect 20748 3490 20804 3502
rect 20860 5460 20916 5470
rect 20860 4338 20916 5404
rect 20860 4286 20862 4338
rect 20914 4286 20916 4338
rect 20748 3220 20804 3230
rect 20748 2994 20804 3164
rect 20860 3108 20916 4286
rect 20860 3042 20916 3052
rect 20748 2942 20750 2994
rect 20802 2942 20804 2994
rect 20748 2930 20804 2942
rect 20972 2772 21028 7196
rect 21308 6690 21364 9660
rect 21420 8372 21476 9884
rect 21532 9716 21588 13694
rect 21644 13412 21700 14812
rect 21756 14642 21812 14654
rect 21756 14590 21758 14642
rect 21810 14590 21812 14642
rect 21756 14532 21812 14590
rect 21756 14466 21812 14476
rect 21756 13636 21812 13646
rect 21756 13542 21812 13580
rect 21644 13356 21812 13412
rect 21532 9650 21588 9660
rect 21644 10052 21700 10062
rect 21644 9044 21700 9996
rect 21644 8978 21700 8988
rect 21644 8820 21700 8830
rect 21420 8316 21588 8372
rect 21420 8148 21476 8158
rect 21420 8054 21476 8092
rect 21420 7588 21476 7598
rect 21420 7474 21476 7532
rect 21420 7422 21422 7474
rect 21474 7422 21476 7474
rect 21420 7410 21476 7422
rect 21308 6638 21310 6690
rect 21362 6638 21364 6690
rect 21308 6626 21364 6638
rect 21420 6802 21476 6814
rect 21420 6750 21422 6802
rect 21474 6750 21476 6802
rect 21420 6692 21476 6750
rect 21420 6626 21476 6636
rect 21084 5124 21140 5134
rect 21084 5122 21364 5124
rect 21084 5070 21086 5122
rect 21138 5070 21364 5122
rect 21084 5068 21364 5070
rect 21084 5058 21140 5068
rect 21308 4340 21364 5068
rect 21532 5122 21588 8316
rect 21644 7362 21700 8764
rect 21756 8596 21812 13356
rect 21868 12964 21924 17612
rect 21980 17602 22036 17612
rect 22092 15148 22148 21980
rect 22316 21028 22372 23324
rect 22428 23156 22484 23166
rect 22428 21252 22484 23100
rect 22540 22372 22596 24220
rect 23100 24052 23156 40348
rect 23436 38668 23492 57820
rect 24464 57260 24728 57270
rect 24520 57204 24568 57260
rect 24624 57204 24672 57260
rect 24464 57194 24728 57204
rect 23804 56476 24068 56486
rect 23860 56420 23908 56476
rect 23964 56420 24012 56476
rect 23804 56410 24068 56420
rect 24464 55692 24728 55702
rect 24520 55636 24568 55692
rect 24624 55636 24672 55692
rect 24464 55626 24728 55636
rect 23660 55188 23716 55198
rect 23548 48020 23604 48030
rect 23548 46562 23604 47964
rect 23548 46510 23550 46562
rect 23602 46510 23604 46562
rect 23548 46498 23604 46510
rect 23660 44548 23716 55132
rect 24780 55188 24836 55198
rect 24780 55094 24836 55132
rect 23804 54908 24068 54918
rect 23860 54852 23908 54908
rect 23964 54852 24012 54908
rect 23804 54842 24068 54852
rect 24464 54124 24728 54134
rect 24520 54068 24568 54124
rect 24624 54068 24672 54124
rect 24464 54058 24728 54068
rect 23804 53340 24068 53350
rect 23860 53284 23908 53340
rect 23964 53284 24012 53340
rect 23804 53274 24068 53284
rect 24464 52556 24728 52566
rect 24520 52500 24568 52556
rect 24624 52500 24672 52556
rect 24464 52490 24728 52500
rect 23804 51772 24068 51782
rect 23860 51716 23908 51772
rect 23964 51716 24012 51772
rect 23804 51706 24068 51716
rect 24464 50988 24728 50998
rect 24520 50932 24568 50988
rect 24624 50932 24672 50988
rect 24464 50922 24728 50932
rect 23804 50204 24068 50214
rect 23860 50148 23908 50204
rect 23964 50148 24012 50204
rect 23804 50138 24068 50148
rect 24464 49420 24728 49430
rect 24520 49364 24568 49420
rect 24624 49364 24672 49420
rect 24464 49354 24728 49364
rect 23804 48636 24068 48646
rect 23860 48580 23908 48636
rect 23964 48580 24012 48636
rect 23804 48570 24068 48580
rect 24464 47852 24728 47862
rect 24520 47796 24568 47852
rect 24624 47796 24672 47852
rect 24464 47786 24728 47796
rect 23804 47068 24068 47078
rect 23860 47012 23908 47068
rect 23964 47012 24012 47068
rect 23804 47002 24068 47012
rect 24464 46284 24728 46294
rect 24520 46228 24568 46284
rect 24624 46228 24672 46284
rect 24464 46218 24728 46228
rect 23804 45500 24068 45510
rect 23860 45444 23908 45500
rect 23964 45444 24012 45500
rect 23804 45434 24068 45444
rect 24892 45332 24948 88732
rect 25004 79604 25060 79614
rect 25004 62356 25060 79548
rect 25004 62290 25060 62300
rect 25116 63924 25172 63934
rect 25116 57540 25172 63868
rect 25116 57474 25172 57484
rect 24892 45266 24948 45276
rect 25004 53060 25060 53070
rect 24464 44716 24728 44726
rect 24520 44660 24568 44716
rect 24624 44660 24672 44716
rect 24464 44650 24728 44660
rect 23324 38612 23492 38668
rect 23548 44492 23716 44548
rect 23548 38668 23604 44492
rect 23804 43932 24068 43942
rect 23860 43876 23908 43932
rect 23964 43876 24012 43932
rect 23804 43866 24068 43876
rect 23660 43538 23716 43550
rect 23660 43486 23662 43538
rect 23714 43486 23716 43538
rect 23660 42196 23716 43486
rect 24464 43148 24728 43158
rect 24520 43092 24568 43148
rect 24624 43092 24672 43148
rect 24464 43082 24728 43092
rect 23804 42364 24068 42374
rect 23860 42308 23908 42364
rect 23964 42308 24012 42364
rect 23804 42298 24068 42308
rect 23660 42140 23828 42196
rect 23660 41970 23716 41982
rect 23660 41918 23662 41970
rect 23714 41918 23716 41970
rect 23660 41636 23716 41918
rect 23660 41570 23716 41580
rect 23772 41188 23828 42140
rect 24464 41580 24728 41590
rect 24520 41524 24568 41580
rect 24624 41524 24672 41580
rect 24464 41514 24728 41524
rect 23772 40964 23828 41132
rect 23660 40908 23828 40964
rect 23660 40404 23716 40908
rect 23804 40796 24068 40806
rect 23860 40740 23908 40796
rect 23964 40740 24012 40796
rect 23804 40730 24068 40740
rect 23660 40310 23716 40348
rect 24464 40012 24728 40022
rect 24520 39956 24568 40012
rect 24624 39956 24672 40012
rect 24464 39946 24728 39956
rect 23804 39228 24068 39238
rect 23860 39172 23908 39228
rect 23964 39172 24012 39228
rect 23804 39162 24068 39172
rect 23548 38612 23716 38668
rect 23212 31892 23268 31902
rect 23212 31798 23268 31836
rect 22876 23996 23156 24052
rect 23212 29092 23268 29102
rect 22764 23714 22820 23726
rect 22764 23662 22766 23714
rect 22818 23662 22820 23714
rect 22764 22708 22820 23662
rect 22764 22642 22820 22652
rect 22540 22306 22596 22316
rect 22764 22372 22820 22382
rect 22876 22372 22932 23996
rect 23212 23878 23268 29036
rect 23324 26908 23380 38612
rect 23660 36706 23716 38612
rect 24464 38444 24728 38454
rect 24520 38388 24568 38444
rect 24624 38388 24672 38444
rect 24464 38378 24728 38388
rect 24332 38276 24388 38286
rect 23804 37660 24068 37670
rect 23860 37604 23908 37660
rect 23964 37604 24012 37660
rect 23804 37594 24068 37604
rect 23660 36654 23662 36706
rect 23714 36654 23716 36706
rect 23660 36642 23716 36654
rect 23996 36596 24052 36606
rect 23996 36502 24052 36540
rect 23804 36092 24068 36102
rect 23860 36036 23908 36092
rect 23964 36036 24012 36092
rect 23804 36026 24068 36036
rect 24108 35700 24164 35710
rect 24108 35698 24276 35700
rect 24108 35646 24110 35698
rect 24162 35646 24276 35698
rect 24108 35644 24276 35646
rect 24108 35634 24164 35644
rect 23436 34916 23492 34926
rect 23772 34916 23828 34926
rect 23436 32786 23492 34860
rect 23660 34914 23828 34916
rect 23660 34862 23774 34914
rect 23826 34862 23828 34914
rect 23660 34860 23828 34862
rect 23660 33460 23716 34860
rect 23772 34850 23828 34860
rect 23804 34524 24068 34534
rect 23860 34468 23908 34524
rect 23964 34468 24012 34524
rect 23804 34458 24068 34468
rect 23996 34132 24052 34142
rect 24220 34132 24276 35644
rect 23996 34130 24276 34132
rect 23996 34078 23998 34130
rect 24050 34078 24276 34130
rect 23996 34076 24276 34078
rect 23772 33460 23828 33470
rect 23660 33404 23772 33460
rect 23772 33346 23828 33404
rect 23772 33294 23774 33346
rect 23826 33294 23828 33346
rect 23772 33282 23828 33294
rect 23996 33124 24052 34076
rect 23436 32734 23438 32786
rect 23490 32734 23492 32786
rect 23436 32722 23492 32734
rect 23660 33068 24052 33124
rect 23660 32788 23716 33068
rect 23804 32956 24068 32966
rect 23860 32900 23908 32956
rect 23964 32900 24012 32956
rect 23804 32890 24068 32900
rect 23660 26908 23716 32732
rect 23804 31388 24068 31398
rect 23860 31332 23908 31388
rect 23964 31332 24012 31388
rect 23804 31322 24068 31332
rect 23804 29820 24068 29830
rect 23860 29764 23908 29820
rect 23964 29764 24012 29820
rect 23804 29754 24068 29764
rect 23804 28252 24068 28262
rect 23860 28196 23908 28252
rect 23964 28196 24012 28252
rect 23804 28186 24068 28196
rect 23324 26852 23492 26908
rect 22988 23822 23268 23878
rect 23324 23826 23380 23838
rect 22988 23044 23044 23822
rect 23324 23774 23326 23826
rect 23378 23774 23380 23826
rect 23212 23714 23268 23726
rect 23212 23662 23214 23714
rect 23266 23662 23268 23714
rect 23212 23604 23268 23662
rect 23212 23538 23268 23548
rect 23324 23380 23380 23774
rect 23100 23324 23380 23380
rect 23436 23380 23492 26852
rect 23548 26852 23716 26908
rect 23548 23938 23604 26852
rect 23804 26684 24068 26694
rect 23860 26628 23908 26684
rect 23964 26628 24012 26684
rect 23804 26618 24068 26628
rect 23804 25116 24068 25126
rect 23860 25060 23908 25116
rect 23964 25060 24012 25116
rect 23804 25050 24068 25060
rect 23548 23886 23550 23938
rect 23602 23886 23604 23938
rect 23548 23874 23604 23886
rect 23804 23548 24068 23558
rect 23860 23492 23908 23548
rect 23964 23492 24012 23548
rect 23804 23482 24068 23492
rect 23436 23324 23604 23380
rect 23100 23154 23156 23324
rect 23100 23102 23102 23154
rect 23154 23102 23156 23154
rect 23100 23090 23156 23102
rect 23212 23156 23268 23194
rect 23212 23090 23268 23100
rect 23324 23154 23380 23166
rect 23324 23102 23326 23154
rect 23378 23102 23380 23154
rect 22988 22978 23044 22988
rect 22764 22370 22932 22372
rect 22764 22318 22766 22370
rect 22818 22318 22932 22370
rect 22764 22316 22932 22318
rect 23100 22932 23156 22942
rect 22540 21812 22596 21822
rect 22540 21718 22596 21756
rect 22764 21588 22820 22316
rect 23100 21810 23156 22876
rect 23212 22930 23268 22942
rect 23212 22878 23214 22930
rect 23266 22878 23268 22930
rect 23212 22820 23268 22878
rect 23212 22754 23268 22764
rect 23100 21758 23102 21810
rect 23154 21758 23156 21810
rect 23100 21746 23156 21758
rect 23324 22370 23380 23102
rect 23436 23156 23492 23166
rect 23436 22594 23492 23100
rect 23548 22932 23604 23324
rect 23660 23156 23716 23166
rect 23884 23156 23940 23166
rect 23660 23154 23940 23156
rect 23660 23102 23662 23154
rect 23714 23102 23886 23154
rect 23938 23102 23940 23154
rect 23660 23100 23940 23102
rect 23660 23090 23716 23100
rect 23884 23090 23940 23100
rect 24220 23042 24276 23054
rect 24220 22990 24222 23042
rect 24274 22990 24276 23042
rect 24108 22932 24164 22942
rect 23548 22876 23716 22932
rect 23436 22542 23438 22594
rect 23490 22542 23492 22594
rect 23436 22530 23492 22542
rect 23548 22708 23604 22718
rect 23548 22372 23604 22652
rect 23324 22318 23326 22370
rect 23378 22318 23380 22370
rect 23324 21812 23380 22318
rect 23324 21746 23380 21756
rect 23436 22370 23604 22372
rect 23436 22318 23550 22370
rect 23602 22318 23604 22370
rect 23436 22316 23604 22318
rect 22764 21522 22820 21532
rect 22988 21588 23044 21598
rect 23436 21588 23492 22316
rect 23548 22306 23604 22316
rect 22988 21586 23492 21588
rect 22988 21534 22990 21586
rect 23042 21534 23492 21586
rect 22988 21532 23492 21534
rect 22988 21522 23044 21532
rect 23660 21476 23716 22876
rect 24108 22838 24164 22876
rect 23772 22260 23828 22270
rect 23772 22166 23828 22204
rect 24220 22148 24276 22990
rect 24220 22082 24276 22092
rect 23804 21980 24068 21990
rect 23860 21924 23908 21980
rect 23964 21924 24012 21980
rect 23804 21914 24068 21924
rect 23436 21420 23716 21476
rect 22428 21196 22932 21252
rect 21868 12898 21924 12908
rect 21980 15092 22148 15148
rect 22204 20972 22372 21028
rect 21868 11954 21924 11966
rect 21868 11902 21870 11954
rect 21922 11902 21924 11954
rect 21868 11844 21924 11902
rect 21868 10498 21924 11788
rect 21868 10446 21870 10498
rect 21922 10446 21924 10498
rect 21868 10434 21924 10446
rect 21868 9826 21924 9838
rect 21868 9774 21870 9826
rect 21922 9774 21924 9826
rect 21868 9268 21924 9774
rect 21980 9380 22036 15092
rect 22204 14980 22260 20972
rect 22652 16212 22708 16222
rect 22092 14924 22260 14980
rect 22316 16210 22708 16212
rect 22316 16158 22654 16210
rect 22706 16158 22708 16210
rect 22316 16156 22708 16158
rect 22092 13636 22148 14924
rect 22204 14756 22260 14766
rect 22204 13746 22260 14700
rect 22316 13972 22372 16156
rect 22652 16146 22708 16156
rect 22764 15092 22820 15102
rect 22652 15090 22820 15092
rect 22652 15038 22766 15090
rect 22818 15038 22820 15090
rect 22652 15036 22820 15038
rect 22428 14532 22484 14542
rect 22652 14532 22708 15036
rect 22764 15026 22820 15036
rect 22428 14530 22708 14532
rect 22428 14478 22430 14530
rect 22482 14478 22708 14530
rect 22428 14476 22708 14478
rect 22764 14530 22820 14542
rect 22764 14478 22766 14530
rect 22818 14478 22820 14530
rect 22428 14466 22484 14476
rect 22316 13906 22372 13916
rect 22204 13694 22206 13746
rect 22258 13694 22260 13746
rect 22204 13682 22260 13694
rect 22764 13746 22820 14478
rect 22764 13694 22766 13746
rect 22818 13694 22820 13746
rect 22092 13570 22148 13580
rect 22540 13076 22596 13086
rect 22540 12982 22596 13020
rect 22428 12180 22484 12190
rect 22316 10610 22372 10622
rect 22316 10558 22318 10610
rect 22370 10558 22372 10610
rect 22204 9828 22260 9838
rect 21980 9314 22036 9324
rect 22092 9826 22260 9828
rect 22092 9774 22206 9826
rect 22258 9774 22260 9826
rect 22092 9772 22260 9774
rect 21868 9202 21924 9212
rect 21756 8530 21812 8540
rect 21868 9044 21924 9054
rect 21644 7310 21646 7362
rect 21698 7310 21700 7362
rect 21644 7298 21700 7310
rect 21756 8370 21812 8382
rect 21756 8318 21758 8370
rect 21810 8318 21812 8370
rect 21756 8036 21812 8318
rect 21756 6132 21812 7980
rect 21868 6132 21924 8988
rect 22092 7252 22148 9772
rect 22204 9762 22260 9772
rect 22316 9156 22372 10558
rect 22428 10052 22484 12124
rect 22428 9986 22484 9996
rect 22428 9828 22484 9838
rect 22764 9828 22820 13694
rect 22428 9826 22820 9828
rect 22428 9774 22430 9826
rect 22482 9774 22820 9826
rect 22428 9772 22820 9774
rect 22428 9762 22484 9772
rect 22876 9492 22932 21196
rect 23212 19908 23268 19918
rect 23100 16100 23156 16110
rect 22988 12852 23044 12862
rect 23100 12852 23156 16044
rect 22988 12850 23156 12852
rect 22988 12798 22990 12850
rect 23042 12798 23156 12850
rect 22988 12796 23156 12798
rect 22988 12180 23044 12796
rect 22988 12114 23044 12124
rect 22876 9436 23156 9492
rect 22764 9380 22820 9390
rect 22428 9268 22484 9278
rect 22428 9174 22484 9212
rect 22316 9090 22372 9100
rect 22316 7476 22372 7486
rect 22316 7474 22596 7476
rect 22316 7422 22318 7474
rect 22370 7422 22596 7474
rect 22316 7420 22596 7422
rect 22316 7410 22372 7420
rect 22092 7196 22372 7252
rect 22092 6692 22148 6702
rect 22316 6692 22372 7196
rect 22428 6692 22484 6702
rect 22316 6690 22484 6692
rect 22316 6638 22430 6690
rect 22482 6638 22484 6690
rect 22316 6636 22484 6638
rect 22092 6598 22148 6636
rect 22204 6468 22260 6478
rect 21868 6076 22036 6132
rect 21756 6066 21812 6076
rect 21532 5070 21534 5122
rect 21586 5070 21588 5122
rect 21532 4564 21588 5070
rect 21532 4498 21588 4508
rect 21868 5908 21924 5918
rect 21868 5794 21924 5852
rect 21868 5742 21870 5794
rect 21922 5742 21924 5794
rect 21308 4284 21588 4340
rect 21196 4226 21252 4238
rect 21196 4174 21198 4226
rect 21250 4174 21252 4226
rect 21196 4116 21252 4174
rect 21196 3892 21252 4060
rect 21196 3826 21252 3836
rect 21420 4116 21476 4126
rect 21420 3778 21476 4060
rect 21420 3726 21422 3778
rect 21474 3726 21476 3778
rect 21420 3714 21476 3726
rect 20972 2706 21028 2716
rect 21084 3556 21140 3566
rect 20188 700 20356 756
rect 20412 1708 20580 1764
rect 20860 1988 20916 1998
rect 19740 420 19796 430
rect 19740 112 19796 364
rect 19964 308 20020 318
rect 19964 112 20020 252
rect 20188 112 20244 700
rect 20412 112 20468 1708
rect 20636 308 20692 318
rect 20636 112 20692 252
rect 20860 112 20916 1932
rect 20972 1764 21028 1774
rect 20972 532 21028 1708
rect 21084 644 21140 3500
rect 21420 2884 21476 2894
rect 21420 2548 21476 2828
rect 21420 1090 21476 2492
rect 21532 2210 21588 4284
rect 21868 4228 21924 5742
rect 21868 4162 21924 4172
rect 21532 2158 21534 2210
rect 21586 2158 21588 2210
rect 21532 2146 21588 2158
rect 21756 2772 21812 2782
rect 21420 1038 21422 1090
rect 21474 1038 21476 1090
rect 21420 1026 21476 1038
rect 21532 1540 21588 1550
rect 21084 588 21364 644
rect 20972 476 21140 532
rect 21084 112 21140 476
rect 21308 112 21364 588
rect 21532 112 21588 1484
rect 21756 1204 21812 2716
rect 21868 2546 21924 2558
rect 21868 2494 21870 2546
rect 21922 2494 21924 2546
rect 21868 2212 21924 2494
rect 21868 2146 21924 2156
rect 21756 112 21812 1148
rect 21980 112 22036 6076
rect 22092 2212 22148 2222
rect 22092 2118 22148 2156
rect 22204 112 22260 6412
rect 22316 5908 22372 5918
rect 22316 5460 22372 5852
rect 22316 5394 22372 5404
rect 22428 5348 22484 6636
rect 22428 5282 22484 5292
rect 22428 5124 22484 5134
rect 22428 5030 22484 5068
rect 22428 4564 22484 4574
rect 22540 4564 22596 7420
rect 22764 4676 22820 9324
rect 22988 8820 23044 8830
rect 22876 8818 23044 8820
rect 22876 8766 22990 8818
rect 23042 8766 23044 8818
rect 22876 8764 23044 8766
rect 22876 7924 22932 8764
rect 22988 8754 23044 8764
rect 22876 7858 22932 7868
rect 22988 8034 23044 8046
rect 22988 7982 22990 8034
rect 23042 7982 23044 8034
rect 22876 7474 22932 7486
rect 22876 7422 22878 7474
rect 22930 7422 22932 7474
rect 22876 7028 22932 7422
rect 22876 6580 22932 6972
rect 22988 6692 23044 7982
rect 22988 6626 23044 6636
rect 22876 6514 22932 6524
rect 22988 6244 23044 6254
rect 22988 6130 23044 6188
rect 22988 6078 22990 6130
rect 23042 6078 23044 6130
rect 22988 6066 23044 6078
rect 22988 5234 23044 5246
rect 22988 5182 22990 5234
rect 23042 5182 23044 5234
rect 22988 5012 23044 5182
rect 22988 4946 23044 4956
rect 22764 4610 22820 4620
rect 22988 4788 23044 4798
rect 22428 4562 22596 4564
rect 22428 4510 22430 4562
rect 22482 4510 22596 4562
rect 22428 4508 22596 4510
rect 22988 4562 23044 4732
rect 22988 4510 22990 4562
rect 23042 4510 23044 4562
rect 22428 4498 22484 4508
rect 22988 4498 23044 4510
rect 22428 4340 22484 4350
rect 22316 2772 22372 2782
rect 22316 2678 22372 2716
rect 22316 978 22372 990
rect 22316 926 22318 978
rect 22370 926 22372 978
rect 22316 532 22372 926
rect 22316 466 22372 476
rect 22428 112 22484 4284
rect 22540 3892 22596 3902
rect 22540 3778 22596 3836
rect 22540 3726 22542 3778
rect 22594 3726 22596 3778
rect 22540 3714 22596 3726
rect 22876 3780 22932 3790
rect 22876 2996 22932 3724
rect 22988 3442 23044 3454
rect 22988 3390 22990 3442
rect 23042 3390 23044 3442
rect 22988 3220 23044 3390
rect 22988 3154 23044 3164
rect 22988 2996 23044 3006
rect 22876 2994 23044 2996
rect 22876 2942 22990 2994
rect 23042 2942 23044 2994
rect 22876 2940 23044 2942
rect 22988 2930 23044 2940
rect 22876 2436 22932 2446
rect 22652 2212 22708 2222
rect 22540 1652 22596 1662
rect 22540 1202 22596 1596
rect 22540 1150 22542 1202
rect 22594 1150 22596 1202
rect 22540 1138 22596 1150
rect 22652 112 22708 2156
rect 22876 112 22932 2380
rect 22988 980 23044 990
rect 22988 886 23044 924
rect 23100 112 23156 9436
rect 23212 6468 23268 19852
rect 23436 15316 23492 21420
rect 23804 20412 24068 20422
rect 23860 20356 23908 20412
rect 23964 20356 24012 20412
rect 23804 20346 24068 20356
rect 23804 18844 24068 18854
rect 23860 18788 23908 18844
rect 23964 18788 24012 18844
rect 23804 18778 24068 18788
rect 23436 15250 23492 15260
rect 23660 18676 23716 18686
rect 23660 14532 23716 18620
rect 23804 17276 24068 17286
rect 23860 17220 23908 17276
rect 23964 17220 24012 17276
rect 23804 17210 24068 17220
rect 23804 15708 24068 15718
rect 23860 15652 23908 15708
rect 23964 15652 24012 15708
rect 23804 15642 24068 15652
rect 23772 14532 23828 14542
rect 23660 14530 23828 14532
rect 23660 14478 23774 14530
rect 23826 14478 23828 14530
rect 23660 14476 23828 14478
rect 23660 13748 23716 14476
rect 23772 14466 23828 14476
rect 23804 14140 24068 14150
rect 23860 14084 23908 14140
rect 23964 14084 24012 14140
rect 23804 14074 24068 14084
rect 23772 13748 23828 13758
rect 23660 13746 23828 13748
rect 23660 13694 23774 13746
rect 23826 13694 23828 13746
rect 23660 13692 23828 13694
rect 23660 11844 23716 13692
rect 23772 13682 23828 13692
rect 23804 12572 24068 12582
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 23804 12506 24068 12516
rect 23436 11788 23716 11844
rect 23324 9828 23380 9838
rect 23436 9828 23492 11788
rect 23324 9826 23492 9828
rect 23324 9774 23326 9826
rect 23378 9774 23492 9826
rect 23324 9772 23492 9774
rect 23324 9762 23380 9772
rect 23212 6402 23268 6412
rect 23436 6690 23492 9772
rect 23660 11396 23716 11406
rect 23660 8260 23716 11340
rect 23804 11004 24068 11014
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 23804 10938 24068 10948
rect 23804 9436 24068 9446
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 23804 9370 24068 9380
rect 24108 8932 24164 8942
rect 24108 8838 24164 8876
rect 23660 8204 24276 8260
rect 23436 6638 23438 6690
rect 23490 6638 23492 6690
rect 23212 6020 23268 6030
rect 23212 3388 23268 5964
rect 23324 5348 23380 5358
rect 23324 5254 23380 5292
rect 23436 5124 23492 6638
rect 23436 5058 23492 5068
rect 23548 8148 23604 8158
rect 23436 4676 23492 4686
rect 23212 3332 23380 3388
rect 23212 2100 23268 2110
rect 23212 2006 23268 2044
rect 23324 1202 23380 3332
rect 23324 1150 23326 1202
rect 23378 1150 23380 1202
rect 23324 1138 23380 1150
rect 23436 980 23492 4620
rect 23548 4228 23604 8092
rect 23804 7868 24068 7878
rect 23660 7812 23716 7822
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 23804 7802 24068 7812
rect 23660 7588 23716 7756
rect 23660 7474 23716 7532
rect 23660 7422 23662 7474
rect 23714 7422 23716 7474
rect 23660 7410 23716 7422
rect 23804 6300 24068 6310
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 23804 6234 24068 6244
rect 24108 6132 24164 6142
rect 24108 5794 24164 6076
rect 24108 5742 24110 5794
rect 24162 5742 24164 5794
rect 24108 5730 24164 5742
rect 23996 5348 24052 5358
rect 23996 5254 24052 5292
rect 23660 5234 23716 5246
rect 23660 5182 23662 5234
rect 23714 5182 23716 5234
rect 23660 4452 23716 5182
rect 23804 4732 24068 4742
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 23804 4666 24068 4676
rect 23660 4386 23716 4396
rect 23772 4340 23828 4350
rect 23548 4172 23716 4228
rect 23548 3780 23604 3790
rect 23548 3686 23604 3724
rect 23660 3388 23716 4172
rect 23772 3556 23828 4284
rect 24108 4228 24164 4238
rect 24108 4134 24164 4172
rect 23772 3490 23828 3500
rect 23884 3666 23940 3678
rect 23884 3614 23886 3666
rect 23938 3614 23940 3666
rect 23324 924 23492 980
rect 23548 3332 23716 3388
rect 23884 3332 23940 3614
rect 23324 112 23380 924
rect 23548 112 23604 3332
rect 23884 3266 23940 3276
rect 23804 3164 24068 3174
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 23804 3098 24068 3108
rect 23660 2996 23716 3006
rect 23660 2436 23716 2940
rect 24108 2548 24164 2558
rect 24108 2454 24164 2492
rect 23660 1986 23716 2380
rect 23660 1934 23662 1986
rect 23714 1934 23716 1986
rect 23660 1922 23716 1934
rect 23804 1596 24068 1606
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 23804 1530 24068 1540
rect 23772 1428 23828 1438
rect 23772 112 23828 1372
rect 23996 1428 24052 1438
rect 24220 1428 24276 8204
rect 24332 5348 24388 38220
rect 24464 36876 24728 36886
rect 24520 36820 24568 36876
rect 24624 36820 24672 36876
rect 24464 36810 24728 36820
rect 24464 35308 24728 35318
rect 24520 35252 24568 35308
rect 24624 35252 24672 35308
rect 24464 35242 24728 35252
rect 24780 35028 24836 35038
rect 24780 34934 24836 34972
rect 24668 34916 24724 34926
rect 24668 34822 24724 34860
rect 24892 34130 24948 34142
rect 24892 34078 24894 34130
rect 24946 34078 24948 34130
rect 24668 34020 24724 34030
rect 24668 33926 24724 33964
rect 24464 33740 24728 33750
rect 24520 33684 24568 33740
rect 24624 33684 24672 33740
rect 24464 33674 24728 33684
rect 24464 32172 24728 32182
rect 24520 32116 24568 32172
rect 24624 32116 24672 32172
rect 24464 32106 24728 32116
rect 24892 31892 24948 34078
rect 24892 31826 24948 31836
rect 24464 30604 24728 30614
rect 24520 30548 24568 30604
rect 24624 30548 24672 30604
rect 24464 30538 24728 30548
rect 24464 29036 24728 29046
rect 24520 28980 24568 29036
rect 24624 28980 24672 29036
rect 24464 28970 24728 28980
rect 24464 27468 24728 27478
rect 24520 27412 24568 27468
rect 24624 27412 24672 27468
rect 24464 27402 24728 27412
rect 24464 25900 24728 25910
rect 24520 25844 24568 25900
rect 24624 25844 24672 25900
rect 24464 25834 24728 25844
rect 24464 24332 24728 24342
rect 24520 24276 24568 24332
rect 24624 24276 24672 24332
rect 24464 24266 24728 24276
rect 24464 22764 24728 22774
rect 24520 22708 24568 22764
rect 24624 22708 24672 22764
rect 24464 22698 24728 22708
rect 24464 21196 24728 21206
rect 24520 21140 24568 21196
rect 24624 21140 24672 21196
rect 24464 21130 24728 21140
rect 24464 19628 24728 19638
rect 24520 19572 24568 19628
rect 24624 19572 24672 19628
rect 24464 19562 24728 19572
rect 25004 18452 25060 53004
rect 25004 18386 25060 18396
rect 24464 18060 24728 18070
rect 24520 18004 24568 18060
rect 24624 18004 24672 18060
rect 24464 17994 24728 18004
rect 24892 16772 24948 16782
rect 24464 16492 24728 16502
rect 24520 16436 24568 16492
rect 24624 16436 24672 16492
rect 24464 16426 24728 16436
rect 24464 14924 24728 14934
rect 24520 14868 24568 14924
rect 24624 14868 24672 14924
rect 24464 14858 24728 14868
rect 24892 14868 24948 16716
rect 25340 15148 25396 110012
rect 25788 109228 25844 112478
rect 25900 111412 25956 113260
rect 26348 113314 26404 113326
rect 26348 113262 26350 113314
rect 26402 113262 26404 113314
rect 26236 112306 26292 112318
rect 26236 112254 26238 112306
rect 26290 112254 26292 112306
rect 26012 111748 26068 111786
rect 26236 111748 26292 112254
rect 26012 111682 26068 111692
rect 26124 111746 26292 111748
rect 26124 111694 26238 111746
rect 26290 111694 26292 111746
rect 26124 111692 26292 111694
rect 25900 111356 26068 111412
rect 25900 110068 25956 110078
rect 25900 109974 25956 110012
rect 26012 109956 26068 111356
rect 26124 110962 26180 111692
rect 26236 111682 26292 111692
rect 26348 111300 26404 113262
rect 26572 113316 26628 113326
rect 26460 112980 26516 112990
rect 26460 112418 26516 112924
rect 26460 112366 26462 112418
rect 26514 112366 26516 112418
rect 26460 112354 26516 112366
rect 26572 111970 26628 113260
rect 27020 113314 27076 113326
rect 27020 113262 27022 113314
rect 27074 113262 27076 113314
rect 27020 112868 27076 113262
rect 27916 113314 27972 113326
rect 27916 113262 27918 113314
rect 27970 113262 27972 113314
rect 27020 112802 27076 112812
rect 27132 113204 27188 113214
rect 26908 112420 26964 112430
rect 26572 111918 26574 111970
rect 26626 111918 26628 111970
rect 26572 111906 26628 111918
rect 26796 112306 26852 112318
rect 26796 112254 26798 112306
rect 26850 112254 26852 112306
rect 26796 111972 26852 112254
rect 26796 111906 26852 111916
rect 26124 110910 26126 110962
rect 26178 110910 26180 110962
rect 26124 110852 26180 110910
rect 26124 110786 26180 110796
rect 26236 111244 26404 111300
rect 26460 111748 26516 111758
rect 26012 109890 26068 109900
rect 25788 109172 25956 109228
rect 25676 96180 25732 96190
rect 25452 92708 25508 92718
rect 25452 92614 25508 92652
rect 25452 35476 25508 35486
rect 25452 34914 25508 35420
rect 25452 34862 25454 34914
rect 25506 34862 25508 34914
rect 25452 34850 25508 34862
rect 25452 34132 25508 34142
rect 25452 34038 25508 34076
rect 24892 14802 24948 14812
rect 25228 15092 25396 15148
rect 24464 13356 24728 13366
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24464 13290 24728 13300
rect 25116 12852 25172 12862
rect 24464 11788 24728 11798
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24464 11722 24728 11732
rect 25004 10388 25060 10398
rect 24464 10220 24728 10230
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24464 10154 24728 10164
rect 24556 9156 24612 9166
rect 24556 9062 24612 9100
rect 24892 9156 24948 9166
rect 24464 8652 24728 8662
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24464 8586 24728 8596
rect 24464 7084 24728 7094
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 24464 7018 24728 7028
rect 24556 5908 24612 5918
rect 24556 5814 24612 5852
rect 24464 5516 24728 5526
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24464 5450 24728 5460
rect 24444 5348 24500 5358
rect 24892 5348 24948 9100
rect 24332 5346 24500 5348
rect 24332 5294 24446 5346
rect 24498 5294 24500 5346
rect 24332 5292 24500 5294
rect 24332 3780 24388 5292
rect 24444 5282 24500 5292
rect 24668 5292 24948 5348
rect 24668 4338 24724 5292
rect 25004 5236 25060 10332
rect 25116 5460 25172 12796
rect 25228 5684 25284 15092
rect 25676 10052 25732 96124
rect 25788 92708 25844 92718
rect 25788 92614 25844 92652
rect 25900 87556 25956 109172
rect 26124 109170 26180 109182
rect 26124 109118 26126 109170
rect 26178 109118 26180 109170
rect 26124 108500 26180 109118
rect 26124 108406 26180 108444
rect 26236 106148 26292 111244
rect 26460 110738 26516 111692
rect 26796 111748 26852 111758
rect 26796 110850 26852 111692
rect 26796 110798 26798 110850
rect 26850 110798 26852 110850
rect 26796 110786 26852 110798
rect 26460 110686 26462 110738
rect 26514 110686 26516 110738
rect 26348 110178 26404 110190
rect 26348 110126 26350 110178
rect 26402 110126 26404 110178
rect 26348 108500 26404 110126
rect 26460 110068 26516 110686
rect 26796 110628 26852 110638
rect 26572 110292 26628 110302
rect 26572 110198 26628 110236
rect 26460 110002 26516 110012
rect 26796 110066 26852 110572
rect 26796 110014 26798 110066
rect 26850 110014 26852 110066
rect 26796 109282 26852 110014
rect 26908 109396 26964 112364
rect 27132 112418 27188 113148
rect 27580 113092 27636 113102
rect 27132 112366 27134 112418
rect 27186 112366 27188 112418
rect 27132 112354 27188 112366
rect 27468 112420 27524 112430
rect 27468 112326 27524 112364
rect 27468 112084 27524 112094
rect 27244 111972 27300 111982
rect 27244 111878 27300 111916
rect 27020 111748 27076 111758
rect 27020 111746 27300 111748
rect 27020 111694 27022 111746
rect 27074 111694 27300 111746
rect 27020 111692 27300 111694
rect 27020 111682 27076 111692
rect 27244 110852 27300 111692
rect 27244 110786 27300 110796
rect 27468 110850 27524 112028
rect 27580 111970 27636 113036
rect 27580 111918 27582 111970
rect 27634 111918 27636 111970
rect 27580 111906 27636 111918
rect 27804 111746 27860 111758
rect 27804 111694 27806 111746
rect 27858 111694 27860 111746
rect 27804 111076 27860 111694
rect 27916 111412 27972 113262
rect 28252 112644 28308 112654
rect 28252 111970 28308 112588
rect 28476 112418 28532 114716
rect 29148 114660 29204 114670
rect 29036 114212 29092 114222
rect 29036 113538 29092 114156
rect 29036 113486 29038 113538
rect 29090 113486 29092 113538
rect 29036 113474 29092 113486
rect 28476 112366 28478 112418
rect 28530 112366 28532 112418
rect 28476 112354 28532 112366
rect 28588 113314 28644 113326
rect 28588 113262 28590 113314
rect 28642 113262 28644 113314
rect 28252 111918 28254 111970
rect 28306 111918 28308 111970
rect 28252 111906 28308 111918
rect 28476 111748 28532 111758
rect 28476 111654 28532 111692
rect 28588 111524 28644 113262
rect 28924 112532 28980 112542
rect 28812 112308 28868 112318
rect 28812 112214 28868 112252
rect 28924 111970 28980 112476
rect 29148 112418 29204 114604
rect 29820 113540 29876 113550
rect 29820 113446 29876 113484
rect 29260 113316 29316 113326
rect 29260 113222 29316 113260
rect 30044 113314 30100 113326
rect 30044 113262 30046 113314
rect 30098 113262 30100 113314
rect 29932 112980 29988 112990
rect 29148 112366 29150 112418
rect 29202 112366 29204 112418
rect 29148 112354 29204 112366
rect 29820 112756 29876 112766
rect 29820 112418 29876 112700
rect 29820 112366 29822 112418
rect 29874 112366 29876 112418
rect 29820 112354 29876 112366
rect 28924 111918 28926 111970
rect 28978 111918 28980 111970
rect 28924 111906 28980 111918
rect 29484 112306 29540 112318
rect 29484 112254 29486 112306
rect 29538 112254 29540 112306
rect 29260 111860 29316 111870
rect 29260 111766 29316 111804
rect 28588 111458 28644 111468
rect 27916 111346 27972 111356
rect 29484 111300 29540 112254
rect 29932 111970 29988 112924
rect 30044 112084 30100 113262
rect 30044 112018 30100 112028
rect 30156 112306 30212 112318
rect 30156 112254 30158 112306
rect 30210 112254 30212 112306
rect 29932 111918 29934 111970
rect 29986 111918 29988 111970
rect 29932 111906 29988 111918
rect 30156 111972 30212 112254
rect 30156 111906 30212 111916
rect 30604 111860 30660 111870
rect 30604 111766 30660 111804
rect 29484 111234 29540 111244
rect 29596 111746 29652 111758
rect 29596 111694 29598 111746
rect 29650 111694 29652 111746
rect 29596 111188 29652 111694
rect 30268 111746 30324 111758
rect 30268 111694 30270 111746
rect 30322 111694 30324 111746
rect 30268 111636 30324 111694
rect 30268 111570 30324 111580
rect 29596 111122 29652 111132
rect 27804 111010 27860 111020
rect 30268 110964 30324 110974
rect 27468 110798 27470 110850
rect 27522 110798 27524 110850
rect 27468 110786 27524 110798
rect 29820 110962 30324 110964
rect 29820 110910 30270 110962
rect 30322 110910 30324 110962
rect 29820 110908 30324 110910
rect 29820 110850 29876 110908
rect 30268 110898 30324 110908
rect 29820 110798 29822 110850
rect 29874 110798 29876 110850
rect 29820 110786 29876 110798
rect 27132 110740 27188 110750
rect 29484 110740 29540 110750
rect 27020 110738 27188 110740
rect 27020 110686 27134 110738
rect 27186 110686 27188 110738
rect 27020 110684 27188 110686
rect 27020 110404 27076 110684
rect 27132 110674 27188 110684
rect 29260 110738 29540 110740
rect 29260 110686 29486 110738
rect 29538 110686 29540 110738
rect 29260 110684 29540 110686
rect 27020 110310 27076 110348
rect 27356 110404 27412 110414
rect 27356 110310 27412 110348
rect 27692 110292 27748 110302
rect 27692 110198 27748 110236
rect 26908 109330 26964 109340
rect 27244 110180 27300 110190
rect 26796 109230 26798 109282
rect 26850 109230 26852 109282
rect 26348 108434 26404 108444
rect 26572 109060 26628 109070
rect 26236 106082 26292 106092
rect 26348 94276 26404 94286
rect 26348 90748 26404 94220
rect 25900 87490 25956 87500
rect 26124 90692 26404 90748
rect 26124 73948 26180 90692
rect 26236 89124 26292 89134
rect 26236 76580 26292 89068
rect 26460 82516 26516 82526
rect 26460 82348 26516 82460
rect 26236 76514 26292 76524
rect 26348 82292 26516 82348
rect 26348 76468 26404 82292
rect 26572 80052 26628 109004
rect 26796 97468 26852 109230
rect 27020 109170 27076 109182
rect 27020 109118 27022 109170
rect 27074 109118 27076 109170
rect 27020 109060 27076 109118
rect 27020 108994 27076 109004
rect 26684 97412 26852 97468
rect 27020 108836 27076 108846
rect 26684 85708 26740 97412
rect 26908 93714 26964 93726
rect 26908 93662 26910 93714
rect 26962 93662 26964 93714
rect 26684 85652 26852 85708
rect 26572 79986 26628 79996
rect 26684 76580 26740 76590
rect 26572 76468 26628 76478
rect 26348 76412 26516 76468
rect 26124 73892 26404 73948
rect 26012 39844 26068 39854
rect 25788 34692 25844 34702
rect 25788 34690 25956 34692
rect 25788 34638 25790 34690
rect 25842 34638 25956 34690
rect 25788 34636 25956 34638
rect 25788 34626 25844 34636
rect 25788 33906 25844 33918
rect 25788 33854 25790 33906
rect 25842 33854 25844 33906
rect 25788 32900 25844 33854
rect 25788 32834 25844 32844
rect 25676 9986 25732 9996
rect 25788 17668 25844 17678
rect 25788 7028 25844 17612
rect 25900 16324 25956 34636
rect 26012 30212 26068 39788
rect 26012 30146 26068 30156
rect 25900 16258 25956 16268
rect 26348 15092 26404 73892
rect 26460 15204 26516 76412
rect 26572 15988 26628 76412
rect 26572 15922 26628 15932
rect 26684 15204 26740 76524
rect 26796 17668 26852 85652
rect 26908 75010 26964 93662
rect 26908 74958 26910 75010
rect 26962 74958 26964 75010
rect 26908 74946 26964 74958
rect 27020 20188 27076 108780
rect 27132 108500 27188 108510
rect 27132 89124 27188 108444
rect 27132 89058 27188 89068
rect 27020 20132 27188 20188
rect 26796 17602 26852 17612
rect 27020 17780 27076 17790
rect 26684 15148 26964 15204
rect 26460 15138 26516 15148
rect 26348 15026 26404 15036
rect 26236 14868 26292 14878
rect 25788 6962 25844 6972
rect 26012 14644 26068 14654
rect 25788 6804 25844 6814
rect 25340 5908 25396 5918
rect 25340 5814 25396 5852
rect 25788 5794 25844 6748
rect 25788 5742 25790 5794
rect 25842 5742 25844 5794
rect 25788 5730 25844 5742
rect 25228 5628 25396 5684
rect 25116 5394 25172 5404
rect 25116 5236 25172 5246
rect 25004 5234 25172 5236
rect 25004 5182 25118 5234
rect 25170 5182 25172 5234
rect 25004 5180 25172 5182
rect 25116 4788 25172 5180
rect 25116 4722 25172 4732
rect 24668 4286 24670 4338
rect 24722 4286 24724 4338
rect 24668 4228 24724 4286
rect 25116 4340 25172 4350
rect 24668 4162 24724 4172
rect 25004 4228 25060 4238
rect 24464 3948 24728 3958
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24464 3882 24728 3892
rect 24556 3780 24612 3790
rect 24332 3778 24612 3780
rect 24332 3726 24558 3778
rect 24610 3726 24612 3778
rect 24332 3724 24612 3726
rect 24556 3714 24612 3724
rect 24892 3780 24948 3818
rect 24892 3714 24948 3724
rect 24556 2996 24612 3006
rect 24556 2882 24612 2940
rect 25004 2996 25060 4172
rect 25116 4226 25172 4284
rect 25116 4174 25118 4226
rect 25170 4174 25172 4226
rect 25116 4162 25172 4174
rect 25228 3780 25284 3790
rect 25228 3722 25284 3724
rect 25228 3670 25230 3722
rect 25282 3670 25284 3722
rect 25228 3658 25284 3670
rect 25004 2930 25060 2940
rect 25228 3220 25284 3230
rect 24556 2830 24558 2882
rect 24610 2830 24612 2882
rect 24556 2818 24612 2830
rect 25116 2546 25172 2558
rect 25116 2494 25118 2546
rect 25170 2494 25172 2546
rect 24464 2380 24728 2390
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24464 2314 24728 2324
rect 24892 2324 24948 2334
rect 24668 2212 24724 2222
rect 24892 2212 24948 2268
rect 24668 2210 24948 2212
rect 24668 2158 24670 2210
rect 24722 2158 24948 2210
rect 24668 2156 24948 2158
rect 24668 2146 24724 2156
rect 25116 1876 25172 2494
rect 25116 1810 25172 1820
rect 25116 1652 25172 1662
rect 23996 1426 24276 1428
rect 23996 1374 23998 1426
rect 24050 1374 24276 1426
rect 23996 1372 24276 1374
rect 24332 1540 24388 1550
rect 23996 1362 24052 1372
rect 23996 1204 24052 1214
rect 23996 112 24052 1148
rect 24332 756 24388 1484
rect 24892 1316 24948 1326
rect 24220 700 24388 756
rect 24464 812 24728 822
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24464 746 24728 756
rect 24220 112 24276 700
rect 24444 644 24500 654
rect 24444 112 24500 588
rect 24668 644 24724 654
rect 24668 112 24724 588
rect 24892 112 24948 1260
rect 25116 112 25172 1596
rect 25228 1090 25284 3164
rect 25228 1038 25230 1090
rect 25282 1038 25284 1090
rect 25228 1026 25284 1038
rect 25340 112 25396 5628
rect 25564 4788 25620 4798
rect 25452 4114 25508 4126
rect 25452 4062 25454 4114
rect 25506 4062 25508 4114
rect 25452 4004 25508 4062
rect 25452 3938 25508 3948
rect 25564 3778 25620 4732
rect 25564 3726 25566 3778
rect 25618 3726 25620 3778
rect 25564 3714 25620 3726
rect 25900 3666 25956 3678
rect 25900 3614 25902 3666
rect 25954 3614 25956 3666
rect 25900 3556 25956 3614
rect 25900 3490 25956 3500
rect 26012 3220 26068 14588
rect 26012 3154 26068 3164
rect 26124 9940 26180 9950
rect 26124 2996 26180 9884
rect 26236 3778 26292 14812
rect 26460 14868 26516 14878
rect 26348 5348 26404 5358
rect 26460 5348 26516 14812
rect 26572 14644 26628 14654
rect 26572 7364 26628 14588
rect 26908 11788 26964 15148
rect 26572 7298 26628 7308
rect 26684 11732 26964 11788
rect 26348 5346 26516 5348
rect 26348 5294 26350 5346
rect 26402 5294 26516 5346
rect 26348 5292 26516 5294
rect 26348 5282 26404 5292
rect 26460 4452 26516 5292
rect 26460 4386 26516 4396
rect 26236 3726 26238 3778
rect 26290 3726 26292 3778
rect 26236 3714 26292 3726
rect 26348 4228 26404 4238
rect 25900 2940 26180 2996
rect 25452 2772 25508 2782
rect 25452 2678 25508 2716
rect 25788 2548 25844 2558
rect 25788 2454 25844 2492
rect 25788 2324 25844 2334
rect 25452 2212 25508 2222
rect 25452 1316 25508 2156
rect 25564 1316 25620 1326
rect 25452 1314 25620 1316
rect 25452 1262 25566 1314
rect 25618 1262 25620 1314
rect 25452 1260 25620 1262
rect 25564 1250 25620 1260
rect 25564 868 25620 878
rect 25564 112 25620 812
rect 25788 112 25844 2268
rect 25900 2098 25956 2940
rect 26124 2772 26180 2782
rect 26348 2772 26404 4172
rect 26572 4116 26628 4126
rect 26572 3778 26628 4060
rect 26684 3892 26740 11732
rect 26908 5796 26964 5806
rect 26908 5702 26964 5740
rect 26684 3826 26740 3836
rect 26572 3726 26574 3778
rect 26626 3726 26628 3778
rect 26572 3714 26628 3726
rect 26796 3556 26852 3566
rect 26796 3462 26852 3500
rect 26684 2772 26740 2782
rect 26348 2770 26740 2772
rect 26348 2718 26686 2770
rect 26738 2718 26740 2770
rect 26348 2716 26740 2718
rect 26124 2678 26180 2716
rect 26684 2706 26740 2716
rect 26460 2546 26516 2558
rect 26460 2494 26462 2546
rect 26514 2494 26516 2546
rect 25900 2046 25902 2098
rect 25954 2046 25956 2098
rect 25900 2034 25956 2046
rect 26348 2212 26404 2222
rect 26236 1876 26292 1886
rect 26236 1782 26292 1820
rect 26012 1652 26068 1662
rect 26012 112 26068 1596
rect 26348 1202 26404 2156
rect 26348 1150 26350 1202
rect 26402 1150 26404 1202
rect 26348 1138 26404 1150
rect 26124 1092 26180 1102
rect 26124 998 26180 1036
rect 5376 0 5488 112
rect 5600 0 5712 112
rect 5824 0 5936 112
rect 6048 0 6160 112
rect 6272 0 6384 112
rect 6496 0 6608 112
rect 6720 0 6832 112
rect 6944 0 7056 112
rect 7168 0 7280 112
rect 7392 0 7504 112
rect 7616 0 7728 112
rect 7840 0 7952 112
rect 8064 0 8176 112
rect 8288 0 8400 112
rect 8512 0 8624 112
rect 8736 0 8848 112
rect 8960 0 9072 112
rect 9184 0 9296 112
rect 9408 0 9520 112
rect 9632 0 9744 112
rect 9856 0 9968 112
rect 10080 0 10192 112
rect 10304 0 10416 112
rect 10528 0 10640 112
rect 10752 0 10864 112
rect 10976 0 11088 112
rect 11200 0 11312 112
rect 11424 0 11536 112
rect 11648 0 11760 112
rect 11872 0 11984 112
rect 12096 0 12208 112
rect 12320 0 12432 112
rect 12544 0 12656 112
rect 12768 0 12880 112
rect 12992 0 13104 112
rect 13216 0 13328 112
rect 13440 0 13552 112
rect 13664 0 13776 112
rect 13888 0 14000 112
rect 14112 0 14224 112
rect 14336 0 14448 112
rect 14560 0 14672 112
rect 14784 0 14896 112
rect 15008 0 15120 112
rect 15232 0 15344 112
rect 15456 0 15568 112
rect 15680 0 15792 112
rect 15904 0 16016 112
rect 16128 0 16240 112
rect 16352 0 16464 112
rect 16576 0 16688 112
rect 16800 0 16912 112
rect 17024 0 17136 112
rect 17248 0 17360 112
rect 17472 0 17584 112
rect 17696 0 17808 112
rect 17920 0 18032 112
rect 18144 0 18256 112
rect 18368 0 18480 112
rect 18592 0 18704 112
rect 18816 0 18928 112
rect 19040 0 19152 112
rect 19264 0 19376 112
rect 19488 0 19600 112
rect 19712 0 19824 112
rect 19936 0 20048 112
rect 20160 0 20272 112
rect 20384 0 20496 112
rect 20608 0 20720 112
rect 20832 0 20944 112
rect 21056 0 21168 112
rect 21280 0 21392 112
rect 21504 0 21616 112
rect 21728 0 21840 112
rect 21952 0 22064 112
rect 22176 0 22288 112
rect 22400 0 22512 112
rect 22624 0 22736 112
rect 22848 0 22960 112
rect 23072 0 23184 112
rect 23296 0 23408 112
rect 23520 0 23632 112
rect 23744 0 23856 112
rect 23968 0 24080 112
rect 24192 0 24304 112
rect 24416 0 24528 112
rect 24640 0 24752 112
rect 24864 0 24976 112
rect 25088 0 25200 112
rect 25312 0 25424 112
rect 25536 0 25648 112
rect 25760 0 25872 112
rect 25984 0 26096 112
rect 26460 84 26516 2494
rect 26796 2100 26852 2110
rect 26796 2006 26852 2044
rect 27020 1986 27076 17724
rect 27132 2772 27188 20132
rect 27244 5124 27300 110124
rect 28476 109060 28532 109070
rect 27356 108388 27412 108398
rect 27356 6916 27412 108332
rect 27804 94388 27860 94398
rect 27692 74786 27748 74798
rect 27692 74734 27694 74786
rect 27746 74734 27748 74786
rect 27692 55300 27748 74734
rect 27692 55234 27748 55244
rect 27356 6850 27412 6860
rect 27692 38164 27748 38174
rect 27692 6580 27748 38108
rect 27804 17892 27860 94332
rect 28028 92708 28084 92718
rect 27916 90356 27972 90366
rect 27916 19460 27972 90300
rect 28028 35140 28084 92652
rect 28028 35074 28084 35084
rect 28140 85652 28196 85662
rect 28140 27972 28196 85596
rect 28252 56308 28308 56318
rect 28252 43708 28308 56252
rect 28364 55300 28420 55310
rect 28364 55206 28420 55244
rect 28252 43652 28420 43708
rect 28140 27906 28196 27916
rect 28252 40964 28308 40974
rect 27916 19394 27972 19404
rect 28028 26852 28084 26862
rect 27804 17826 27860 17836
rect 27692 6514 27748 6524
rect 27804 15204 27860 15214
rect 27244 5058 27300 5068
rect 27468 6468 27524 6478
rect 27356 4900 27412 4910
rect 27132 2716 27300 2772
rect 27020 1934 27022 1986
rect 27074 1934 27076 1986
rect 27020 1922 27076 1934
rect 27132 2546 27188 2558
rect 27132 2494 27134 2546
rect 27186 2494 27188 2546
rect 27132 1988 27188 2494
rect 27132 1922 27188 1932
rect 27244 1204 27300 2716
rect 27356 2770 27412 4844
rect 27356 2718 27358 2770
rect 27410 2718 27412 2770
rect 27356 2706 27412 2718
rect 27468 2324 27524 6412
rect 27244 1138 27300 1148
rect 27356 2268 27524 2324
rect 26796 978 26852 990
rect 26796 926 26798 978
rect 26850 926 26852 978
rect 26796 196 26852 926
rect 27132 980 27188 990
rect 27356 980 27412 2268
rect 27804 2210 27860 15148
rect 28028 11620 28084 26796
rect 28028 11554 28084 11564
rect 28252 9268 28308 40908
rect 28364 24724 28420 43652
rect 28364 24658 28420 24668
rect 28252 9202 28308 9212
rect 28476 8428 28532 109004
rect 29260 98980 29316 110684
rect 29484 110674 29540 110684
rect 30604 110740 30660 110750
rect 30604 110646 30660 110684
rect 30604 110290 30660 110302
rect 30604 110238 30606 110290
rect 30658 110238 30660 110290
rect 30268 110180 30324 110190
rect 29820 110178 30324 110180
rect 29820 110126 30270 110178
rect 30322 110126 30324 110178
rect 29820 110124 30324 110126
rect 29484 109508 29540 109518
rect 29484 109394 29540 109452
rect 29484 109342 29486 109394
rect 29538 109342 29540 109394
rect 29484 109330 29540 109342
rect 29820 109282 29876 110124
rect 30268 110114 30324 110124
rect 30604 109620 30660 110238
rect 30604 109554 30660 109564
rect 29820 109230 29822 109282
rect 29874 109230 29876 109282
rect 29820 109218 29876 109230
rect 29820 108724 29876 108734
rect 30268 108724 30324 108734
rect 29820 108722 30324 108724
rect 29820 108670 29822 108722
rect 29874 108670 30270 108722
rect 30322 108670 30324 108722
rect 29820 108668 30324 108670
rect 29820 108658 29876 108668
rect 30268 108658 30324 108668
rect 30380 108724 30436 108734
rect 29596 108610 29652 108622
rect 29596 108558 29598 108610
rect 29650 108558 29652 108610
rect 29484 106034 29540 106046
rect 29484 105982 29486 106034
rect 29538 105982 29540 106034
rect 29484 102508 29540 105982
rect 29596 106036 29652 108558
rect 30380 107826 30436 108668
rect 30604 108722 30660 108734
rect 30604 108670 30606 108722
rect 30658 108670 30660 108722
rect 30604 108500 30660 108670
rect 30604 108434 30660 108444
rect 30380 107774 30382 107826
rect 30434 107774 30436 107826
rect 30380 107762 30436 107774
rect 30604 107602 30660 107614
rect 30604 107550 30606 107602
rect 30658 107550 30660 107602
rect 30604 107380 30660 107550
rect 30604 107314 30660 107324
rect 30604 107154 30660 107166
rect 30604 107102 30606 107154
rect 30658 107102 30660 107154
rect 30268 107044 30324 107054
rect 29820 107042 30324 107044
rect 29820 106990 30270 107042
rect 30322 106990 30324 107042
rect 29820 106988 30324 106990
rect 29820 106146 29876 106988
rect 30268 106978 30324 106988
rect 30604 106260 30660 107102
rect 30604 106194 30660 106204
rect 29820 106094 29822 106146
rect 29874 106094 29876 106146
rect 29820 106082 29876 106094
rect 29596 105970 29652 105980
rect 30268 105588 30324 105598
rect 30268 105494 30324 105532
rect 30604 105586 30660 105598
rect 30604 105534 30606 105586
rect 30658 105534 30660 105586
rect 30604 105140 30660 105534
rect 30604 105074 30660 105084
rect 30268 104466 30324 104478
rect 30268 104414 30270 104466
rect 30322 104414 30324 104466
rect 30268 104132 30324 104414
rect 30268 104066 30324 104076
rect 30604 104466 30660 104478
rect 30604 104414 30606 104466
rect 30658 104414 30660 104466
rect 30604 104020 30660 104414
rect 30604 103954 30660 103964
rect 30268 102900 30324 102910
rect 30268 102806 30324 102844
rect 30604 102900 30660 102910
rect 30604 102806 30660 102844
rect 29372 102452 29540 102508
rect 30268 102452 30324 102462
rect 29372 99092 29428 102452
rect 30268 102358 30324 102396
rect 30604 102450 30660 102462
rect 30604 102398 30606 102450
rect 30658 102398 30660 102450
rect 30604 101780 30660 102398
rect 30604 101714 30660 101724
rect 29820 100882 29876 100894
rect 29820 100830 29822 100882
rect 29874 100830 29876 100882
rect 29484 100772 29540 100782
rect 29820 100772 29876 100830
rect 30604 100882 30660 100894
rect 30604 100830 30606 100882
rect 30658 100830 30660 100882
rect 30268 100772 30324 100782
rect 29820 100770 30324 100772
rect 29820 100718 30270 100770
rect 30322 100718 30324 100770
rect 29820 100716 30324 100718
rect 29484 100678 29540 100716
rect 30268 100706 30324 100716
rect 30604 100660 30660 100830
rect 30604 100594 30660 100604
rect 30268 99764 30324 99774
rect 30268 99670 30324 99708
rect 30604 99762 30660 99774
rect 30604 99710 30606 99762
rect 30658 99710 30660 99762
rect 30604 99540 30660 99710
rect 30604 99474 30660 99484
rect 30268 99316 30324 99326
rect 30268 99222 30324 99260
rect 30604 99314 30660 99326
rect 30604 99262 30606 99314
rect 30658 99262 30660 99314
rect 29372 99026 29428 99036
rect 29260 98914 29316 98924
rect 30604 98420 30660 99262
rect 30604 98354 30660 98364
rect 29820 97748 29876 97758
rect 30268 97748 30324 97758
rect 29820 97746 30324 97748
rect 29820 97694 29822 97746
rect 29874 97694 30270 97746
rect 30322 97694 30324 97746
rect 29820 97692 30324 97694
rect 29820 97682 29876 97692
rect 30268 97682 30324 97692
rect 30604 97746 30660 97758
rect 30604 97694 30606 97746
rect 30658 97694 30660 97746
rect 29484 97634 29540 97646
rect 29484 97582 29486 97634
rect 29538 97582 29540 97634
rect 29484 96852 29540 97582
rect 30604 97300 30660 97694
rect 30604 97234 30660 97244
rect 29484 96786 29540 96796
rect 29484 96628 29540 96638
rect 30268 96628 30324 96638
rect 29484 96290 29540 96572
rect 29484 96238 29486 96290
rect 29538 96238 29540 96290
rect 29484 96226 29540 96238
rect 29820 96626 30324 96628
rect 29820 96574 30270 96626
rect 30322 96574 30324 96626
rect 29820 96572 30324 96574
rect 29820 96290 29876 96572
rect 30268 96562 30324 96572
rect 30604 96626 30660 96638
rect 30604 96574 30606 96626
rect 30658 96574 30660 96626
rect 29820 96238 29822 96290
rect 29874 96238 29876 96290
rect 29820 96226 29876 96238
rect 30604 96180 30660 96574
rect 30604 96114 30660 96124
rect 30380 95284 30436 95294
rect 30268 95058 30324 95070
rect 30268 95006 30270 95058
rect 30322 95006 30324 95058
rect 30268 94724 30324 95006
rect 30268 94658 30324 94668
rect 30380 94498 30436 95228
rect 30604 95060 30660 95070
rect 30604 94966 30660 95004
rect 30380 94446 30382 94498
rect 30434 94446 30436 94498
rect 30380 94434 30436 94446
rect 30604 94610 30660 94622
rect 30604 94558 30606 94610
rect 30658 94558 30660 94610
rect 30604 93940 30660 94558
rect 30604 93874 30660 93884
rect 30268 93492 30324 93502
rect 30268 93154 30324 93436
rect 30268 93102 30270 93154
rect 30322 93102 30324 93154
rect 30268 93090 30324 93102
rect 30604 93042 30660 93054
rect 30604 92990 30606 93042
rect 30658 92990 30660 93042
rect 30604 92820 30660 92990
rect 30604 92754 30660 92764
rect 30268 91924 30324 91934
rect 30268 91830 30324 91868
rect 30604 91922 30660 91934
rect 30604 91870 30606 91922
rect 30658 91870 30660 91922
rect 30604 91700 30660 91870
rect 30604 91634 30660 91644
rect 30604 91474 30660 91486
rect 30604 91422 30606 91474
rect 30658 91422 30660 91474
rect 30268 91362 30324 91374
rect 30268 91310 30270 91362
rect 30322 91310 30324 91362
rect 30268 90468 30324 91310
rect 30604 90580 30660 91422
rect 30604 90514 30660 90524
rect 30268 90402 30324 90412
rect 30268 89908 30324 89918
rect 30268 89814 30324 89852
rect 30604 89906 30660 89918
rect 30604 89854 30606 89906
rect 30658 89854 30660 89906
rect 30604 89460 30660 89854
rect 30604 89394 30660 89404
rect 30268 88788 30324 88798
rect 29820 88786 30324 88788
rect 29820 88734 30270 88786
rect 30322 88734 30324 88786
rect 29820 88732 30324 88734
rect 29820 88450 29876 88732
rect 30268 88722 30324 88732
rect 30604 88786 30660 88798
rect 30604 88734 30606 88786
rect 30658 88734 30660 88786
rect 29820 88398 29822 88450
rect 29874 88398 29876 88450
rect 29820 88386 29876 88398
rect 30604 88340 30660 88734
rect 30604 88274 30660 88284
rect 29484 88228 29540 88238
rect 29372 88226 29540 88228
rect 29372 88174 29486 88226
rect 29538 88174 29540 88226
rect 29372 88172 29540 88174
rect 29372 77812 29428 88172
rect 29484 88162 29540 88172
rect 30268 87444 30324 87454
rect 30268 87350 30324 87388
rect 30604 87220 30660 87230
rect 30604 87126 30660 87164
rect 30604 86770 30660 86782
rect 30604 86718 30606 86770
rect 30658 86718 30660 86770
rect 30268 86658 30324 86670
rect 30268 86606 30270 86658
rect 30322 86606 30324 86658
rect 30268 85764 30324 86606
rect 30604 86100 30660 86718
rect 30604 86034 30660 86044
rect 30268 85698 30324 85708
rect 30268 85204 30324 85214
rect 30268 85110 30324 85148
rect 30604 85202 30660 85214
rect 30604 85150 30606 85202
rect 30658 85150 30660 85202
rect 30604 84980 30660 85150
rect 30604 84914 30660 84924
rect 30268 84084 30324 84094
rect 30268 83990 30324 84028
rect 30604 84082 30660 84094
rect 30604 84030 30606 84082
rect 30658 84030 30660 84082
rect 30604 83860 30660 84030
rect 30604 83794 30660 83804
rect 30604 83634 30660 83646
rect 30604 83582 30606 83634
rect 30658 83582 30660 83634
rect 30268 83522 30324 83534
rect 30268 83470 30270 83522
rect 30322 83470 30324 83522
rect 30268 82628 30324 83470
rect 30604 82740 30660 83582
rect 30604 82674 30660 82684
rect 30268 82562 30324 82572
rect 29820 82068 29876 82078
rect 30268 82068 30324 82078
rect 29820 82066 30324 82068
rect 29820 82014 29822 82066
rect 29874 82014 30270 82066
rect 30322 82014 30324 82066
rect 29820 82012 30324 82014
rect 29820 82002 29876 82012
rect 30268 82002 30324 82012
rect 30604 82066 30660 82078
rect 30604 82014 30606 82066
rect 30658 82014 30660 82066
rect 29484 81956 29540 81966
rect 29484 81862 29540 81900
rect 30604 81620 30660 82014
rect 30604 81554 30660 81564
rect 30268 80948 30324 80958
rect 29820 80946 30324 80948
rect 29820 80894 30270 80946
rect 30322 80894 30324 80946
rect 29820 80892 30324 80894
rect 29820 80610 29876 80892
rect 30268 80882 30324 80892
rect 30604 80946 30660 80958
rect 30604 80894 30606 80946
rect 30658 80894 30660 80946
rect 29820 80558 29822 80610
rect 29874 80558 29876 80610
rect 29820 80546 29876 80558
rect 30604 80500 30660 80894
rect 30604 80434 30660 80444
rect 29484 80386 29540 80398
rect 29484 80334 29486 80386
rect 29538 80334 29540 80386
rect 29484 79716 29540 80334
rect 29484 79650 29540 79660
rect 29484 79378 29540 79390
rect 29484 79326 29486 79378
rect 29538 79326 29540 79378
rect 29484 78932 29540 79326
rect 29820 79380 29876 79390
rect 30268 79380 30324 79390
rect 29820 79378 30324 79380
rect 29820 79326 29822 79378
rect 29874 79326 30270 79378
rect 30322 79326 30324 79378
rect 29820 79324 30324 79326
rect 29820 79314 29876 79324
rect 30268 79314 30324 79324
rect 30604 79380 30660 79390
rect 30604 79286 30660 79324
rect 29484 78866 29540 78876
rect 30604 78930 30660 78942
rect 30604 78878 30606 78930
rect 30658 78878 30660 78930
rect 30268 78820 30324 78830
rect 29820 78818 30324 78820
rect 29820 78766 30270 78818
rect 30322 78766 30324 78818
rect 29820 78764 30324 78766
rect 29484 77924 29540 77934
rect 29484 77830 29540 77868
rect 29820 77922 29876 78764
rect 30268 78754 30324 78764
rect 30604 78260 30660 78878
rect 30604 78194 30660 78204
rect 29820 77870 29822 77922
rect 29874 77870 29876 77922
rect 29820 77858 29876 77870
rect 29372 77746 29428 77756
rect 30268 74676 30324 74686
rect 30268 74582 30324 74620
rect 30604 74676 30660 74686
rect 30604 74582 30660 74620
rect 30604 74226 30660 74238
rect 30604 74174 30606 74226
rect 30658 74174 30660 74226
rect 30268 74116 30324 74126
rect 30268 74022 30324 74060
rect 30604 73556 30660 74174
rect 30604 73490 30660 73500
rect 30604 72658 30660 72670
rect 30604 72606 30606 72658
rect 30658 72606 30660 72658
rect 30268 72548 30324 72558
rect 29820 72546 30324 72548
rect 29820 72494 30270 72546
rect 30322 72494 30324 72546
rect 29820 72492 30324 72494
rect 29820 71202 29876 72492
rect 30268 72482 30324 72492
rect 30604 72436 30660 72606
rect 30604 72370 30660 72380
rect 29820 71150 29822 71202
rect 29874 71150 29876 71202
rect 29820 71138 29876 71150
rect 30380 71762 30436 71774
rect 30380 71710 30382 71762
rect 30434 71710 30436 71762
rect 29484 70980 29540 70990
rect 30268 70980 30324 70990
rect 29484 70886 29540 70924
rect 29820 70978 30324 70980
rect 29820 70926 30270 70978
rect 30322 70926 30324 70978
rect 29820 70924 30324 70926
rect 29820 68514 29876 70924
rect 30268 70914 30324 70924
rect 30268 69412 30324 69422
rect 29820 68462 29822 68514
rect 29874 68462 29876 68514
rect 29820 68450 29876 68462
rect 29932 69410 30324 69412
rect 29932 69358 30270 69410
rect 30322 69358 30324 69410
rect 29932 69356 30324 69358
rect 28700 68404 28756 68414
rect 28700 58212 28756 68348
rect 29484 68404 29540 68414
rect 29484 68310 29540 68348
rect 29820 68068 29876 68078
rect 29932 68068 29988 69356
rect 30268 69346 30324 69356
rect 29820 68066 29988 68068
rect 29820 68014 29822 68066
rect 29874 68014 29988 68066
rect 29820 68012 29988 68014
rect 30268 68402 30324 68414
rect 30268 68350 30270 68402
rect 30322 68350 30324 68402
rect 29820 68002 29876 68012
rect 29596 67842 29652 67854
rect 29596 67790 29598 67842
rect 29650 67790 29652 67842
rect 29596 67228 29652 67790
rect 29596 67172 29764 67228
rect 29484 63700 29540 63710
rect 29148 63698 29540 63700
rect 29148 63646 29486 63698
rect 29538 63646 29540 63698
rect 29148 63644 29540 63646
rect 28700 58146 28756 58156
rect 28812 63140 28868 63150
rect 28812 48132 28868 63084
rect 29148 55468 29204 63644
rect 29484 63634 29540 63644
rect 29484 63140 29540 63150
rect 29484 63046 29540 63084
rect 29596 61570 29652 61582
rect 29596 61518 29598 61570
rect 29650 61518 29652 61570
rect 29484 60562 29540 60574
rect 29484 60510 29486 60562
rect 29538 60510 29540 60562
rect 29484 60340 29540 60510
rect 29260 60284 29540 60340
rect 29260 56644 29316 60284
rect 29596 60228 29652 61518
rect 29596 60162 29652 60172
rect 29484 60002 29540 60014
rect 29484 59950 29486 60002
rect 29538 59950 29540 60002
rect 29484 59444 29540 59950
rect 29708 59780 29764 67172
rect 30268 66500 30324 68350
rect 30380 67228 30436 71710
rect 30604 71538 30660 71550
rect 30604 71486 30606 71538
rect 30658 71486 30660 71538
rect 30604 71316 30660 71486
rect 30604 71250 30660 71260
rect 30604 71090 30660 71102
rect 30604 71038 30606 71090
rect 30658 71038 30660 71090
rect 30604 70196 30660 71038
rect 30604 70130 30660 70140
rect 30604 69522 30660 69534
rect 30604 69470 30606 69522
rect 30658 69470 30660 69522
rect 30604 69076 30660 69470
rect 30604 69010 30660 69020
rect 30604 68402 30660 68414
rect 30604 68350 30606 68402
rect 30658 68350 30660 68402
rect 30604 67956 30660 68350
rect 30604 67890 30660 67900
rect 30380 67172 30548 67228
rect 30268 66434 30324 66444
rect 30380 67058 30436 67070
rect 30380 67006 30382 67058
rect 30434 67006 30436 67058
rect 30268 66276 30324 66286
rect 29820 66274 30324 66276
rect 29820 66222 30270 66274
rect 30322 66222 30324 66274
rect 29820 66220 30324 66222
rect 29820 63810 29876 66220
rect 30268 66210 30324 66220
rect 30380 64820 30436 67006
rect 30380 64754 30436 64764
rect 30268 64708 30324 64718
rect 29820 63758 29822 63810
rect 29874 63758 29876 63810
rect 29820 63746 29876 63758
rect 29932 64706 30324 64708
rect 29932 64654 30270 64706
rect 30322 64654 30324 64706
rect 29932 64652 30324 64654
rect 29820 63364 29876 63374
rect 29932 63364 29988 64652
rect 30268 64642 30324 64652
rect 30492 63924 30548 67172
rect 30604 66836 30660 66846
rect 30604 66742 30660 66780
rect 30604 66386 30660 66398
rect 30604 66334 30606 66386
rect 30658 66334 30660 66386
rect 30604 65716 30660 66334
rect 30604 65650 30660 65660
rect 30604 64818 30660 64830
rect 30604 64766 30606 64818
rect 30658 64766 30660 64818
rect 30604 64596 30660 64766
rect 30604 64530 30660 64540
rect 30492 63858 30548 63868
rect 30268 63700 30324 63710
rect 29820 63362 29988 63364
rect 29820 63310 29822 63362
rect 29874 63310 29988 63362
rect 29820 63308 29988 63310
rect 30044 63698 30324 63700
rect 30044 63646 30270 63698
rect 30322 63646 30324 63698
rect 30044 63644 30324 63646
rect 29820 63298 29876 63308
rect 30044 62692 30100 63644
rect 30268 63634 30324 63644
rect 30604 63698 30660 63710
rect 30604 63646 30606 63698
rect 30658 63646 30660 63698
rect 30604 63476 30660 63646
rect 30604 63410 30660 63420
rect 30604 63250 30660 63262
rect 30604 63198 30606 63250
rect 30658 63198 30660 63250
rect 30268 63140 30324 63150
rect 29820 62636 30100 62692
rect 30156 63138 30324 63140
rect 30156 63086 30270 63138
rect 30322 63086 30324 63138
rect 30156 63084 30324 63086
rect 29820 61794 29876 62636
rect 30156 61796 30212 63084
rect 30268 63074 30324 63084
rect 30604 62356 30660 63198
rect 30604 62290 30660 62300
rect 29820 61742 29822 61794
rect 29874 61742 29876 61794
rect 29820 61730 29876 61742
rect 29932 61740 30212 61796
rect 29932 61572 29988 61740
rect 30604 61682 30660 61694
rect 30604 61630 30606 61682
rect 30658 61630 30660 61682
rect 30268 61572 30324 61582
rect 29820 61516 29988 61572
rect 30044 61570 30324 61572
rect 30044 61518 30270 61570
rect 30322 61518 30324 61570
rect 30044 61516 30324 61518
rect 29820 60674 29876 61516
rect 30044 60676 30100 61516
rect 30268 61506 30324 61516
rect 30604 61236 30660 61630
rect 30604 61170 30660 61180
rect 29820 60622 29822 60674
rect 29874 60622 29876 60674
rect 29820 60610 29876 60622
rect 29932 60620 30100 60676
rect 29820 60228 29876 60238
rect 29932 60228 29988 60620
rect 30268 60564 30324 60574
rect 29820 60226 29988 60228
rect 29820 60174 29822 60226
rect 29874 60174 29988 60226
rect 29820 60172 29988 60174
rect 30044 60562 30324 60564
rect 30044 60510 30270 60562
rect 30322 60510 30324 60562
rect 30044 60508 30324 60510
rect 29820 60162 29876 60172
rect 29708 59714 29764 59724
rect 30044 59556 30100 60508
rect 30268 60498 30324 60508
rect 30604 60562 30660 60574
rect 30604 60510 30606 60562
rect 30658 60510 30660 60562
rect 30604 60116 30660 60510
rect 30604 60050 30660 60060
rect 29484 59378 29540 59388
rect 29820 59500 30100 59556
rect 29820 58658 29876 59500
rect 30268 58996 30324 59006
rect 29820 58606 29822 58658
rect 29874 58606 29876 58658
rect 29820 58594 29876 58606
rect 29932 58994 30324 58996
rect 29932 58942 30270 58994
rect 30322 58942 30324 58994
rect 29932 58940 30324 58942
rect 29484 58434 29540 58446
rect 29484 58382 29486 58434
rect 29538 58382 29540 58434
rect 29484 57764 29540 58382
rect 29484 57698 29540 57708
rect 29820 57540 29876 57550
rect 29932 57540 29988 58940
rect 30268 58930 30324 58940
rect 30604 58996 30660 59006
rect 30604 58902 30660 58940
rect 30604 58546 30660 58558
rect 30604 58494 30606 58546
rect 30658 58494 30660 58546
rect 29820 57538 29988 57540
rect 29820 57486 29822 57538
rect 29874 57486 29988 57538
rect 29820 57484 29988 57486
rect 30268 58434 30324 58446
rect 30268 58382 30270 58434
rect 30322 58382 30324 58434
rect 29820 57474 29876 57484
rect 29260 56578 29316 56588
rect 29484 57426 29540 57438
rect 29484 57374 29486 57426
rect 29538 57374 29540 57426
rect 29148 55412 29428 55468
rect 29372 50708 29428 55412
rect 29484 51940 29540 57374
rect 30268 56084 30324 58382
rect 30604 57876 30660 58494
rect 30604 57810 30660 57820
rect 30604 56978 30660 56990
rect 30604 56926 30606 56978
rect 30658 56926 30660 56978
rect 30268 56018 30324 56028
rect 30380 56866 30436 56878
rect 30380 56814 30382 56866
rect 30434 56814 30436 56866
rect 30268 55858 30324 55870
rect 30268 55806 30270 55858
rect 30322 55806 30324 55858
rect 30268 55468 30324 55806
rect 30380 55524 30436 56814
rect 30604 56756 30660 56926
rect 30604 56690 30660 56700
rect 30604 55858 30660 55870
rect 30604 55806 30606 55858
rect 30658 55806 30660 55858
rect 30604 55636 30660 55806
rect 30604 55570 30660 55580
rect 30492 55524 30548 55534
rect 30380 55522 30548 55524
rect 30380 55470 30494 55522
rect 30546 55470 30548 55522
rect 30380 55468 30548 55470
rect 29932 55412 30324 55468
rect 30492 55458 30548 55468
rect 29932 53732 29988 55412
rect 30156 55300 30212 55310
rect 29932 53666 29988 53676
rect 30044 55298 30212 55300
rect 30044 55246 30158 55298
rect 30210 55246 30212 55298
rect 30044 55244 30212 55246
rect 29484 51874 29540 51884
rect 29372 50642 29428 50652
rect 30044 48356 30100 55244
rect 30156 55234 30212 55244
rect 30604 54516 30660 54526
rect 30604 54402 30660 54460
rect 30604 54350 30606 54402
rect 30658 54350 30660 54402
rect 30604 54338 30660 54350
rect 30268 54292 30324 54302
rect 30156 54290 30324 54292
rect 30156 54238 30270 54290
rect 30322 54238 30324 54290
rect 30156 54236 30324 54238
rect 30156 53508 30212 54236
rect 30268 54226 30324 54236
rect 30604 53842 30660 53854
rect 30604 53790 30606 53842
rect 30658 53790 30660 53842
rect 30156 53442 30212 53452
rect 30380 53730 30436 53742
rect 30380 53678 30382 53730
rect 30434 53678 30436 53730
rect 30268 52722 30324 52734
rect 30268 52670 30270 52722
rect 30322 52670 30324 52722
rect 30268 52276 30324 52670
rect 30380 52724 30436 53678
rect 30604 53396 30660 53790
rect 30604 53330 30660 53340
rect 30380 52658 30436 52668
rect 30604 52722 30660 52734
rect 30604 52670 30606 52722
rect 30658 52670 30660 52722
rect 30268 52210 30324 52220
rect 30604 52276 30660 52670
rect 30604 52210 30660 52220
rect 30268 51156 30324 51166
rect 30268 51062 30324 51100
rect 30604 51156 30660 51166
rect 30604 51062 30660 51100
rect 30604 50706 30660 50718
rect 30604 50654 30606 50706
rect 30658 50654 30660 50706
rect 30380 50594 30436 50606
rect 30380 50542 30382 50594
rect 30434 50542 30436 50594
rect 30380 49140 30436 50542
rect 30604 50036 30660 50654
rect 30604 49970 30660 49980
rect 30380 49074 30436 49084
rect 30492 49700 30548 49710
rect 30044 48290 30100 48300
rect 30268 49026 30324 49038
rect 30268 48974 30270 49026
rect 30322 48974 30324 49026
rect 30268 48244 30324 48974
rect 30268 48178 30324 48188
rect 28812 48066 28868 48076
rect 30268 48020 30324 48030
rect 30268 47926 30324 47964
rect 30268 47460 30324 47470
rect 30268 47366 30324 47404
rect 30268 45892 30324 45902
rect 29820 45890 30324 45892
rect 29820 45838 30270 45890
rect 30322 45838 30324 45890
rect 29820 45836 30324 45838
rect 29708 45332 29764 45342
rect 29484 44884 29540 44894
rect 29484 44790 29540 44828
rect 29596 44322 29652 44334
rect 29596 44270 29598 44322
rect 29650 44270 29652 44322
rect 29484 43316 29540 43326
rect 29148 43314 29540 43316
rect 29148 43262 29486 43314
rect 29538 43262 29540 43314
rect 29148 43260 29540 43262
rect 29148 29204 29204 43260
rect 29484 43250 29540 43260
rect 29484 41748 29540 41758
rect 29372 41746 29540 41748
rect 29372 41694 29486 41746
rect 29538 41694 29540 41746
rect 29372 41692 29540 41694
rect 29372 30772 29428 41692
rect 29484 41682 29540 41692
rect 29484 41186 29540 41198
rect 29484 41134 29486 41186
rect 29538 41134 29540 41186
rect 29484 40516 29540 41134
rect 29484 40450 29540 40460
rect 29484 40178 29540 40190
rect 29484 40126 29486 40178
rect 29538 40126 29540 40178
rect 29484 39508 29540 40126
rect 29484 39442 29540 39452
rect 29484 38052 29540 38062
rect 29484 35588 29540 37996
rect 29596 36708 29652 44270
rect 29596 36642 29652 36652
rect 29708 35700 29764 45276
rect 29820 44994 29876 45836
rect 30268 45826 30324 45836
rect 29820 44942 29822 44994
rect 29874 44942 29876 44994
rect 29820 44930 29876 44942
rect 30268 44884 30324 44894
rect 29932 44882 30324 44884
rect 29932 44830 30270 44882
rect 30322 44830 30324 44882
rect 29932 44828 30324 44830
rect 29820 44548 29876 44558
rect 29932 44548 29988 44828
rect 30268 44818 30324 44828
rect 29820 44546 29988 44548
rect 29820 44494 29822 44546
rect 29874 44494 29988 44546
rect 29820 44492 29988 44494
rect 29820 44482 29876 44492
rect 29820 43316 29876 43326
rect 30268 43316 30324 43326
rect 29820 43314 30324 43316
rect 29820 43262 29822 43314
rect 29874 43262 30270 43314
rect 30322 43262 30324 43314
rect 29820 43260 30324 43262
rect 29820 43250 29876 43260
rect 30268 43250 30324 43260
rect 30380 42868 30436 42878
rect 30268 42756 30324 42766
rect 29820 42754 30324 42756
rect 29820 42702 30270 42754
rect 30322 42702 30324 42754
rect 29820 42700 30324 42702
rect 29820 41858 29876 42700
rect 30268 42690 30324 42700
rect 29820 41806 29822 41858
rect 29874 41806 29876 41858
rect 29820 41794 29876 41806
rect 29820 41300 29876 41310
rect 30268 41300 30324 41310
rect 29820 41298 30324 41300
rect 29820 41246 29822 41298
rect 29874 41246 30270 41298
rect 30322 41246 30324 41298
rect 29820 41244 30324 41246
rect 29820 41234 29876 41244
rect 30268 41234 30324 41244
rect 30268 40404 30324 40414
rect 29820 40402 30324 40404
rect 29820 40350 30270 40402
rect 30322 40350 30324 40402
rect 29820 40348 30324 40350
rect 29820 40290 29876 40348
rect 30268 40338 30324 40348
rect 29820 40238 29822 40290
rect 29874 40238 29876 40290
rect 29820 40226 29876 40238
rect 30268 36596 30324 36606
rect 29708 35644 30212 35700
rect 29484 35532 29876 35588
rect 29596 33234 29652 33246
rect 29596 33182 29598 33234
rect 29650 33182 29652 33234
rect 29596 32676 29652 33182
rect 29596 32610 29652 32620
rect 29708 33122 29764 33134
rect 29708 33070 29710 33122
rect 29762 33070 29764 33122
rect 29708 31948 29764 33070
rect 29372 30706 29428 30716
rect 29484 31892 29764 31948
rect 29148 29138 29204 29148
rect 29484 25060 29540 31892
rect 29596 27860 29652 27870
rect 29596 27766 29652 27804
rect 29708 27748 29764 27758
rect 29708 27654 29764 27692
rect 29820 27300 29876 35532
rect 30156 32004 30212 35644
rect 30268 35698 30324 36540
rect 30268 35646 30270 35698
rect 30322 35646 30324 35698
rect 30268 35634 30324 35646
rect 30268 35140 30324 35150
rect 30268 35046 30324 35084
rect 30268 34356 30324 34366
rect 30268 34130 30324 34300
rect 30268 34078 30270 34130
rect 30322 34078 30324 34130
rect 30268 34066 30324 34078
rect 30380 33908 30436 42812
rect 30268 33852 30436 33908
rect 30268 33124 30324 33852
rect 30380 33348 30436 33358
rect 30492 33348 30548 49644
rect 30604 49138 30660 49150
rect 30604 49086 30606 49138
rect 30658 49086 30660 49138
rect 30604 48916 30660 49086
rect 30604 48850 30660 48860
rect 30604 48018 30660 48030
rect 30604 47966 30606 48018
rect 30658 47966 30660 48018
rect 30604 47796 30660 47966
rect 30604 47730 30660 47740
rect 30604 47570 30660 47582
rect 30604 47518 30606 47570
rect 30658 47518 30660 47570
rect 30604 46676 30660 47518
rect 30604 46610 30660 46620
rect 30604 46002 30660 46014
rect 30604 45950 30606 46002
rect 30658 45950 30660 46002
rect 30604 45556 30660 45950
rect 30604 45490 30660 45500
rect 30604 44882 30660 44894
rect 30604 44830 30606 44882
rect 30658 44830 30660 44882
rect 30604 44436 30660 44830
rect 30604 44370 30660 44380
rect 30604 43316 30660 43326
rect 30604 43222 30660 43260
rect 30604 42866 30660 42878
rect 30604 42814 30606 42866
rect 30658 42814 30660 42866
rect 30604 42196 30660 42814
rect 30604 42130 30660 42140
rect 30604 41298 30660 41310
rect 30604 41246 30606 41298
rect 30658 41246 30660 41298
rect 30604 41076 30660 41246
rect 30604 41010 30660 41020
rect 30604 40178 30660 40190
rect 30604 40126 30606 40178
rect 30658 40126 30660 40178
rect 30604 39956 30660 40126
rect 30604 39890 30660 39900
rect 31276 37828 31332 37838
rect 30604 35474 30660 35486
rect 30604 35422 30606 35474
rect 30658 35422 30660 35474
rect 30604 35252 30660 35422
rect 30604 35186 30660 35196
rect 30604 35026 30660 35038
rect 30604 34974 30606 35026
rect 30658 34974 30660 35026
rect 30604 34356 30660 34974
rect 30604 34290 30660 34300
rect 30604 33908 30660 33918
rect 30604 33906 30772 33908
rect 30604 33854 30606 33906
rect 30658 33854 30772 33906
rect 30604 33852 30772 33854
rect 30604 33842 30660 33852
rect 30380 33346 30548 33348
rect 30380 33294 30382 33346
rect 30434 33294 30548 33346
rect 30380 33292 30548 33294
rect 30604 33458 30660 33470
rect 30604 33406 30606 33458
rect 30658 33406 30660 33458
rect 30380 33282 30436 33292
rect 30268 33068 30548 33124
rect 30380 32900 30436 32910
rect 30268 32004 30324 32014
rect 30156 32002 30324 32004
rect 30156 31950 30270 32002
rect 30322 31950 30324 32002
rect 30156 31948 30324 31950
rect 30268 31938 30324 31948
rect 30380 30994 30436 32844
rect 30380 30942 30382 30994
rect 30434 30942 30436 30994
rect 30380 30930 30436 30942
rect 30156 30884 30212 30894
rect 30156 29428 30212 30828
rect 30268 30212 30324 30222
rect 30268 30118 30324 30156
rect 30268 29428 30324 29438
rect 30156 29426 30324 29428
rect 30156 29374 30270 29426
rect 30322 29374 30324 29426
rect 30156 29372 30324 29374
rect 30268 29362 30324 29372
rect 30268 28756 30324 28766
rect 30268 28662 30324 28700
rect 30268 27972 30324 27982
rect 30268 27858 30324 27916
rect 30268 27806 30270 27858
rect 30322 27806 30324 27858
rect 30268 27794 30324 27806
rect 30268 27300 30324 27310
rect 29820 27298 30324 27300
rect 29820 27246 30270 27298
rect 30322 27246 30324 27298
rect 29820 27244 30324 27246
rect 30268 27234 30324 27244
rect 30268 25732 30324 25742
rect 30268 25638 30324 25676
rect 30492 25284 30548 33068
rect 30604 32564 30660 33406
rect 30716 33460 30772 33852
rect 30716 33394 30772 33404
rect 30604 32498 30660 32508
rect 30604 31890 30660 31902
rect 30604 31838 30606 31890
rect 30658 31838 30660 31890
rect 30604 31668 30660 31838
rect 30604 31602 30660 31612
rect 30604 30772 30660 30782
rect 30604 30678 30660 30716
rect 30604 30322 30660 30334
rect 30604 30270 30606 30322
rect 30658 30270 30660 30322
rect 30604 29876 30660 30270
rect 30604 29810 30660 29820
rect 30604 29202 30660 29214
rect 30604 29150 30606 29202
rect 30658 29150 30660 29202
rect 30604 28980 30660 29150
rect 30604 28914 30660 28924
rect 30604 28754 30660 28766
rect 30604 28702 30606 28754
rect 30658 28702 30660 28754
rect 30604 28084 30660 28702
rect 30604 28018 30660 28028
rect 30604 27636 30660 27646
rect 30604 27634 30772 27636
rect 30604 27582 30606 27634
rect 30658 27582 30772 27634
rect 30604 27580 30772 27582
rect 30604 27570 30660 27580
rect 30604 27186 30660 27198
rect 30604 27134 30606 27186
rect 30658 27134 30660 27186
rect 30604 26292 30660 27134
rect 30716 27188 30772 27580
rect 30716 27122 30772 27132
rect 30604 26226 30660 26236
rect 30604 25618 30660 25630
rect 30604 25566 30606 25618
rect 30658 25566 30660 25618
rect 30604 25396 30660 25566
rect 30604 25330 30660 25340
rect 29484 24994 29540 25004
rect 30380 25228 30548 25284
rect 30268 24724 30324 24734
rect 30268 24630 30324 24668
rect 30268 24052 30324 24062
rect 30268 23958 30324 23996
rect 30268 23380 30324 23390
rect 30268 23154 30324 23324
rect 30268 23102 30270 23154
rect 30322 23102 30324 23154
rect 30268 23090 30324 23102
rect 30268 22596 30324 22606
rect 30268 22502 30324 22540
rect 30268 21364 30324 21374
rect 30156 21362 30324 21364
rect 30156 21310 30270 21362
rect 30322 21310 30324 21362
rect 30156 21308 30324 21310
rect 30156 20692 30212 21308
rect 30268 21298 30324 21308
rect 30268 20804 30324 20814
rect 30268 20710 30324 20748
rect 30156 20626 30212 20636
rect 30268 19460 30324 19470
rect 30268 19366 30324 19404
rect 30268 18452 30324 18462
rect 30268 18358 30324 18396
rect 30268 17892 30324 17902
rect 30268 17798 30324 17836
rect 30268 16660 30324 16670
rect 30156 16604 30268 16660
rect 30156 13858 30212 16604
rect 30268 16566 30324 16604
rect 30268 16324 30324 16334
rect 30268 16230 30324 16268
rect 30380 15314 30436 25228
rect 30380 15262 30382 15314
rect 30434 15262 30436 15314
rect 30380 15250 30436 15262
rect 30492 25060 30548 25070
rect 30268 14756 30324 14766
rect 30268 14662 30324 14700
rect 30156 13806 30158 13858
rect 30210 13806 30212 13858
rect 30156 13794 30212 13806
rect 30268 13188 30324 13198
rect 30268 13094 30324 13132
rect 30380 12180 30436 12190
rect 30492 12180 30548 25004
rect 30604 24500 30660 24510
rect 30604 24406 30660 24444
rect 30604 24050 30660 24062
rect 30604 23998 30606 24050
rect 30658 23998 30660 24050
rect 30604 23604 30660 23998
rect 30604 23538 30660 23548
rect 30604 22930 30660 22942
rect 30604 22878 30606 22930
rect 30658 22878 30660 22930
rect 30604 22708 30660 22878
rect 30604 22642 30660 22652
rect 30604 22482 30660 22494
rect 30604 22430 30606 22482
rect 30658 22430 30660 22482
rect 30604 21812 30660 22430
rect 30604 21746 30660 21756
rect 30604 21364 30660 21374
rect 30604 21362 30772 21364
rect 30604 21310 30606 21362
rect 30658 21310 30772 21362
rect 30604 21308 30772 21310
rect 30604 21298 30660 21308
rect 30604 20914 30660 20926
rect 30604 20862 30606 20914
rect 30658 20862 30660 20914
rect 30604 20020 30660 20862
rect 30716 20916 30772 21308
rect 30716 20850 30772 20860
rect 30604 19954 30660 19964
rect 30604 19346 30660 19358
rect 30604 19294 30606 19346
rect 30658 19294 30660 19346
rect 30604 19124 30660 19294
rect 30604 19058 30660 19068
rect 30604 18228 30660 18238
rect 30604 18134 30660 18172
rect 30604 17778 30660 17790
rect 30604 17726 30606 17778
rect 30658 17726 30660 17778
rect 30604 17332 30660 17726
rect 30604 17266 30660 17276
rect 30604 16658 30660 16670
rect 30604 16606 30606 16658
rect 30658 16606 30660 16658
rect 30604 16436 30660 16606
rect 30604 16370 30660 16380
rect 30604 16210 30660 16222
rect 30604 16158 30606 16210
rect 30658 16158 30660 16210
rect 30604 15540 30660 16158
rect 30604 15474 30660 15484
rect 30604 15092 30660 15102
rect 30604 15090 30772 15092
rect 30604 15038 30606 15090
rect 30658 15038 30772 15090
rect 30604 15036 30772 15038
rect 30604 15026 30660 15036
rect 30604 14642 30660 14654
rect 30604 14590 30606 14642
rect 30658 14590 30660 14642
rect 30604 13748 30660 14590
rect 30716 14644 30772 15036
rect 30716 14578 30772 14588
rect 30604 13682 30660 13692
rect 30604 13074 30660 13086
rect 30604 13022 30606 13074
rect 30658 13022 30660 13074
rect 30604 12852 30660 13022
rect 30604 12786 30660 12796
rect 30380 12178 30548 12180
rect 30380 12126 30382 12178
rect 30434 12126 30548 12178
rect 30380 12124 30548 12126
rect 30380 12114 30436 12124
rect 30604 11956 30660 11966
rect 30604 11862 30660 11900
rect 30268 11620 30324 11630
rect 30268 11526 30324 11564
rect 30604 11506 30660 11518
rect 30604 11454 30606 11506
rect 30658 11454 30660 11506
rect 30604 11060 30660 11454
rect 30604 10994 30660 11004
rect 27804 2158 27806 2210
rect 27858 2158 27860 2210
rect 27804 2146 27860 2158
rect 28364 8372 28532 8428
rect 27132 978 27412 980
rect 27132 926 27134 978
rect 27186 926 27412 978
rect 27132 924 27412 926
rect 27468 2098 27524 2110
rect 27468 2046 27470 2098
rect 27522 2046 27524 2098
rect 27132 914 27188 924
rect 27468 532 27524 2046
rect 28140 2098 28196 2110
rect 28140 2046 28142 2098
rect 28194 2046 28196 2098
rect 28140 1764 28196 2046
rect 28140 1698 28196 1708
rect 28364 1652 28420 8372
rect 31276 7476 31332 37772
rect 31500 27748 31556 27758
rect 31388 15316 31444 15326
rect 31388 8372 31444 15260
rect 31500 10164 31556 27692
rect 31500 10098 31556 10108
rect 31388 8306 31444 8316
rect 31276 7410 31332 7420
rect 29260 5684 29316 5694
rect 28476 3332 28532 3342
rect 28476 2210 28532 3276
rect 28476 2158 28478 2210
rect 28530 2158 28532 2210
rect 28476 2146 28532 2158
rect 28364 1586 28420 1596
rect 28588 1428 28644 1438
rect 27692 1316 27748 1326
rect 27692 1090 27748 1260
rect 28028 1204 28084 1214
rect 28028 1110 28084 1148
rect 28588 1202 28644 1372
rect 28588 1150 28590 1202
rect 28642 1150 28644 1202
rect 28588 1138 28644 1150
rect 29260 1202 29316 5628
rect 29260 1150 29262 1202
rect 29314 1150 29316 1202
rect 29260 1138 29316 1150
rect 27692 1038 27694 1090
rect 27746 1038 27748 1090
rect 27692 1026 27748 1038
rect 28364 1092 28420 1102
rect 28364 998 28420 1036
rect 27468 466 27524 476
rect 29036 978 29092 990
rect 29036 926 29038 978
rect 29090 926 29092 978
rect 29036 308 29092 926
rect 29036 242 29092 252
rect 26796 130 26852 140
rect 26460 18 26516 28
<< via2 >>
rect 140 114156 196 114212
rect 4844 114156 4900 114212
rect 1932 113932 1988 113988
rect 812 113708 868 113764
rect 588 111916 644 111972
rect 588 110908 644 110964
rect 1484 113538 1540 113540
rect 1484 113486 1486 113538
rect 1486 113486 1538 113538
rect 1538 113486 1540 113538
rect 1484 113484 1540 113486
rect 1260 113314 1316 113316
rect 1260 113262 1262 113314
rect 1262 113262 1314 113314
rect 1314 113262 1316 113314
rect 1260 113260 1316 113262
rect 1484 113148 1540 113204
rect 812 111804 868 111860
rect 476 108332 532 108388
rect 364 106204 420 106260
rect 140 96460 196 96516
rect 252 99932 308 99988
rect 140 85708 196 85764
rect 252 83692 308 83748
rect 476 97804 532 97860
rect 476 92764 532 92820
rect 588 100492 644 100548
rect 1820 112306 1876 112308
rect 1820 112254 1822 112306
rect 1822 112254 1874 112306
rect 1874 112254 1876 112306
rect 1820 112252 1876 112254
rect 1708 112140 1764 112196
rect 1596 111858 1652 111860
rect 1596 111806 1598 111858
rect 1598 111806 1650 111858
rect 1650 111806 1652 111858
rect 1596 111804 1652 111806
rect 1260 111634 1316 111636
rect 1260 111582 1262 111634
rect 1262 111582 1314 111634
rect 1314 111582 1316 111634
rect 1260 111580 1316 111582
rect 1484 111468 1540 111524
rect 1148 109452 1204 109508
rect 1484 110796 1540 110852
rect 1260 107996 1316 108052
rect 924 104860 980 104916
rect 1596 110908 1652 110964
rect 4464 113706 4520 113708
rect 4464 113654 4466 113706
rect 4466 113654 4518 113706
rect 4518 113654 4520 113706
rect 4464 113652 4520 113654
rect 4568 113706 4624 113708
rect 4568 113654 4570 113706
rect 4570 113654 4622 113706
rect 4622 113654 4624 113706
rect 4568 113652 4624 113654
rect 4672 113706 4728 113708
rect 4672 113654 4674 113706
rect 4674 113654 4726 113706
rect 4726 113654 4728 113706
rect 4672 113652 4728 113654
rect 5404 113820 5460 113876
rect 5180 113596 5236 113652
rect 1596 107324 1652 107380
rect 1372 106540 1428 106596
rect 1260 106258 1316 106260
rect 1260 106206 1262 106258
rect 1262 106206 1314 106258
rect 1314 106206 1316 106258
rect 1260 106204 1316 106206
rect 1036 103180 1092 103236
rect 812 102172 868 102228
rect 1036 102844 1092 102900
rect 700 98476 756 98532
rect 1148 102284 1204 102340
rect 1260 104860 1316 104916
rect 1372 104524 1428 104580
rect 1372 103906 1428 103908
rect 1372 103854 1374 103906
rect 1374 103854 1426 103906
rect 1426 103854 1428 103906
rect 1372 103852 1428 103854
rect 1036 101164 1092 101220
rect 1260 100716 1316 100772
rect 1260 100546 1316 100548
rect 1260 100494 1262 100546
rect 1262 100494 1314 100546
rect 1314 100494 1316 100546
rect 1260 100492 1316 100494
rect 1260 99986 1316 99988
rect 1260 99934 1262 99986
rect 1262 99934 1314 99986
rect 1314 99934 1316 99986
rect 1260 99932 1316 99934
rect 1372 98812 1428 98868
rect 588 90636 644 90692
rect 364 83244 420 83300
rect 588 90300 644 90356
rect 1036 92652 1092 92708
rect 1260 96236 1316 96292
rect 1260 94556 1316 94612
rect 812 91196 868 91252
rect 1596 106540 1652 106596
rect 1820 109676 1876 109732
rect 1820 106204 1876 106260
rect 1932 106316 1988 106372
rect 1596 104636 1652 104692
rect 1708 104578 1764 104580
rect 1708 104526 1710 104578
rect 1710 104526 1762 104578
rect 1762 104526 1764 104578
rect 1708 104524 1764 104526
rect 1596 104018 1652 104020
rect 1596 103966 1598 104018
rect 1598 103966 1650 104018
rect 1650 103966 1652 104018
rect 1596 103964 1652 103966
rect 1596 102732 1652 102788
rect 2268 109004 2324 109060
rect 2716 111580 2772 111636
rect 2828 110908 2884 110964
rect 2268 107660 2324 107716
rect 2380 106876 2436 106932
rect 2156 106428 2212 106484
rect 2380 106428 2436 106484
rect 2156 106258 2212 106260
rect 2156 106206 2158 106258
rect 2158 106206 2210 106258
rect 2210 106206 2212 106258
rect 2156 106204 2212 106206
rect 2156 105868 2212 105924
rect 2044 105420 2100 105476
rect 2156 104076 2212 104132
rect 1708 102450 1764 102452
rect 1708 102398 1710 102450
rect 1710 102398 1762 102450
rect 1762 102398 1764 102450
rect 1708 102396 1764 102398
rect 1932 103404 1988 103460
rect 2156 99596 2212 99652
rect 2380 102844 2436 102900
rect 2380 100994 2436 100996
rect 2380 100942 2382 100994
rect 2382 100942 2434 100994
rect 2434 100942 2436 100994
rect 2380 100940 2436 100942
rect 2268 98812 2324 98868
rect 2380 100716 2436 100772
rect 2380 98588 2436 98644
rect 2380 98252 2436 98308
rect 2268 98194 2324 98196
rect 2268 98142 2270 98194
rect 2270 98142 2322 98194
rect 2322 98142 2324 98194
rect 2268 98140 2324 98142
rect 1708 97858 1764 97860
rect 1708 97806 1710 97858
rect 1710 97806 1762 97858
rect 1762 97806 1764 97858
rect 1708 97804 1764 97806
rect 2156 96908 2212 96964
rect 1596 96796 1652 96852
rect 2156 96348 2212 96404
rect 1708 96178 1764 96180
rect 1708 96126 1710 96178
rect 1710 96126 1762 96178
rect 1762 96126 1764 96178
rect 1708 96124 1764 96126
rect 1484 95788 1540 95844
rect 1708 95900 1764 95956
rect 1484 95282 1540 95284
rect 1484 95230 1486 95282
rect 1486 95230 1538 95282
rect 1538 95230 1540 95282
rect 1484 95228 1540 95230
rect 1484 94332 1540 94388
rect 1596 92988 1652 93044
rect 1260 91250 1316 91252
rect 1260 91198 1262 91250
rect 1262 91198 1314 91250
rect 1314 91198 1316 91250
rect 1260 91196 1316 91198
rect 1148 90354 1204 90356
rect 1148 90302 1150 90354
rect 1150 90302 1202 90354
rect 1202 90302 1204 90354
rect 1148 90300 1204 90302
rect 1036 88956 1092 89012
rect 1148 90076 1204 90132
rect 1148 87164 1204 87220
rect 700 86716 756 86772
rect 1036 85762 1092 85764
rect 1036 85710 1038 85762
rect 1038 85710 1090 85762
rect 1090 85710 1092 85762
rect 1036 85708 1092 85710
rect 588 79996 644 80052
rect 700 85596 756 85652
rect 588 79772 644 79828
rect 1484 91196 1540 91252
rect 1484 90636 1540 90692
rect 1932 95676 1988 95732
rect 1820 94668 1876 94724
rect 1932 94444 1988 94500
rect 2156 94332 2212 94388
rect 2044 94220 2100 94276
rect 2156 94108 2212 94164
rect 2044 93042 2100 93044
rect 2044 92990 2046 93042
rect 2046 92990 2098 93042
rect 2098 92990 2100 93042
rect 2044 92988 2100 92990
rect 2604 109004 2660 109060
rect 3164 113372 3220 113428
rect 5516 113426 5572 113428
rect 5516 113374 5518 113426
rect 5518 113374 5570 113426
rect 5570 113374 5572 113426
rect 5516 113372 5572 113374
rect 3164 111468 3220 111524
rect 3388 113260 3444 113316
rect 3804 112922 3860 112924
rect 3804 112870 3806 112922
rect 3806 112870 3858 112922
rect 3858 112870 3860 112922
rect 3804 112868 3860 112870
rect 3908 112922 3964 112924
rect 3908 112870 3910 112922
rect 3910 112870 3962 112922
rect 3962 112870 3964 112922
rect 3908 112868 3964 112870
rect 4012 112922 4068 112924
rect 4012 112870 4014 112922
rect 4014 112870 4066 112922
rect 4066 112870 4068 112922
rect 4012 112868 4068 112870
rect 3500 111634 3556 111636
rect 3500 111582 3502 111634
rect 3502 111582 3554 111634
rect 3554 111582 3556 111634
rect 3500 111580 3556 111582
rect 3388 110348 3444 110404
rect 2940 109676 2996 109732
rect 3276 109900 3332 109956
rect 2940 107996 2996 108052
rect 2716 106428 2772 106484
rect 2828 106204 2884 106260
rect 2940 106428 2996 106484
rect 2604 105868 2660 105924
rect 2716 106092 2772 106148
rect 2716 105196 2772 105252
rect 2604 104188 2660 104244
rect 2604 104018 2660 104020
rect 2604 103966 2606 104018
rect 2606 103966 2658 104018
rect 2658 103966 2660 104018
rect 2604 103964 2660 103966
rect 2940 102114 2996 102116
rect 2940 102062 2942 102114
rect 2942 102062 2994 102114
rect 2994 102062 2996 102114
rect 2940 102060 2996 102062
rect 2940 101724 2996 101780
rect 2828 100770 2884 100772
rect 2828 100718 2830 100770
rect 2830 100718 2882 100770
rect 2882 100718 2884 100770
rect 2828 100716 2884 100718
rect 2940 100156 2996 100212
rect 2604 98252 2660 98308
rect 2828 99484 2884 99540
rect 2828 98140 2884 98196
rect 2380 93660 2436 93716
rect 2716 96850 2772 96852
rect 2716 96798 2718 96850
rect 2718 96798 2770 96850
rect 2770 96798 2772 96850
rect 2716 96796 2772 96798
rect 2940 96348 2996 96404
rect 3804 111354 3860 111356
rect 3804 111302 3806 111354
rect 3806 111302 3858 111354
rect 3858 111302 3860 111354
rect 3804 111300 3860 111302
rect 3908 111354 3964 111356
rect 3908 111302 3910 111354
rect 3910 111302 3962 111354
rect 3962 111302 3964 111354
rect 3908 111300 3964 111302
rect 4012 111354 4068 111356
rect 4012 111302 4014 111354
rect 4014 111302 4066 111354
rect 4066 111302 4068 111354
rect 4012 111300 4068 111302
rect 3724 111020 3780 111076
rect 4060 110738 4116 110740
rect 4060 110686 4062 110738
rect 4062 110686 4114 110738
rect 4114 110686 4116 110738
rect 4060 110684 4116 110686
rect 3948 110460 4004 110516
rect 3948 110124 4004 110180
rect 3500 109340 3556 109396
rect 3804 109786 3860 109788
rect 3804 109734 3806 109786
rect 3806 109734 3858 109786
rect 3858 109734 3860 109786
rect 3804 109732 3860 109734
rect 3908 109786 3964 109788
rect 3908 109734 3910 109786
rect 3910 109734 3962 109786
rect 3962 109734 3964 109786
rect 3908 109732 3964 109734
rect 4012 109786 4068 109788
rect 4012 109734 4014 109786
rect 4014 109734 4066 109786
rect 4066 109734 4068 109786
rect 4012 109732 4068 109734
rect 4956 112588 5012 112644
rect 4844 112364 4900 112420
rect 4464 112138 4520 112140
rect 4464 112086 4466 112138
rect 4466 112086 4518 112138
rect 4518 112086 4520 112138
rect 4464 112084 4520 112086
rect 4568 112138 4624 112140
rect 4568 112086 4570 112138
rect 4570 112086 4622 112138
rect 4622 112086 4624 112138
rect 4568 112084 4624 112086
rect 4672 112138 4728 112140
rect 4672 112086 4674 112138
rect 4674 112086 4726 112138
rect 4726 112086 4728 112138
rect 4672 112084 4728 112086
rect 4284 111132 4340 111188
rect 4396 111916 4452 111972
rect 4844 111020 4900 111076
rect 4844 110684 4900 110740
rect 4464 110570 4520 110572
rect 4284 110460 4340 110516
rect 4464 110518 4466 110570
rect 4466 110518 4518 110570
rect 4518 110518 4520 110570
rect 4464 110516 4520 110518
rect 4568 110570 4624 110572
rect 4568 110518 4570 110570
rect 4570 110518 4622 110570
rect 4622 110518 4624 110570
rect 4568 110516 4624 110518
rect 4672 110570 4728 110572
rect 4672 110518 4674 110570
rect 4674 110518 4726 110570
rect 4726 110518 4728 110570
rect 4672 110516 4728 110518
rect 4284 109788 4340 109844
rect 4396 110236 4452 110292
rect 3836 109340 3892 109396
rect 3724 109282 3780 109284
rect 3724 109230 3726 109282
rect 3726 109230 3778 109282
rect 3778 109230 3780 109282
rect 3724 109228 3780 109230
rect 3612 108668 3668 108724
rect 3276 108556 3332 108612
rect 3948 108892 4004 108948
rect 4620 109564 4676 109620
rect 4172 109004 4228 109060
rect 4464 109002 4520 109004
rect 4464 108950 4466 109002
rect 4466 108950 4518 109002
rect 4518 108950 4520 109002
rect 4464 108948 4520 108950
rect 4568 109002 4624 109004
rect 4568 108950 4570 109002
rect 4570 108950 4622 109002
rect 4622 108950 4624 109002
rect 4568 108948 4624 108950
rect 4672 109002 4728 109004
rect 4672 108950 4674 109002
rect 4674 108950 4726 109002
rect 4726 108950 4728 109002
rect 4672 108948 4728 108950
rect 5516 112476 5572 112532
rect 5068 112306 5124 112308
rect 5068 112254 5070 112306
rect 5070 112254 5122 112306
rect 5122 112254 5124 112306
rect 5068 112252 5124 112254
rect 5068 111858 5124 111860
rect 5068 111806 5070 111858
rect 5070 111806 5122 111858
rect 5122 111806 5124 111858
rect 5068 111804 5124 111806
rect 5852 113820 5908 113876
rect 5852 113426 5908 113428
rect 5852 113374 5854 113426
rect 5854 113374 5906 113426
rect 5906 113374 5908 113426
rect 5852 113372 5908 113374
rect 6300 113932 6356 113988
rect 6076 113260 6132 113316
rect 6076 112812 6132 112868
rect 6300 112476 6356 112532
rect 5740 112306 5796 112308
rect 5740 112254 5742 112306
rect 5742 112254 5794 112306
rect 5794 112254 5796 112306
rect 5740 112252 5796 112254
rect 5404 111356 5460 111412
rect 5516 110962 5572 110964
rect 5516 110910 5518 110962
rect 5518 110910 5570 110962
rect 5570 110910 5572 110962
rect 5516 110908 5572 110910
rect 5404 110572 5460 110628
rect 5292 109954 5348 109956
rect 5292 109902 5294 109954
rect 5294 109902 5346 109954
rect 5346 109902 5348 109954
rect 5292 109900 5348 109902
rect 5628 110066 5684 110068
rect 5628 110014 5630 110066
rect 5630 110014 5682 110066
rect 5682 110014 5684 110066
rect 5628 110012 5684 110014
rect 5740 109900 5796 109956
rect 5404 109788 5460 109844
rect 5404 109452 5460 109508
rect 4844 108892 4900 108948
rect 4956 109340 5012 109396
rect 4060 108780 4116 108836
rect 4844 108668 4900 108724
rect 3388 108332 3444 108388
rect 3500 107996 3556 108052
rect 3500 107772 3556 107828
rect 3804 108218 3860 108220
rect 3804 108166 3806 108218
rect 3806 108166 3858 108218
rect 3858 108166 3860 108218
rect 3804 108164 3860 108166
rect 3908 108218 3964 108220
rect 3908 108166 3910 108218
rect 3910 108166 3962 108218
rect 3962 108166 3964 108218
rect 3908 108164 3964 108166
rect 4012 108218 4068 108220
rect 4012 108166 4014 108218
rect 4014 108166 4066 108218
rect 4066 108166 4068 108218
rect 4012 108164 4068 108166
rect 4620 108444 4676 108500
rect 4732 108220 4788 108276
rect 4396 107548 4452 107604
rect 4464 107434 4520 107436
rect 4464 107382 4466 107434
rect 4466 107382 4518 107434
rect 4518 107382 4520 107434
rect 4464 107380 4520 107382
rect 4568 107434 4624 107436
rect 4568 107382 4570 107434
rect 4570 107382 4622 107434
rect 4622 107382 4624 107434
rect 4568 107380 4624 107382
rect 4672 107434 4728 107436
rect 4672 107382 4674 107434
rect 4674 107382 4726 107434
rect 4726 107382 4728 107434
rect 4672 107380 4728 107382
rect 3500 107100 3556 107156
rect 3388 106764 3444 106820
rect 3276 105980 3332 106036
rect 3164 105196 3220 105252
rect 3612 106988 3668 107044
rect 4732 107042 4788 107044
rect 4732 106990 4734 107042
rect 4734 106990 4786 107042
rect 4786 106990 4788 107042
rect 4732 106988 4788 106990
rect 4620 106876 4676 106932
rect 3804 106650 3860 106652
rect 3804 106598 3806 106650
rect 3806 106598 3858 106650
rect 3858 106598 3860 106650
rect 3804 106596 3860 106598
rect 3908 106650 3964 106652
rect 3908 106598 3910 106650
rect 3910 106598 3962 106650
rect 3962 106598 3964 106650
rect 3908 106596 3964 106598
rect 4012 106650 4068 106652
rect 4012 106598 4014 106650
rect 4014 106598 4066 106650
rect 4066 106598 4068 106650
rect 4012 106596 4068 106598
rect 3612 106258 3668 106260
rect 3612 106206 3614 106258
rect 3614 106206 3666 106258
rect 3666 106206 3668 106258
rect 3612 106204 3668 106206
rect 4508 106316 4564 106372
rect 4172 105980 4228 106036
rect 4060 105756 4116 105812
rect 3836 105420 3892 105476
rect 4060 105420 4116 105476
rect 4396 105980 4452 106036
rect 4284 105868 4340 105924
rect 4464 105866 4520 105868
rect 4464 105814 4466 105866
rect 4466 105814 4518 105866
rect 4518 105814 4520 105866
rect 4464 105812 4520 105814
rect 4568 105866 4624 105868
rect 4568 105814 4570 105866
rect 4570 105814 4622 105866
rect 4622 105814 4624 105866
rect 4568 105812 4624 105814
rect 4672 105866 4728 105868
rect 4672 105814 4674 105866
rect 4674 105814 4726 105866
rect 4726 105814 4728 105866
rect 4672 105812 4728 105814
rect 4508 105196 4564 105252
rect 3804 105082 3860 105084
rect 3804 105030 3806 105082
rect 3806 105030 3858 105082
rect 3858 105030 3860 105082
rect 3804 105028 3860 105030
rect 3908 105082 3964 105084
rect 3908 105030 3910 105082
rect 3910 105030 3962 105082
rect 3962 105030 3964 105082
rect 3908 105028 3964 105030
rect 4012 105082 4068 105084
rect 4012 105030 4014 105082
rect 4014 105030 4066 105082
rect 4066 105030 4068 105082
rect 4012 105028 4068 105030
rect 4060 104748 4116 104804
rect 3724 104578 3780 104580
rect 3724 104526 3726 104578
rect 3726 104526 3778 104578
rect 3778 104526 3780 104578
rect 3724 104524 3780 104526
rect 4732 105586 4788 105588
rect 4732 105534 4734 105586
rect 4734 105534 4786 105586
rect 4786 105534 4788 105586
rect 4732 105532 4788 105534
rect 4620 104748 4676 104804
rect 4172 104412 4228 104468
rect 4172 104076 4228 104132
rect 3276 102396 3332 102452
rect 3804 103514 3860 103516
rect 3804 103462 3806 103514
rect 3806 103462 3858 103514
rect 3858 103462 3860 103514
rect 3804 103460 3860 103462
rect 3908 103514 3964 103516
rect 3908 103462 3910 103514
rect 3910 103462 3962 103514
rect 3962 103462 3964 103514
rect 3908 103460 3964 103462
rect 4012 103514 4068 103516
rect 4012 103462 4014 103514
rect 4014 103462 4066 103514
rect 4066 103462 4068 103514
rect 4012 103460 4068 103462
rect 3724 103292 3780 103348
rect 3948 103180 4004 103236
rect 3836 103068 3892 103124
rect 3836 102732 3892 102788
rect 4060 102732 4116 102788
rect 3804 101946 3860 101948
rect 3804 101894 3806 101946
rect 3806 101894 3858 101946
rect 3858 101894 3860 101946
rect 3804 101892 3860 101894
rect 3908 101946 3964 101948
rect 3908 101894 3910 101946
rect 3910 101894 3962 101946
rect 3962 101894 3964 101946
rect 3908 101892 3964 101894
rect 4012 101946 4068 101948
rect 4012 101894 4014 101946
rect 4014 101894 4066 101946
rect 4066 101894 4068 101946
rect 4012 101892 4068 101894
rect 4060 100940 4116 100996
rect 3836 100770 3892 100772
rect 3836 100718 3838 100770
rect 3838 100718 3890 100770
rect 3890 100718 3892 100770
rect 3836 100716 3892 100718
rect 3612 100492 3668 100548
rect 3804 100378 3860 100380
rect 3804 100326 3806 100378
rect 3806 100326 3858 100378
rect 3858 100326 3860 100378
rect 3804 100324 3860 100326
rect 3908 100378 3964 100380
rect 3908 100326 3910 100378
rect 3910 100326 3962 100378
rect 3962 100326 3964 100378
rect 3908 100324 3964 100326
rect 4012 100378 4068 100380
rect 4012 100326 4014 100378
rect 4014 100326 4066 100378
rect 4066 100326 4068 100378
rect 4012 100324 4068 100326
rect 4060 100044 4116 100100
rect 3164 99484 3220 99540
rect 3276 99260 3332 99316
rect 3164 99202 3220 99204
rect 3164 99150 3166 99202
rect 3166 99150 3218 99202
rect 3218 99150 3220 99202
rect 3164 99148 3220 99150
rect 3612 99596 3668 99652
rect 3164 96236 3220 96292
rect 2716 95900 2772 95956
rect 2828 95228 2884 95284
rect 2716 95116 2772 95172
rect 2268 92092 2324 92148
rect 1708 90076 1764 90132
rect 2380 91420 2436 91476
rect 1820 87554 1876 87556
rect 1820 87502 1822 87554
rect 1822 87502 1874 87554
rect 1874 87502 1876 87554
rect 1820 87500 1876 87502
rect 1708 87052 1764 87108
rect 1372 86492 1428 86548
rect 1484 86716 1540 86772
rect 1260 86268 1316 86324
rect 700 78876 756 78932
rect 812 80892 868 80948
rect 588 76972 644 77028
rect 140 76524 196 76580
rect 252 76748 308 76804
rect 28 75404 84 75460
rect 1148 84924 1204 84980
rect 1148 84028 1204 84084
rect 1596 86770 1652 86772
rect 1596 86718 1598 86770
rect 1598 86718 1650 86770
rect 1650 86718 1652 86770
rect 1596 86716 1652 86718
rect 1484 85596 1540 85652
rect 1596 86492 1652 86548
rect 1484 85372 1540 85428
rect 1372 84700 1428 84756
rect 1484 84028 1540 84084
rect 924 80780 980 80836
rect 1148 82012 1204 82068
rect 1036 80220 1092 80276
rect 1260 79436 1316 79492
rect 924 79100 980 79156
rect 1036 76748 1092 76804
rect 924 76636 980 76692
rect 924 75404 980 75460
rect 812 75180 868 75236
rect 140 69356 196 69412
rect 252 74172 308 74228
rect 140 68012 196 68068
rect 140 67788 196 67844
rect 252 66668 308 66724
rect 364 68348 420 68404
rect 140 63084 196 63140
rect 252 65996 308 66052
rect 364 62636 420 62692
rect 476 67900 532 67956
rect 1036 74226 1092 74228
rect 1036 74174 1038 74226
rect 1038 74174 1090 74226
rect 1090 74174 1092 74226
rect 1036 74172 1092 74174
rect 1260 78146 1316 78148
rect 1260 78094 1262 78146
rect 1262 78094 1314 78146
rect 1314 78094 1316 78146
rect 1260 78092 1316 78094
rect 1932 86268 1988 86324
rect 1820 84978 1876 84980
rect 1820 84926 1822 84978
rect 1822 84926 1874 84978
rect 1874 84926 1876 84978
rect 1820 84924 1876 84926
rect 2156 87330 2212 87332
rect 2156 87278 2158 87330
rect 2158 87278 2210 87330
rect 2210 87278 2212 87330
rect 2156 87276 2212 87278
rect 2268 89180 2324 89236
rect 2044 85372 2100 85428
rect 2044 85036 2100 85092
rect 1820 83692 1876 83748
rect 1932 83356 1988 83412
rect 1708 82684 1764 82740
rect 1484 82012 1540 82068
rect 1484 78988 1540 79044
rect 1596 82236 1652 82292
rect 1372 76242 1428 76244
rect 1372 76190 1374 76242
rect 1374 76190 1426 76242
rect 1426 76190 1428 76242
rect 1372 76188 1428 76190
rect 1484 75852 1540 75908
rect 1260 75628 1316 75684
rect 1260 75404 1316 75460
rect 1372 74114 1428 74116
rect 1372 74062 1374 74114
rect 1374 74062 1426 74114
rect 1426 74062 1428 74114
rect 1372 74060 1428 74062
rect 1260 73948 1316 74004
rect 1148 72380 1204 72436
rect 588 67116 644 67172
rect 476 62188 532 62244
rect 588 66780 644 66836
rect 700 65772 756 65828
rect 924 70476 980 70532
rect 1036 68572 1092 68628
rect 1036 68402 1092 68404
rect 1036 68350 1038 68402
rect 1038 68350 1090 68402
rect 1090 68350 1092 68402
rect 1036 68348 1092 68350
rect 1036 67954 1092 67956
rect 1036 67902 1038 67954
rect 1038 67902 1090 67954
rect 1090 67902 1092 67954
rect 1036 67900 1092 67902
rect 1260 71484 1316 71540
rect 1484 71036 1540 71092
rect 1372 70700 1428 70756
rect 1260 70588 1316 70644
rect 1484 70588 1540 70644
rect 1260 70364 1316 70420
rect 1372 69410 1428 69412
rect 1372 69358 1374 69410
rect 1374 69358 1426 69410
rect 1426 69358 1428 69410
rect 1372 69356 1428 69358
rect 1260 69244 1316 69300
rect 2268 85260 2324 85316
rect 2380 85372 2436 85428
rect 2268 84924 2324 84980
rect 2156 84082 2212 84084
rect 2156 84030 2158 84082
rect 2158 84030 2210 84082
rect 2210 84030 2212 84082
rect 2156 84028 2212 84030
rect 2828 91420 2884 91476
rect 2716 91084 2772 91140
rect 2716 90076 2772 90132
rect 2604 89570 2660 89572
rect 2604 89518 2606 89570
rect 2606 89518 2658 89570
rect 2658 89518 2660 89570
rect 2604 89516 2660 89518
rect 2716 89180 2772 89236
rect 2604 89010 2660 89012
rect 2604 88958 2606 89010
rect 2606 88958 2658 89010
rect 2658 88958 2660 89010
rect 2604 88956 2660 88958
rect 3052 91084 3108 91140
rect 3836 98924 3892 98980
rect 3804 98810 3860 98812
rect 3804 98758 3806 98810
rect 3806 98758 3858 98810
rect 3858 98758 3860 98810
rect 3804 98756 3860 98758
rect 3908 98810 3964 98812
rect 3908 98758 3910 98810
rect 3910 98758 3962 98810
rect 3962 98758 3964 98810
rect 3908 98756 3964 98758
rect 4012 98810 4068 98812
rect 4012 98758 4014 98810
rect 4014 98758 4066 98810
rect 4066 98758 4068 98810
rect 4012 98756 4068 98758
rect 4464 104298 4520 104300
rect 4464 104246 4466 104298
rect 4466 104246 4518 104298
rect 4518 104246 4520 104298
rect 4464 104244 4520 104246
rect 4568 104298 4624 104300
rect 4568 104246 4570 104298
rect 4570 104246 4622 104298
rect 4622 104246 4624 104298
rect 4568 104244 4624 104246
rect 4672 104298 4728 104300
rect 4672 104246 4674 104298
rect 4674 104246 4726 104298
rect 4726 104246 4728 104298
rect 4672 104244 4728 104246
rect 4844 104188 4900 104244
rect 4396 103794 4452 103796
rect 4396 103742 4398 103794
rect 4398 103742 4450 103794
rect 4450 103742 4452 103794
rect 4396 103740 4452 103742
rect 4396 103010 4452 103012
rect 4396 102958 4398 103010
rect 4398 102958 4450 103010
rect 4450 102958 4452 103010
rect 4396 102956 4452 102958
rect 4732 102844 4788 102900
rect 4464 102730 4520 102732
rect 4464 102678 4466 102730
rect 4466 102678 4518 102730
rect 4518 102678 4520 102730
rect 4464 102676 4520 102678
rect 4568 102730 4624 102732
rect 4568 102678 4570 102730
rect 4570 102678 4622 102730
rect 4622 102678 4624 102730
rect 4568 102676 4624 102678
rect 4672 102730 4728 102732
rect 4672 102678 4674 102730
rect 4674 102678 4726 102730
rect 4726 102678 4728 102730
rect 4672 102676 4728 102678
rect 4396 101442 4452 101444
rect 4396 101390 4398 101442
rect 4398 101390 4450 101442
rect 4450 101390 4452 101442
rect 4396 101388 4452 101390
rect 4844 101388 4900 101444
rect 4464 101162 4520 101164
rect 4464 101110 4466 101162
rect 4466 101110 4518 101162
rect 4518 101110 4520 101162
rect 4464 101108 4520 101110
rect 4568 101162 4624 101164
rect 4568 101110 4570 101162
rect 4570 101110 4622 101162
rect 4622 101110 4624 101162
rect 4568 101108 4624 101110
rect 4672 101162 4728 101164
rect 4672 101110 4674 101162
rect 4674 101110 4726 101162
rect 4726 101110 4728 101162
rect 4672 101108 4728 101110
rect 4732 99820 4788 99876
rect 4464 99594 4520 99596
rect 4464 99542 4466 99594
rect 4466 99542 4518 99594
rect 4518 99542 4520 99594
rect 4464 99540 4520 99542
rect 4568 99594 4624 99596
rect 4568 99542 4570 99594
rect 4570 99542 4622 99594
rect 4622 99542 4624 99594
rect 4568 99540 4624 99542
rect 4672 99594 4728 99596
rect 4672 99542 4674 99594
rect 4674 99542 4726 99594
rect 4726 99542 4728 99594
rect 4672 99540 4728 99542
rect 4284 99372 4340 99428
rect 4396 99314 4452 99316
rect 4396 99262 4398 99314
rect 4398 99262 4450 99314
rect 4450 99262 4452 99314
rect 4396 99260 4452 99262
rect 4284 98924 4340 98980
rect 4172 98306 4228 98308
rect 4172 98254 4174 98306
rect 4174 98254 4226 98306
rect 4226 98254 4228 98306
rect 4172 98252 4228 98254
rect 4396 98700 4452 98756
rect 4732 98364 4788 98420
rect 4396 98252 4452 98308
rect 5740 109282 5796 109284
rect 5740 109230 5742 109282
rect 5742 109230 5794 109282
rect 5794 109230 5796 109282
rect 5740 109228 5796 109230
rect 5292 109116 5348 109172
rect 5068 108780 5124 108836
rect 5180 107826 5236 107828
rect 5180 107774 5182 107826
rect 5182 107774 5234 107826
rect 5234 107774 5236 107826
rect 5180 107772 5236 107774
rect 5628 108610 5684 108612
rect 5628 108558 5630 108610
rect 5630 108558 5682 108610
rect 5682 108558 5684 108610
rect 5628 108556 5684 108558
rect 5516 107884 5572 107940
rect 5404 107154 5460 107156
rect 5404 107102 5406 107154
rect 5406 107102 5458 107154
rect 5458 107102 5460 107154
rect 5404 107100 5460 107102
rect 5740 107884 5796 107940
rect 5068 103292 5124 103348
rect 5068 102396 5124 102452
rect 6636 113036 6692 113092
rect 5516 106652 5572 106708
rect 5292 105196 5348 105252
rect 5404 106540 5460 106596
rect 5292 104972 5348 105028
rect 5292 102898 5348 102900
rect 5292 102846 5294 102898
rect 5294 102846 5346 102898
rect 5346 102846 5348 102898
rect 5292 102844 5348 102846
rect 5516 106092 5572 106148
rect 5404 102508 5460 102564
rect 5516 105196 5572 105252
rect 5292 101948 5348 102004
rect 5180 101836 5236 101892
rect 5404 101442 5460 101444
rect 5404 101390 5406 101442
rect 5406 101390 5458 101442
rect 5458 101390 5460 101442
rect 5404 101388 5460 101390
rect 5292 101276 5348 101332
rect 5740 105868 5796 105924
rect 5740 103516 5796 103572
rect 5740 103292 5796 103348
rect 6860 112476 6916 112532
rect 6188 110460 6244 110516
rect 6412 111132 6468 111188
rect 6860 110962 6916 110964
rect 6860 110910 6862 110962
rect 6862 110910 6914 110962
rect 6914 110910 6916 110962
rect 6860 110908 6916 110910
rect 6412 110460 6468 110516
rect 6412 110124 6468 110180
rect 6076 108220 6132 108276
rect 6636 110460 6692 110516
rect 6636 109900 6692 109956
rect 6300 108108 6356 108164
rect 6076 107436 6132 107492
rect 5628 102898 5684 102900
rect 5628 102846 5630 102898
rect 5630 102846 5682 102898
rect 5682 102846 5684 102898
rect 5628 102844 5684 102846
rect 6300 107938 6356 107940
rect 6300 107886 6302 107938
rect 6302 107886 6354 107938
rect 6354 107886 6356 107938
rect 6300 107884 6356 107886
rect 6076 104188 6132 104244
rect 5964 103964 6020 104020
rect 6300 106540 6356 106596
rect 6412 107548 6468 107604
rect 6412 103964 6468 104020
rect 6300 103292 6356 103348
rect 6188 103068 6244 103124
rect 6412 102620 6468 102676
rect 5740 101388 5796 101444
rect 5852 102396 5908 102452
rect 5852 102172 5908 102228
rect 6748 108668 6804 108724
rect 6860 108556 6916 108612
rect 6748 106652 6804 106708
rect 6636 105868 6692 105924
rect 7084 113148 7140 113204
rect 7420 112924 7476 112980
rect 7196 112588 7252 112644
rect 7084 109340 7140 109396
rect 7084 108780 7140 108836
rect 7196 108444 7252 108500
rect 7084 107660 7140 107716
rect 6972 106034 7028 106036
rect 6972 105982 6974 106034
rect 6974 105982 7026 106034
rect 7026 105982 7028 106034
rect 6972 105980 7028 105982
rect 6972 105756 7028 105812
rect 6972 105586 7028 105588
rect 6972 105534 6974 105586
rect 6974 105534 7026 105586
rect 7026 105534 7028 105586
rect 6972 105532 7028 105534
rect 6860 104972 6916 105028
rect 6972 104524 7028 104580
rect 7308 107548 7364 107604
rect 7308 107100 7364 107156
rect 7196 106092 7252 106148
rect 7308 106876 7364 106932
rect 7644 111804 7700 111860
rect 7532 111020 7588 111076
rect 7756 111746 7812 111748
rect 7756 111694 7758 111746
rect 7758 111694 7810 111746
rect 7810 111694 7812 111746
rect 7756 111692 7812 111694
rect 8092 113484 8148 113540
rect 7980 113090 8036 113092
rect 7980 113038 7982 113090
rect 7982 113038 8034 113090
rect 8034 113038 8036 113090
rect 7980 113036 8036 113038
rect 8092 112700 8148 112756
rect 7980 112306 8036 112308
rect 7980 112254 7982 112306
rect 7982 112254 8034 112306
rect 8034 112254 8036 112306
rect 7980 112252 8036 112254
rect 7980 111468 8036 111524
rect 7980 110908 8036 110964
rect 8092 109394 8148 109396
rect 8092 109342 8094 109394
rect 8094 109342 8146 109394
rect 8146 109342 8148 109394
rect 8092 109340 8148 109342
rect 7868 108444 7924 108500
rect 7756 108108 7812 108164
rect 7868 107714 7924 107716
rect 7868 107662 7870 107714
rect 7870 107662 7922 107714
rect 7922 107662 7924 107714
rect 7868 107660 7924 107662
rect 7756 106930 7812 106932
rect 7756 106878 7758 106930
rect 7758 106878 7810 106930
rect 7810 106878 7812 106930
rect 7756 106876 7812 106878
rect 7644 106258 7700 106260
rect 7644 106206 7646 106258
rect 7646 106206 7698 106258
rect 7698 106206 7700 106258
rect 7644 106204 7700 106206
rect 7532 105980 7588 106036
rect 7420 104412 7476 104468
rect 7308 104300 7364 104356
rect 6748 103740 6804 103796
rect 6636 103628 6692 103684
rect 6748 103122 6804 103124
rect 6748 103070 6750 103122
rect 6750 103070 6802 103122
rect 6802 103070 6804 103122
rect 6748 103068 6804 103070
rect 7084 104018 7140 104020
rect 7084 103966 7086 104018
rect 7086 103966 7138 104018
rect 7138 103966 7140 104018
rect 7084 103964 7140 103966
rect 7308 103852 7364 103908
rect 6076 102284 6132 102340
rect 5516 101164 5572 101220
rect 5516 100492 5572 100548
rect 5180 100268 5236 100324
rect 5628 100380 5684 100436
rect 6076 101388 6132 101444
rect 6076 101164 6132 101220
rect 5852 99596 5908 99652
rect 5068 98812 5124 98868
rect 5180 98924 5236 98980
rect 4956 98252 5012 98308
rect 4060 97746 4116 97748
rect 4060 97694 4062 97746
rect 4062 97694 4114 97746
rect 4114 97694 4116 97746
rect 4060 97692 4116 97694
rect 4464 98026 4520 98028
rect 4464 97974 4466 98026
rect 4466 97974 4518 98026
rect 4518 97974 4520 98026
rect 4464 97972 4520 97974
rect 4568 98026 4624 98028
rect 4568 97974 4570 98026
rect 4570 97974 4622 98026
rect 4622 97974 4624 98026
rect 4568 97972 4624 97974
rect 4672 98026 4728 98028
rect 4672 97974 4674 98026
rect 4674 97974 4726 98026
rect 4726 97974 4728 98026
rect 4672 97972 4728 97974
rect 4508 97804 4564 97860
rect 3804 97242 3860 97244
rect 3804 97190 3806 97242
rect 3806 97190 3858 97242
rect 3858 97190 3860 97242
rect 3804 97188 3860 97190
rect 3908 97242 3964 97244
rect 3908 97190 3910 97242
rect 3910 97190 3962 97242
rect 3962 97190 3964 97242
rect 3908 97188 3964 97190
rect 4012 97242 4068 97244
rect 4012 97190 4014 97242
rect 4014 97190 4066 97242
rect 4066 97190 4068 97242
rect 4012 97188 4068 97190
rect 3500 96908 3556 96964
rect 4508 97468 4564 97524
rect 4844 97468 4900 97524
rect 3500 95900 3556 95956
rect 3612 95676 3668 95732
rect 3804 95674 3860 95676
rect 3804 95622 3806 95674
rect 3806 95622 3858 95674
rect 3858 95622 3860 95674
rect 3804 95620 3860 95622
rect 3908 95674 3964 95676
rect 3908 95622 3910 95674
rect 3910 95622 3962 95674
rect 3962 95622 3964 95674
rect 3908 95620 3964 95622
rect 4012 95674 4068 95676
rect 4012 95622 4014 95674
rect 4014 95622 4066 95674
rect 4066 95622 4068 95674
rect 4012 95620 4068 95622
rect 4172 95282 4228 95284
rect 4172 95230 4174 95282
rect 4174 95230 4226 95282
rect 4226 95230 4228 95282
rect 4172 95228 4228 95230
rect 4060 95116 4116 95172
rect 3388 94332 3444 94388
rect 4060 94498 4116 94500
rect 4060 94446 4062 94498
rect 4062 94446 4114 94498
rect 4114 94446 4116 94498
rect 4060 94444 4116 94446
rect 3612 93996 3668 94052
rect 3804 94106 3860 94108
rect 3804 94054 3806 94106
rect 3806 94054 3858 94106
rect 3858 94054 3860 94106
rect 3804 94052 3860 94054
rect 3908 94106 3964 94108
rect 3908 94054 3910 94106
rect 3910 94054 3962 94106
rect 3962 94054 3964 94106
rect 3908 94052 3964 94054
rect 4012 94106 4068 94108
rect 4012 94054 4014 94106
rect 4014 94054 4066 94106
rect 4066 94054 4068 94106
rect 4012 94052 4068 94054
rect 3276 93772 3332 93828
rect 3500 93772 3556 93828
rect 3948 93714 4004 93716
rect 3948 93662 3950 93714
rect 3950 93662 4002 93714
rect 4002 93662 4004 93714
rect 3948 93660 4004 93662
rect 3804 92538 3860 92540
rect 3804 92486 3806 92538
rect 3806 92486 3858 92538
rect 3858 92486 3860 92538
rect 3804 92484 3860 92486
rect 3908 92538 3964 92540
rect 3908 92486 3910 92538
rect 3910 92486 3962 92538
rect 3962 92486 3964 92538
rect 3908 92484 3964 92486
rect 4012 92538 4068 92540
rect 4012 92486 4014 92538
rect 4014 92486 4066 92538
rect 4066 92486 4068 92538
rect 4012 92484 4068 92486
rect 3276 90972 3332 91028
rect 3164 90524 3220 90580
rect 3164 89628 3220 89684
rect 3052 89516 3108 89572
rect 3164 88956 3220 89012
rect 2716 87500 2772 87556
rect 2604 87164 2660 87220
rect 2604 86828 2660 86884
rect 2716 86716 2772 86772
rect 2716 86156 2772 86212
rect 2604 85596 2660 85652
rect 2604 85090 2660 85092
rect 2604 85038 2606 85090
rect 2606 85038 2658 85090
rect 2658 85038 2660 85090
rect 2604 85036 2660 85038
rect 2492 84924 2548 84980
rect 2380 83634 2436 83636
rect 2380 83582 2382 83634
rect 2382 83582 2434 83634
rect 2434 83582 2436 83634
rect 2380 83580 2436 83582
rect 2268 82460 2324 82516
rect 2156 82236 2212 82292
rect 2044 82124 2100 82180
rect 2156 81788 2212 81844
rect 2828 85202 2884 85204
rect 2828 85150 2830 85202
rect 2830 85150 2882 85202
rect 2882 85150 2884 85202
rect 2828 85148 2884 85150
rect 2828 84306 2884 84308
rect 2828 84254 2830 84306
rect 2830 84254 2882 84306
rect 2882 84254 2884 84306
rect 2828 84252 2884 84254
rect 2828 82738 2884 82740
rect 2828 82686 2830 82738
rect 2830 82686 2882 82738
rect 2882 82686 2884 82738
rect 2828 82684 2884 82686
rect 2044 80332 2100 80388
rect 1932 79996 1988 80052
rect 1932 79436 1988 79492
rect 1708 78876 1764 78932
rect 1708 78540 1764 78596
rect 1932 78204 1988 78260
rect 1820 78092 1876 78148
rect 2044 77532 2100 77588
rect 1932 75740 1988 75796
rect 2492 80498 2548 80500
rect 2492 80446 2494 80498
rect 2494 80446 2546 80498
rect 2546 80446 2548 80498
rect 2492 80444 2548 80446
rect 2380 80386 2436 80388
rect 2380 80334 2382 80386
rect 2382 80334 2434 80386
rect 2434 80334 2436 80386
rect 2380 80332 2436 80334
rect 2156 77196 2212 77252
rect 2268 80108 2324 80164
rect 2156 76524 2212 76580
rect 2492 79324 2548 79380
rect 2380 78652 2436 78708
rect 2380 77250 2436 77252
rect 2380 77198 2382 77250
rect 2382 77198 2434 77250
rect 2434 77198 2436 77250
rect 2380 77196 2436 77198
rect 2380 76354 2436 76356
rect 2380 76302 2382 76354
rect 2382 76302 2434 76354
rect 2434 76302 2436 76354
rect 2380 76300 2436 76302
rect 2716 82236 2772 82292
rect 3276 88114 3332 88116
rect 3276 88062 3278 88114
rect 3278 88062 3330 88114
rect 3330 88062 3332 88114
rect 3276 88060 3332 88062
rect 3804 90970 3860 90972
rect 3804 90918 3806 90970
rect 3806 90918 3858 90970
rect 3858 90918 3860 90970
rect 3804 90916 3860 90918
rect 3908 90970 3964 90972
rect 3908 90918 3910 90970
rect 3910 90918 3962 90970
rect 3962 90918 3964 90970
rect 3908 90916 3964 90918
rect 4012 90970 4068 90972
rect 4012 90918 4014 90970
rect 4014 90918 4066 90970
rect 4066 90918 4068 90970
rect 4012 90916 4068 90918
rect 4060 90300 4116 90356
rect 3724 89740 3780 89796
rect 3804 89402 3860 89404
rect 3804 89350 3806 89402
rect 3806 89350 3858 89402
rect 3858 89350 3860 89402
rect 3804 89348 3860 89350
rect 3908 89402 3964 89404
rect 3908 89350 3910 89402
rect 3910 89350 3962 89402
rect 3962 89350 3964 89402
rect 3908 89348 3964 89350
rect 4012 89402 4068 89404
rect 4012 89350 4014 89402
rect 4014 89350 4066 89402
rect 4066 89350 4068 89402
rect 4012 89348 4068 89350
rect 3612 88226 3668 88228
rect 3612 88174 3614 88226
rect 3614 88174 3666 88226
rect 3666 88174 3668 88226
rect 3612 88172 3668 88174
rect 4464 96458 4520 96460
rect 4464 96406 4466 96458
rect 4466 96406 4518 96458
rect 4518 96406 4520 96458
rect 4464 96404 4520 96406
rect 4568 96458 4624 96460
rect 4568 96406 4570 96458
rect 4570 96406 4622 96458
rect 4622 96406 4624 96458
rect 4568 96404 4624 96406
rect 4672 96458 4728 96460
rect 4672 96406 4674 96458
rect 4674 96406 4726 96458
rect 4726 96406 4728 96458
rect 4672 96404 4728 96406
rect 4956 96348 5012 96404
rect 4620 95900 4676 95956
rect 4620 95116 4676 95172
rect 4464 94890 4520 94892
rect 4464 94838 4466 94890
rect 4466 94838 4518 94890
rect 4518 94838 4520 94890
rect 4464 94836 4520 94838
rect 4568 94890 4624 94892
rect 4568 94838 4570 94890
rect 4570 94838 4622 94890
rect 4622 94838 4624 94890
rect 4568 94836 4624 94838
rect 4672 94890 4728 94892
rect 4672 94838 4674 94890
rect 4674 94838 4726 94890
rect 4726 94838 4728 94890
rect 4672 94836 4728 94838
rect 4396 94668 4452 94724
rect 4844 94556 4900 94612
rect 4844 94108 4900 94164
rect 4464 93322 4520 93324
rect 4464 93270 4466 93322
rect 4466 93270 4518 93322
rect 4518 93270 4520 93322
rect 4464 93268 4520 93270
rect 4568 93322 4624 93324
rect 4568 93270 4570 93322
rect 4570 93270 4622 93322
rect 4622 93270 4624 93322
rect 4568 93268 4624 93270
rect 4672 93322 4728 93324
rect 4672 93270 4674 93322
rect 4674 93270 4726 93322
rect 4726 93270 4728 93322
rect 4672 93268 4728 93270
rect 5068 92876 5124 92932
rect 4956 92652 5012 92708
rect 4844 92428 4900 92484
rect 4464 91754 4520 91756
rect 4464 91702 4466 91754
rect 4466 91702 4518 91754
rect 4518 91702 4520 91754
rect 4464 91700 4520 91702
rect 4568 91754 4624 91756
rect 4568 91702 4570 91754
rect 4570 91702 4622 91754
rect 4622 91702 4624 91754
rect 4568 91700 4624 91702
rect 4672 91754 4728 91756
rect 4672 91702 4674 91754
rect 4674 91702 4726 91754
rect 4726 91702 4728 91754
rect 4672 91700 4728 91702
rect 4620 91474 4676 91476
rect 4620 91422 4622 91474
rect 4622 91422 4674 91474
rect 4674 91422 4676 91474
rect 4620 91420 4676 91422
rect 4464 90186 4520 90188
rect 4464 90134 4466 90186
rect 4466 90134 4518 90186
rect 4518 90134 4520 90186
rect 4464 90132 4520 90134
rect 4568 90186 4624 90188
rect 4568 90134 4570 90186
rect 4570 90134 4622 90186
rect 4622 90134 4624 90186
rect 4568 90132 4624 90134
rect 4672 90186 4728 90188
rect 4672 90134 4674 90186
rect 4674 90134 4726 90186
rect 4726 90134 4728 90186
rect 4672 90132 4728 90134
rect 4172 89068 4228 89124
rect 3724 88060 3780 88116
rect 4060 88060 4116 88116
rect 3804 87834 3860 87836
rect 3804 87782 3806 87834
rect 3806 87782 3858 87834
rect 3858 87782 3860 87834
rect 3804 87780 3860 87782
rect 3908 87834 3964 87836
rect 3908 87782 3910 87834
rect 3910 87782 3962 87834
rect 3962 87782 3964 87834
rect 3908 87780 3964 87782
rect 4012 87834 4068 87836
rect 4012 87782 4014 87834
rect 4014 87782 4066 87834
rect 4066 87782 4068 87834
rect 4012 87780 4068 87782
rect 3388 87612 3444 87668
rect 3164 85650 3220 85652
rect 3164 85598 3166 85650
rect 3166 85598 3218 85650
rect 3218 85598 3220 85650
rect 3164 85596 3220 85598
rect 3164 84476 3220 84532
rect 3500 85090 3556 85092
rect 3500 85038 3502 85090
rect 3502 85038 3554 85090
rect 3554 85038 3556 85090
rect 3500 85036 3556 85038
rect 3276 84252 3332 84308
rect 3052 82684 3108 82740
rect 3164 84028 3220 84084
rect 3052 81676 3108 81732
rect 2828 79378 2884 79380
rect 2828 79326 2830 79378
rect 2830 79326 2882 79378
rect 2882 79326 2884 79378
rect 2828 79324 2884 79326
rect 2716 78092 2772 78148
rect 2940 78652 2996 78708
rect 2716 76860 2772 76916
rect 2268 75628 2324 75684
rect 2604 76636 2660 76692
rect 2156 75516 2212 75572
rect 2268 74844 2324 74900
rect 2044 73164 2100 73220
rect 1820 72828 1876 72884
rect 2044 72716 2100 72772
rect 1820 72380 1876 72436
rect 2268 73500 2324 73556
rect 2156 72380 2212 72436
rect 2268 72604 2324 72660
rect 2044 71820 2100 71876
rect 1932 70812 1988 70868
rect 1708 70140 1764 70196
rect 1820 70588 1876 70644
rect 1708 69580 1764 69636
rect 1148 67228 1204 67284
rect 2156 71484 2212 71540
rect 2492 75516 2548 75572
rect 2492 72716 2548 72772
rect 3276 81730 3332 81732
rect 3276 81678 3278 81730
rect 3278 81678 3330 81730
rect 3330 81678 3332 81730
rect 3276 81676 3332 81678
rect 3388 81564 3444 81620
rect 3164 80108 3220 80164
rect 3388 79324 3444 79380
rect 4464 88618 4520 88620
rect 4464 88566 4466 88618
rect 4466 88566 4518 88618
rect 4518 88566 4520 88618
rect 4464 88564 4520 88566
rect 4568 88618 4624 88620
rect 4568 88566 4570 88618
rect 4570 88566 4622 88618
rect 4622 88566 4624 88618
rect 4568 88564 4624 88566
rect 4672 88618 4728 88620
rect 4672 88566 4674 88618
rect 4674 88566 4726 88618
rect 4726 88566 4728 88618
rect 4672 88564 4728 88566
rect 5292 98588 5348 98644
rect 5292 98364 5348 98420
rect 5292 98140 5348 98196
rect 5292 96460 5348 96516
rect 5964 99148 6020 99204
rect 5740 98306 5796 98308
rect 5740 98254 5742 98306
rect 5742 98254 5794 98306
rect 5794 98254 5796 98306
rect 5740 98252 5796 98254
rect 5516 96962 5572 96964
rect 5516 96910 5518 96962
rect 5518 96910 5570 96962
rect 5570 96910 5572 96962
rect 5516 96908 5572 96910
rect 6188 100492 6244 100548
rect 6188 99596 6244 99652
rect 6188 97692 6244 97748
rect 6076 97468 6132 97524
rect 5740 96460 5796 96516
rect 5292 92652 5348 92708
rect 5740 94668 5796 94724
rect 6076 95340 6132 95396
rect 6412 101500 6468 101556
rect 6412 98812 6468 98868
rect 6636 101164 6692 101220
rect 7196 102284 7252 102340
rect 8540 113708 8596 113764
rect 8316 109116 8372 109172
rect 8428 111580 8484 111636
rect 8316 106930 8372 106932
rect 8316 106878 8318 106930
rect 8318 106878 8370 106930
rect 8370 106878 8372 106930
rect 8316 106876 8372 106878
rect 8540 112252 8596 112308
rect 8988 114268 9044 114324
rect 9100 114380 9156 114436
rect 9212 114044 9268 114100
rect 9100 112306 9156 112308
rect 9100 112254 9102 112306
rect 9102 112254 9154 112306
rect 9154 112254 9156 112306
rect 9100 112252 9156 112254
rect 8764 111580 8820 111636
rect 8876 112028 8932 112084
rect 9324 112924 9380 112980
rect 9884 114716 9940 114772
rect 9660 113932 9716 113988
rect 10220 114156 10276 114212
rect 10556 114380 10612 114436
rect 10332 113596 10388 113652
rect 10220 113036 10276 113092
rect 10108 112588 10164 112644
rect 10220 112476 10276 112532
rect 9660 112028 9716 112084
rect 8876 110460 8932 110516
rect 8652 109228 8708 109284
rect 8540 106764 8596 106820
rect 8428 106204 8484 106260
rect 8092 105532 8148 105588
rect 8316 105868 8372 105924
rect 8092 104972 8148 105028
rect 8092 104412 8148 104468
rect 6636 100604 6692 100660
rect 6524 98028 6580 98084
rect 6412 97580 6468 97636
rect 6412 97244 6468 97300
rect 6524 97804 6580 97860
rect 6412 96460 6468 96516
rect 6412 96124 6468 96180
rect 6972 98700 7028 98756
rect 6860 98194 6916 98196
rect 6860 98142 6862 98194
rect 6862 98142 6914 98194
rect 6914 98142 6916 98194
rect 6860 98140 6916 98142
rect 7084 97468 7140 97524
rect 6636 96908 6692 96964
rect 6748 96066 6804 96068
rect 6748 96014 6750 96066
rect 6750 96014 6802 96066
rect 6802 96014 6804 96066
rect 6748 96012 6804 96014
rect 6636 95170 6692 95172
rect 6636 95118 6638 95170
rect 6638 95118 6690 95170
rect 6690 95118 6692 95170
rect 6636 95116 6692 95118
rect 5404 92428 5460 92484
rect 5516 93996 5572 94052
rect 4956 91420 5012 91476
rect 5404 92258 5460 92260
rect 5404 92206 5406 92258
rect 5406 92206 5458 92258
rect 5458 92206 5460 92258
rect 5404 92204 5460 92206
rect 4956 91250 5012 91252
rect 4956 91198 4958 91250
rect 4958 91198 5010 91250
rect 5010 91198 5012 91250
rect 4956 91196 5012 91198
rect 5740 93714 5796 93716
rect 5740 93662 5742 93714
rect 5742 93662 5794 93714
rect 5794 93662 5796 93714
rect 5740 93660 5796 93662
rect 5740 93436 5796 93492
rect 5628 92930 5684 92932
rect 5628 92878 5630 92930
rect 5630 92878 5682 92930
rect 5682 92878 5684 92930
rect 5628 92876 5684 92878
rect 5740 92428 5796 92484
rect 5740 91980 5796 92036
rect 5404 90188 5460 90244
rect 5068 88956 5124 89012
rect 4284 87388 4340 87444
rect 4464 87050 4520 87052
rect 4464 86998 4466 87050
rect 4466 86998 4518 87050
rect 4518 86998 4520 87050
rect 4464 86996 4520 86998
rect 4568 87050 4624 87052
rect 4568 86998 4570 87050
rect 4570 86998 4622 87050
rect 4622 86998 4624 87050
rect 4568 86996 4624 86998
rect 4672 87050 4728 87052
rect 4672 86998 4674 87050
rect 4674 86998 4726 87050
rect 4726 86998 4728 87050
rect 4672 86996 4728 86998
rect 3948 86828 4004 86884
rect 3724 86658 3780 86660
rect 3724 86606 3726 86658
rect 3726 86606 3778 86658
rect 3778 86606 3780 86658
rect 3724 86604 3780 86606
rect 3948 86492 4004 86548
rect 3804 86266 3860 86268
rect 3804 86214 3806 86266
rect 3806 86214 3858 86266
rect 3858 86214 3860 86266
rect 3804 86212 3860 86214
rect 3908 86266 3964 86268
rect 3908 86214 3910 86266
rect 3910 86214 3962 86266
rect 3962 86214 3964 86266
rect 3908 86212 3964 86214
rect 4012 86266 4068 86268
rect 4012 86214 4014 86266
rect 4014 86214 4066 86266
rect 4066 86214 4068 86266
rect 4012 86212 4068 86214
rect 3948 86044 4004 86100
rect 3836 84812 3892 84868
rect 4284 85650 4340 85652
rect 4284 85598 4286 85650
rect 4286 85598 4338 85650
rect 4338 85598 4340 85650
rect 4284 85596 4340 85598
rect 4464 85482 4520 85484
rect 4464 85430 4466 85482
rect 4466 85430 4518 85482
rect 4518 85430 4520 85482
rect 4464 85428 4520 85430
rect 4568 85482 4624 85484
rect 4568 85430 4570 85482
rect 4570 85430 4622 85482
rect 4622 85430 4624 85482
rect 4568 85428 4624 85430
rect 4672 85482 4728 85484
rect 4672 85430 4674 85482
rect 4674 85430 4726 85482
rect 4726 85430 4728 85482
rect 4672 85428 4728 85430
rect 3804 84698 3860 84700
rect 3804 84646 3806 84698
rect 3806 84646 3858 84698
rect 3858 84646 3860 84698
rect 3804 84644 3860 84646
rect 3908 84698 3964 84700
rect 3908 84646 3910 84698
rect 3910 84646 3962 84698
rect 3962 84646 3964 84698
rect 3908 84644 3964 84646
rect 4012 84698 4068 84700
rect 4012 84646 4014 84698
rect 4014 84646 4066 84698
rect 4066 84646 4068 84698
rect 4012 84644 4068 84646
rect 4172 84306 4228 84308
rect 4172 84254 4174 84306
rect 4174 84254 4226 84306
rect 4226 84254 4228 84306
rect 4172 84252 4228 84254
rect 3948 83468 4004 83524
rect 3804 83130 3860 83132
rect 3804 83078 3806 83130
rect 3806 83078 3858 83130
rect 3858 83078 3860 83130
rect 3804 83076 3860 83078
rect 3908 83130 3964 83132
rect 3908 83078 3910 83130
rect 3910 83078 3962 83130
rect 3962 83078 3964 83130
rect 3908 83076 3964 83078
rect 4012 83130 4068 83132
rect 4012 83078 4014 83130
rect 4014 83078 4066 83130
rect 4066 83078 4068 83130
rect 4012 83076 4068 83078
rect 3724 82066 3780 82068
rect 3724 82014 3726 82066
rect 3726 82014 3778 82066
rect 3778 82014 3780 82066
rect 3724 82012 3780 82014
rect 4844 84252 4900 84308
rect 4396 84028 4452 84084
rect 4464 83914 4520 83916
rect 4464 83862 4466 83914
rect 4466 83862 4518 83914
rect 4518 83862 4520 83914
rect 4464 83860 4520 83862
rect 4568 83914 4624 83916
rect 4568 83862 4570 83914
rect 4570 83862 4622 83914
rect 4622 83862 4624 83914
rect 4568 83860 4624 83862
rect 4672 83914 4728 83916
rect 4672 83862 4674 83914
rect 4674 83862 4726 83914
rect 4726 83862 4728 83914
rect 4672 83860 4728 83862
rect 5292 87948 5348 88004
rect 5740 90860 5796 90916
rect 6188 94444 6244 94500
rect 6188 93660 6244 93716
rect 5964 93324 6020 93380
rect 5964 92818 6020 92820
rect 5964 92766 5966 92818
rect 5966 92766 6018 92818
rect 6018 92766 6020 92818
rect 5964 92764 6020 92766
rect 6076 92540 6132 92596
rect 5964 92428 6020 92484
rect 6188 91420 6244 91476
rect 6188 90188 6244 90244
rect 6300 94108 6356 94164
rect 6636 92930 6692 92932
rect 6636 92878 6638 92930
rect 6638 92878 6690 92930
rect 6690 92878 6692 92930
rect 6636 92876 6692 92878
rect 6748 92540 6804 92596
rect 7084 95564 7140 95620
rect 7084 95394 7140 95396
rect 7084 95342 7086 95394
rect 7086 95342 7138 95394
rect 7138 95342 7140 95394
rect 7084 95340 7140 95342
rect 7084 94498 7140 94500
rect 7084 94446 7086 94498
rect 7086 94446 7138 94498
rect 7138 94446 7140 94498
rect 7084 94444 7140 94446
rect 6972 94220 7028 94276
rect 7084 93212 7140 93268
rect 7084 92540 7140 92596
rect 6636 92034 6692 92036
rect 6636 91982 6638 92034
rect 6638 91982 6690 92034
rect 6690 91982 6692 92034
rect 6636 91980 6692 91982
rect 6524 91868 6580 91924
rect 6524 91420 6580 91476
rect 6524 91084 6580 91140
rect 5852 89292 5908 89348
rect 6188 89292 6244 89348
rect 5404 86604 5460 86660
rect 5292 85932 5348 85988
rect 5068 83580 5124 83636
rect 3612 81676 3668 81732
rect 3804 81562 3860 81564
rect 3804 81510 3806 81562
rect 3806 81510 3858 81562
rect 3858 81510 3860 81562
rect 3804 81508 3860 81510
rect 3908 81562 3964 81564
rect 3908 81510 3910 81562
rect 3910 81510 3962 81562
rect 3962 81510 3964 81562
rect 3908 81508 3964 81510
rect 4012 81562 4068 81564
rect 4012 81510 4014 81562
rect 4014 81510 4066 81562
rect 4066 81510 4068 81562
rect 4012 81508 4068 81510
rect 4464 82346 4520 82348
rect 4464 82294 4466 82346
rect 4466 82294 4518 82346
rect 4518 82294 4520 82346
rect 4464 82292 4520 82294
rect 4568 82346 4624 82348
rect 4568 82294 4570 82346
rect 4570 82294 4622 82346
rect 4622 82294 4624 82346
rect 4568 82292 4624 82294
rect 4672 82346 4728 82348
rect 4672 82294 4674 82346
rect 4674 82294 4726 82346
rect 4726 82294 4728 82346
rect 4672 82292 4728 82294
rect 4508 81676 4564 81732
rect 4172 81228 4228 81284
rect 3948 80946 4004 80948
rect 3948 80894 3950 80946
rect 3950 80894 4002 80946
rect 4002 80894 4004 80946
rect 3948 80892 4004 80894
rect 3612 80386 3668 80388
rect 3612 80334 3614 80386
rect 3614 80334 3666 80386
rect 3666 80334 3668 80386
rect 3612 80332 3668 80334
rect 4508 80892 4564 80948
rect 5068 82012 5124 82068
rect 5404 83916 5460 83972
rect 5292 82684 5348 82740
rect 5292 82348 5348 82404
rect 4844 81452 4900 81508
rect 4464 80778 4520 80780
rect 4464 80726 4466 80778
rect 4466 80726 4518 80778
rect 4518 80726 4520 80778
rect 4464 80724 4520 80726
rect 4568 80778 4624 80780
rect 4568 80726 4570 80778
rect 4570 80726 4622 80778
rect 4622 80726 4624 80778
rect 4568 80724 4624 80726
rect 4672 80778 4728 80780
rect 4672 80726 4674 80778
rect 4674 80726 4726 80778
rect 4726 80726 4728 80778
rect 4672 80724 4728 80726
rect 3804 79994 3860 79996
rect 3804 79942 3806 79994
rect 3806 79942 3858 79994
rect 3858 79942 3860 79994
rect 3804 79940 3860 79942
rect 3908 79994 3964 79996
rect 3908 79942 3910 79994
rect 3910 79942 3962 79994
rect 3962 79942 3964 79994
rect 3908 79940 3964 79942
rect 4012 79994 4068 79996
rect 4012 79942 4014 79994
rect 4014 79942 4066 79994
rect 4066 79942 4068 79994
rect 4012 79940 4068 79942
rect 3500 78316 3556 78372
rect 4060 79100 4116 79156
rect 3948 78764 4004 78820
rect 3804 78426 3860 78428
rect 3804 78374 3806 78426
rect 3806 78374 3858 78426
rect 3858 78374 3860 78426
rect 3804 78372 3860 78374
rect 3908 78426 3964 78428
rect 3908 78374 3910 78426
rect 3910 78374 3962 78426
rect 3962 78374 3964 78426
rect 3908 78372 3964 78374
rect 4012 78426 4068 78428
rect 4012 78374 4014 78426
rect 4014 78374 4066 78426
rect 4066 78374 4068 78426
rect 4012 78372 4068 78374
rect 4172 78316 4228 78372
rect 3052 77868 3108 77924
rect 3052 77532 3108 77588
rect 3388 77868 3444 77924
rect 3276 77810 3332 77812
rect 3276 77758 3278 77810
rect 3278 77758 3330 77810
rect 3330 77758 3332 77810
rect 3276 77756 3332 77758
rect 2940 75682 2996 75684
rect 2940 75630 2942 75682
rect 2942 75630 2994 75682
rect 2994 75630 2996 75682
rect 2940 75628 2996 75630
rect 2940 74732 2996 74788
rect 3164 76860 3220 76916
rect 3164 76412 3220 76468
rect 3388 77196 3444 77252
rect 3612 77810 3668 77812
rect 3612 77758 3614 77810
rect 3614 77758 3666 77810
rect 3666 77758 3668 77810
rect 3612 77756 3668 77758
rect 4464 79210 4520 79212
rect 4464 79158 4466 79210
rect 4466 79158 4518 79210
rect 4518 79158 4520 79210
rect 4464 79156 4520 79158
rect 4568 79210 4624 79212
rect 4568 79158 4570 79210
rect 4570 79158 4622 79210
rect 4622 79158 4624 79210
rect 4568 79156 4624 79158
rect 4672 79210 4728 79212
rect 4672 79158 4674 79210
rect 4674 79158 4726 79210
rect 4726 79158 4728 79210
rect 4672 79156 4728 79158
rect 4172 77756 4228 77812
rect 5068 80668 5124 80724
rect 4956 79772 5012 79828
rect 4464 77642 4520 77644
rect 4464 77590 4466 77642
rect 4466 77590 4518 77642
rect 4518 77590 4520 77642
rect 4464 77588 4520 77590
rect 4568 77642 4624 77644
rect 4568 77590 4570 77642
rect 4570 77590 4622 77642
rect 4622 77590 4624 77642
rect 4568 77588 4624 77590
rect 4672 77642 4728 77644
rect 4672 77590 4674 77642
rect 4674 77590 4726 77642
rect 4726 77590 4728 77642
rect 4672 77588 4728 77590
rect 3948 77308 4004 77364
rect 4844 77308 4900 77364
rect 4396 77084 4452 77140
rect 4172 76972 4228 77028
rect 3804 76858 3860 76860
rect 3804 76806 3806 76858
rect 3806 76806 3858 76858
rect 3858 76806 3860 76858
rect 3804 76804 3860 76806
rect 3908 76858 3964 76860
rect 3908 76806 3910 76858
rect 3910 76806 3962 76858
rect 3962 76806 3964 76858
rect 3908 76804 3964 76806
rect 4012 76858 4068 76860
rect 4012 76806 4014 76858
rect 4014 76806 4066 76858
rect 4066 76806 4068 76858
rect 4012 76804 4068 76806
rect 2604 72492 2660 72548
rect 2940 73276 2996 73332
rect 2044 70476 2100 70532
rect 2828 72492 2884 72548
rect 2268 70978 2324 70980
rect 2268 70926 2270 70978
rect 2270 70926 2322 70978
rect 2322 70926 2324 70978
rect 2268 70924 2324 70926
rect 2044 70140 2100 70196
rect 924 66892 980 66948
rect 1148 66834 1204 66836
rect 1148 66782 1150 66834
rect 1150 66782 1202 66834
rect 1202 66782 1204 66834
rect 1148 66780 1204 66782
rect 1932 68626 1988 68628
rect 1932 68574 1934 68626
rect 1934 68574 1986 68626
rect 1986 68574 1988 68626
rect 1932 68572 1988 68574
rect 1372 68012 1428 68068
rect 1820 68066 1876 68068
rect 1820 68014 1822 68066
rect 1822 68014 1874 68066
rect 1874 68014 1876 68066
rect 1820 68012 1876 68014
rect 1820 67228 1876 67284
rect 1484 66946 1540 66948
rect 1484 66894 1486 66946
rect 1486 66894 1538 66946
rect 1538 66894 1540 66946
rect 1484 66892 1540 66894
rect 1260 66332 1316 66388
rect 812 63980 868 64036
rect 1260 64092 1316 64148
rect 588 61964 644 62020
rect 1372 63308 1428 63364
rect 1596 66444 1652 66500
rect 1820 66332 1876 66388
rect 2492 70588 2548 70644
rect 2604 70812 2660 70868
rect 2492 69916 2548 69972
rect 2156 67564 2212 67620
rect 2044 66668 2100 66724
rect 2156 66556 2212 66612
rect 2156 66220 2212 66276
rect 1932 65602 1988 65604
rect 1932 65550 1934 65602
rect 1934 65550 1986 65602
rect 1986 65550 1988 65602
rect 1932 65548 1988 65550
rect 1596 64540 1652 64596
rect 1708 63980 1764 64036
rect 1820 63084 1876 63140
rect 700 61292 756 61348
rect 700 60844 756 60900
rect 1148 62076 1204 62132
rect 2044 62354 2100 62356
rect 2044 62302 2046 62354
rect 2046 62302 2098 62354
rect 2098 62302 2100 62354
rect 2044 62300 2100 62302
rect 1932 62188 1988 62244
rect 2380 67004 2436 67060
rect 2492 66892 2548 66948
rect 2828 70812 2884 70868
rect 3052 72770 3108 72772
rect 3052 72718 3054 72770
rect 3054 72718 3106 72770
rect 3106 72718 3108 72770
rect 3052 72716 3108 72718
rect 2940 70924 2996 70980
rect 2828 69970 2884 69972
rect 2828 69918 2830 69970
rect 2830 69918 2882 69970
rect 2882 69918 2884 69970
rect 2828 69916 2884 69918
rect 3276 70700 3332 70756
rect 2940 69244 2996 69300
rect 2940 68572 2996 68628
rect 3052 66946 3108 66948
rect 3052 66894 3054 66946
rect 3054 66894 3106 66946
rect 3106 66894 3108 66946
rect 3052 66892 3108 66894
rect 2716 66332 2772 66388
rect 3052 66556 3108 66612
rect 2492 64988 2548 65044
rect 2380 63810 2436 63812
rect 2380 63758 2382 63810
rect 2382 63758 2434 63810
rect 2434 63758 2436 63810
rect 2380 63756 2436 63758
rect 812 60396 868 60452
rect 924 59948 980 60004
rect 2156 61794 2212 61796
rect 2156 61742 2158 61794
rect 2158 61742 2210 61794
rect 2210 61742 2212 61794
rect 2156 61740 2212 61742
rect 1372 61682 1428 61684
rect 1372 61630 1374 61682
rect 1374 61630 1426 61682
rect 1426 61630 1428 61682
rect 1372 61628 1428 61630
rect 1820 61682 1876 61684
rect 1820 61630 1822 61682
rect 1822 61630 1874 61682
rect 1874 61630 1876 61682
rect 1820 61628 1876 61630
rect 1484 61404 1540 61460
rect 1372 60562 1428 60564
rect 1372 60510 1374 60562
rect 1374 60510 1426 60562
rect 1426 60510 1428 60562
rect 1372 60508 1428 60510
rect 1036 59500 1092 59556
rect 1596 61292 1652 61348
rect 924 58604 980 58660
rect 2828 64988 2884 65044
rect 2716 62300 2772 62356
rect 2828 63868 2884 63924
rect 2940 63362 2996 63364
rect 2940 63310 2942 63362
rect 2942 63310 2994 63362
rect 2994 63310 2996 63362
rect 2940 63308 2996 63310
rect 2940 63084 2996 63140
rect 3948 75628 4004 75684
rect 4172 75404 4228 75460
rect 3804 75290 3860 75292
rect 3804 75238 3806 75290
rect 3806 75238 3858 75290
rect 3858 75238 3860 75290
rect 3804 75236 3860 75238
rect 3908 75290 3964 75292
rect 3908 75238 3910 75290
rect 3910 75238 3962 75290
rect 3962 75238 3964 75290
rect 3908 75236 3964 75238
rect 4012 75290 4068 75292
rect 4012 75238 4014 75290
rect 4014 75238 4066 75290
rect 4066 75238 4068 75290
rect 4012 75236 4068 75238
rect 3836 74844 3892 74900
rect 3836 74620 3892 74676
rect 4060 74508 4116 74564
rect 3948 74396 4004 74452
rect 3836 74172 3892 74228
rect 3612 73948 3668 74004
rect 3804 73722 3860 73724
rect 3804 73670 3806 73722
rect 3806 73670 3858 73722
rect 3858 73670 3860 73722
rect 3804 73668 3860 73670
rect 3908 73722 3964 73724
rect 3908 73670 3910 73722
rect 3910 73670 3962 73722
rect 3962 73670 3964 73722
rect 3908 73668 3964 73670
rect 4012 73722 4068 73724
rect 4012 73670 4014 73722
rect 4014 73670 4066 73722
rect 4066 73670 4068 73722
rect 4012 73668 4068 73670
rect 4464 76074 4520 76076
rect 4464 76022 4466 76074
rect 4466 76022 4518 76074
rect 4518 76022 4520 76074
rect 4464 76020 4520 76022
rect 4568 76074 4624 76076
rect 4568 76022 4570 76074
rect 4570 76022 4622 76074
rect 4622 76022 4624 76074
rect 4568 76020 4624 76022
rect 4672 76074 4728 76076
rect 4672 76022 4674 76074
rect 4674 76022 4726 76074
rect 4726 76022 4728 76074
rect 4672 76020 4728 76022
rect 4284 75068 4340 75124
rect 4396 74956 4452 75012
rect 4284 74844 4340 74900
rect 4464 74506 4520 74508
rect 4464 74454 4466 74506
rect 4466 74454 4518 74506
rect 4518 74454 4520 74506
rect 4464 74452 4520 74454
rect 4568 74506 4624 74508
rect 4568 74454 4570 74506
rect 4570 74454 4622 74506
rect 4622 74454 4624 74506
rect 4568 74452 4624 74454
rect 4672 74506 4728 74508
rect 4672 74454 4674 74506
rect 4674 74454 4726 74506
rect 4726 74454 4728 74506
rect 4672 74452 4728 74454
rect 4284 74060 4340 74116
rect 5068 77308 5124 77364
rect 5404 81676 5460 81732
rect 5628 84028 5684 84084
rect 5628 82796 5684 82852
rect 6860 90300 6916 90356
rect 7084 91586 7140 91588
rect 7084 91534 7086 91586
rect 7086 91534 7138 91586
rect 7138 91534 7140 91586
rect 7084 91532 7140 91534
rect 6636 89010 6692 89012
rect 6636 88958 6638 89010
rect 6638 88958 6690 89010
rect 6690 88958 6692 89010
rect 6636 88956 6692 88958
rect 6860 88898 6916 88900
rect 6860 88846 6862 88898
rect 6862 88846 6914 88898
rect 6914 88846 6916 88898
rect 6860 88844 6916 88846
rect 6300 87554 6356 87556
rect 6300 87502 6302 87554
rect 6302 87502 6354 87554
rect 6354 87502 6356 87554
rect 6300 87500 6356 87502
rect 5852 84252 5908 84308
rect 5964 84028 6020 84084
rect 6188 87276 6244 87332
rect 6188 85820 6244 85876
rect 5852 83244 5908 83300
rect 5852 82850 5908 82852
rect 5852 82798 5854 82850
rect 5854 82798 5906 82850
rect 5906 82798 5908 82850
rect 5852 82796 5908 82798
rect 5740 80668 5796 80724
rect 5852 80108 5908 80164
rect 5404 79324 5460 79380
rect 5292 77308 5348 77364
rect 5404 78316 5460 78372
rect 5404 78092 5460 78148
rect 5180 77196 5236 77252
rect 5068 76300 5124 76356
rect 4956 75404 5012 75460
rect 5068 74114 5124 74116
rect 5068 74062 5070 74114
rect 5070 74062 5122 74114
rect 5122 74062 5124 74114
rect 5068 74060 5124 74062
rect 4956 73218 5012 73220
rect 4956 73166 4958 73218
rect 4958 73166 5010 73218
rect 5010 73166 5012 73218
rect 4956 73164 5012 73166
rect 4464 72938 4520 72940
rect 4464 72886 4466 72938
rect 4466 72886 4518 72938
rect 4518 72886 4520 72938
rect 4464 72884 4520 72886
rect 4568 72938 4624 72940
rect 4568 72886 4570 72938
rect 4570 72886 4622 72938
rect 4622 72886 4624 72938
rect 4568 72884 4624 72886
rect 4672 72938 4728 72940
rect 4672 72886 4674 72938
rect 4674 72886 4726 72938
rect 4726 72886 4728 72938
rect 4672 72884 4728 72886
rect 4396 72492 4452 72548
rect 3804 72154 3860 72156
rect 3804 72102 3806 72154
rect 3806 72102 3858 72154
rect 3858 72102 3860 72154
rect 3804 72100 3860 72102
rect 3908 72154 3964 72156
rect 3908 72102 3910 72154
rect 3910 72102 3962 72154
rect 3962 72102 3964 72154
rect 3908 72100 3964 72102
rect 4012 72154 4068 72156
rect 4012 72102 4014 72154
rect 4014 72102 4066 72154
rect 4066 72102 4068 72154
rect 4012 72100 4068 72102
rect 4284 71762 4340 71764
rect 4284 71710 4286 71762
rect 4286 71710 4338 71762
rect 4338 71710 4340 71762
rect 4284 71708 4340 71710
rect 5180 73052 5236 73108
rect 5292 72716 5348 72772
rect 5068 72546 5124 72548
rect 5068 72494 5070 72546
rect 5070 72494 5122 72546
rect 5122 72494 5124 72546
rect 5068 72492 5124 72494
rect 5180 71820 5236 71876
rect 4464 71370 4520 71372
rect 4464 71318 4466 71370
rect 4466 71318 4518 71370
rect 4518 71318 4520 71370
rect 4464 71316 4520 71318
rect 4568 71370 4624 71372
rect 4568 71318 4570 71370
rect 4570 71318 4622 71370
rect 4622 71318 4624 71370
rect 4568 71316 4624 71318
rect 4672 71370 4728 71372
rect 4672 71318 4674 71370
rect 4674 71318 4726 71370
rect 4726 71318 4728 71370
rect 4672 71316 4728 71318
rect 3500 70978 3556 70980
rect 3500 70926 3502 70978
rect 3502 70926 3554 70978
rect 3554 70926 3556 70978
rect 3500 70924 3556 70926
rect 3500 70588 3556 70644
rect 4508 70978 4564 70980
rect 4508 70926 4510 70978
rect 4510 70926 4562 70978
rect 4562 70926 4564 70978
rect 4508 70924 4564 70926
rect 3804 70586 3860 70588
rect 3804 70534 3806 70586
rect 3806 70534 3858 70586
rect 3858 70534 3860 70586
rect 3804 70532 3860 70534
rect 3908 70586 3964 70588
rect 3908 70534 3910 70586
rect 3910 70534 3962 70586
rect 3962 70534 3964 70586
rect 3908 70532 3964 70534
rect 4012 70586 4068 70588
rect 4012 70534 4014 70586
rect 4014 70534 4066 70586
rect 4066 70534 4068 70586
rect 4012 70532 4068 70534
rect 4284 70476 4340 70532
rect 3388 69244 3444 69300
rect 3836 69132 3892 69188
rect 3804 69018 3860 69020
rect 3804 68966 3806 69018
rect 3806 68966 3858 69018
rect 3858 68966 3860 69018
rect 3804 68964 3860 68966
rect 3908 69018 3964 69020
rect 3908 68966 3910 69018
rect 3910 68966 3962 69018
rect 3962 68966 3964 69018
rect 3908 68964 3964 68966
rect 4012 69018 4068 69020
rect 4012 68966 4014 69018
rect 4014 68966 4066 69018
rect 4066 68966 4068 69018
rect 4012 68964 4068 68966
rect 4464 69802 4520 69804
rect 4464 69750 4466 69802
rect 4466 69750 4518 69802
rect 4518 69750 4520 69802
rect 4464 69748 4520 69750
rect 4568 69802 4624 69804
rect 4568 69750 4570 69802
rect 4570 69750 4622 69802
rect 4622 69750 4624 69802
rect 4568 69748 4624 69750
rect 4672 69802 4728 69804
rect 4672 69750 4674 69802
rect 4674 69750 4726 69802
rect 4726 69750 4728 69802
rect 4672 69748 4728 69750
rect 4172 68796 4228 68852
rect 3388 67228 3444 67284
rect 3948 67676 4004 67732
rect 3804 67450 3860 67452
rect 3804 67398 3806 67450
rect 3806 67398 3858 67450
rect 3858 67398 3860 67450
rect 3804 67396 3860 67398
rect 3908 67450 3964 67452
rect 3908 67398 3910 67450
rect 3910 67398 3962 67450
rect 3962 67398 3964 67450
rect 3908 67396 3964 67398
rect 4012 67450 4068 67452
rect 4012 67398 4014 67450
rect 4014 67398 4066 67450
rect 4066 67398 4068 67450
rect 4012 67396 4068 67398
rect 4844 68460 4900 68516
rect 4956 70924 5012 70980
rect 5292 71260 5348 71316
rect 5628 78204 5684 78260
rect 5628 77868 5684 77924
rect 5852 79324 5908 79380
rect 5852 76860 5908 76916
rect 6412 86940 6468 86996
rect 6748 86828 6804 86884
rect 6748 86156 6804 86212
rect 6412 85148 6468 85204
rect 6524 85596 6580 85652
rect 6300 84140 6356 84196
rect 7084 90748 7140 90804
rect 7308 100716 7364 100772
rect 7420 100492 7476 100548
rect 7308 98700 7364 98756
rect 7644 100268 7700 100324
rect 8540 104524 8596 104580
rect 8988 108892 9044 108948
rect 9212 110290 9268 110292
rect 9212 110238 9214 110290
rect 9214 110238 9266 110290
rect 9266 110238 9268 110290
rect 9212 110236 9268 110238
rect 8876 108610 8932 108612
rect 8876 108558 8878 108610
rect 8878 108558 8930 108610
rect 8930 108558 8932 108610
rect 8876 108556 8932 108558
rect 9212 108834 9268 108836
rect 9212 108782 9214 108834
rect 9214 108782 9266 108834
rect 9266 108782 9268 108834
rect 9212 108780 9268 108782
rect 9100 108444 9156 108500
rect 8876 106930 8932 106932
rect 8876 106878 8878 106930
rect 8878 106878 8930 106930
rect 8930 106878 8932 106930
rect 8876 106876 8932 106878
rect 9324 108108 9380 108164
rect 9436 111804 9492 111860
rect 9324 107826 9380 107828
rect 9324 107774 9326 107826
rect 9326 107774 9378 107826
rect 9378 107774 9380 107826
rect 9324 107772 9380 107774
rect 9100 105756 9156 105812
rect 10332 111804 10388 111860
rect 10220 111692 10276 111748
rect 9996 110402 10052 110404
rect 9996 110350 9998 110402
rect 9998 110350 10050 110402
rect 10050 110350 10052 110402
rect 9996 110348 10052 110350
rect 10332 110178 10388 110180
rect 10332 110126 10334 110178
rect 10334 110126 10386 110178
rect 10386 110126 10388 110178
rect 10332 110124 10388 110126
rect 9884 109394 9940 109396
rect 9884 109342 9886 109394
rect 9886 109342 9938 109394
rect 9938 109342 9940 109394
rect 9884 109340 9940 109342
rect 10220 109900 10276 109956
rect 9548 109116 9604 109172
rect 9548 108892 9604 108948
rect 9548 106930 9604 106932
rect 9548 106878 9550 106930
rect 9550 106878 9602 106930
rect 9602 106878 9604 106930
rect 9548 106876 9604 106878
rect 10668 112476 10724 112532
rect 10556 111746 10612 111748
rect 10556 111694 10558 111746
rect 10558 111694 10610 111746
rect 10610 111694 10612 111746
rect 10556 111692 10612 111694
rect 10780 112140 10836 112196
rect 10892 111970 10948 111972
rect 10892 111918 10894 111970
rect 10894 111918 10946 111970
rect 10946 111918 10948 111970
rect 10892 111916 10948 111918
rect 10892 111356 10948 111412
rect 10668 111020 10724 111076
rect 10556 110962 10612 110964
rect 10556 110910 10558 110962
rect 10558 110910 10610 110962
rect 10610 110910 10612 110962
rect 10556 110908 10612 110910
rect 9996 108668 10052 108724
rect 9884 108610 9940 108612
rect 9884 108558 9886 108610
rect 9886 108558 9938 108610
rect 9938 108558 9940 108610
rect 9884 108556 9940 108558
rect 9884 107884 9940 107940
rect 9772 107826 9828 107828
rect 9772 107774 9774 107826
rect 9774 107774 9826 107826
rect 9826 107774 9828 107826
rect 9772 107772 9828 107774
rect 10556 108892 10612 108948
rect 10892 110684 10948 110740
rect 10780 109170 10836 109172
rect 10780 109118 10782 109170
rect 10782 109118 10834 109170
rect 10834 109118 10836 109170
rect 10780 109116 10836 109118
rect 11116 112476 11172 112532
rect 11340 112364 11396 112420
rect 11228 111634 11284 111636
rect 11228 111582 11230 111634
rect 11230 111582 11282 111634
rect 11282 111582 11284 111634
rect 11228 111580 11284 111582
rect 11228 109900 11284 109956
rect 10668 108332 10724 108388
rect 9996 107772 10052 107828
rect 10444 107714 10500 107716
rect 10444 107662 10446 107714
rect 10446 107662 10498 107714
rect 10498 107662 10500 107714
rect 10444 107660 10500 107662
rect 9996 106146 10052 106148
rect 9996 106094 9998 106146
rect 9998 106094 10050 106146
rect 10050 106094 10052 106146
rect 9996 106092 10052 106094
rect 11004 107826 11060 107828
rect 11004 107774 11006 107826
rect 11006 107774 11058 107826
rect 11058 107774 11060 107826
rect 11004 107772 11060 107774
rect 10780 106930 10836 106932
rect 10780 106878 10782 106930
rect 10782 106878 10834 106930
rect 10834 106878 10836 106930
rect 10780 106876 10836 106878
rect 11564 113426 11620 113428
rect 11564 113374 11566 113426
rect 11566 113374 11618 113426
rect 11618 113374 11620 113426
rect 11564 113372 11620 113374
rect 11900 114380 11956 114436
rect 12124 114156 12180 114212
rect 12348 113820 12404 113876
rect 12460 114492 12516 114548
rect 11900 113708 11956 113764
rect 11676 112700 11732 112756
rect 11564 112418 11620 112420
rect 11564 112366 11566 112418
rect 11566 112366 11618 112418
rect 11618 112366 11620 112418
rect 11564 112364 11620 112366
rect 12572 113596 12628 113652
rect 12236 113036 12292 113092
rect 11900 112476 11956 112532
rect 12012 112924 12068 112980
rect 11900 112028 11956 112084
rect 12124 112588 12180 112644
rect 13020 113484 13076 113540
rect 13244 113036 13300 113092
rect 12796 112924 12852 112980
rect 11564 110908 11620 110964
rect 12236 112028 12292 112084
rect 12236 111132 12292 111188
rect 11564 110460 11620 110516
rect 12460 112028 12516 112084
rect 12236 110348 12292 110404
rect 12124 109282 12180 109284
rect 12124 109230 12126 109282
rect 12126 109230 12178 109282
rect 12178 109230 12180 109282
rect 12124 109228 12180 109230
rect 11340 107100 11396 107156
rect 11676 109116 11732 109172
rect 8876 103292 8932 103348
rect 8204 100716 8260 100772
rect 8652 102284 8708 102340
rect 8652 100492 8708 100548
rect 8988 102396 9044 102452
rect 8092 99932 8148 99988
rect 7532 98812 7588 98868
rect 8204 98978 8260 98980
rect 8204 98926 8206 98978
rect 8206 98926 8258 98978
rect 8258 98926 8260 98978
rect 8204 98924 8260 98926
rect 8092 98812 8148 98868
rect 7308 97692 7364 97748
rect 7420 98418 7476 98420
rect 7420 98366 7422 98418
rect 7422 98366 7474 98418
rect 7474 98366 7476 98418
rect 7420 98364 7476 98366
rect 7420 97580 7476 97636
rect 7980 98306 8036 98308
rect 7980 98254 7982 98306
rect 7982 98254 8034 98306
rect 8034 98254 8036 98306
rect 7980 98252 8036 98254
rect 7644 97468 7700 97524
rect 7420 97132 7476 97188
rect 7308 96348 7364 96404
rect 7308 95564 7364 95620
rect 7756 97356 7812 97412
rect 8204 97634 8260 97636
rect 8204 97582 8206 97634
rect 8206 97582 8258 97634
rect 8258 97582 8260 97634
rect 8204 97580 8260 97582
rect 8092 97468 8148 97524
rect 8204 96796 8260 96852
rect 8428 97244 8484 97300
rect 7196 89906 7252 89908
rect 7196 89854 7198 89906
rect 7198 89854 7250 89906
rect 7250 89854 7252 89906
rect 7196 89852 7252 89854
rect 7420 90636 7476 90692
rect 7084 87500 7140 87556
rect 7084 86716 7140 86772
rect 6748 82124 6804 82180
rect 6860 84140 6916 84196
rect 6412 81564 6468 81620
rect 6188 80780 6244 80836
rect 6748 81228 6804 81284
rect 6412 81004 6468 81060
rect 6636 81058 6692 81060
rect 6636 81006 6638 81058
rect 6638 81006 6690 81058
rect 6690 81006 6692 81058
rect 6636 81004 6692 81006
rect 6636 80780 6692 80836
rect 6076 80220 6132 80276
rect 6188 80108 6244 80164
rect 6076 78652 6132 78708
rect 6076 78316 6132 78372
rect 5740 76412 5796 76468
rect 5964 76242 6020 76244
rect 5964 76190 5966 76242
rect 5966 76190 6018 76242
rect 6018 76190 6020 76242
rect 5964 76188 6020 76190
rect 5852 75740 5908 75796
rect 6188 75852 6244 75908
rect 5628 74284 5684 74340
rect 6188 75628 6244 75684
rect 5628 71148 5684 71204
rect 5068 70700 5124 70756
rect 5292 70588 5348 70644
rect 5180 68908 5236 68964
rect 4464 68234 4520 68236
rect 4464 68182 4466 68234
rect 4466 68182 4518 68234
rect 4518 68182 4520 68234
rect 4464 68180 4520 68182
rect 4568 68234 4624 68236
rect 4568 68182 4570 68234
rect 4570 68182 4622 68234
rect 4622 68182 4624 68234
rect 4568 68180 4624 68182
rect 4672 68234 4728 68236
rect 4672 68182 4674 68234
rect 4674 68182 4726 68234
rect 4726 68182 4728 68234
rect 4672 68180 4728 68182
rect 4508 67842 4564 67844
rect 4508 67790 4510 67842
rect 4510 67790 4562 67842
rect 4562 67790 4564 67842
rect 4508 67788 4564 67790
rect 4284 66834 4340 66836
rect 4284 66782 4286 66834
rect 4286 66782 4338 66834
rect 4338 66782 4340 66834
rect 4284 66780 4340 66782
rect 4464 66666 4520 66668
rect 4464 66614 4466 66666
rect 4466 66614 4518 66666
rect 4518 66614 4520 66666
rect 4464 66612 4520 66614
rect 4568 66666 4624 66668
rect 4568 66614 4570 66666
rect 4570 66614 4622 66666
rect 4622 66614 4624 66666
rect 4568 66612 4624 66614
rect 4672 66666 4728 66668
rect 4672 66614 4674 66666
rect 4674 66614 4726 66666
rect 4726 66614 4728 66666
rect 4672 66612 4728 66614
rect 3612 66386 3668 66388
rect 3612 66334 3614 66386
rect 3614 66334 3666 66386
rect 3666 66334 3668 66386
rect 3612 66332 3668 66334
rect 3948 66274 4004 66276
rect 3948 66222 3950 66274
rect 3950 66222 4002 66274
rect 4002 66222 4004 66274
rect 3948 66220 4004 66222
rect 3804 65882 3860 65884
rect 3804 65830 3806 65882
rect 3806 65830 3858 65882
rect 3858 65830 3860 65882
rect 3804 65828 3860 65830
rect 3908 65882 3964 65884
rect 3908 65830 3910 65882
rect 3910 65830 3962 65882
rect 3962 65830 3964 65882
rect 3908 65828 3964 65830
rect 4012 65882 4068 65884
rect 4012 65830 4014 65882
rect 4014 65830 4066 65882
rect 4066 65830 4068 65882
rect 4012 65828 4068 65830
rect 4396 65490 4452 65492
rect 4396 65438 4398 65490
rect 4398 65438 4450 65490
rect 4450 65438 4452 65490
rect 4396 65436 4452 65438
rect 5404 70252 5460 70308
rect 5852 75068 5908 75124
rect 6524 80498 6580 80500
rect 6524 80446 6526 80498
rect 6526 80446 6578 80498
rect 6578 80446 6580 80498
rect 6524 80444 6580 80446
rect 6412 79324 6468 79380
rect 6748 79490 6804 79492
rect 6748 79438 6750 79490
rect 6750 79438 6802 79490
rect 6802 79438 6804 79490
rect 6748 79436 6804 79438
rect 6412 77868 6468 77924
rect 6972 83468 7028 83524
rect 7308 86828 7364 86884
rect 7756 91922 7812 91924
rect 7756 91870 7758 91922
rect 7758 91870 7810 91922
rect 7810 91870 7812 91922
rect 7756 91868 7812 91870
rect 8540 95564 8596 95620
rect 8652 97580 8708 97636
rect 8540 94780 8596 94836
rect 8204 94444 8260 94500
rect 8428 93884 8484 93940
rect 8316 93212 8372 93268
rect 8316 92876 8372 92932
rect 8204 92316 8260 92372
rect 7980 92204 8036 92260
rect 8540 92988 8596 93044
rect 8316 91868 8372 91924
rect 8204 91586 8260 91588
rect 8204 91534 8206 91586
rect 8206 91534 8258 91586
rect 8258 91534 8260 91586
rect 8204 91532 8260 91534
rect 7532 89682 7588 89684
rect 7532 89630 7534 89682
rect 7534 89630 7586 89682
rect 7586 89630 7588 89682
rect 7532 89628 7588 89630
rect 7868 89570 7924 89572
rect 7868 89518 7870 89570
rect 7870 89518 7922 89570
rect 7922 89518 7924 89570
rect 7868 89516 7924 89518
rect 7420 84588 7476 84644
rect 7532 84252 7588 84308
rect 8092 89292 8148 89348
rect 8092 85260 8148 85316
rect 8540 91868 8596 91924
rect 8204 84812 8260 84868
rect 8092 84028 8148 84084
rect 7868 83916 7924 83972
rect 7084 82348 7140 82404
rect 7084 82124 7140 82180
rect 7196 80444 7252 80500
rect 6636 77474 6692 77476
rect 6636 77422 6638 77474
rect 6638 77422 6690 77474
rect 6690 77422 6692 77474
rect 6636 77420 6692 77422
rect 6636 76748 6692 76804
rect 6636 76578 6692 76580
rect 6636 76526 6638 76578
rect 6638 76526 6690 76578
rect 6690 76526 6692 76578
rect 6636 76524 6692 76526
rect 6524 75852 6580 75908
rect 6636 75740 6692 75796
rect 5852 72940 5908 72996
rect 5852 71820 5908 71876
rect 6076 71874 6132 71876
rect 6076 71822 6078 71874
rect 6078 71822 6130 71874
rect 6130 71822 6132 71874
rect 6076 71820 6132 71822
rect 6860 78092 6916 78148
rect 6524 74620 6580 74676
rect 7196 79324 7252 79380
rect 7868 82012 7924 82068
rect 7308 78876 7364 78932
rect 7420 81340 7476 81396
rect 7084 78428 7140 78484
rect 7084 77980 7140 78036
rect 6972 76524 7028 76580
rect 6524 73388 6580 73444
rect 6300 72658 6356 72660
rect 6300 72606 6302 72658
rect 6302 72606 6354 72658
rect 6354 72606 6356 72658
rect 6300 72604 6356 72606
rect 6412 71762 6468 71764
rect 6412 71710 6414 71762
rect 6414 71710 6466 71762
rect 6466 71710 6468 71762
rect 6412 71708 6468 71710
rect 6300 71596 6356 71652
rect 6300 71372 6356 71428
rect 5852 70812 5908 70868
rect 5740 69132 5796 69188
rect 5628 68684 5684 68740
rect 4956 67954 5012 67956
rect 4956 67902 4958 67954
rect 4958 67902 5010 67954
rect 5010 67902 5012 67954
rect 4956 67900 5012 67902
rect 5292 67842 5348 67844
rect 5292 67790 5294 67842
rect 5294 67790 5346 67842
rect 5346 67790 5348 67842
rect 5292 67788 5348 67790
rect 5404 66780 5460 66836
rect 5180 66220 5236 66276
rect 4464 65098 4520 65100
rect 4464 65046 4466 65098
rect 4466 65046 4518 65098
rect 4518 65046 4520 65098
rect 4464 65044 4520 65046
rect 4568 65098 4624 65100
rect 4568 65046 4570 65098
rect 4570 65046 4622 65098
rect 4622 65046 4624 65098
rect 4568 65044 4624 65046
rect 4672 65098 4728 65100
rect 4672 65046 4674 65098
rect 4674 65046 4726 65098
rect 4726 65046 4728 65098
rect 4672 65044 4728 65046
rect 4956 64876 5012 64932
rect 3948 64428 4004 64484
rect 4284 64706 4340 64708
rect 4284 64654 4286 64706
rect 4286 64654 4338 64706
rect 4338 64654 4340 64706
rect 4284 64652 4340 64654
rect 3804 64314 3860 64316
rect 3804 64262 3806 64314
rect 3806 64262 3858 64314
rect 3858 64262 3860 64314
rect 3804 64260 3860 64262
rect 3908 64314 3964 64316
rect 3908 64262 3910 64314
rect 3910 64262 3962 64314
rect 3962 64262 3964 64314
rect 3908 64260 3964 64262
rect 4012 64314 4068 64316
rect 4012 64262 4014 64314
rect 4014 64262 4066 64314
rect 4066 64262 4068 64314
rect 4012 64260 4068 64262
rect 4172 63980 4228 64036
rect 3500 63922 3556 63924
rect 3500 63870 3502 63922
rect 3502 63870 3554 63922
rect 3554 63870 3556 63922
rect 3500 63868 3556 63870
rect 3164 63084 3220 63140
rect 3388 62860 3444 62916
rect 4956 64540 5012 64596
rect 5068 64316 5124 64372
rect 5180 64764 5236 64820
rect 4464 63530 4520 63532
rect 4464 63478 4466 63530
rect 4466 63478 4518 63530
rect 4518 63478 4520 63530
rect 4464 63476 4520 63478
rect 4568 63530 4624 63532
rect 4568 63478 4570 63530
rect 4570 63478 4622 63530
rect 4622 63478 4624 63530
rect 4568 63476 4624 63478
rect 4672 63530 4728 63532
rect 4672 63478 4674 63530
rect 4674 63478 4726 63530
rect 4726 63478 4728 63530
rect 4672 63476 4728 63478
rect 5292 63308 5348 63364
rect 4172 62860 4228 62916
rect 3804 62746 3860 62748
rect 3804 62694 3806 62746
rect 3806 62694 3858 62746
rect 3858 62694 3860 62746
rect 3804 62692 3860 62694
rect 3908 62746 3964 62748
rect 3908 62694 3910 62746
rect 3910 62694 3962 62746
rect 3962 62694 3964 62746
rect 3908 62692 3964 62694
rect 4012 62746 4068 62748
rect 4012 62694 4014 62746
rect 4014 62694 4066 62746
rect 4066 62694 4068 62746
rect 4012 62692 4068 62694
rect 3612 61852 3668 61908
rect 4172 62636 4228 62692
rect 3500 61682 3556 61684
rect 3500 61630 3502 61682
rect 3502 61630 3554 61682
rect 3554 61630 3556 61682
rect 3500 61628 3556 61630
rect 2156 60674 2212 60676
rect 2156 60622 2158 60674
rect 2158 60622 2210 60674
rect 2210 60622 2212 60674
rect 2156 60620 2212 60622
rect 1820 60562 1876 60564
rect 1820 60510 1822 60562
rect 1822 60510 1874 60562
rect 1874 60510 1876 60562
rect 1820 60508 1876 60510
rect 2380 59948 2436 60004
rect 2604 59836 2660 59892
rect 3804 61178 3860 61180
rect 3804 61126 3806 61178
rect 3806 61126 3858 61178
rect 3858 61126 3860 61178
rect 3804 61124 3860 61126
rect 3908 61178 3964 61180
rect 3908 61126 3910 61178
rect 3910 61126 3962 61178
rect 3962 61126 3964 61178
rect 3908 61124 3964 61126
rect 4012 61178 4068 61180
rect 4012 61126 4014 61178
rect 4014 61126 4066 61178
rect 4066 61126 4068 61178
rect 4012 61124 4068 61126
rect 3164 60562 3220 60564
rect 3164 60510 3166 60562
rect 3166 60510 3218 60562
rect 3218 60510 3220 60562
rect 3164 60508 3220 60510
rect 4956 62412 5012 62468
rect 5292 62242 5348 62244
rect 5292 62190 5294 62242
rect 5294 62190 5346 62242
rect 5346 62190 5348 62242
rect 5292 62188 5348 62190
rect 4284 62076 4340 62132
rect 4464 61962 4520 61964
rect 4464 61910 4466 61962
rect 4466 61910 4518 61962
rect 4518 61910 4520 61962
rect 4464 61908 4520 61910
rect 4568 61962 4624 61964
rect 4568 61910 4570 61962
rect 4570 61910 4622 61962
rect 4622 61910 4624 61962
rect 4568 61908 4624 61910
rect 4672 61962 4728 61964
rect 4672 61910 4674 61962
rect 4674 61910 4726 61962
rect 4726 61910 4728 61962
rect 4672 61908 4728 61910
rect 5068 61964 5124 62020
rect 4620 61570 4676 61572
rect 4620 61518 4622 61570
rect 4622 61518 4674 61570
rect 4674 61518 4676 61570
rect 4620 61516 4676 61518
rect 5404 61570 5460 61572
rect 5404 61518 5406 61570
rect 5406 61518 5458 61570
rect 5458 61518 5460 61570
rect 5404 61516 5460 61518
rect 4464 60394 4520 60396
rect 4464 60342 4466 60394
rect 4466 60342 4518 60394
rect 4518 60342 4520 60394
rect 4464 60340 4520 60342
rect 4568 60394 4624 60396
rect 4568 60342 4570 60394
rect 4570 60342 4622 60394
rect 4622 60342 4624 60394
rect 4568 60340 4624 60342
rect 4672 60394 4728 60396
rect 4672 60342 4674 60394
rect 4674 60342 4726 60394
rect 4726 60342 4728 60394
rect 4672 60340 4728 60342
rect 5180 60226 5236 60228
rect 5180 60174 5182 60226
rect 5182 60174 5234 60226
rect 5234 60174 5236 60226
rect 5180 60172 5236 60174
rect 3612 59890 3668 59892
rect 3612 59838 3614 59890
rect 3614 59838 3666 59890
rect 3666 59838 3668 59890
rect 3612 59836 3668 59838
rect 1372 58994 1428 58996
rect 1372 58942 1374 58994
rect 1374 58942 1426 58994
rect 1426 58942 1428 58994
rect 1372 58940 1428 58942
rect 1820 58994 1876 58996
rect 1820 58942 1822 58994
rect 1822 58942 1874 58994
rect 1874 58942 1876 58994
rect 1820 58940 1876 58942
rect 1372 58658 1428 58660
rect 1372 58606 1374 58658
rect 1374 58606 1426 58658
rect 1426 58606 1428 58658
rect 1372 58604 1428 58606
rect 1036 58156 1092 58212
rect 1260 56700 1316 56756
rect 252 41356 308 41412
rect 1148 50818 1204 50820
rect 1148 50766 1150 50818
rect 1150 50766 1202 50818
rect 1202 50766 1204 50818
rect 1148 50764 1204 50766
rect 812 50652 868 50708
rect 700 45836 756 45892
rect 700 40908 756 40964
rect 252 31612 308 31668
rect 364 29596 420 29652
rect 364 26236 420 26292
rect 1036 49980 1092 50036
rect 1260 49868 1316 49924
rect 1596 58716 1652 58772
rect 1036 48300 1092 48356
rect 1148 49532 1204 49588
rect 1484 53900 1540 53956
rect 2044 58434 2100 58436
rect 2044 58382 2046 58434
rect 2046 58382 2098 58434
rect 2098 58382 2100 58434
rect 2044 58380 2100 58382
rect 1708 57708 1764 57764
rect 1932 58044 1988 58100
rect 1932 55356 1988 55412
rect 1596 52780 1652 52836
rect 1820 54908 1876 54964
rect 1484 52668 1540 52724
rect 1484 50706 1540 50708
rect 1484 50654 1486 50706
rect 1486 50654 1538 50706
rect 1538 50654 1540 50706
rect 1484 50652 1540 50654
rect 1372 48524 1428 48580
rect 1596 48412 1652 48468
rect 1708 48300 1764 48356
rect 1484 46732 1540 46788
rect 1708 46508 1764 46564
rect 2156 54626 2212 54628
rect 2156 54574 2158 54626
rect 2158 54574 2210 54626
rect 2210 54574 2212 54626
rect 2156 54572 2212 54574
rect 2044 50594 2100 50596
rect 2044 50542 2046 50594
rect 2046 50542 2098 50594
rect 2098 50542 2100 50594
rect 2044 50540 2100 50542
rect 2268 49250 2324 49252
rect 2268 49198 2270 49250
rect 2270 49198 2322 49250
rect 2322 49198 2324 49250
rect 2268 49196 2324 49198
rect 1932 49026 1988 49028
rect 1932 48974 1934 49026
rect 1934 48974 1986 49026
rect 1986 48974 1988 49026
rect 1932 48972 1988 48974
rect 2156 48466 2212 48468
rect 2156 48414 2158 48466
rect 2158 48414 2210 48466
rect 2210 48414 2212 48466
rect 2156 48412 2212 48414
rect 2268 48076 2324 48132
rect 2044 47964 2100 48020
rect 1932 47570 1988 47572
rect 1932 47518 1934 47570
rect 1934 47518 1986 47570
rect 1986 47518 1988 47570
rect 1932 47516 1988 47518
rect 2268 47740 2324 47796
rect 1820 46060 1876 46116
rect 2268 47516 2324 47572
rect 1596 45836 1652 45892
rect 1148 45388 1204 45444
rect 1260 44156 1316 44212
rect 1260 43596 1316 43652
rect 364 19852 420 19908
rect 924 40796 980 40852
rect 588 19740 644 19796
rect 476 12796 532 12852
rect 364 11900 420 11956
rect 252 9884 308 9940
rect 252 5628 308 5684
rect 476 5292 532 5348
rect 364 4172 420 4228
rect 1148 39340 1204 39396
rect 1260 39506 1316 39508
rect 1260 39454 1262 39506
rect 1262 39454 1314 39506
rect 1314 39454 1316 39506
rect 1260 39452 1316 39454
rect 1708 45388 1764 45444
rect 1596 44828 1652 44884
rect 1484 44604 1540 44660
rect 1484 44044 1540 44100
rect 1708 44716 1764 44772
rect 1596 41580 1652 41636
rect 3804 59610 3860 59612
rect 3804 59558 3806 59610
rect 3806 59558 3858 59610
rect 3858 59558 3860 59610
rect 3804 59556 3860 59558
rect 3908 59610 3964 59612
rect 3908 59558 3910 59610
rect 3910 59558 3962 59610
rect 3962 59558 3964 59610
rect 3908 59556 3964 59558
rect 4012 59610 4068 59612
rect 4012 59558 4014 59610
rect 4014 59558 4066 59610
rect 4066 59558 4068 59610
rect 4012 59556 4068 59558
rect 2492 59106 2548 59108
rect 2492 59054 2494 59106
rect 2494 59054 2546 59106
rect 2546 59054 2548 59106
rect 2492 59052 2548 59054
rect 2828 59106 2884 59108
rect 2828 59054 2830 59106
rect 2830 59054 2882 59106
rect 2882 59054 2884 59106
rect 2828 59052 2884 59054
rect 4464 58826 4520 58828
rect 4464 58774 4466 58826
rect 4466 58774 4518 58826
rect 4518 58774 4520 58826
rect 4464 58772 4520 58774
rect 4568 58826 4624 58828
rect 4568 58774 4570 58826
rect 4570 58774 4622 58826
rect 4622 58774 4624 58826
rect 4568 58772 4624 58774
rect 4672 58826 4728 58828
rect 4672 58774 4674 58826
rect 4674 58774 4726 58826
rect 4726 58774 4728 58826
rect 4672 58772 4728 58774
rect 3804 58042 3860 58044
rect 3804 57990 3806 58042
rect 3806 57990 3858 58042
rect 3858 57990 3860 58042
rect 3804 57988 3860 57990
rect 3908 58042 3964 58044
rect 3908 57990 3910 58042
rect 3910 57990 3962 58042
rect 3962 57990 3964 58042
rect 3908 57988 3964 57990
rect 4012 58042 4068 58044
rect 4012 57990 4014 58042
rect 4014 57990 4066 58042
rect 4066 57990 4068 58042
rect 4012 57988 4068 57990
rect 4464 57258 4520 57260
rect 4464 57206 4466 57258
rect 4466 57206 4518 57258
rect 4518 57206 4520 57258
rect 4464 57204 4520 57206
rect 4568 57258 4624 57260
rect 4568 57206 4570 57258
rect 4570 57206 4622 57258
rect 4622 57206 4624 57258
rect 4568 57204 4624 57206
rect 4672 57258 4728 57260
rect 4672 57206 4674 57258
rect 4674 57206 4726 57258
rect 4726 57206 4728 57258
rect 4672 57204 4728 57206
rect 2940 56700 2996 56756
rect 2492 55804 2548 55860
rect 4396 56754 4452 56756
rect 4396 56702 4398 56754
rect 4398 56702 4450 56754
rect 4450 56702 4452 56754
rect 4396 56700 4452 56702
rect 3804 56474 3860 56476
rect 3804 56422 3806 56474
rect 3806 56422 3858 56474
rect 3858 56422 3860 56474
rect 3804 56420 3860 56422
rect 3908 56474 3964 56476
rect 3908 56422 3910 56474
rect 3910 56422 3962 56474
rect 3962 56422 3964 56474
rect 3908 56420 3964 56422
rect 4012 56474 4068 56476
rect 4012 56422 4014 56474
rect 4014 56422 4066 56474
rect 4066 56422 4068 56474
rect 4012 56420 4068 56422
rect 3500 56252 3556 56308
rect 2940 54572 2996 54628
rect 2492 53452 2548 53508
rect 2492 50652 2548 50708
rect 3276 55804 3332 55860
rect 4396 56140 4452 56196
rect 4844 56588 4900 56644
rect 4464 55690 4520 55692
rect 4464 55638 4466 55690
rect 4466 55638 4518 55690
rect 4518 55638 4520 55690
rect 4464 55636 4520 55638
rect 4568 55690 4624 55692
rect 4568 55638 4570 55690
rect 4570 55638 4622 55690
rect 4622 55638 4624 55690
rect 4568 55636 4624 55638
rect 4672 55690 4728 55692
rect 4672 55638 4674 55690
rect 4674 55638 4726 55690
rect 4726 55638 4728 55690
rect 4672 55636 4728 55638
rect 4620 55298 4676 55300
rect 4620 55246 4622 55298
rect 4622 55246 4674 55298
rect 4674 55246 4676 55298
rect 4620 55244 4676 55246
rect 3804 54906 3860 54908
rect 3804 54854 3806 54906
rect 3806 54854 3858 54906
rect 3858 54854 3860 54906
rect 3804 54852 3860 54854
rect 3908 54906 3964 54908
rect 3908 54854 3910 54906
rect 3910 54854 3962 54906
rect 3962 54854 3964 54906
rect 3908 54852 3964 54854
rect 4012 54906 4068 54908
rect 4012 54854 4014 54906
rect 4014 54854 4066 54906
rect 4066 54854 4068 54906
rect 4012 54852 4068 54854
rect 3724 54738 3780 54740
rect 3724 54686 3726 54738
rect 3726 54686 3778 54738
rect 3778 54686 3780 54738
rect 3724 54684 3780 54686
rect 4464 54122 4520 54124
rect 4464 54070 4466 54122
rect 4466 54070 4518 54122
rect 4518 54070 4520 54122
rect 4464 54068 4520 54070
rect 4568 54122 4624 54124
rect 4568 54070 4570 54122
rect 4570 54070 4622 54122
rect 4622 54070 4624 54122
rect 4568 54068 4624 54070
rect 4672 54122 4728 54124
rect 4672 54070 4674 54122
rect 4674 54070 4726 54122
rect 4726 54070 4728 54122
rect 4672 54068 4728 54070
rect 3500 53452 3556 53508
rect 4620 53506 4676 53508
rect 4620 53454 4622 53506
rect 4622 53454 4674 53506
rect 4674 53454 4676 53506
rect 4620 53452 4676 53454
rect 3804 53338 3860 53340
rect 3804 53286 3806 53338
rect 3806 53286 3858 53338
rect 3858 53286 3860 53338
rect 3804 53284 3860 53286
rect 3908 53338 3964 53340
rect 3908 53286 3910 53338
rect 3910 53286 3962 53338
rect 3962 53286 3964 53338
rect 3908 53284 3964 53286
rect 4012 53338 4068 53340
rect 4012 53286 4014 53338
rect 4014 53286 4066 53338
rect 4066 53286 4068 53338
rect 4012 53284 4068 53286
rect 4284 52722 4340 52724
rect 4284 52670 4286 52722
rect 4286 52670 4338 52722
rect 4338 52670 4340 52722
rect 4284 52668 4340 52670
rect 4464 52554 4520 52556
rect 4464 52502 4466 52554
rect 4466 52502 4518 52554
rect 4518 52502 4520 52554
rect 4464 52500 4520 52502
rect 4568 52554 4624 52556
rect 4568 52502 4570 52554
rect 4570 52502 4622 52554
rect 4622 52502 4624 52554
rect 4568 52500 4624 52502
rect 4672 52554 4728 52556
rect 4672 52502 4674 52554
rect 4674 52502 4726 52554
rect 4726 52502 4728 52554
rect 4672 52500 4728 52502
rect 3052 52108 3108 52164
rect 2828 50540 2884 50596
rect 2604 49980 2660 50036
rect 2716 48914 2772 48916
rect 2716 48862 2718 48914
rect 2718 48862 2770 48914
rect 2770 48862 2772 48914
rect 2716 48860 2772 48862
rect 2604 48076 2660 48132
rect 2716 48636 2772 48692
rect 2492 47964 2548 48020
rect 3276 49980 3332 50036
rect 4508 52386 4564 52388
rect 4508 52334 4510 52386
rect 4510 52334 4562 52386
rect 4562 52334 4564 52386
rect 4508 52332 4564 52334
rect 4844 52220 4900 52276
rect 5068 55410 5124 55412
rect 5068 55358 5070 55410
rect 5070 55358 5122 55410
rect 5122 55358 5124 55410
rect 5068 55356 5124 55358
rect 3804 51770 3860 51772
rect 3804 51718 3806 51770
rect 3806 51718 3858 51770
rect 3858 51718 3860 51770
rect 3804 51716 3860 51718
rect 3908 51770 3964 51772
rect 3908 51718 3910 51770
rect 3910 51718 3962 51770
rect 3962 51718 3964 51770
rect 3908 51716 3964 51718
rect 4012 51770 4068 51772
rect 4012 51718 4014 51770
rect 4014 51718 4066 51770
rect 4066 51718 4068 51770
rect 4012 51716 4068 51718
rect 5404 54684 5460 54740
rect 5292 53452 5348 53508
rect 3388 51212 3444 51268
rect 2940 49532 2996 49588
rect 3276 49084 3332 49140
rect 2828 48300 2884 48356
rect 2716 47458 2772 47460
rect 2716 47406 2718 47458
rect 2718 47406 2770 47458
rect 2770 47406 2772 47458
rect 2716 47404 2772 47406
rect 2716 47180 2772 47236
rect 3276 48524 3332 48580
rect 2940 47516 2996 47572
rect 3052 47964 3108 48020
rect 4284 51154 4340 51156
rect 4284 51102 4286 51154
rect 4286 51102 4338 51154
rect 4338 51102 4340 51154
rect 4284 51100 4340 51102
rect 4464 50986 4520 50988
rect 4464 50934 4466 50986
rect 4466 50934 4518 50986
rect 4518 50934 4520 50986
rect 4464 50932 4520 50934
rect 4568 50986 4624 50988
rect 4568 50934 4570 50986
rect 4570 50934 4622 50986
rect 4622 50934 4624 50986
rect 4568 50932 4624 50934
rect 4672 50986 4728 50988
rect 4672 50934 4674 50986
rect 4674 50934 4726 50986
rect 4726 50934 4728 50986
rect 4672 50932 4728 50934
rect 5068 50818 5124 50820
rect 5068 50766 5070 50818
rect 5070 50766 5122 50818
rect 5122 50766 5124 50818
rect 5068 50764 5124 50766
rect 4956 50594 5012 50596
rect 4956 50542 4958 50594
rect 4958 50542 5010 50594
rect 5010 50542 5012 50594
rect 4956 50540 5012 50542
rect 4060 50482 4116 50484
rect 4060 50430 4062 50482
rect 4062 50430 4114 50482
rect 4114 50430 4116 50482
rect 4060 50428 4116 50430
rect 5964 68796 6020 68852
rect 6188 68124 6244 68180
rect 5964 66556 6020 66612
rect 6076 67564 6132 67620
rect 5964 66332 6020 66388
rect 5852 66274 5908 66276
rect 5852 66222 5854 66274
rect 5854 66222 5906 66274
rect 5906 66222 5908 66274
rect 5852 66220 5908 66222
rect 5852 65602 5908 65604
rect 5852 65550 5854 65602
rect 5854 65550 5906 65602
rect 5906 65550 5908 65602
rect 5852 65548 5908 65550
rect 6076 65884 6132 65940
rect 5740 64652 5796 64708
rect 5628 63644 5684 63700
rect 5628 63196 5684 63252
rect 5740 63138 5796 63140
rect 5740 63086 5742 63138
rect 5742 63086 5794 63138
rect 5794 63086 5796 63138
rect 5740 63084 5796 63086
rect 5628 61964 5684 62020
rect 6076 62412 6132 62468
rect 5964 62354 6020 62356
rect 5964 62302 5966 62354
rect 5966 62302 6018 62354
rect 6018 62302 6020 62354
rect 5964 62300 6020 62302
rect 6076 61794 6132 61796
rect 6076 61742 6078 61794
rect 6078 61742 6130 61794
rect 6130 61742 6132 61794
rect 6076 61740 6132 61742
rect 5964 60172 6020 60228
rect 5852 59890 5908 59892
rect 5852 59838 5854 59890
rect 5854 59838 5906 59890
rect 5906 59838 5908 59890
rect 5852 59836 5908 59838
rect 6636 72604 6692 72660
rect 6636 72268 6692 72324
rect 6860 73948 6916 74004
rect 7420 77756 7476 77812
rect 7868 79548 7924 79604
rect 8092 81228 8148 81284
rect 8092 79212 8148 79268
rect 7980 78428 8036 78484
rect 7868 78034 7924 78036
rect 7868 77982 7870 78034
rect 7870 77982 7922 78034
rect 7922 77982 7924 78034
rect 7868 77980 7924 77982
rect 7756 77532 7812 77588
rect 7868 77756 7924 77812
rect 7532 77084 7588 77140
rect 7084 75906 7140 75908
rect 7084 75854 7086 75906
rect 7086 75854 7138 75906
rect 7138 75854 7140 75906
rect 7084 75852 7140 75854
rect 7644 76354 7700 76356
rect 7644 76302 7646 76354
rect 7646 76302 7698 76354
rect 7698 76302 7700 76354
rect 7644 76300 7700 76302
rect 7532 74338 7588 74340
rect 7532 74286 7534 74338
rect 7534 74286 7586 74338
rect 7586 74286 7588 74338
rect 7532 74284 7588 74286
rect 7420 74172 7476 74228
rect 7084 73836 7140 73892
rect 7196 73724 7252 73780
rect 7420 73612 7476 73668
rect 7196 72828 7252 72884
rect 6748 69580 6804 69636
rect 6860 70812 6916 70868
rect 6524 68796 6580 68852
rect 6636 69132 6692 69188
rect 6524 67116 6580 67172
rect 6300 65884 6356 65940
rect 6412 66220 6468 66276
rect 6300 65100 6356 65156
rect 6300 63644 6356 63700
rect 6524 65548 6580 65604
rect 6524 63084 6580 63140
rect 6412 62354 6468 62356
rect 6412 62302 6414 62354
rect 6414 62302 6466 62354
rect 6466 62302 6468 62354
rect 6412 62300 6468 62302
rect 6524 62860 6580 62916
rect 6636 62242 6692 62244
rect 6636 62190 6638 62242
rect 6638 62190 6690 62242
rect 6690 62190 6692 62242
rect 6636 62188 6692 62190
rect 6636 60674 6692 60676
rect 6636 60622 6638 60674
rect 6638 60622 6690 60674
rect 6690 60622 6692 60674
rect 6636 60620 6692 60622
rect 6300 60114 6356 60116
rect 6300 60062 6302 60114
rect 6302 60062 6354 60114
rect 6354 60062 6356 60114
rect 6300 60060 6356 60062
rect 5852 56194 5908 56196
rect 5852 56142 5854 56194
rect 5854 56142 5906 56194
rect 5906 56142 5908 56194
rect 5852 56140 5908 56142
rect 5628 54684 5684 54740
rect 5740 55356 5796 55412
rect 5516 53228 5572 53284
rect 5628 51996 5684 52052
rect 5516 51100 5572 51156
rect 5628 50428 5684 50484
rect 3804 50202 3860 50204
rect 3804 50150 3806 50202
rect 3806 50150 3858 50202
rect 3858 50150 3860 50202
rect 3804 50148 3860 50150
rect 3908 50202 3964 50204
rect 3908 50150 3910 50202
rect 3910 50150 3962 50202
rect 3962 50150 3964 50202
rect 3908 50148 3964 50150
rect 4012 50202 4068 50204
rect 4012 50150 4014 50202
rect 4014 50150 4066 50202
rect 4066 50150 4068 50202
rect 4012 50148 4068 50150
rect 4956 49868 5012 49924
rect 4464 49418 4520 49420
rect 4464 49366 4466 49418
rect 4466 49366 4518 49418
rect 4518 49366 4520 49418
rect 4464 49364 4520 49366
rect 4568 49418 4624 49420
rect 4568 49366 4570 49418
rect 4570 49366 4622 49418
rect 4622 49366 4624 49418
rect 4568 49364 4624 49366
rect 4672 49418 4728 49420
rect 4672 49366 4674 49418
rect 4674 49366 4726 49418
rect 4726 49366 4728 49418
rect 4672 49364 4728 49366
rect 3724 48972 3780 49028
rect 3612 48748 3668 48804
rect 3804 48634 3860 48636
rect 3804 48582 3806 48634
rect 3806 48582 3858 48634
rect 3858 48582 3860 48634
rect 3804 48580 3860 48582
rect 3908 48634 3964 48636
rect 3908 48582 3910 48634
rect 3910 48582 3962 48634
rect 3962 48582 3964 48634
rect 3908 48580 3964 48582
rect 4012 48634 4068 48636
rect 4012 48582 4014 48634
rect 4014 48582 4066 48634
rect 4066 48582 4068 48634
rect 4012 48580 4068 48582
rect 3612 48300 3668 48356
rect 3500 48188 3556 48244
rect 3164 47180 3220 47236
rect 2940 46620 2996 46676
rect 2156 45612 2212 45668
rect 1932 42642 1988 42644
rect 1932 42590 1934 42642
rect 1934 42590 1986 42642
rect 1986 42590 1988 42642
rect 1932 42588 1988 42590
rect 2044 43538 2100 43540
rect 2044 43486 2046 43538
rect 2046 43486 2098 43538
rect 2098 43486 2100 43538
rect 2044 43484 2100 43486
rect 1708 39452 1764 39508
rect 1596 39340 1652 39396
rect 1484 37324 1540 37380
rect 1484 36482 1540 36484
rect 1484 36430 1486 36482
rect 1486 36430 1538 36482
rect 1538 36430 1540 36482
rect 1484 36428 1540 36430
rect 1148 35810 1204 35812
rect 1148 35758 1150 35810
rect 1150 35758 1202 35810
rect 1202 35758 1204 35810
rect 1148 35756 1204 35758
rect 1036 35196 1092 35252
rect 1148 32786 1204 32788
rect 1148 32734 1150 32786
rect 1150 32734 1202 32786
rect 1202 32734 1204 32786
rect 1148 32732 1204 32734
rect 1372 32172 1428 32228
rect 1260 28588 1316 28644
rect 1148 27970 1204 27972
rect 1148 27918 1150 27970
rect 1150 27918 1202 27970
rect 1202 27918 1204 27970
rect 1148 27916 1204 27918
rect 1148 25228 1204 25284
rect 812 23324 868 23380
rect 700 17388 756 17444
rect 812 22988 868 23044
rect 1036 21308 1092 21364
rect 924 20412 980 20468
rect 1260 24722 1316 24724
rect 1260 24670 1262 24722
rect 1262 24670 1314 24722
rect 1314 24670 1316 24722
rect 1260 24668 1316 24670
rect 2828 44882 2884 44884
rect 2828 44830 2830 44882
rect 2830 44830 2882 44882
rect 2882 44830 2884 44882
rect 2828 44828 2884 44830
rect 2156 41746 2212 41748
rect 2156 41694 2158 41746
rect 2158 41694 2210 41746
rect 2210 41694 2212 41746
rect 2156 41692 2212 41694
rect 2604 41580 2660 41636
rect 2044 40290 2100 40292
rect 2044 40238 2046 40290
rect 2046 40238 2098 40290
rect 2098 40238 2100 40290
rect 2044 40236 2100 40238
rect 1932 38162 1988 38164
rect 1932 38110 1934 38162
rect 1934 38110 1986 38162
rect 1986 38110 1988 38162
rect 1932 38108 1988 38110
rect 2380 40572 2436 40628
rect 2940 42028 2996 42084
rect 2940 41020 2996 41076
rect 2828 40236 2884 40292
rect 2828 38668 2884 38724
rect 3500 46732 3556 46788
rect 3724 48242 3780 48244
rect 3724 48190 3726 48242
rect 3726 48190 3778 48242
rect 3778 48190 3780 48242
rect 3724 48188 3780 48190
rect 4060 47964 4116 48020
rect 3724 47570 3780 47572
rect 3724 47518 3726 47570
rect 3726 47518 3778 47570
rect 3778 47518 3780 47570
rect 3724 47516 3780 47518
rect 3612 47292 3668 47348
rect 3388 44828 3444 44884
rect 3164 41804 3220 41860
rect 3388 41580 3444 41636
rect 3276 41468 3332 41524
rect 3388 41132 3444 41188
rect 3276 40402 3332 40404
rect 3276 40350 3278 40402
rect 3278 40350 3330 40402
rect 3330 40350 3332 40402
rect 3276 40348 3332 40350
rect 1932 37266 1988 37268
rect 1932 37214 1934 37266
rect 1934 37214 1986 37266
rect 1986 37214 1988 37266
rect 1932 37212 1988 37214
rect 1820 36988 1876 37044
rect 1708 34748 1764 34804
rect 1708 32732 1764 32788
rect 1820 32172 1876 32228
rect 2268 36316 2324 36372
rect 2044 34524 2100 34580
rect 1708 31836 1764 31892
rect 2044 33740 2100 33796
rect 1596 30380 1652 30436
rect 1708 30940 1764 30996
rect 1484 28812 1540 28868
rect 1932 31666 1988 31668
rect 1932 31614 1934 31666
rect 1934 31614 1986 31666
rect 1986 31614 1988 31666
rect 1932 31612 1988 31614
rect 2156 33628 2212 33684
rect 2156 33458 2212 33460
rect 2156 33406 2158 33458
rect 2158 33406 2210 33458
rect 2210 33406 2212 33458
rect 2156 33404 2212 33406
rect 2492 37212 2548 37268
rect 2716 37378 2772 37380
rect 2716 37326 2718 37378
rect 2718 37326 2770 37378
rect 2770 37326 2772 37378
rect 2716 37324 2772 37326
rect 2604 36316 2660 36372
rect 2716 35196 2772 35252
rect 3052 37826 3108 37828
rect 3052 37774 3054 37826
rect 3054 37774 3106 37826
rect 3106 37774 3108 37826
rect 3052 37772 3108 37774
rect 3164 37042 3220 37044
rect 3164 36990 3166 37042
rect 3166 36990 3218 37042
rect 3218 36990 3220 37042
rect 3164 36988 3220 36990
rect 2380 34242 2436 34244
rect 2380 34190 2382 34242
rect 2382 34190 2434 34242
rect 2434 34190 2436 34242
rect 2380 34188 2436 34190
rect 2380 33740 2436 33796
rect 2940 34188 2996 34244
rect 2828 32396 2884 32452
rect 2492 31836 2548 31892
rect 2156 31612 2212 31668
rect 2268 31724 2324 31780
rect 2716 31778 2772 31780
rect 2716 31726 2718 31778
rect 2718 31726 2770 31778
rect 2770 31726 2772 31778
rect 2716 31724 2772 31726
rect 2716 31500 2772 31556
rect 2044 31052 2100 31108
rect 1820 29148 1876 29204
rect 2044 29932 2100 29988
rect 1708 28642 1764 28644
rect 1708 28590 1710 28642
rect 1710 28590 1762 28642
rect 1762 28590 1764 28642
rect 1708 28588 1764 28590
rect 1484 27916 1540 27972
rect 2268 29314 2324 29316
rect 2268 29262 2270 29314
rect 2270 29262 2322 29314
rect 2322 29262 2324 29314
rect 2268 29260 2324 29262
rect 2156 28866 2212 28868
rect 2156 28814 2158 28866
rect 2158 28814 2210 28866
rect 2210 28814 2212 28866
rect 2156 28812 2212 28814
rect 1932 27692 1988 27748
rect 1260 23660 1316 23716
rect 1372 21698 1428 21700
rect 1372 21646 1374 21698
rect 1374 21646 1426 21698
rect 1426 21646 1428 21698
rect 1372 21644 1428 21646
rect 1260 20300 1316 20356
rect 1708 26460 1764 26516
rect 1596 26178 1652 26180
rect 1596 26126 1598 26178
rect 1598 26126 1650 26178
rect 1650 26126 1652 26178
rect 1596 26124 1652 26126
rect 2156 27356 2212 27412
rect 1932 26460 1988 26516
rect 2492 30380 2548 30436
rect 2492 30044 2548 30100
rect 2492 29484 2548 29540
rect 2492 27692 2548 27748
rect 1820 25228 1876 25284
rect 1932 26236 1988 26292
rect 1708 24668 1764 24724
rect 2156 25506 2212 25508
rect 2156 25454 2158 25506
rect 2158 25454 2210 25506
rect 2210 25454 2212 25506
rect 2156 25452 2212 25454
rect 2492 26908 2548 26964
rect 2716 29538 2772 29540
rect 2716 29486 2718 29538
rect 2718 29486 2770 29538
rect 2770 29486 2772 29538
rect 2716 29484 2772 29486
rect 2940 31890 2996 31892
rect 2940 31838 2942 31890
rect 2942 31838 2994 31890
rect 2994 31838 2996 31890
rect 2940 31836 2996 31838
rect 3388 36428 3444 36484
rect 3500 41020 3556 41076
rect 4464 47850 4520 47852
rect 4464 47798 4466 47850
rect 4466 47798 4518 47850
rect 4518 47798 4520 47850
rect 4464 47796 4520 47798
rect 4568 47850 4624 47852
rect 4568 47798 4570 47850
rect 4570 47798 4622 47850
rect 4622 47798 4624 47850
rect 4568 47796 4624 47798
rect 4672 47850 4728 47852
rect 4672 47798 4674 47850
rect 4674 47798 4726 47850
rect 4726 47798 4728 47850
rect 4672 47796 4728 47798
rect 4172 47404 4228 47460
rect 3804 47066 3860 47068
rect 3804 47014 3806 47066
rect 3806 47014 3858 47066
rect 3858 47014 3860 47066
rect 3804 47012 3860 47014
rect 3908 47066 3964 47068
rect 3908 47014 3910 47066
rect 3910 47014 3962 47066
rect 3962 47014 3964 47066
rect 3908 47012 3964 47014
rect 4012 47066 4068 47068
rect 4012 47014 4014 47066
rect 4014 47014 4066 47066
rect 4066 47014 4068 47066
rect 4012 47012 4068 47014
rect 3804 45498 3860 45500
rect 3804 45446 3806 45498
rect 3806 45446 3858 45498
rect 3858 45446 3860 45498
rect 3804 45444 3860 45446
rect 3908 45498 3964 45500
rect 3908 45446 3910 45498
rect 3910 45446 3962 45498
rect 3962 45446 3964 45498
rect 3908 45444 3964 45446
rect 4012 45498 4068 45500
rect 4012 45446 4014 45498
rect 4014 45446 4066 45498
rect 4066 45446 4068 45498
rect 4012 45444 4068 45446
rect 3804 43930 3860 43932
rect 3804 43878 3806 43930
rect 3806 43878 3858 43930
rect 3858 43878 3860 43930
rect 3804 43876 3860 43878
rect 3908 43930 3964 43932
rect 3908 43878 3910 43930
rect 3910 43878 3962 43930
rect 3962 43878 3964 43930
rect 3908 43876 3964 43878
rect 4012 43930 4068 43932
rect 4012 43878 4014 43930
rect 4014 43878 4066 43930
rect 4066 43878 4068 43930
rect 4012 43876 4068 43878
rect 5292 49532 5348 49588
rect 4956 48748 5012 48804
rect 5068 48860 5124 48916
rect 4844 47068 4900 47124
rect 5068 46956 5124 47012
rect 4956 46732 5012 46788
rect 4464 46282 4520 46284
rect 4464 46230 4466 46282
rect 4466 46230 4518 46282
rect 4518 46230 4520 46282
rect 4464 46228 4520 46230
rect 4568 46282 4624 46284
rect 4568 46230 4570 46282
rect 4570 46230 4622 46282
rect 4622 46230 4624 46282
rect 4568 46228 4624 46230
rect 4672 46282 4728 46284
rect 4672 46230 4674 46282
rect 4674 46230 4726 46282
rect 4726 46230 4728 46282
rect 4672 46228 4728 46230
rect 4844 45836 4900 45892
rect 4396 45500 4452 45556
rect 5068 45612 5124 45668
rect 4956 45388 5012 45444
rect 4464 44714 4520 44716
rect 4464 44662 4466 44714
rect 4466 44662 4518 44714
rect 4518 44662 4520 44714
rect 4464 44660 4520 44662
rect 4568 44714 4624 44716
rect 4568 44662 4570 44714
rect 4570 44662 4622 44714
rect 4622 44662 4624 44714
rect 4568 44660 4624 44662
rect 4672 44714 4728 44716
rect 4672 44662 4674 44714
rect 4674 44662 4726 44714
rect 4726 44662 4728 44714
rect 4672 44660 4728 44662
rect 4284 43484 4340 43540
rect 4956 43708 5012 43764
rect 4464 43146 4520 43148
rect 4464 43094 4466 43146
rect 4466 43094 4518 43146
rect 4518 43094 4520 43146
rect 4464 43092 4520 43094
rect 4568 43146 4624 43148
rect 4568 43094 4570 43146
rect 4570 43094 4622 43146
rect 4622 43094 4624 43146
rect 4568 43092 4624 43094
rect 4672 43146 4728 43148
rect 4672 43094 4674 43146
rect 4674 43094 4726 43146
rect 4726 43094 4728 43146
rect 4672 43092 4728 43094
rect 3804 42362 3860 42364
rect 3804 42310 3806 42362
rect 3806 42310 3858 42362
rect 3858 42310 3860 42362
rect 3804 42308 3860 42310
rect 3908 42362 3964 42364
rect 3908 42310 3910 42362
rect 3910 42310 3962 42362
rect 3962 42310 3964 42362
rect 3908 42308 3964 42310
rect 4012 42362 4068 42364
rect 4012 42310 4014 42362
rect 4014 42310 4066 42362
rect 4066 42310 4068 42362
rect 4012 42308 4068 42310
rect 4172 41970 4228 41972
rect 4172 41918 4174 41970
rect 4174 41918 4226 41970
rect 4226 41918 4228 41970
rect 4172 41916 4228 41918
rect 4172 41356 4228 41412
rect 4396 41916 4452 41972
rect 4284 41804 4340 41860
rect 3804 40794 3860 40796
rect 3804 40742 3806 40794
rect 3806 40742 3858 40794
rect 3858 40742 3860 40794
rect 3804 40740 3860 40742
rect 3908 40794 3964 40796
rect 3908 40742 3910 40794
rect 3910 40742 3962 40794
rect 3962 40742 3964 40794
rect 3908 40740 3964 40742
rect 4012 40794 4068 40796
rect 4012 40742 4014 40794
rect 4014 40742 4066 40794
rect 4066 40742 4068 40794
rect 4012 40740 4068 40742
rect 3804 39226 3860 39228
rect 3804 39174 3806 39226
rect 3806 39174 3858 39226
rect 3858 39174 3860 39226
rect 3804 39172 3860 39174
rect 3908 39226 3964 39228
rect 3908 39174 3910 39226
rect 3910 39174 3962 39226
rect 3962 39174 3964 39226
rect 3908 39172 3964 39174
rect 4012 39226 4068 39228
rect 4012 39174 4014 39226
rect 4014 39174 4066 39226
rect 4066 39174 4068 39226
rect 4012 39172 4068 39174
rect 4956 41970 5012 41972
rect 4956 41918 4958 41970
rect 4958 41918 5010 41970
rect 5010 41918 5012 41970
rect 4956 41916 5012 41918
rect 4464 41578 4520 41580
rect 4464 41526 4466 41578
rect 4466 41526 4518 41578
rect 4518 41526 4520 41578
rect 4464 41524 4520 41526
rect 4568 41578 4624 41580
rect 4568 41526 4570 41578
rect 4570 41526 4622 41578
rect 4622 41526 4624 41578
rect 4568 41524 4624 41526
rect 4672 41578 4728 41580
rect 4672 41526 4674 41578
rect 4674 41526 4726 41578
rect 4726 41526 4728 41578
rect 4672 41524 4728 41526
rect 4396 41410 4452 41412
rect 4396 41358 4398 41410
rect 4398 41358 4450 41410
rect 4450 41358 4452 41410
rect 4396 41356 4452 41358
rect 4844 41186 4900 41188
rect 4844 41134 4846 41186
rect 4846 41134 4898 41186
rect 4898 41134 4900 41186
rect 4844 41132 4900 41134
rect 5068 41692 5124 41748
rect 4464 40010 4520 40012
rect 4464 39958 4466 40010
rect 4466 39958 4518 40010
rect 4518 39958 4520 40010
rect 4464 39956 4520 39958
rect 4568 40010 4624 40012
rect 4568 39958 4570 40010
rect 4570 39958 4622 40010
rect 4622 39958 4624 40010
rect 4568 39956 4624 39958
rect 4672 40010 4728 40012
rect 4672 39958 4674 40010
rect 4674 39958 4726 40010
rect 4726 39958 4728 40010
rect 4672 39956 4728 39958
rect 4956 40236 5012 40292
rect 5404 47458 5460 47460
rect 5404 47406 5406 47458
rect 5406 47406 5458 47458
rect 5458 47406 5460 47458
rect 5404 47404 5460 47406
rect 5292 45836 5348 45892
rect 5292 45500 5348 45556
rect 5852 49026 5908 49028
rect 5852 48974 5854 49026
rect 5854 48974 5906 49026
rect 5906 48974 5908 49026
rect 5852 48972 5908 48974
rect 6076 50594 6132 50596
rect 6076 50542 6078 50594
rect 6078 50542 6130 50594
rect 6130 50542 6132 50594
rect 6076 50540 6132 50542
rect 6636 56866 6692 56868
rect 6636 56814 6638 56866
rect 6638 56814 6690 56866
rect 6690 56814 6692 56866
rect 6636 56812 6692 56814
rect 6972 70700 7028 70756
rect 7420 72322 7476 72324
rect 7420 72270 7422 72322
rect 7422 72270 7474 72322
rect 7474 72270 7476 72322
rect 7420 72268 7476 72270
rect 7756 73276 7812 73332
rect 8428 83804 8484 83860
rect 8316 82738 8372 82740
rect 8316 82686 8318 82738
rect 8318 82686 8370 82738
rect 8370 82686 8372 82738
rect 8316 82684 8372 82686
rect 8316 82460 8372 82516
rect 8316 82236 8372 82292
rect 8540 82124 8596 82180
rect 8540 81004 8596 81060
rect 9660 104466 9716 104468
rect 9660 104414 9662 104466
rect 9662 104414 9714 104466
rect 9714 104414 9716 104466
rect 9660 104412 9716 104414
rect 9772 103740 9828 103796
rect 9324 103122 9380 103124
rect 9324 103070 9326 103122
rect 9326 103070 9378 103122
rect 9378 103070 9380 103122
rect 9324 103068 9380 103070
rect 9660 102508 9716 102564
rect 9548 100828 9604 100884
rect 9436 100156 9492 100212
rect 9548 100492 9604 100548
rect 9324 99986 9380 99988
rect 9324 99934 9326 99986
rect 9326 99934 9378 99986
rect 9378 99934 9380 99986
rect 9324 99932 9380 99934
rect 9548 99820 9604 99876
rect 9660 99596 9716 99652
rect 9660 99260 9716 99316
rect 9212 97580 9268 97636
rect 9548 98140 9604 98196
rect 8764 94780 8820 94836
rect 8876 95676 8932 95732
rect 8876 93996 8932 94052
rect 8764 93436 8820 93492
rect 8988 95228 9044 95284
rect 9100 94892 9156 94948
rect 8876 93042 8932 93044
rect 8876 92990 8878 93042
rect 8878 92990 8930 93042
rect 8930 92990 8932 93042
rect 8876 92988 8932 92990
rect 8764 92876 8820 92932
rect 9324 93884 9380 93940
rect 9324 93436 9380 93492
rect 9548 95282 9604 95284
rect 9548 95230 9550 95282
rect 9550 95230 9602 95282
rect 9602 95230 9604 95282
rect 9548 95228 9604 95230
rect 9884 100770 9940 100772
rect 9884 100718 9886 100770
rect 9886 100718 9938 100770
rect 9938 100718 9940 100770
rect 9884 100716 9940 100718
rect 10108 103628 10164 103684
rect 10556 102898 10612 102900
rect 10556 102846 10558 102898
rect 10558 102846 10610 102898
rect 10610 102846 10612 102898
rect 10556 102844 10612 102846
rect 10668 102508 10724 102564
rect 10780 105980 10836 106036
rect 10780 103628 10836 103684
rect 10444 101836 10500 101892
rect 10108 101442 10164 101444
rect 10108 101390 10110 101442
rect 10110 101390 10162 101442
rect 10162 101390 10164 101442
rect 10108 101388 10164 101390
rect 10108 101052 10164 101108
rect 9996 100156 10052 100212
rect 9884 99708 9940 99764
rect 10332 100828 10388 100884
rect 10332 100156 10388 100212
rect 10220 99932 10276 99988
rect 10108 98476 10164 98532
rect 9996 97356 10052 97412
rect 9884 95228 9940 95284
rect 9996 95564 10052 95620
rect 9548 93602 9604 93604
rect 9548 93550 9550 93602
rect 9550 93550 9602 93602
rect 9602 93550 9604 93602
rect 9548 93548 9604 93550
rect 9324 92316 9380 92372
rect 8764 91868 8820 91924
rect 8988 89010 9044 89012
rect 8988 88958 8990 89010
rect 8990 88958 9042 89010
rect 9042 88958 9044 89010
rect 8988 88956 9044 88958
rect 8988 88732 9044 88788
rect 8876 85708 8932 85764
rect 8988 85036 9044 85092
rect 8876 84306 8932 84308
rect 8876 84254 8878 84306
rect 8878 84254 8930 84306
rect 8930 84254 8932 84306
rect 8876 84252 8932 84254
rect 8876 83634 8932 83636
rect 8876 83582 8878 83634
rect 8878 83582 8930 83634
rect 8930 83582 8932 83634
rect 8876 83580 8932 83582
rect 8876 83356 8932 83412
rect 8764 82796 8820 82852
rect 8652 79772 8708 79828
rect 9100 84588 9156 84644
rect 9436 92204 9492 92260
rect 9324 89852 9380 89908
rect 9324 88956 9380 89012
rect 9212 83522 9268 83524
rect 9212 83470 9214 83522
rect 9214 83470 9266 83522
rect 9266 83470 9268 83522
rect 9212 83468 9268 83470
rect 9100 81340 9156 81396
rect 9212 83244 9268 83300
rect 8764 79602 8820 79604
rect 8764 79550 8766 79602
rect 8766 79550 8818 79602
rect 8818 79550 8820 79602
rect 8764 79548 8820 79550
rect 8428 79436 8484 79492
rect 9100 79772 9156 79828
rect 9436 87276 9492 87332
rect 9436 85932 9492 85988
rect 9660 92930 9716 92932
rect 9660 92878 9662 92930
rect 9662 92878 9714 92930
rect 9714 92878 9716 92930
rect 9660 92876 9716 92878
rect 9660 92204 9716 92260
rect 10108 95340 10164 95396
rect 10668 100156 10724 100212
rect 10668 99986 10724 99988
rect 10668 99934 10670 99986
rect 10670 99934 10722 99986
rect 10722 99934 10724 99986
rect 10668 99932 10724 99934
rect 10556 99708 10612 99764
rect 11004 104748 11060 104804
rect 10892 102226 10948 102228
rect 10892 102174 10894 102226
rect 10894 102174 10946 102226
rect 10946 102174 10948 102226
rect 10892 102172 10948 102174
rect 11116 104466 11172 104468
rect 11116 104414 11118 104466
rect 11118 104414 11170 104466
rect 11170 104414 11172 104466
rect 11116 104412 11172 104414
rect 11788 107324 11844 107380
rect 11564 106428 11620 106484
rect 11788 106540 11844 106596
rect 11452 104748 11508 104804
rect 11340 104412 11396 104468
rect 11004 102060 11060 102116
rect 11004 101052 11060 101108
rect 11452 103852 11508 103908
rect 11116 100828 11172 100884
rect 11228 103628 11284 103684
rect 11676 104412 11732 104468
rect 12012 107548 12068 107604
rect 11900 104076 11956 104132
rect 11676 103852 11732 103908
rect 13692 113426 13748 113428
rect 13692 113374 13694 113426
rect 13694 113374 13746 113426
rect 13746 113374 13748 113426
rect 13692 113372 13748 113374
rect 13468 112028 13524 112084
rect 12908 111020 12964 111076
rect 13132 111804 13188 111860
rect 12460 110460 12516 110516
rect 13020 110684 13076 110740
rect 12908 110066 12964 110068
rect 12908 110014 12910 110066
rect 12910 110014 12962 110066
rect 12962 110014 12964 110066
rect 12908 110012 12964 110014
rect 12908 109676 12964 109732
rect 13020 109452 13076 109508
rect 12908 109004 12964 109060
rect 12796 107548 12852 107604
rect 12684 107266 12740 107268
rect 12684 107214 12686 107266
rect 12686 107214 12738 107266
rect 12738 107214 12740 107266
rect 12684 107212 12740 107214
rect 12348 104524 12404 104580
rect 13692 111804 13748 111860
rect 13692 111580 13748 111636
rect 13244 111356 13300 111412
rect 13244 110124 13300 110180
rect 13580 110962 13636 110964
rect 13580 110910 13582 110962
rect 13582 110910 13634 110962
rect 13634 110910 13636 110962
rect 13580 110908 13636 110910
rect 13692 110796 13748 110852
rect 13580 110684 13636 110740
rect 13244 109564 13300 109620
rect 13468 109506 13524 109508
rect 13468 109454 13470 109506
rect 13470 109454 13522 109506
rect 13522 109454 13524 109506
rect 13468 109452 13524 109454
rect 13244 109004 13300 109060
rect 13580 108220 13636 108276
rect 13468 107826 13524 107828
rect 13468 107774 13470 107826
rect 13470 107774 13522 107826
rect 13522 107774 13524 107826
rect 13468 107772 13524 107774
rect 13356 107436 13412 107492
rect 13132 107324 13188 107380
rect 12012 103852 12068 103908
rect 11900 103794 11956 103796
rect 11900 103742 11902 103794
rect 11902 103742 11954 103794
rect 11954 103742 11956 103794
rect 11900 103740 11956 103742
rect 11676 103628 11732 103684
rect 12124 103628 12180 103684
rect 11564 103180 11620 103236
rect 12908 106764 12964 106820
rect 13020 106428 13076 106484
rect 13020 106258 13076 106260
rect 13020 106206 13022 106258
rect 13022 106206 13074 106258
rect 13074 106206 13076 106258
rect 13020 106204 13076 106206
rect 13356 106540 13412 106596
rect 13244 106204 13300 106260
rect 13132 105980 13188 106036
rect 13468 105980 13524 106036
rect 13132 105756 13188 105812
rect 13468 105532 13524 105588
rect 13468 104636 13524 104692
rect 13692 107714 13748 107716
rect 13692 107662 13694 107714
rect 13694 107662 13746 107714
rect 13746 107662 13748 107714
rect 13692 107660 13748 107662
rect 14140 113372 14196 113428
rect 14140 112700 14196 112756
rect 14700 113538 14756 113540
rect 14700 113486 14702 113538
rect 14702 113486 14754 113538
rect 14754 113486 14756 113538
rect 14700 113484 14756 113486
rect 14588 113372 14644 113428
rect 14588 113148 14644 113204
rect 14364 112588 14420 112644
rect 14476 112700 14532 112756
rect 14028 111244 14084 111300
rect 14476 111580 14532 111636
rect 15036 113484 15092 113540
rect 14812 112588 14868 112644
rect 14924 111858 14980 111860
rect 14924 111806 14926 111858
rect 14926 111806 14978 111858
rect 14978 111806 14980 111858
rect 14924 111804 14980 111806
rect 14252 110908 14308 110964
rect 14924 111580 14980 111636
rect 13916 110684 13972 110740
rect 13916 110460 13972 110516
rect 14028 110012 14084 110068
rect 14252 109900 14308 109956
rect 13916 109340 13972 109396
rect 13916 108610 13972 108612
rect 13916 108558 13918 108610
rect 13918 108558 13970 108610
rect 13970 108558 13972 108610
rect 13916 108556 13972 108558
rect 14028 108108 14084 108164
rect 13804 107548 13860 107604
rect 13916 107884 13972 107940
rect 14140 107772 14196 107828
rect 14028 107436 14084 107492
rect 13804 105644 13860 105700
rect 12908 103740 12964 103796
rect 13132 103682 13188 103684
rect 13132 103630 13134 103682
rect 13134 103630 13186 103682
rect 13186 103630 13188 103682
rect 13132 103628 13188 103630
rect 12908 103234 12964 103236
rect 12908 103182 12910 103234
rect 12910 103182 12962 103234
rect 12962 103182 12964 103234
rect 12908 103180 12964 103182
rect 11452 103068 11508 103124
rect 11676 103068 11732 103124
rect 11340 101052 11396 101108
rect 11228 99820 11284 99876
rect 11340 99708 11396 99764
rect 11452 99932 11508 99988
rect 11564 99372 11620 99428
rect 11004 98588 11060 98644
rect 11228 98588 11284 98644
rect 11676 99148 11732 99204
rect 10332 97244 10388 97300
rect 10556 97692 10612 97748
rect 10444 96626 10500 96628
rect 10444 96574 10446 96626
rect 10446 96574 10498 96626
rect 10498 96574 10500 96626
rect 10444 96572 10500 96574
rect 10332 96012 10388 96068
rect 10444 95676 10500 95732
rect 10892 96796 10948 96852
rect 11340 97356 11396 97412
rect 11564 96850 11620 96852
rect 11564 96798 11566 96850
rect 11566 96798 11618 96850
rect 11618 96798 11620 96850
rect 11564 96796 11620 96798
rect 11452 96290 11508 96292
rect 11452 96238 11454 96290
rect 11454 96238 11506 96290
rect 11506 96238 11508 96290
rect 11452 96236 11508 96238
rect 10780 95340 10836 95396
rect 9996 94108 10052 94164
rect 10332 94780 10388 94836
rect 10220 94274 10276 94276
rect 10220 94222 10222 94274
rect 10222 94222 10274 94274
rect 10274 94222 10276 94274
rect 10220 94220 10276 94222
rect 10444 93884 10500 93940
rect 10332 92988 10388 93044
rect 9660 90188 9716 90244
rect 9660 89122 9716 89124
rect 9660 89070 9662 89122
rect 9662 89070 9714 89122
rect 9714 89070 9716 89122
rect 9660 89068 9716 89070
rect 10220 90412 10276 90468
rect 10108 89906 10164 89908
rect 10108 89854 10110 89906
rect 10110 89854 10162 89906
rect 10162 89854 10164 89906
rect 10108 89852 10164 89854
rect 9660 84306 9716 84308
rect 9660 84254 9662 84306
rect 9662 84254 9714 84306
rect 9714 84254 9716 84306
rect 9660 84252 9716 84254
rect 9660 84028 9716 84084
rect 9884 88284 9940 88340
rect 9884 84140 9940 84196
rect 9996 86716 10052 86772
rect 9884 83746 9940 83748
rect 9884 83694 9886 83746
rect 9886 83694 9938 83746
rect 9938 83694 9940 83746
rect 9884 83692 9940 83694
rect 9772 83356 9828 83412
rect 9884 83468 9940 83524
rect 9324 81900 9380 81956
rect 9324 81452 9380 81508
rect 9660 81004 9716 81060
rect 8428 79100 8484 79156
rect 8316 78876 8372 78932
rect 8316 78092 8372 78148
rect 8540 78988 8596 79044
rect 8540 77756 8596 77812
rect 8092 76188 8148 76244
rect 8204 75682 8260 75684
rect 8204 75630 8206 75682
rect 8206 75630 8258 75682
rect 8258 75630 8260 75682
rect 8204 75628 8260 75630
rect 8204 75180 8260 75236
rect 8428 77532 8484 77588
rect 7980 74114 8036 74116
rect 7980 74062 7982 74114
rect 7982 74062 8034 74114
rect 8034 74062 8036 74114
rect 7980 74060 8036 74062
rect 8204 73388 8260 73444
rect 7756 72492 7812 72548
rect 7756 71484 7812 71540
rect 7756 71036 7812 71092
rect 8316 73164 8372 73220
rect 8092 72268 8148 72324
rect 7868 69916 7924 69972
rect 8092 71484 8148 71540
rect 8092 70082 8148 70084
rect 8092 70030 8094 70082
rect 8094 70030 8146 70082
rect 8146 70030 8148 70082
rect 8092 70028 8148 70030
rect 7308 69186 7364 69188
rect 7308 69134 7310 69186
rect 7310 69134 7362 69186
rect 7362 69134 7364 69186
rect 7308 69132 7364 69134
rect 7308 68796 7364 68852
rect 7756 68514 7812 68516
rect 7756 68462 7758 68514
rect 7758 68462 7810 68514
rect 7810 68462 7812 68514
rect 7756 68460 7812 68462
rect 7084 67228 7140 67284
rect 7644 67340 7700 67396
rect 6972 67170 7028 67172
rect 6972 67118 6974 67170
rect 6974 67118 7026 67170
rect 7026 67118 7028 67170
rect 6972 67116 7028 67118
rect 6972 66780 7028 66836
rect 7308 67004 7364 67060
rect 7308 66668 7364 66724
rect 6972 61516 7028 61572
rect 7532 64540 7588 64596
rect 7420 62914 7476 62916
rect 7420 62862 7422 62914
rect 7422 62862 7474 62914
rect 7474 62862 7476 62914
rect 7420 62860 7476 62862
rect 7644 63756 7700 63812
rect 7196 58492 7252 58548
rect 7756 57820 7812 57876
rect 6860 56252 6916 56308
rect 6636 56140 6692 56196
rect 6524 55298 6580 55300
rect 6524 55246 6526 55298
rect 6526 55246 6578 55298
rect 6578 55246 6580 55298
rect 6524 55244 6580 55246
rect 6636 54796 6692 54852
rect 6300 54348 6356 54404
rect 6300 53900 6356 53956
rect 6636 53788 6692 53844
rect 6300 53116 6356 53172
rect 6412 52668 6468 52724
rect 6188 48860 6244 48916
rect 5964 48188 6020 48244
rect 6412 47964 6468 48020
rect 6748 53730 6804 53732
rect 6748 53678 6750 53730
rect 6750 53678 6802 53730
rect 6802 53678 6804 53730
rect 6748 53676 6804 53678
rect 6636 52556 6692 52612
rect 6972 53676 7028 53732
rect 6972 52946 7028 52948
rect 6972 52894 6974 52946
rect 6974 52894 7026 52946
rect 7026 52894 7028 52946
rect 6972 52892 7028 52894
rect 6636 52108 6692 52164
rect 6636 49532 6692 49588
rect 6860 52162 6916 52164
rect 6860 52110 6862 52162
rect 6862 52110 6914 52162
rect 6914 52110 6916 52162
rect 6860 52108 6916 52110
rect 6748 48972 6804 49028
rect 6860 51212 6916 51268
rect 6860 50876 6916 50932
rect 6636 48242 6692 48244
rect 6636 48190 6638 48242
rect 6638 48190 6690 48242
rect 6690 48190 6692 48242
rect 6636 48188 6692 48190
rect 6076 47346 6132 47348
rect 6076 47294 6078 47346
rect 6078 47294 6130 47346
rect 6130 47294 6132 47346
rect 6076 47292 6132 47294
rect 5852 46674 5908 46676
rect 5852 46622 5854 46674
rect 5854 46622 5906 46674
rect 5906 46622 5908 46674
rect 5852 46620 5908 46622
rect 5852 45388 5908 45444
rect 5516 44994 5572 44996
rect 5516 44942 5518 44994
rect 5518 44942 5570 44994
rect 5570 44942 5572 44994
rect 5516 44940 5572 44942
rect 5628 44882 5684 44884
rect 5628 44830 5630 44882
rect 5630 44830 5682 44882
rect 5682 44830 5684 44882
rect 5628 44828 5684 44830
rect 6188 45500 6244 45556
rect 5964 45164 6020 45220
rect 6076 44994 6132 44996
rect 6076 44942 6078 44994
rect 6078 44942 6130 44994
rect 6130 44942 6132 44994
rect 6076 44940 6132 44942
rect 5740 43036 5796 43092
rect 5852 42924 5908 42980
rect 6524 47570 6580 47572
rect 6524 47518 6526 47570
rect 6526 47518 6578 47570
rect 6578 47518 6580 47570
rect 6524 47516 6580 47518
rect 6636 47292 6692 47348
rect 6748 46956 6804 47012
rect 6076 42140 6132 42196
rect 5852 42028 5908 42084
rect 5740 41970 5796 41972
rect 5740 41918 5742 41970
rect 5742 41918 5794 41970
rect 5794 41918 5796 41970
rect 5740 41916 5796 41918
rect 5292 41356 5348 41412
rect 5628 41186 5684 41188
rect 5628 41134 5630 41186
rect 5630 41134 5682 41186
rect 5682 41134 5684 41186
rect 5628 41132 5684 41134
rect 5180 40402 5236 40404
rect 5180 40350 5182 40402
rect 5182 40350 5234 40402
rect 5234 40350 5236 40402
rect 5180 40348 5236 40350
rect 4956 39618 5012 39620
rect 4956 39566 4958 39618
rect 4958 39566 5010 39618
rect 5010 39566 5012 39618
rect 4956 39564 5012 39566
rect 4844 38780 4900 38836
rect 4284 38668 4340 38724
rect 4464 38442 4520 38444
rect 4464 38390 4466 38442
rect 4466 38390 4518 38442
rect 4518 38390 4520 38442
rect 4464 38388 4520 38390
rect 4568 38442 4624 38444
rect 4568 38390 4570 38442
rect 4570 38390 4622 38442
rect 4622 38390 4624 38442
rect 4568 38388 4624 38390
rect 4672 38442 4728 38444
rect 4672 38390 4674 38442
rect 4674 38390 4726 38442
rect 4726 38390 4728 38442
rect 4672 38388 4728 38390
rect 5180 38220 5236 38276
rect 3804 37658 3860 37660
rect 3804 37606 3806 37658
rect 3806 37606 3858 37658
rect 3858 37606 3860 37658
rect 3804 37604 3860 37606
rect 3908 37658 3964 37660
rect 3908 37606 3910 37658
rect 3910 37606 3962 37658
rect 3962 37606 3964 37658
rect 3908 37604 3964 37606
rect 4012 37658 4068 37660
rect 4012 37606 4014 37658
rect 4014 37606 4066 37658
rect 4066 37606 4068 37658
rect 4012 37604 4068 37606
rect 5404 39228 5460 39284
rect 5964 41746 6020 41748
rect 5964 41694 5966 41746
rect 5966 41694 6018 41746
rect 6018 41694 6020 41746
rect 5964 41692 6020 41694
rect 6188 39788 6244 39844
rect 6076 39452 6132 39508
rect 6188 38780 6244 38836
rect 5516 38556 5572 38612
rect 6076 38722 6132 38724
rect 6076 38670 6078 38722
rect 6078 38670 6130 38722
rect 6130 38670 6132 38722
rect 6076 38668 6132 38670
rect 5292 37772 5348 37828
rect 5740 38444 5796 38500
rect 5180 37212 5236 37268
rect 4464 36874 4520 36876
rect 4464 36822 4466 36874
rect 4466 36822 4518 36874
rect 4518 36822 4520 36874
rect 4464 36820 4520 36822
rect 4568 36874 4624 36876
rect 4568 36822 4570 36874
rect 4570 36822 4622 36874
rect 4622 36822 4624 36874
rect 4568 36820 4624 36822
rect 4672 36874 4728 36876
rect 4672 36822 4674 36874
rect 4674 36822 4726 36874
rect 4726 36822 4728 36874
rect 4672 36820 4728 36822
rect 4284 36652 4340 36708
rect 3804 36090 3860 36092
rect 3804 36038 3806 36090
rect 3806 36038 3858 36090
rect 3858 36038 3860 36090
rect 3804 36036 3860 36038
rect 3908 36090 3964 36092
rect 3908 36038 3910 36090
rect 3910 36038 3962 36090
rect 3962 36038 3964 36090
rect 3908 36036 3964 36038
rect 4012 36090 4068 36092
rect 4012 36038 4014 36090
rect 4014 36038 4066 36090
rect 4066 36038 4068 36090
rect 4012 36036 4068 36038
rect 3500 35756 3556 35812
rect 3052 31724 3108 31780
rect 3164 35196 3220 35252
rect 2940 31612 2996 31668
rect 3948 35196 4004 35252
rect 3388 34972 3444 35028
rect 3948 34972 4004 35028
rect 2380 24220 2436 24276
rect 2716 24220 2772 24276
rect 1596 22988 1652 23044
rect 2268 24108 2324 24164
rect 1596 20860 1652 20916
rect 1708 20972 1764 21028
rect 1708 20412 1764 20468
rect 1148 20130 1204 20132
rect 1148 20078 1150 20130
rect 1150 20078 1202 20130
rect 1202 20078 1204 20130
rect 1148 20076 1204 20078
rect 1596 20300 1652 20356
rect 1260 19346 1316 19348
rect 1260 19294 1262 19346
rect 1262 19294 1314 19346
rect 1314 19294 1316 19346
rect 1260 19292 1316 19294
rect 1932 23826 1988 23828
rect 1932 23774 1934 23826
rect 1934 23774 1986 23826
rect 1986 23774 1988 23826
rect 1932 23772 1988 23774
rect 2044 21420 2100 21476
rect 2156 21644 2212 21700
rect 2156 20412 2212 20468
rect 1932 20076 1988 20132
rect 1932 19404 1988 19460
rect 2156 19794 2212 19796
rect 2156 19742 2158 19794
rect 2158 19742 2210 19794
rect 2210 19742 2212 19794
rect 2156 19740 2212 19742
rect 2716 23660 2772 23716
rect 2604 22482 2660 22484
rect 2604 22430 2606 22482
rect 2606 22430 2658 22482
rect 2658 22430 2660 22482
rect 2604 22428 2660 22430
rect 2604 21644 2660 21700
rect 2716 21532 2772 21588
rect 2940 24050 2996 24052
rect 2940 23998 2942 24050
rect 2942 23998 2994 24050
rect 2994 23998 2996 24050
rect 2940 23996 2996 23998
rect 3836 34748 3892 34804
rect 5628 37772 5684 37828
rect 6076 38444 6132 38500
rect 5852 37660 5908 37716
rect 5628 37324 5684 37380
rect 4508 35756 4564 35812
rect 5516 36988 5572 37044
rect 5180 35756 5236 35812
rect 4464 35306 4520 35308
rect 4464 35254 4466 35306
rect 4466 35254 4518 35306
rect 4518 35254 4520 35306
rect 4464 35252 4520 35254
rect 4568 35306 4624 35308
rect 4568 35254 4570 35306
rect 4570 35254 4622 35306
rect 4622 35254 4624 35306
rect 4568 35252 4624 35254
rect 4672 35306 4728 35308
rect 4672 35254 4674 35306
rect 4674 35254 4726 35306
rect 4726 35254 4728 35306
rect 4672 35252 4728 35254
rect 4172 34636 4228 34692
rect 3804 34522 3860 34524
rect 3612 34412 3668 34468
rect 3804 34470 3806 34522
rect 3806 34470 3858 34522
rect 3858 34470 3860 34522
rect 3804 34468 3860 34470
rect 3908 34522 3964 34524
rect 3908 34470 3910 34522
rect 3910 34470 3962 34522
rect 3962 34470 3964 34522
rect 3908 34468 3964 34470
rect 4012 34522 4068 34524
rect 4012 34470 4014 34522
rect 4014 34470 4066 34522
rect 4066 34470 4068 34522
rect 4012 34468 4068 34470
rect 3500 34076 3556 34132
rect 3724 34076 3780 34132
rect 4172 33852 4228 33908
rect 3948 33740 4004 33796
rect 4732 34914 4788 34916
rect 4732 34862 4734 34914
rect 4734 34862 4786 34914
rect 4786 34862 4788 34914
rect 4732 34860 4788 34862
rect 4464 33738 4520 33740
rect 4464 33686 4466 33738
rect 4466 33686 4518 33738
rect 4518 33686 4520 33738
rect 4464 33684 4520 33686
rect 4568 33738 4624 33740
rect 4568 33686 4570 33738
rect 4570 33686 4622 33738
rect 4622 33686 4624 33738
rect 4568 33684 4624 33686
rect 4672 33738 4728 33740
rect 4672 33686 4674 33738
rect 4674 33686 4726 33738
rect 4726 33686 4728 33738
rect 4672 33684 4728 33686
rect 4284 33516 4340 33572
rect 3612 33458 3668 33460
rect 3612 33406 3614 33458
rect 3614 33406 3666 33458
rect 3666 33406 3668 33458
rect 3612 33404 3668 33406
rect 3388 33346 3444 33348
rect 3388 33294 3390 33346
rect 3390 33294 3442 33346
rect 3442 33294 3444 33346
rect 3388 33292 3444 33294
rect 4284 33346 4340 33348
rect 4284 33294 4286 33346
rect 4286 33294 4338 33346
rect 4338 33294 4340 33346
rect 4284 33292 4340 33294
rect 5068 34802 5124 34804
rect 5068 34750 5070 34802
rect 5070 34750 5122 34802
rect 5122 34750 5124 34802
rect 5068 34748 5124 34750
rect 5292 34748 5348 34804
rect 5516 34914 5572 34916
rect 5516 34862 5518 34914
rect 5518 34862 5570 34914
rect 5570 34862 5572 34914
rect 5516 34860 5572 34862
rect 5404 34636 5460 34692
rect 5068 34076 5124 34132
rect 4956 33852 5012 33908
rect 3804 32954 3860 32956
rect 3804 32902 3806 32954
rect 3806 32902 3858 32954
rect 3858 32902 3860 32954
rect 3804 32900 3860 32902
rect 3908 32954 3964 32956
rect 3908 32902 3910 32954
rect 3910 32902 3962 32954
rect 3962 32902 3964 32954
rect 3908 32900 3964 32902
rect 4012 32954 4068 32956
rect 4012 32902 4014 32954
rect 4014 32902 4066 32954
rect 4066 32902 4068 32954
rect 4012 32900 4068 32902
rect 4464 32170 4520 32172
rect 4464 32118 4466 32170
rect 4466 32118 4518 32170
rect 4518 32118 4520 32170
rect 4464 32116 4520 32118
rect 4568 32170 4624 32172
rect 4568 32118 4570 32170
rect 4570 32118 4622 32170
rect 4622 32118 4624 32170
rect 4568 32116 4624 32118
rect 4672 32170 4728 32172
rect 4672 32118 4674 32170
rect 4674 32118 4726 32170
rect 4726 32118 4728 32170
rect 4672 32116 4728 32118
rect 4844 31836 4900 31892
rect 3804 31386 3860 31388
rect 3804 31334 3806 31386
rect 3806 31334 3858 31386
rect 3858 31334 3860 31386
rect 3804 31332 3860 31334
rect 3908 31386 3964 31388
rect 3908 31334 3910 31386
rect 3910 31334 3962 31386
rect 3962 31334 3964 31386
rect 3908 31332 3964 31334
rect 4012 31386 4068 31388
rect 4012 31334 4014 31386
rect 4014 31334 4066 31386
rect 4066 31334 4068 31386
rect 4012 31332 4068 31334
rect 4464 30602 4520 30604
rect 4464 30550 4466 30602
rect 4466 30550 4518 30602
rect 4518 30550 4520 30602
rect 4464 30548 4520 30550
rect 4568 30602 4624 30604
rect 4568 30550 4570 30602
rect 4570 30550 4622 30602
rect 4622 30550 4624 30602
rect 4568 30548 4624 30550
rect 4672 30602 4728 30604
rect 4672 30550 4674 30602
rect 4674 30550 4726 30602
rect 4726 30550 4728 30602
rect 4672 30548 4728 30550
rect 3612 30380 3668 30436
rect 3388 29932 3444 29988
rect 3276 27858 3332 27860
rect 3276 27806 3278 27858
rect 3278 27806 3330 27858
rect 3330 27806 3332 27858
rect 3276 27804 3332 27806
rect 3164 26012 3220 26068
rect 3164 25228 3220 25284
rect 3164 22930 3220 22932
rect 3164 22878 3166 22930
rect 3166 22878 3218 22930
rect 3218 22878 3220 22930
rect 3164 22876 3220 22878
rect 4172 30156 4228 30212
rect 3804 29818 3860 29820
rect 3804 29766 3806 29818
rect 3806 29766 3858 29818
rect 3858 29766 3860 29818
rect 3804 29764 3860 29766
rect 3908 29818 3964 29820
rect 3908 29766 3910 29818
rect 3910 29766 3962 29818
rect 3962 29766 3964 29818
rect 3908 29764 3964 29766
rect 4012 29818 4068 29820
rect 4012 29766 4014 29818
rect 4014 29766 4066 29818
rect 4066 29766 4068 29818
rect 4012 29764 4068 29766
rect 3804 28250 3860 28252
rect 3804 28198 3806 28250
rect 3806 28198 3858 28250
rect 3858 28198 3860 28250
rect 3804 28196 3860 28198
rect 3908 28250 3964 28252
rect 3908 28198 3910 28250
rect 3910 28198 3962 28250
rect 3962 28198 3964 28250
rect 3908 28196 3964 28198
rect 4012 28250 4068 28252
rect 4012 28198 4014 28250
rect 4014 28198 4066 28250
rect 4066 28198 4068 28250
rect 4012 28196 4068 28198
rect 3948 27804 4004 27860
rect 3724 27244 3780 27300
rect 3948 27020 4004 27076
rect 4172 27020 4228 27076
rect 3804 26682 3860 26684
rect 3804 26630 3806 26682
rect 3806 26630 3858 26682
rect 3858 26630 3860 26682
rect 3804 26628 3860 26630
rect 3908 26682 3964 26684
rect 3908 26630 3910 26682
rect 3910 26630 3962 26682
rect 3962 26630 3964 26682
rect 3908 26628 3964 26630
rect 4012 26682 4068 26684
rect 4012 26630 4014 26682
rect 4014 26630 4066 26682
rect 4066 26630 4068 26682
rect 4012 26628 4068 26630
rect 4172 26348 4228 26404
rect 3724 25676 3780 25732
rect 5068 33292 5124 33348
rect 4956 30156 5012 30212
rect 5068 30380 5124 30436
rect 4464 29034 4520 29036
rect 4464 28982 4466 29034
rect 4466 28982 4518 29034
rect 4518 28982 4520 29034
rect 4464 28980 4520 28982
rect 4568 29034 4624 29036
rect 4568 28982 4570 29034
rect 4570 28982 4622 29034
rect 4622 28982 4624 29034
rect 4568 28980 4624 28982
rect 4672 29034 4728 29036
rect 4672 28982 4674 29034
rect 4674 28982 4726 29034
rect 4726 28982 4728 29034
rect 4672 28980 4728 28982
rect 4464 27466 4520 27468
rect 4464 27414 4466 27466
rect 4466 27414 4518 27466
rect 4518 27414 4520 27466
rect 4464 27412 4520 27414
rect 4568 27466 4624 27468
rect 4568 27414 4570 27466
rect 4570 27414 4622 27466
rect 4622 27414 4624 27466
rect 4568 27412 4624 27414
rect 4672 27466 4728 27468
rect 4672 27414 4674 27466
rect 4674 27414 4726 27466
rect 4726 27414 4728 27466
rect 4672 27412 4728 27414
rect 4508 27074 4564 27076
rect 4508 27022 4510 27074
rect 4510 27022 4562 27074
rect 4562 27022 4564 27074
rect 4508 27020 4564 27022
rect 5180 26796 5236 26852
rect 5740 37100 5796 37156
rect 6076 37660 6132 37716
rect 6188 37772 6244 37828
rect 5628 34076 5684 34132
rect 5964 37548 6020 37604
rect 5628 33852 5684 33908
rect 5516 33516 5572 33572
rect 5852 35084 5908 35140
rect 5852 34636 5908 34692
rect 6524 45890 6580 45892
rect 6524 45838 6526 45890
rect 6526 45838 6578 45890
rect 6578 45838 6580 45890
rect 6524 45836 6580 45838
rect 6636 45612 6692 45668
rect 7084 50594 7140 50596
rect 7084 50542 7086 50594
rect 7086 50542 7138 50594
rect 7138 50542 7140 50594
rect 7084 50540 7140 50542
rect 6972 49644 7028 49700
rect 6972 47292 7028 47348
rect 7084 48636 7140 48692
rect 7084 48130 7140 48132
rect 7084 48078 7086 48130
rect 7086 48078 7138 48130
rect 7138 48078 7140 48130
rect 7084 48076 7140 48078
rect 6972 47068 7028 47124
rect 7532 53564 7588 53620
rect 7420 49586 7476 49588
rect 7420 49534 7422 49586
rect 7422 49534 7474 49586
rect 7474 49534 7476 49586
rect 7420 49532 7476 49534
rect 7980 68348 8036 68404
rect 8204 69580 8260 69636
rect 8316 72380 8372 72436
rect 8092 68012 8148 68068
rect 7980 63362 8036 63364
rect 7980 63310 7982 63362
rect 7982 63310 8034 63362
rect 8034 63310 8036 63362
rect 7980 63308 8036 63310
rect 8316 64764 8372 64820
rect 8204 64706 8260 64708
rect 8204 64654 8206 64706
rect 8206 64654 8258 64706
rect 8258 64654 8260 64706
rect 8204 64652 8260 64654
rect 8204 64146 8260 64148
rect 8204 64094 8206 64146
rect 8206 64094 8258 64146
rect 8258 64094 8260 64146
rect 8204 64092 8260 64094
rect 8540 75628 8596 75684
rect 9100 78204 9156 78260
rect 9436 79378 9492 79380
rect 9436 79326 9438 79378
rect 9438 79326 9490 79378
rect 9490 79326 9492 79378
rect 9436 79324 9492 79326
rect 9548 78930 9604 78932
rect 9548 78878 9550 78930
rect 9550 78878 9602 78930
rect 9602 78878 9604 78930
rect 9548 78876 9604 78878
rect 9324 78540 9380 78596
rect 8988 77644 9044 77700
rect 8876 76466 8932 76468
rect 8876 76414 8878 76466
rect 8878 76414 8930 76466
rect 8930 76414 8932 76466
rect 8876 76412 8932 76414
rect 8876 72828 8932 72884
rect 9884 79996 9940 80052
rect 10220 86380 10276 86436
rect 10108 84700 10164 84756
rect 10108 84364 10164 84420
rect 11116 95282 11172 95284
rect 11116 95230 11118 95282
rect 11118 95230 11170 95282
rect 11170 95230 11172 95282
rect 11116 95228 11172 95230
rect 10780 93996 10836 94052
rect 10892 94556 10948 94612
rect 11004 94108 11060 94164
rect 10780 93714 10836 93716
rect 10780 93662 10782 93714
rect 10782 93662 10834 93714
rect 10834 93662 10836 93714
rect 10780 93660 10836 93662
rect 10668 93212 10724 93268
rect 10780 93324 10836 93380
rect 10892 92930 10948 92932
rect 10892 92878 10894 92930
rect 10894 92878 10946 92930
rect 10946 92878 10948 92930
rect 10892 92876 10948 92878
rect 10892 91474 10948 91476
rect 10892 91422 10894 91474
rect 10894 91422 10946 91474
rect 10946 91422 10948 91474
rect 10892 91420 10948 91422
rect 10556 89068 10612 89124
rect 10556 84364 10612 84420
rect 10332 83522 10388 83524
rect 10332 83470 10334 83522
rect 10334 83470 10386 83522
rect 10386 83470 10388 83522
rect 10332 83468 10388 83470
rect 10220 82684 10276 82740
rect 10108 82460 10164 82516
rect 10108 82124 10164 82180
rect 10332 82460 10388 82516
rect 9660 78428 9716 78484
rect 9436 78146 9492 78148
rect 9436 78094 9438 78146
rect 9438 78094 9490 78146
rect 9490 78094 9492 78146
rect 9436 78092 9492 78094
rect 9548 77980 9604 78036
rect 9660 77644 9716 77700
rect 9772 77868 9828 77924
rect 9548 77532 9604 77588
rect 9436 77420 9492 77476
rect 9324 77196 9380 77252
rect 9548 77250 9604 77252
rect 9548 77198 9550 77250
rect 9550 77198 9602 77250
rect 9602 77198 9604 77250
rect 9548 77196 9604 77198
rect 10332 80892 10388 80948
rect 10220 80444 10276 80500
rect 10108 79324 10164 79380
rect 10108 78204 10164 78260
rect 9884 76412 9940 76468
rect 9884 74060 9940 74116
rect 9548 73836 9604 73892
rect 9324 73500 9380 73556
rect 9324 73052 9380 73108
rect 9212 72828 9268 72884
rect 9100 72322 9156 72324
rect 9100 72270 9102 72322
rect 9102 72270 9154 72322
rect 9154 72270 9156 72322
rect 9100 72268 9156 72270
rect 8988 71820 9044 71876
rect 8876 71372 8932 71428
rect 9436 72492 9492 72548
rect 9772 73330 9828 73332
rect 9772 73278 9774 73330
rect 9774 73278 9826 73330
rect 9826 73278 9828 73330
rect 9772 73276 9828 73278
rect 11900 99372 11956 99428
rect 11788 97916 11844 97972
rect 12684 102396 12740 102452
rect 12460 101836 12516 101892
rect 12348 100828 12404 100884
rect 12124 99986 12180 99988
rect 12124 99934 12126 99986
rect 12126 99934 12178 99986
rect 12178 99934 12180 99986
rect 12124 99932 12180 99934
rect 12124 97244 12180 97300
rect 11676 96124 11732 96180
rect 11228 93660 11284 93716
rect 11564 93714 11620 93716
rect 11564 93662 11566 93714
rect 11566 93662 11618 93714
rect 11618 93662 11620 93714
rect 11564 93660 11620 93662
rect 12012 96796 12068 96852
rect 12236 94668 12292 94724
rect 11900 94556 11956 94612
rect 11676 92988 11732 93044
rect 11788 92652 11844 92708
rect 11900 93660 11956 93716
rect 11900 92428 11956 92484
rect 11116 90354 11172 90356
rect 11116 90302 11118 90354
rect 11118 90302 11170 90354
rect 11170 90302 11172 90354
rect 11116 90300 11172 90302
rect 12124 91362 12180 91364
rect 12124 91310 12126 91362
rect 12126 91310 12178 91362
rect 12178 91310 12180 91362
rect 12124 91308 12180 91310
rect 11900 90860 11956 90916
rect 11676 90188 11732 90244
rect 11228 89570 11284 89572
rect 11228 89518 11230 89570
rect 11230 89518 11282 89570
rect 11282 89518 11284 89570
rect 11228 89516 11284 89518
rect 11788 89516 11844 89572
rect 11116 88956 11172 89012
rect 11452 88338 11508 88340
rect 11452 88286 11454 88338
rect 11454 88286 11506 88338
rect 11506 88286 11508 88338
rect 11452 88284 11508 88286
rect 11452 87500 11508 87556
rect 11004 87276 11060 87332
rect 11228 87388 11284 87444
rect 11564 87388 11620 87444
rect 11340 86828 11396 86884
rect 11004 86658 11060 86660
rect 11004 86606 11006 86658
rect 11006 86606 11058 86658
rect 11058 86606 11060 86658
rect 11004 86604 11060 86606
rect 11340 86268 11396 86324
rect 11004 86044 11060 86100
rect 10892 85260 10948 85316
rect 11004 82908 11060 82964
rect 11116 85932 11172 85988
rect 11228 85202 11284 85204
rect 11228 85150 11230 85202
rect 11230 85150 11282 85202
rect 11282 85150 11284 85202
rect 11228 85148 11284 85150
rect 10556 82460 10612 82516
rect 11004 82348 11060 82404
rect 11116 81900 11172 81956
rect 11228 84588 11284 84644
rect 10668 81452 10724 81508
rect 10556 80108 10612 80164
rect 10444 79772 10500 79828
rect 10780 80946 10836 80948
rect 10780 80894 10782 80946
rect 10782 80894 10834 80946
rect 10834 80894 10836 80946
rect 10780 80892 10836 80894
rect 10892 79884 10948 79940
rect 10332 79324 10388 79380
rect 10780 78652 10836 78708
rect 11340 84418 11396 84420
rect 11340 84366 11342 84418
rect 11342 84366 11394 84418
rect 11394 84366 11396 84418
rect 11340 84364 11396 84366
rect 11452 84924 11508 84980
rect 11228 80556 11284 80612
rect 11340 83132 11396 83188
rect 11228 78876 11284 78932
rect 10892 78316 10948 78372
rect 11228 78652 11284 78708
rect 11228 78316 11284 78372
rect 10444 78204 10500 78260
rect 10220 76300 10276 76356
rect 11452 79884 11508 79940
rect 11452 79660 11508 79716
rect 11452 79042 11508 79044
rect 11452 78990 11454 79042
rect 11454 78990 11506 79042
rect 11506 78990 11508 79042
rect 11452 78988 11508 78990
rect 11452 78594 11508 78596
rect 11452 78542 11454 78594
rect 11454 78542 11506 78594
rect 11506 78542 11508 78594
rect 11452 78540 11508 78542
rect 11340 78204 11396 78260
rect 11788 86658 11844 86660
rect 11788 86606 11790 86658
rect 11790 86606 11842 86658
rect 11842 86606 11844 86658
rect 11788 86604 11844 86606
rect 12124 90524 12180 90580
rect 12236 90076 12292 90132
rect 12012 85820 12068 85876
rect 12572 99148 12628 99204
rect 13244 101836 13300 101892
rect 12908 101500 12964 101556
rect 13132 100156 13188 100212
rect 12908 99202 12964 99204
rect 12908 99150 12910 99202
rect 12910 99150 12962 99202
rect 12962 99150 12964 99202
rect 12908 99148 12964 99150
rect 13020 98588 13076 98644
rect 13020 97468 13076 97524
rect 12460 96066 12516 96068
rect 12460 96014 12462 96066
rect 12462 96014 12514 96066
rect 12514 96014 12516 96066
rect 12460 96012 12516 96014
rect 12460 90748 12516 90804
rect 12684 97244 12740 97300
rect 12908 97244 12964 97300
rect 12796 97020 12852 97076
rect 12684 91532 12740 91588
rect 12908 96236 12964 96292
rect 12908 92428 12964 92484
rect 13356 100156 13412 100212
rect 13468 102396 13524 102452
rect 13804 105308 13860 105364
rect 13692 105196 13748 105252
rect 13692 103740 13748 103796
rect 13804 103292 13860 103348
rect 13692 102508 13748 102564
rect 14028 106428 14084 106484
rect 13580 101554 13636 101556
rect 13580 101502 13582 101554
rect 13582 101502 13634 101554
rect 13634 101502 13636 101554
rect 13580 101500 13636 101502
rect 13468 99820 13524 99876
rect 13244 95788 13300 95844
rect 13580 101276 13636 101332
rect 13692 100828 13748 100884
rect 13468 96124 13524 96180
rect 13132 93660 13188 93716
rect 13468 93996 13524 94052
rect 13916 102450 13972 102452
rect 13916 102398 13918 102450
rect 13918 102398 13970 102450
rect 13970 102398 13972 102450
rect 13916 102396 13972 102398
rect 14588 110908 14644 110964
rect 14476 110684 14532 110740
rect 14476 109340 14532 109396
rect 15148 113260 15204 113316
rect 15372 114156 15428 114212
rect 15260 112588 15316 112644
rect 15372 113260 15428 113316
rect 15036 111356 15092 111412
rect 15148 110962 15204 110964
rect 15148 110910 15150 110962
rect 15150 110910 15202 110962
rect 15202 110910 15204 110962
rect 15148 110908 15204 110910
rect 15036 109564 15092 109620
rect 15260 108892 15316 108948
rect 15036 107660 15092 107716
rect 14700 107548 14756 107604
rect 14364 107436 14420 107492
rect 14812 107436 14868 107492
rect 14588 106930 14644 106932
rect 14588 106878 14590 106930
rect 14590 106878 14642 106930
rect 14642 106878 14644 106930
rect 14588 106876 14644 106878
rect 14364 105196 14420 105252
rect 14252 104972 14308 105028
rect 14700 103794 14756 103796
rect 14700 103742 14702 103794
rect 14702 103742 14754 103794
rect 14754 103742 14756 103794
rect 14700 103740 14756 103742
rect 14140 103180 14196 103236
rect 14140 101612 14196 101668
rect 14028 100828 14084 100884
rect 13916 100156 13972 100212
rect 14140 99932 14196 99988
rect 14028 99372 14084 99428
rect 14252 100716 14308 100772
rect 14588 102338 14644 102340
rect 14588 102286 14590 102338
rect 14590 102286 14642 102338
rect 14642 102286 14644 102338
rect 14588 102284 14644 102286
rect 14476 100156 14532 100212
rect 14364 98028 14420 98084
rect 13692 96850 13748 96852
rect 13692 96798 13694 96850
rect 13694 96798 13746 96850
rect 13746 96798 13748 96850
rect 13692 96796 13748 96798
rect 13468 93436 13524 93492
rect 13580 93212 13636 93268
rect 13580 92876 13636 92932
rect 13020 90636 13076 90692
rect 13244 91308 13300 91364
rect 12796 90466 12852 90468
rect 12796 90414 12798 90466
rect 12798 90414 12850 90466
rect 12850 90414 12852 90466
rect 12796 90412 12852 90414
rect 13132 90466 13188 90468
rect 13132 90414 13134 90466
rect 13134 90414 13186 90466
rect 13186 90414 13188 90466
rect 13132 90412 13188 90414
rect 12572 89906 12628 89908
rect 12572 89854 12574 89906
rect 12574 89854 12626 89906
rect 12626 89854 12628 89906
rect 12572 89852 12628 89854
rect 13468 90300 13524 90356
rect 13580 90188 13636 90244
rect 13356 90076 13412 90132
rect 13916 96908 13972 96964
rect 13916 96236 13972 96292
rect 14028 95788 14084 95844
rect 14140 95170 14196 95172
rect 14140 95118 14142 95170
rect 14142 95118 14194 95170
rect 14194 95118 14196 95170
rect 14140 95116 14196 95118
rect 13916 94332 13972 94388
rect 13916 94108 13972 94164
rect 14140 93996 14196 94052
rect 14028 93324 14084 93380
rect 13916 92428 13972 92484
rect 14028 91196 14084 91252
rect 13804 91084 13860 91140
rect 13916 90300 13972 90356
rect 13692 89740 13748 89796
rect 13020 89122 13076 89124
rect 13020 89070 13022 89122
rect 13022 89070 13074 89122
rect 13074 89070 13076 89122
rect 13020 89068 13076 89070
rect 13356 88620 13412 88676
rect 12684 88172 12740 88228
rect 13244 88226 13300 88228
rect 13244 88174 13246 88226
rect 13246 88174 13298 88226
rect 13298 88174 13300 88226
rect 13244 88172 13300 88174
rect 12460 86770 12516 86772
rect 12460 86718 12462 86770
rect 12462 86718 12514 86770
rect 12514 86718 12516 86770
rect 12460 86716 12516 86718
rect 11676 78930 11732 78932
rect 11676 78878 11678 78930
rect 11678 78878 11730 78930
rect 11730 78878 11732 78930
rect 11676 78876 11732 78878
rect 11676 78652 11732 78708
rect 10556 77868 10612 77924
rect 10556 76076 10612 76132
rect 10668 74060 10724 74116
rect 10220 73442 10276 73444
rect 10220 73390 10222 73442
rect 10222 73390 10274 73442
rect 10274 73390 10276 73442
rect 10220 73388 10276 73390
rect 10668 73890 10724 73892
rect 10668 73838 10670 73890
rect 10670 73838 10722 73890
rect 10722 73838 10724 73890
rect 10668 73836 10724 73838
rect 10556 73612 10612 73668
rect 10892 77196 10948 77252
rect 11676 77308 11732 77364
rect 10892 76354 10948 76356
rect 10892 76302 10894 76354
rect 10894 76302 10946 76354
rect 10946 76302 10948 76354
rect 10892 76300 10948 76302
rect 11228 76300 11284 76356
rect 11004 75068 11060 75124
rect 10780 73500 10836 73556
rect 11452 74060 11508 74116
rect 10780 73218 10836 73220
rect 10780 73166 10782 73218
rect 10782 73166 10834 73218
rect 10834 73166 10836 73218
rect 10780 73164 10836 73166
rect 9324 72434 9380 72436
rect 9324 72382 9326 72434
rect 9326 72382 9378 72434
rect 9378 72382 9380 72434
rect 9324 72380 9380 72382
rect 9772 72380 9828 72436
rect 10108 72380 10164 72436
rect 10108 72156 10164 72212
rect 9100 70476 9156 70532
rect 8876 69244 8932 69300
rect 8652 67116 8708 67172
rect 8988 67004 9044 67060
rect 9436 68402 9492 68404
rect 9436 68350 9438 68402
rect 9438 68350 9490 68402
rect 9490 68350 9492 68402
rect 9436 68348 9492 68350
rect 9772 70754 9828 70756
rect 9772 70702 9774 70754
rect 9774 70702 9826 70754
rect 9826 70702 9828 70754
rect 9772 70700 9828 70702
rect 9772 69916 9828 69972
rect 9324 67564 9380 67620
rect 8540 65436 8596 65492
rect 8876 65548 8932 65604
rect 8428 63756 8484 63812
rect 8764 63980 8820 64036
rect 9324 65490 9380 65492
rect 9324 65438 9326 65490
rect 9326 65438 9378 65490
rect 9378 65438 9380 65490
rect 9324 65436 9380 65438
rect 9548 67004 9604 67060
rect 9660 66780 9716 66836
rect 9996 69970 10052 69972
rect 9996 69918 9998 69970
rect 9998 69918 10050 69970
rect 10050 69918 10052 69970
rect 9996 69916 10052 69918
rect 9996 69468 10052 69524
rect 9996 68908 10052 68964
rect 9884 67004 9940 67060
rect 9996 67116 10052 67172
rect 8988 61740 9044 61796
rect 8764 59724 8820 59780
rect 8316 58716 8372 58772
rect 8540 57708 8596 57764
rect 8092 56812 8148 56868
rect 8988 56924 9044 56980
rect 7644 50540 7700 50596
rect 7980 54460 8036 54516
rect 9212 64988 9268 65044
rect 9324 64706 9380 64708
rect 9324 64654 9326 64706
rect 9326 64654 9378 64706
rect 9378 64654 9380 64706
rect 9324 64652 9380 64654
rect 9996 64988 10052 65044
rect 9996 64818 10052 64820
rect 9996 64766 9998 64818
rect 9998 64766 10050 64818
rect 10050 64766 10052 64818
rect 9996 64764 10052 64766
rect 9548 63868 9604 63924
rect 9324 63810 9380 63812
rect 9324 63758 9326 63810
rect 9326 63758 9378 63810
rect 9378 63758 9380 63810
rect 9324 63756 9380 63758
rect 9884 63756 9940 63812
rect 9884 63420 9940 63476
rect 9212 61404 9268 61460
rect 9436 61740 9492 61796
rect 9548 61068 9604 61124
rect 9996 62524 10052 62580
rect 9996 61852 10052 61908
rect 9884 59948 9940 60004
rect 9436 59836 9492 59892
rect 9436 59164 9492 59220
rect 10108 59836 10164 59892
rect 9324 58716 9380 58772
rect 10108 58716 10164 58772
rect 9996 58156 10052 58212
rect 9548 56924 9604 56980
rect 8764 54514 8820 54516
rect 8764 54462 8766 54514
rect 8766 54462 8818 54514
rect 8818 54462 8820 54514
rect 8764 54460 8820 54462
rect 8204 53788 8260 53844
rect 8092 52946 8148 52948
rect 8092 52894 8094 52946
rect 8094 52894 8146 52946
rect 8146 52894 8148 52946
rect 8092 52892 8148 52894
rect 7532 48636 7588 48692
rect 7756 48972 7812 49028
rect 7196 48300 7252 48356
rect 7196 47516 7252 47572
rect 7532 46956 7588 47012
rect 7868 48188 7924 48244
rect 7756 46562 7812 46564
rect 7756 46510 7758 46562
rect 7758 46510 7810 46562
rect 7810 46510 7812 46562
rect 7756 46508 7812 46510
rect 7084 46002 7140 46004
rect 7084 45950 7086 46002
rect 7086 45950 7138 46002
rect 7138 45950 7140 46002
rect 7084 45948 7140 45950
rect 6860 45106 6916 45108
rect 6860 45054 6862 45106
rect 6862 45054 6914 45106
rect 6914 45054 6916 45106
rect 6860 45052 6916 45054
rect 7084 44434 7140 44436
rect 7084 44382 7086 44434
rect 7086 44382 7138 44434
rect 7138 44382 7140 44434
rect 7084 44380 7140 44382
rect 6860 43036 6916 43092
rect 6412 41244 6468 41300
rect 6300 37660 6356 37716
rect 6412 40124 6468 40180
rect 6188 36540 6244 36596
rect 6076 35420 6132 35476
rect 6188 35698 6244 35700
rect 6188 35646 6190 35698
rect 6190 35646 6242 35698
rect 6242 35646 6244 35698
rect 6188 35644 6244 35646
rect 6188 35084 6244 35140
rect 6076 35026 6132 35028
rect 6076 34974 6078 35026
rect 6078 34974 6130 35026
rect 6130 34974 6132 35026
rect 6076 34972 6132 34974
rect 6188 34860 6244 34916
rect 7532 45164 7588 45220
rect 7196 42924 7252 42980
rect 7196 42700 7252 42756
rect 7196 42476 7252 42532
rect 7308 41804 7364 41860
rect 6860 39564 6916 39620
rect 6412 36428 6468 36484
rect 6524 39116 6580 39172
rect 6860 38668 6916 38724
rect 6860 37772 6916 37828
rect 6636 36652 6692 36708
rect 6636 34860 6692 34916
rect 7308 40012 7364 40068
rect 7084 39116 7140 39172
rect 7196 37826 7252 37828
rect 7196 37774 7198 37826
rect 7198 37774 7250 37826
rect 7250 37774 7252 37826
rect 7196 37772 7252 37774
rect 7308 37100 7364 37156
rect 7420 37548 7476 37604
rect 7756 43260 7812 43316
rect 7756 42140 7812 42196
rect 7532 37324 7588 37380
rect 7196 36988 7252 37044
rect 7532 36988 7588 37044
rect 7308 36594 7364 36596
rect 7308 36542 7310 36594
rect 7310 36542 7362 36594
rect 7362 36542 7364 36594
rect 7308 36540 7364 36542
rect 7196 35868 7252 35924
rect 4464 25898 4520 25900
rect 4464 25846 4466 25898
rect 4466 25846 4518 25898
rect 4518 25846 4520 25898
rect 4464 25844 4520 25846
rect 4568 25898 4624 25900
rect 4568 25846 4570 25898
rect 4570 25846 4622 25898
rect 4622 25846 4624 25898
rect 4568 25844 4624 25846
rect 4672 25898 4728 25900
rect 4672 25846 4674 25898
rect 4674 25846 4726 25898
rect 4726 25846 4728 25898
rect 4672 25844 4728 25846
rect 5404 29260 5460 29316
rect 3612 25228 3668 25284
rect 3804 25114 3860 25116
rect 3612 25004 3668 25060
rect 3804 25062 3806 25114
rect 3806 25062 3858 25114
rect 3858 25062 3860 25114
rect 3804 25060 3860 25062
rect 3908 25114 3964 25116
rect 3908 25062 3910 25114
rect 3910 25062 3962 25114
rect 3962 25062 3964 25114
rect 3908 25060 3964 25062
rect 4012 25114 4068 25116
rect 4012 25062 4014 25114
rect 4014 25062 4066 25114
rect 4066 25062 4068 25114
rect 4284 25116 4340 25172
rect 4012 25060 4068 25062
rect 4508 25676 4564 25732
rect 4956 25564 5012 25620
rect 4508 25452 4564 25508
rect 3612 24556 3668 24612
rect 3388 24108 3444 24164
rect 3388 21644 3444 21700
rect 4060 23772 4116 23828
rect 4172 23884 4228 23940
rect 3804 23546 3860 23548
rect 3804 23494 3806 23546
rect 3806 23494 3858 23546
rect 3858 23494 3860 23546
rect 3804 23492 3860 23494
rect 3908 23546 3964 23548
rect 3908 23494 3910 23546
rect 3910 23494 3962 23546
rect 3962 23494 3964 23546
rect 3908 23492 3964 23494
rect 4012 23546 4068 23548
rect 4012 23494 4014 23546
rect 4014 23494 4066 23546
rect 4066 23494 4068 23546
rect 4012 23492 4068 23494
rect 4060 22652 4116 22708
rect 4060 22204 4116 22260
rect 3804 21978 3860 21980
rect 3804 21926 3806 21978
rect 3806 21926 3858 21978
rect 3858 21926 3860 21978
rect 3804 21924 3860 21926
rect 3908 21978 3964 21980
rect 3908 21926 3910 21978
rect 3910 21926 3962 21978
rect 3962 21926 3964 21978
rect 3908 21924 3964 21926
rect 4012 21978 4068 21980
rect 4012 21926 4014 21978
rect 4014 21926 4066 21978
rect 4066 21926 4068 21978
rect 4012 21924 4068 21926
rect 2604 20636 2660 20692
rect 2044 19180 2100 19236
rect 1596 18396 1652 18452
rect 1484 16716 1540 16772
rect 1708 18060 1764 18116
rect 812 15148 868 15204
rect 1036 15484 1092 15540
rect 924 14588 980 14644
rect 700 13244 756 13300
rect 812 12124 868 12180
rect 812 10332 868 10388
rect 700 8204 756 8260
rect 812 10108 868 10164
rect 2156 18338 2212 18340
rect 2156 18286 2158 18338
rect 2158 18286 2210 18338
rect 2210 18286 2212 18338
rect 2156 18284 2212 18286
rect 1820 17836 1876 17892
rect 2268 17612 2324 17668
rect 2156 17500 2212 17556
rect 1260 15426 1316 15428
rect 1260 15374 1262 15426
rect 1262 15374 1314 15426
rect 1314 15374 1316 15426
rect 1260 15372 1316 15374
rect 1932 15372 1988 15428
rect 1372 15260 1428 15316
rect 1260 14700 1316 14756
rect 1260 10780 1316 10836
rect 1260 10332 1316 10388
rect 1596 15202 1652 15204
rect 1596 15150 1598 15202
rect 1598 15150 1650 15202
rect 1650 15150 1652 15202
rect 1596 15148 1652 15150
rect 1820 14924 1876 14980
rect 1484 14812 1540 14868
rect 1708 14700 1764 14756
rect 1596 11564 1652 11620
rect 2044 14588 2100 14644
rect 2268 14476 2324 14532
rect 2268 13746 2324 13748
rect 2268 13694 2270 13746
rect 2270 13694 2322 13746
rect 2322 13694 2324 13746
rect 2268 13692 2324 13694
rect 2268 12908 2324 12964
rect 1820 11004 1876 11060
rect 1932 10892 1988 10948
rect 2044 11116 2100 11172
rect 1820 10108 1876 10164
rect 1932 10668 1988 10724
rect 1820 9212 1876 9268
rect 1036 8092 1092 8148
rect 1036 5346 1092 5348
rect 1036 5294 1038 5346
rect 1038 5294 1090 5346
rect 1090 5294 1092 5346
rect 1036 5292 1092 5294
rect 1036 4226 1092 4228
rect 1036 4174 1038 4226
rect 1038 4174 1090 4226
rect 1090 4174 1092 4226
rect 1036 4172 1092 4174
rect 1260 8540 1316 8596
rect 1484 8428 1540 8484
rect 1372 8258 1428 8260
rect 1372 8206 1374 8258
rect 1374 8206 1426 8258
rect 1426 8206 1428 8258
rect 1372 8204 1428 8206
rect 1372 6690 1428 6692
rect 1372 6638 1374 6690
rect 1374 6638 1426 6690
rect 1426 6638 1428 6690
rect 1372 6636 1428 6638
rect 1372 5346 1428 5348
rect 1372 5294 1374 5346
rect 1374 5294 1426 5346
rect 1426 5294 1428 5346
rect 1372 5292 1428 5294
rect 1372 4338 1428 4340
rect 1372 4286 1374 4338
rect 1374 4286 1426 4338
rect 1426 4286 1428 4338
rect 1372 4284 1428 4286
rect 2492 16268 2548 16324
rect 2492 13692 2548 13748
rect 2380 11228 2436 11284
rect 2492 12460 2548 12516
rect 2268 10050 2324 10052
rect 2268 9998 2270 10050
rect 2270 9998 2322 10050
rect 2322 9998 2324 10050
rect 2268 9996 2324 9998
rect 1708 6412 1764 6468
rect 1820 6300 1876 6356
rect 1708 5068 1764 5124
rect 1708 4226 1764 4228
rect 1708 4174 1710 4226
rect 1710 4174 1762 4226
rect 1762 4174 1764 4226
rect 1708 4172 1764 4174
rect 2268 7362 2324 7364
rect 2268 7310 2270 7362
rect 2270 7310 2322 7362
rect 2322 7310 2324 7362
rect 2268 7308 2324 7310
rect 2156 6690 2212 6692
rect 2156 6638 2158 6690
rect 2158 6638 2210 6690
rect 2210 6638 2212 6690
rect 2156 6636 2212 6638
rect 2380 6636 2436 6692
rect 2268 6188 2324 6244
rect 2156 5628 2212 5684
rect 2044 5346 2100 5348
rect 2044 5294 2046 5346
rect 2046 5294 2098 5346
rect 2098 5294 2100 5346
rect 2044 5292 2100 5294
rect 1932 4284 1988 4340
rect 2044 4396 2100 4452
rect 2044 3778 2100 3780
rect 2044 3726 2046 3778
rect 2046 3726 2098 3778
rect 2098 3726 2100 3778
rect 2044 3724 2100 3726
rect 1596 3276 1652 3332
rect 924 1820 980 1876
rect 924 700 980 756
rect 2716 19740 2772 19796
rect 2716 19234 2772 19236
rect 2716 19182 2718 19234
rect 2718 19182 2770 19234
rect 2770 19182 2772 19234
rect 2716 19180 2772 19182
rect 2716 18284 2772 18340
rect 2716 18060 2772 18116
rect 2716 17164 2772 17220
rect 2716 15484 2772 15540
rect 3164 20636 3220 20692
rect 2940 13634 2996 13636
rect 2940 13582 2942 13634
rect 2942 13582 2994 13634
rect 2994 13582 2996 13634
rect 2940 13580 2996 13582
rect 4060 21362 4116 21364
rect 4060 21310 4062 21362
rect 4062 21310 4114 21362
rect 4114 21310 4116 21362
rect 4060 21308 4116 21310
rect 4464 24330 4520 24332
rect 4464 24278 4466 24330
rect 4466 24278 4518 24330
rect 4518 24278 4520 24330
rect 4464 24276 4520 24278
rect 4568 24330 4624 24332
rect 4568 24278 4570 24330
rect 4570 24278 4622 24330
rect 4622 24278 4624 24330
rect 4568 24276 4624 24278
rect 4672 24330 4728 24332
rect 4672 24278 4674 24330
rect 4674 24278 4726 24330
rect 4726 24278 4728 24330
rect 4672 24276 4728 24278
rect 4396 23772 4452 23828
rect 4396 22988 4452 23044
rect 4464 22762 4520 22764
rect 4464 22710 4466 22762
rect 4466 22710 4518 22762
rect 4518 22710 4520 22762
rect 4464 22708 4520 22710
rect 4568 22762 4624 22764
rect 4568 22710 4570 22762
rect 4570 22710 4622 22762
rect 4622 22710 4624 22762
rect 4568 22708 4624 22710
rect 4672 22762 4728 22764
rect 4672 22710 4674 22762
rect 4674 22710 4726 22762
rect 4726 22710 4728 22762
rect 4672 22708 4728 22710
rect 4956 23938 5012 23940
rect 4956 23886 4958 23938
rect 4958 23886 5010 23938
rect 5010 23886 5012 23938
rect 4956 23884 5012 23886
rect 4956 23324 5012 23380
rect 4844 22092 4900 22148
rect 4464 21194 4520 21196
rect 4464 21142 4466 21194
rect 4466 21142 4518 21194
rect 4518 21142 4520 21194
rect 4464 21140 4520 21142
rect 4568 21194 4624 21196
rect 4568 21142 4570 21194
rect 4570 21142 4622 21194
rect 4622 21142 4624 21194
rect 4568 21140 4624 21142
rect 4672 21194 4728 21196
rect 4672 21142 4674 21194
rect 4674 21142 4726 21194
rect 4726 21142 4728 21194
rect 4672 21140 4728 21142
rect 4172 20972 4228 21028
rect 4396 20972 4452 21028
rect 3804 20410 3860 20412
rect 3804 20358 3806 20410
rect 3806 20358 3858 20410
rect 3858 20358 3860 20410
rect 3804 20356 3860 20358
rect 3908 20410 3964 20412
rect 3908 20358 3910 20410
rect 3910 20358 3962 20410
rect 3962 20358 3964 20410
rect 3908 20356 3964 20358
rect 4012 20410 4068 20412
rect 4012 20358 4014 20410
rect 4014 20358 4066 20410
rect 4066 20358 4068 20410
rect 4012 20356 4068 20358
rect 3612 20188 3668 20244
rect 3500 19740 3556 19796
rect 3388 19180 3444 19236
rect 3276 17836 3332 17892
rect 3164 17276 3220 17332
rect 3276 17164 3332 17220
rect 3388 17388 3444 17444
rect 3276 16940 3332 16996
rect 3276 16322 3332 16324
rect 3276 16270 3278 16322
rect 3278 16270 3330 16322
rect 3330 16270 3332 16322
rect 3276 16268 3332 16270
rect 3948 19234 4004 19236
rect 3948 19182 3950 19234
rect 3950 19182 4002 19234
rect 4002 19182 4004 19234
rect 3948 19180 4004 19182
rect 3612 19068 3668 19124
rect 4172 20018 4228 20020
rect 4172 19966 4174 20018
rect 4174 19966 4226 20018
rect 4226 19966 4228 20018
rect 4172 19964 4228 19966
rect 4060 18956 4116 19012
rect 3804 18842 3860 18844
rect 3804 18790 3806 18842
rect 3806 18790 3858 18842
rect 3858 18790 3860 18842
rect 3804 18788 3860 18790
rect 3908 18842 3964 18844
rect 3908 18790 3910 18842
rect 3910 18790 3962 18842
rect 3962 18790 3964 18842
rect 3908 18788 3964 18790
rect 4012 18842 4068 18844
rect 4012 18790 4014 18842
rect 4014 18790 4066 18842
rect 4066 18790 4068 18842
rect 4012 18788 4068 18790
rect 4172 18450 4228 18452
rect 4172 18398 4174 18450
rect 4174 18398 4226 18450
rect 4226 18398 4228 18450
rect 4172 18396 4228 18398
rect 4732 20524 4788 20580
rect 4396 20188 4452 20244
rect 4464 19626 4520 19628
rect 4464 19574 4466 19626
rect 4466 19574 4518 19626
rect 4518 19574 4520 19626
rect 4464 19572 4520 19574
rect 4568 19626 4624 19628
rect 4568 19574 4570 19626
rect 4570 19574 4622 19626
rect 4622 19574 4624 19626
rect 4568 19572 4624 19574
rect 4672 19626 4728 19628
rect 4672 19574 4674 19626
rect 4674 19574 4726 19626
rect 4726 19574 4728 19626
rect 4672 19572 4728 19574
rect 4464 18058 4520 18060
rect 4464 18006 4466 18058
rect 4466 18006 4518 18058
rect 4518 18006 4520 18058
rect 4464 18004 4520 18006
rect 4568 18058 4624 18060
rect 4568 18006 4570 18058
rect 4570 18006 4622 18058
rect 4622 18006 4624 18058
rect 4568 18004 4624 18006
rect 4672 18058 4728 18060
rect 4672 18006 4674 18058
rect 4674 18006 4726 18058
rect 4726 18006 4728 18058
rect 4672 18004 4728 18006
rect 4956 21084 5012 21140
rect 5292 25676 5348 25732
rect 5180 25618 5236 25620
rect 5180 25566 5182 25618
rect 5182 25566 5234 25618
rect 5234 25566 5236 25618
rect 5180 25564 5236 25566
rect 5180 25116 5236 25172
rect 5180 23772 5236 23828
rect 5068 20524 5124 20580
rect 5180 22988 5236 23044
rect 4956 20188 5012 20244
rect 5740 30210 5796 30212
rect 5740 30158 5742 30210
rect 5742 30158 5794 30210
rect 5794 30158 5796 30210
rect 5740 30156 5796 30158
rect 5628 28252 5684 28308
rect 5628 25676 5684 25732
rect 5740 25564 5796 25620
rect 5628 25452 5684 25508
rect 5628 22930 5684 22932
rect 5628 22878 5630 22930
rect 5630 22878 5682 22930
rect 5682 22878 5684 22930
rect 5628 22876 5684 22878
rect 5404 21644 5460 21700
rect 5404 20018 5460 20020
rect 5404 19966 5406 20018
rect 5406 19966 5458 20018
rect 5458 19966 5460 20018
rect 5404 19964 5460 19966
rect 5068 19628 5124 19684
rect 4956 18226 5012 18228
rect 4956 18174 4958 18226
rect 4958 18174 5010 18226
rect 5010 18174 5012 18226
rect 4956 18172 5012 18174
rect 3612 17724 3668 17780
rect 3948 17554 4004 17556
rect 3948 17502 3950 17554
rect 3950 17502 4002 17554
rect 4002 17502 4004 17554
rect 3948 17500 4004 17502
rect 3804 17274 3860 17276
rect 3804 17222 3806 17274
rect 3806 17222 3858 17274
rect 3858 17222 3860 17274
rect 3804 17220 3860 17222
rect 3908 17274 3964 17276
rect 3908 17222 3910 17274
rect 3910 17222 3962 17274
rect 3962 17222 3964 17274
rect 3908 17220 3964 17222
rect 4012 17274 4068 17276
rect 4012 17222 4014 17274
rect 4014 17222 4066 17274
rect 4066 17222 4068 17274
rect 4012 17220 4068 17222
rect 4284 17778 4340 17780
rect 4284 17726 4286 17778
rect 4286 17726 4338 17778
rect 4338 17726 4340 17778
rect 4284 17724 4340 17726
rect 4284 17164 4340 17220
rect 4844 16828 4900 16884
rect 4464 16490 4520 16492
rect 4464 16438 4466 16490
rect 4466 16438 4518 16490
rect 4518 16438 4520 16490
rect 4464 16436 4520 16438
rect 4568 16490 4624 16492
rect 4568 16438 4570 16490
rect 4570 16438 4622 16490
rect 4622 16438 4624 16490
rect 4568 16436 4624 16438
rect 4672 16490 4728 16492
rect 4672 16438 4674 16490
rect 4674 16438 4726 16490
rect 4726 16438 4728 16490
rect 4672 16436 4728 16438
rect 3612 16156 3668 16212
rect 3804 15706 3860 15708
rect 3804 15654 3806 15706
rect 3806 15654 3858 15706
rect 3858 15654 3860 15706
rect 3804 15652 3860 15654
rect 3908 15706 3964 15708
rect 3908 15654 3910 15706
rect 3910 15654 3962 15706
rect 3962 15654 3964 15706
rect 3908 15652 3964 15654
rect 4012 15706 4068 15708
rect 4012 15654 4014 15706
rect 4014 15654 4066 15706
rect 4066 15654 4068 15706
rect 4012 15652 4068 15654
rect 4284 16098 4340 16100
rect 4284 16046 4286 16098
rect 4286 16046 4338 16098
rect 4338 16046 4340 16098
rect 4284 16044 4340 16046
rect 4172 15372 4228 15428
rect 4060 15260 4116 15316
rect 2828 12796 2884 12852
rect 3164 13804 3220 13860
rect 2828 11228 2884 11284
rect 2716 10780 2772 10836
rect 2716 10220 2772 10276
rect 2492 5068 2548 5124
rect 2604 10108 2660 10164
rect 2716 9042 2772 9044
rect 2716 8990 2718 9042
rect 2718 8990 2770 9042
rect 2770 8990 2772 9042
rect 2716 8988 2772 8990
rect 2828 7644 2884 7700
rect 2940 8652 2996 8708
rect 2716 5682 2772 5684
rect 2716 5630 2718 5682
rect 2718 5630 2770 5682
rect 2770 5630 2772 5682
rect 2716 5628 2772 5630
rect 2716 5346 2772 5348
rect 2716 5294 2718 5346
rect 2718 5294 2770 5346
rect 2770 5294 2772 5346
rect 2716 5292 2772 5294
rect 2716 4620 2772 4676
rect 2604 4172 2660 4228
rect 3500 13746 3556 13748
rect 3500 13694 3502 13746
rect 3502 13694 3554 13746
rect 3554 13694 3556 13746
rect 3500 13692 3556 13694
rect 3388 13522 3444 13524
rect 3388 13470 3390 13522
rect 3390 13470 3442 13522
rect 3442 13470 3444 13522
rect 3388 13468 3444 13470
rect 3724 14642 3780 14644
rect 3724 14590 3726 14642
rect 3726 14590 3778 14642
rect 3778 14590 3780 14642
rect 3724 14588 3780 14590
rect 3836 14530 3892 14532
rect 3836 14478 3838 14530
rect 3838 14478 3890 14530
rect 3890 14478 3892 14530
rect 3836 14476 3892 14478
rect 3804 14138 3860 14140
rect 3804 14086 3806 14138
rect 3806 14086 3858 14138
rect 3858 14086 3860 14138
rect 3804 14084 3860 14086
rect 3908 14138 3964 14140
rect 3908 14086 3910 14138
rect 3910 14086 3962 14138
rect 3962 14086 3964 14138
rect 3908 14084 3964 14086
rect 4012 14138 4068 14140
rect 4012 14086 4014 14138
rect 4014 14086 4066 14138
rect 4066 14086 4068 14138
rect 4012 14084 4068 14086
rect 4060 13804 4116 13860
rect 3948 13692 4004 13748
rect 3500 12124 3556 12180
rect 3276 10892 3332 10948
rect 3500 10780 3556 10836
rect 3804 12570 3860 12572
rect 3804 12518 3806 12570
rect 3806 12518 3858 12570
rect 3858 12518 3860 12570
rect 3804 12516 3860 12518
rect 3908 12570 3964 12572
rect 3908 12518 3910 12570
rect 3910 12518 3962 12570
rect 3962 12518 3964 12570
rect 3908 12516 3964 12518
rect 4012 12570 4068 12572
rect 4012 12518 4014 12570
rect 4014 12518 4066 12570
rect 4066 12518 4068 12570
rect 4012 12516 4068 12518
rect 5852 25228 5908 25284
rect 5852 23826 5908 23828
rect 5852 23774 5854 23826
rect 5854 23774 5906 23826
rect 5906 23774 5908 23826
rect 5852 23772 5908 23774
rect 6188 31052 6244 31108
rect 6076 30716 6132 30772
rect 6188 29314 6244 29316
rect 6188 29262 6190 29314
rect 6190 29262 6242 29314
rect 6242 29262 6244 29314
rect 6188 29260 6244 29262
rect 6412 32732 6468 32788
rect 6972 34300 7028 34356
rect 6860 32338 6916 32340
rect 6860 32286 6862 32338
rect 6862 32286 6914 32338
rect 6914 32286 6916 32338
rect 6860 32284 6916 32286
rect 6636 31948 6692 32004
rect 6748 30994 6804 30996
rect 6748 30942 6750 30994
rect 6750 30942 6802 30994
rect 6802 30942 6804 30994
rect 6748 30940 6804 30942
rect 6524 30268 6580 30324
rect 6636 30210 6692 30212
rect 6636 30158 6638 30210
rect 6638 30158 6690 30210
rect 6690 30158 6692 30210
rect 6636 30156 6692 30158
rect 6188 26460 6244 26516
rect 6300 28812 6356 28868
rect 6636 27746 6692 27748
rect 6636 27694 6638 27746
rect 6638 27694 6690 27746
rect 6690 27694 6692 27746
rect 6636 27692 6692 27694
rect 7084 33068 7140 33124
rect 7420 35420 7476 35476
rect 7196 31948 7252 32004
rect 7532 34860 7588 34916
rect 7196 30940 7252 30996
rect 7420 34412 7476 34468
rect 7420 32060 7476 32116
rect 7644 34300 7700 34356
rect 7532 31164 7588 31220
rect 7420 31106 7476 31108
rect 7420 31054 7422 31106
rect 7422 31054 7474 31106
rect 7474 31054 7476 31106
rect 7420 31052 7476 31054
rect 9212 52946 9268 52948
rect 9212 52894 9214 52946
rect 9214 52894 9266 52946
rect 9266 52894 9268 52946
rect 9212 52892 9268 52894
rect 9100 52108 9156 52164
rect 8540 51436 8596 51492
rect 9324 51436 9380 51492
rect 8764 50988 8820 51044
rect 8204 45890 8260 45892
rect 8204 45838 8206 45890
rect 8206 45838 8258 45890
rect 8258 45838 8260 45890
rect 8204 45836 8260 45838
rect 8204 45106 8260 45108
rect 8204 45054 8206 45106
rect 8206 45054 8258 45106
rect 8258 45054 8260 45106
rect 8204 45052 8260 45054
rect 8092 44828 8148 44884
rect 7980 44492 8036 44548
rect 8092 44380 8148 44436
rect 7980 42140 8036 42196
rect 7868 41020 7924 41076
rect 7980 40684 8036 40740
rect 7980 40460 8036 40516
rect 7868 37548 7924 37604
rect 7868 37154 7924 37156
rect 7868 37102 7870 37154
rect 7870 37102 7922 37154
rect 7922 37102 7924 37154
rect 7868 37100 7924 37102
rect 7868 36652 7924 36708
rect 7868 34354 7924 34356
rect 7868 34302 7870 34354
rect 7870 34302 7922 34354
rect 7922 34302 7924 34354
rect 7868 34300 7924 34302
rect 8316 44268 8372 44324
rect 8204 43484 8260 43540
rect 10108 56978 10164 56980
rect 10108 56926 10110 56978
rect 10110 56926 10162 56978
rect 10162 56926 10164 56978
rect 10108 56924 10164 56926
rect 9660 56812 9716 56868
rect 10332 72770 10388 72772
rect 10332 72718 10334 72770
rect 10334 72718 10386 72770
rect 10386 72718 10388 72770
rect 10332 72716 10388 72718
rect 10332 72546 10388 72548
rect 10332 72494 10334 72546
rect 10334 72494 10386 72546
rect 10386 72494 10388 72546
rect 10332 72492 10388 72494
rect 10780 72492 10836 72548
rect 10444 70700 10500 70756
rect 10556 69020 10612 69076
rect 10444 64092 10500 64148
rect 10332 63868 10388 63924
rect 10444 62860 10500 62916
rect 10668 67228 10724 67284
rect 10892 71650 10948 71652
rect 10892 71598 10894 71650
rect 10894 71598 10946 71650
rect 10946 71598 10948 71650
rect 10892 71596 10948 71598
rect 11340 73836 11396 73892
rect 11228 73218 11284 73220
rect 11228 73166 11230 73218
rect 11230 73166 11282 73218
rect 11282 73166 11284 73218
rect 11228 73164 11284 73166
rect 11340 72940 11396 72996
rect 11004 71090 11060 71092
rect 11004 71038 11006 71090
rect 11006 71038 11058 71090
rect 11058 71038 11060 71090
rect 11004 71036 11060 71038
rect 11116 72828 11172 72884
rect 11452 72716 11508 72772
rect 11340 71874 11396 71876
rect 11340 71822 11342 71874
rect 11342 71822 11394 71874
rect 11394 71822 11396 71874
rect 11340 71820 11396 71822
rect 11340 69020 11396 69076
rect 11228 67788 11284 67844
rect 11116 67228 11172 67284
rect 10892 66892 10948 66948
rect 10780 64034 10836 64036
rect 10780 63982 10782 64034
rect 10782 63982 10834 64034
rect 10834 63982 10836 64034
rect 10780 63980 10836 63982
rect 11004 64540 11060 64596
rect 10892 63644 10948 63700
rect 10556 61292 10612 61348
rect 10556 61068 10612 61124
rect 10892 62466 10948 62468
rect 10892 62414 10894 62466
rect 10894 62414 10946 62466
rect 10946 62414 10948 62466
rect 10892 62412 10948 62414
rect 10780 60620 10836 60676
rect 11004 61852 11060 61908
rect 11116 61570 11172 61572
rect 11116 61518 11118 61570
rect 11118 61518 11170 61570
rect 11170 61518 11172 61570
rect 11116 61516 11172 61518
rect 10780 59388 10836 59444
rect 10332 58716 10388 58772
rect 10668 57932 10724 57988
rect 10444 56866 10500 56868
rect 10444 56814 10446 56866
rect 10446 56814 10498 56866
rect 10498 56814 10500 56866
rect 10444 56812 10500 56814
rect 9884 56082 9940 56084
rect 9884 56030 9886 56082
rect 9886 56030 9938 56082
rect 9938 56030 9940 56082
rect 9884 56028 9940 56030
rect 10332 56028 10388 56084
rect 8876 50204 8932 50260
rect 8988 49644 9044 49700
rect 9884 53788 9940 53844
rect 9772 53564 9828 53620
rect 10108 52834 10164 52836
rect 10108 52782 10110 52834
rect 10110 52782 10162 52834
rect 10162 52782 10164 52834
rect 10108 52780 10164 52782
rect 9772 52444 9828 52500
rect 9660 52332 9716 52388
rect 9772 52220 9828 52276
rect 9660 48748 9716 48804
rect 9548 48524 9604 48580
rect 9324 48412 9380 48468
rect 9212 47628 9268 47684
rect 8876 47180 8932 47236
rect 8988 46674 9044 46676
rect 8988 46622 8990 46674
rect 8990 46622 9042 46674
rect 9042 46622 9044 46674
rect 8988 46620 9044 46622
rect 9212 47292 9268 47348
rect 8652 43260 8708 43316
rect 8652 41970 8708 41972
rect 8652 41918 8654 41970
rect 8654 41918 8706 41970
rect 8706 41918 8708 41970
rect 8652 41916 8708 41918
rect 8428 40626 8484 40628
rect 8428 40574 8430 40626
rect 8430 40574 8482 40626
rect 8482 40574 8484 40626
rect 8428 40572 8484 40574
rect 8204 39394 8260 39396
rect 8204 39342 8206 39394
rect 8206 39342 8258 39394
rect 8258 39342 8260 39394
rect 8204 39340 8260 39342
rect 8316 39116 8372 39172
rect 8316 36482 8372 36484
rect 8316 36430 8318 36482
rect 8318 36430 8370 36482
rect 8370 36430 8372 36482
rect 8316 36428 8372 36430
rect 8876 45388 8932 45444
rect 9100 45890 9156 45892
rect 9100 45838 9102 45890
rect 9102 45838 9154 45890
rect 9154 45838 9156 45890
rect 9100 45836 9156 45838
rect 9100 44322 9156 44324
rect 9100 44270 9102 44322
rect 9102 44270 9154 44322
rect 9154 44270 9156 44322
rect 9100 44268 9156 44270
rect 10108 51996 10164 52052
rect 10220 52332 10276 52388
rect 9884 51772 9940 51828
rect 11228 57932 11284 57988
rect 11004 56924 11060 56980
rect 11004 56028 11060 56084
rect 11228 56082 11284 56084
rect 11228 56030 11230 56082
rect 11230 56030 11282 56082
rect 11282 56030 11284 56082
rect 11228 56028 11284 56030
rect 10444 51436 10500 51492
rect 10332 51324 10388 51380
rect 9884 50988 9940 51044
rect 10332 50428 10388 50484
rect 9996 48914 10052 48916
rect 9996 48862 9998 48914
rect 9998 48862 10050 48914
rect 10050 48862 10052 48914
rect 9996 48860 10052 48862
rect 10220 49644 10276 49700
rect 10220 48860 10276 48916
rect 10108 48636 10164 48692
rect 9884 48076 9940 48132
rect 10108 48412 10164 48468
rect 10220 48018 10276 48020
rect 10220 47966 10222 48018
rect 10222 47966 10274 48018
rect 10274 47966 10276 48018
rect 10220 47964 10276 47966
rect 9884 46508 9940 46564
rect 9660 46114 9716 46116
rect 9660 46062 9662 46114
rect 9662 46062 9714 46114
rect 9714 46062 9716 46114
rect 9660 46060 9716 46062
rect 9660 44828 9716 44884
rect 9884 44882 9940 44884
rect 9884 44830 9886 44882
rect 9886 44830 9938 44882
rect 9938 44830 9940 44882
rect 9884 44828 9940 44830
rect 9772 44380 9828 44436
rect 9324 44098 9380 44100
rect 9324 44046 9326 44098
rect 9326 44046 9378 44098
rect 9378 44046 9380 44098
rect 9324 44044 9380 44046
rect 9324 43820 9380 43876
rect 9772 43708 9828 43764
rect 9324 42924 9380 42980
rect 8988 42082 9044 42084
rect 8988 42030 8990 42082
rect 8990 42030 9042 42082
rect 9042 42030 9044 42082
rect 8988 42028 9044 42030
rect 9660 42476 9716 42532
rect 9324 42364 9380 42420
rect 9212 41858 9268 41860
rect 9212 41806 9214 41858
rect 9214 41806 9266 41858
rect 9266 41806 9268 41858
rect 9212 41804 9268 41806
rect 8876 38444 8932 38500
rect 8652 36316 8708 36372
rect 8092 34914 8148 34916
rect 8092 34862 8094 34914
rect 8094 34862 8146 34914
rect 8146 34862 8148 34914
rect 8092 34860 8148 34862
rect 8652 35420 8708 35476
rect 8764 37884 8820 37940
rect 8428 34860 8484 34916
rect 7980 33516 8036 33572
rect 8316 33516 8372 33572
rect 8092 33292 8148 33348
rect 7868 33234 7924 33236
rect 7868 33182 7870 33234
rect 7870 33182 7922 33234
rect 7922 33182 7924 33234
rect 7868 33180 7924 33182
rect 7980 32786 8036 32788
rect 7980 32734 7982 32786
rect 7982 32734 8034 32786
rect 8034 32734 8036 32786
rect 7980 32732 8036 32734
rect 7084 30434 7140 30436
rect 7084 30382 7086 30434
rect 7086 30382 7138 30434
rect 7138 30382 7140 30434
rect 7084 30380 7140 30382
rect 7308 30268 7364 30324
rect 6972 28700 7028 28756
rect 6748 27244 6804 27300
rect 6972 26572 7028 26628
rect 6524 25900 6580 25956
rect 6188 23884 6244 23940
rect 6412 22876 6468 22932
rect 5852 22092 5908 22148
rect 6188 22204 6244 22260
rect 5964 20636 6020 20692
rect 5852 19740 5908 19796
rect 5964 19292 6020 19348
rect 5516 18620 5572 18676
rect 5740 18956 5796 19012
rect 5628 18226 5684 18228
rect 5628 18174 5630 18226
rect 5630 18174 5682 18226
rect 5682 18174 5684 18226
rect 5628 18172 5684 18174
rect 5964 18060 6020 18116
rect 5292 17388 5348 17444
rect 5404 17612 5460 17668
rect 5404 17052 5460 17108
rect 5516 17500 5572 17556
rect 5516 16098 5572 16100
rect 5516 16046 5518 16098
rect 5518 16046 5570 16098
rect 5570 16046 5572 16098
rect 5516 16044 5572 16046
rect 4396 15372 4452 15428
rect 4844 15932 4900 15988
rect 4620 15148 4676 15204
rect 4464 14922 4520 14924
rect 4464 14870 4466 14922
rect 4466 14870 4518 14922
rect 4518 14870 4520 14922
rect 4464 14868 4520 14870
rect 4568 14922 4624 14924
rect 4568 14870 4570 14922
rect 4570 14870 4622 14922
rect 4622 14870 4624 14922
rect 4568 14868 4624 14870
rect 4672 14922 4728 14924
rect 4672 14870 4674 14922
rect 4674 14870 4726 14922
rect 4726 14870 4728 14922
rect 4672 14868 4728 14870
rect 4396 14530 4452 14532
rect 4396 14478 4398 14530
rect 4398 14478 4450 14530
rect 4450 14478 4452 14530
rect 4396 14476 4452 14478
rect 4284 14028 4340 14084
rect 4396 14140 4452 14196
rect 5068 15596 5124 15652
rect 5180 14924 5236 14980
rect 5068 14642 5124 14644
rect 5068 14590 5070 14642
rect 5070 14590 5122 14642
rect 5122 14590 5124 14642
rect 5068 14588 5124 14590
rect 4732 14140 4788 14196
rect 4844 14028 4900 14084
rect 4172 12124 4228 12180
rect 4284 13468 4340 13524
rect 4464 13354 4520 13356
rect 4464 13302 4466 13354
rect 4466 13302 4518 13354
rect 4518 13302 4520 13354
rect 4464 13300 4520 13302
rect 4568 13354 4624 13356
rect 4568 13302 4570 13354
rect 4570 13302 4622 13354
rect 4622 13302 4624 13354
rect 4568 13300 4624 13302
rect 4672 13354 4728 13356
rect 4672 13302 4674 13354
rect 4674 13302 4726 13354
rect 4726 13302 4728 13354
rect 4672 13300 4728 13302
rect 4732 12572 4788 12628
rect 4396 12460 4452 12516
rect 4464 11786 4520 11788
rect 4464 11734 4466 11786
rect 4466 11734 4518 11786
rect 4518 11734 4520 11786
rect 4464 11732 4520 11734
rect 4568 11786 4624 11788
rect 4568 11734 4570 11786
rect 4570 11734 4622 11786
rect 4622 11734 4624 11786
rect 4568 11732 4624 11734
rect 4672 11786 4728 11788
rect 4672 11734 4674 11786
rect 4674 11734 4726 11786
rect 4726 11734 4728 11786
rect 4672 11732 4728 11734
rect 4284 11564 4340 11620
rect 3804 11002 3860 11004
rect 3804 10950 3806 11002
rect 3806 10950 3858 11002
rect 3858 10950 3860 11002
rect 3804 10948 3860 10950
rect 3908 11002 3964 11004
rect 3908 10950 3910 11002
rect 3910 10950 3962 11002
rect 3962 10950 3964 11002
rect 3908 10948 3964 10950
rect 4012 11002 4068 11004
rect 4012 10950 4014 11002
rect 4014 10950 4066 11002
rect 4066 10950 4068 11002
rect 4012 10948 4068 10950
rect 3612 10668 3668 10724
rect 3164 10444 3220 10500
rect 3948 10498 4004 10500
rect 3948 10446 3950 10498
rect 3950 10446 4002 10498
rect 4002 10446 4004 10498
rect 3948 10444 4004 10446
rect 3164 9996 3220 10052
rect 3804 9434 3860 9436
rect 3804 9382 3806 9434
rect 3806 9382 3858 9434
rect 3858 9382 3860 9434
rect 3804 9380 3860 9382
rect 3908 9434 3964 9436
rect 3908 9382 3910 9434
rect 3910 9382 3962 9434
rect 3962 9382 3964 9434
rect 3908 9380 3964 9382
rect 4012 9434 4068 9436
rect 4012 9382 4014 9434
rect 4014 9382 4066 9434
rect 4066 9382 4068 9434
rect 4012 9380 4068 9382
rect 5068 13074 5124 13076
rect 5068 13022 5070 13074
rect 5070 13022 5122 13074
rect 5122 13022 5124 13074
rect 5068 13020 5124 13022
rect 4956 12236 5012 12292
rect 5292 13916 5348 13972
rect 5404 13580 5460 13636
rect 5292 11954 5348 11956
rect 5292 11902 5294 11954
rect 5294 11902 5346 11954
rect 5346 11902 5348 11954
rect 5292 11900 5348 11902
rect 4956 11394 5012 11396
rect 4956 11342 4958 11394
rect 4958 11342 5010 11394
rect 5010 11342 5012 11394
rect 4956 11340 5012 11342
rect 4844 11116 4900 11172
rect 4620 11004 4676 11060
rect 4464 10218 4520 10220
rect 4464 10166 4466 10218
rect 4466 10166 4518 10218
rect 4518 10166 4520 10218
rect 4464 10164 4520 10166
rect 4568 10218 4624 10220
rect 4568 10166 4570 10218
rect 4570 10166 4622 10218
rect 4622 10166 4624 10218
rect 4568 10164 4624 10166
rect 4672 10218 4728 10220
rect 4672 10166 4674 10218
rect 4674 10166 4726 10218
rect 4726 10166 4728 10218
rect 4672 10164 4728 10166
rect 4732 9996 4788 10052
rect 4732 9436 4788 9492
rect 4844 9660 4900 9716
rect 4396 9100 4452 9156
rect 3276 8540 3332 8596
rect 3948 8988 4004 9044
rect 3500 8258 3556 8260
rect 3500 8206 3502 8258
rect 3502 8206 3554 8258
rect 3554 8206 3556 8258
rect 3500 8204 3556 8206
rect 4284 8876 4340 8932
rect 3388 7698 3444 7700
rect 3388 7646 3390 7698
rect 3390 7646 3442 7698
rect 3442 7646 3444 7698
rect 3388 7644 3444 7646
rect 3388 6690 3444 6692
rect 3388 6638 3390 6690
rect 3390 6638 3442 6690
rect 3442 6638 3444 6690
rect 3388 6636 3444 6638
rect 3052 5628 3108 5684
rect 3388 5964 3444 6020
rect 3164 4956 3220 5012
rect 2268 3500 2324 3556
rect 1708 2156 1764 2212
rect 1820 2492 1876 2548
rect 2156 1932 2212 1988
rect 3164 3500 3220 3556
rect 3388 2994 3444 2996
rect 3388 2942 3390 2994
rect 3390 2942 3442 2994
rect 3442 2942 3444 2994
rect 3388 2940 3444 2942
rect 3388 2604 3444 2660
rect 2492 2268 2548 2324
rect 1820 1708 1876 1764
rect 3388 1708 3444 1764
rect 2268 1372 2324 1428
rect 3804 7866 3860 7868
rect 3804 7814 3806 7866
rect 3806 7814 3858 7866
rect 3858 7814 3860 7866
rect 3804 7812 3860 7814
rect 3908 7866 3964 7868
rect 3908 7814 3910 7866
rect 3910 7814 3962 7866
rect 3962 7814 3964 7866
rect 3908 7812 3964 7814
rect 4012 7866 4068 7868
rect 4012 7814 4014 7866
rect 4014 7814 4066 7866
rect 4066 7814 4068 7866
rect 4012 7812 4068 7814
rect 3948 6748 4004 6804
rect 4060 6636 4116 6692
rect 3804 6298 3860 6300
rect 3804 6246 3806 6298
rect 3806 6246 3858 6298
rect 3858 6246 3860 6298
rect 3804 6244 3860 6246
rect 3908 6298 3964 6300
rect 3908 6246 3910 6298
rect 3910 6246 3962 6298
rect 3962 6246 3964 6298
rect 3908 6244 3964 6246
rect 4012 6298 4068 6300
rect 4012 6246 4014 6298
rect 4014 6246 4066 6298
rect 4066 6246 4068 6298
rect 4012 6244 4068 6246
rect 3836 5906 3892 5908
rect 3836 5854 3838 5906
rect 3838 5854 3890 5906
rect 3890 5854 3892 5906
rect 3836 5852 3892 5854
rect 4172 5122 4228 5124
rect 4172 5070 4174 5122
rect 4174 5070 4226 5122
rect 4226 5070 4228 5122
rect 4172 5068 4228 5070
rect 3804 4730 3860 4732
rect 3804 4678 3806 4730
rect 3806 4678 3858 4730
rect 3858 4678 3860 4730
rect 3804 4676 3860 4678
rect 3908 4730 3964 4732
rect 3908 4678 3910 4730
rect 3910 4678 3962 4730
rect 3962 4678 3964 4730
rect 3908 4676 3964 4678
rect 4012 4730 4068 4732
rect 4012 4678 4014 4730
rect 4014 4678 4066 4730
rect 4066 4678 4068 4730
rect 4012 4676 4068 4678
rect 4464 8650 4520 8652
rect 4464 8598 4466 8650
rect 4466 8598 4518 8650
rect 4518 8598 4520 8650
rect 4464 8596 4520 8598
rect 4568 8650 4624 8652
rect 4568 8598 4570 8650
rect 4570 8598 4622 8650
rect 4622 8598 4624 8650
rect 4568 8596 4624 8598
rect 4672 8650 4728 8652
rect 4672 8598 4674 8650
rect 4674 8598 4726 8650
rect 4726 8598 4728 8650
rect 4672 8596 4728 8598
rect 4732 7756 4788 7812
rect 5404 11564 5460 11620
rect 5740 17612 5796 17668
rect 5964 16492 6020 16548
rect 5852 16380 5908 16436
rect 6188 19068 6244 19124
rect 6188 17948 6244 18004
rect 6188 17500 6244 17556
rect 5852 14364 5908 14420
rect 6076 15148 6132 15204
rect 6188 15090 6244 15092
rect 6188 15038 6190 15090
rect 6190 15038 6242 15090
rect 6242 15038 6244 15090
rect 6188 15036 6244 15038
rect 5964 13468 6020 13524
rect 5740 12908 5796 12964
rect 5852 12572 5908 12628
rect 6300 13580 6356 13636
rect 6076 11900 6132 11956
rect 6188 12236 6244 12292
rect 6076 11564 6132 11620
rect 5740 11282 5796 11284
rect 5740 11230 5742 11282
rect 5742 11230 5794 11282
rect 5794 11230 5796 11282
rect 5740 11228 5796 11230
rect 5628 10444 5684 10500
rect 5516 9996 5572 10052
rect 5068 8988 5124 9044
rect 5292 9042 5348 9044
rect 5292 8990 5294 9042
rect 5294 8990 5346 9042
rect 5346 8990 5348 9042
rect 5292 8988 5348 8990
rect 4956 8428 5012 8484
rect 4956 8204 5012 8260
rect 4956 7868 5012 7924
rect 4464 7082 4520 7084
rect 4464 7030 4466 7082
rect 4466 7030 4518 7082
rect 4518 7030 4520 7082
rect 4464 7028 4520 7030
rect 4568 7082 4624 7084
rect 4568 7030 4570 7082
rect 4570 7030 4622 7082
rect 4622 7030 4624 7082
rect 4568 7028 4624 7030
rect 4672 7082 4728 7084
rect 4672 7030 4674 7082
rect 4674 7030 4726 7082
rect 4726 7030 4728 7082
rect 4672 7028 4728 7030
rect 4732 6860 4788 6916
rect 5964 10498 6020 10500
rect 5964 10446 5966 10498
rect 5966 10446 6018 10498
rect 6018 10446 6020 10498
rect 5964 10444 6020 10446
rect 6076 11228 6132 11284
rect 5964 10050 6020 10052
rect 5964 9998 5966 10050
rect 5966 9998 6018 10050
rect 6018 9998 6020 10050
rect 5964 9996 6020 9998
rect 6300 12178 6356 12180
rect 6300 12126 6302 12178
rect 6302 12126 6354 12178
rect 6354 12126 6356 12178
rect 6300 12124 6356 12126
rect 6636 25452 6692 25508
rect 6748 24946 6804 24948
rect 6748 24894 6750 24946
rect 6750 24894 6802 24946
rect 6802 24894 6804 24946
rect 6748 24892 6804 24894
rect 6860 24108 6916 24164
rect 7196 25900 7252 25956
rect 7868 32060 7924 32116
rect 7532 30156 7588 30212
rect 7532 28812 7588 28868
rect 7532 26908 7588 26964
rect 7420 26572 7476 26628
rect 7308 24556 7364 24612
rect 7532 24668 7588 24724
rect 7420 24162 7476 24164
rect 7420 24110 7422 24162
rect 7422 24110 7474 24162
rect 7474 24110 7476 24162
rect 7420 24108 7476 24110
rect 6748 23378 6804 23380
rect 6748 23326 6750 23378
rect 6750 23326 6802 23378
rect 6802 23326 6804 23378
rect 6748 23324 6804 23326
rect 6860 22428 6916 22484
rect 6636 22258 6692 22260
rect 6636 22206 6638 22258
rect 6638 22206 6690 22258
rect 6690 22206 6692 22258
rect 6636 22204 6692 22206
rect 7084 22316 7140 22372
rect 6748 20018 6804 20020
rect 6748 19966 6750 20018
rect 6750 19966 6802 20018
rect 6802 19966 6804 20018
rect 6748 19964 6804 19966
rect 7308 22092 7364 22148
rect 7308 21196 7364 21252
rect 7308 20802 7364 20804
rect 7308 20750 7310 20802
rect 7310 20750 7362 20802
rect 7362 20750 7364 20802
rect 7308 20748 7364 20750
rect 8204 29986 8260 29988
rect 8204 29934 8206 29986
rect 8206 29934 8258 29986
rect 8258 29934 8260 29986
rect 8204 29932 8260 29934
rect 7868 28252 7924 28308
rect 7756 27020 7812 27076
rect 7644 23548 7700 23604
rect 7980 24892 8036 24948
rect 8092 26012 8148 26068
rect 8428 33292 8484 33348
rect 8428 33068 8484 33124
rect 8652 31052 8708 31108
rect 8428 29260 8484 29316
rect 8428 28700 8484 28756
rect 8540 27916 8596 27972
rect 8652 29932 8708 29988
rect 9212 36988 9268 37044
rect 9212 35420 9268 35476
rect 9100 35026 9156 35028
rect 9100 34974 9102 35026
rect 9102 34974 9154 35026
rect 9154 34974 9156 35026
rect 9100 34972 9156 34974
rect 8988 34300 9044 34356
rect 9212 32732 9268 32788
rect 9100 31052 9156 31108
rect 8988 30268 9044 30324
rect 9548 41692 9604 41748
rect 9436 38556 9492 38612
rect 9436 37938 9492 37940
rect 9436 37886 9438 37938
rect 9438 37886 9490 37938
rect 9490 37886 9492 37938
rect 9436 37884 9492 37886
rect 9436 37266 9492 37268
rect 9436 37214 9438 37266
rect 9438 37214 9490 37266
rect 9490 37214 9492 37266
rect 9436 37212 9492 37214
rect 10220 46732 10276 46788
rect 10220 46172 10276 46228
rect 10108 46060 10164 46116
rect 9996 43260 10052 43316
rect 10892 54402 10948 54404
rect 10892 54350 10894 54402
rect 10894 54350 10946 54402
rect 10946 54350 10948 54402
rect 10892 54348 10948 54350
rect 10892 53788 10948 53844
rect 10892 53228 10948 53284
rect 10780 52220 10836 52276
rect 10668 51772 10724 51828
rect 10892 52162 10948 52164
rect 10892 52110 10894 52162
rect 10894 52110 10946 52162
rect 10946 52110 10948 52162
rect 10892 52108 10948 52110
rect 10668 51212 10724 51268
rect 10780 50988 10836 51044
rect 10556 49644 10612 49700
rect 10444 49308 10500 49364
rect 10668 48748 10724 48804
rect 10444 47964 10500 48020
rect 10780 48242 10836 48244
rect 10780 48190 10782 48242
rect 10782 48190 10834 48242
rect 10834 48190 10836 48242
rect 10780 48188 10836 48190
rect 11116 51324 11172 51380
rect 11004 50876 11060 50932
rect 11004 50540 11060 50596
rect 11004 49756 11060 49812
rect 10444 46732 10500 46788
rect 11004 48412 11060 48468
rect 10332 45778 10388 45780
rect 10332 45726 10334 45778
rect 10334 45726 10386 45778
rect 10386 45726 10388 45778
rect 10332 45724 10388 45726
rect 10220 45052 10276 45108
rect 10444 45388 10500 45444
rect 10892 46844 10948 46900
rect 11004 46508 11060 46564
rect 11228 50764 11284 50820
rect 11228 50594 11284 50596
rect 11228 50542 11230 50594
rect 11230 50542 11282 50594
rect 11282 50542 11284 50594
rect 11228 50540 11284 50542
rect 11676 75068 11732 75124
rect 11900 84476 11956 84532
rect 12796 87724 12852 87780
rect 12460 85090 12516 85092
rect 12460 85038 12462 85090
rect 12462 85038 12514 85090
rect 12514 85038 12516 85090
rect 12460 85036 12516 85038
rect 12348 84252 12404 84308
rect 12460 84812 12516 84868
rect 11900 82348 11956 82404
rect 12012 83244 12068 83300
rect 12460 83132 12516 83188
rect 12012 82572 12068 82628
rect 12348 81116 12404 81172
rect 12236 80892 12292 80948
rect 12124 79490 12180 79492
rect 12124 79438 12126 79490
rect 12126 79438 12178 79490
rect 12178 79438 12180 79490
rect 12124 79436 12180 79438
rect 12012 78876 12068 78932
rect 12012 78428 12068 78484
rect 13132 87612 13188 87668
rect 12796 85372 12852 85428
rect 13692 88338 13748 88340
rect 13692 88286 13694 88338
rect 13694 88286 13746 88338
rect 13746 88286 13748 88338
rect 13692 88284 13748 88286
rect 13804 88060 13860 88116
rect 13468 86658 13524 86660
rect 13468 86606 13470 86658
rect 13470 86606 13522 86658
rect 13522 86606 13524 86658
rect 13468 86604 13524 86606
rect 13580 86156 13636 86212
rect 13580 85932 13636 85988
rect 13468 85820 13524 85876
rect 13244 85260 13300 85316
rect 13244 85090 13300 85092
rect 13244 85038 13246 85090
rect 13246 85038 13298 85090
rect 13298 85038 13300 85090
rect 13244 85036 13300 85038
rect 13132 84364 13188 84420
rect 13020 84194 13076 84196
rect 13020 84142 13022 84194
rect 13022 84142 13074 84194
rect 13074 84142 13076 84194
rect 13020 84140 13076 84142
rect 12572 78988 12628 79044
rect 12796 83804 12852 83860
rect 13020 83692 13076 83748
rect 13020 82460 13076 82516
rect 12908 82012 12964 82068
rect 13020 81340 13076 81396
rect 12908 81170 12964 81172
rect 12908 81118 12910 81170
rect 12910 81118 12962 81170
rect 12962 81118 12964 81170
rect 12908 81116 12964 81118
rect 12908 80610 12964 80612
rect 12908 80558 12910 80610
rect 12910 80558 12962 80610
rect 12962 80558 12964 80610
rect 12908 80556 12964 80558
rect 12908 79436 12964 79492
rect 12348 78876 12404 78932
rect 12236 78594 12292 78596
rect 12236 78542 12238 78594
rect 12238 78542 12290 78594
rect 12290 78542 12292 78594
rect 12236 78540 12292 78542
rect 12348 78316 12404 78372
rect 12572 78594 12628 78596
rect 12572 78542 12574 78594
rect 12574 78542 12626 78594
rect 12626 78542 12628 78594
rect 12572 78540 12628 78542
rect 12236 78146 12292 78148
rect 12236 78094 12238 78146
rect 12238 78094 12290 78146
rect 12290 78094 12292 78146
rect 12236 78092 12292 78094
rect 11900 76524 11956 76580
rect 12124 76466 12180 76468
rect 12124 76414 12126 76466
rect 12126 76414 12178 76466
rect 12178 76414 12180 76466
rect 12124 76412 12180 76414
rect 12348 75740 12404 75796
rect 12236 75516 12292 75572
rect 12124 74898 12180 74900
rect 12124 74846 12126 74898
rect 12126 74846 12178 74898
rect 12178 74846 12180 74898
rect 12124 74844 12180 74846
rect 12012 74732 12068 74788
rect 11788 73948 11844 74004
rect 11676 72828 11732 72884
rect 11788 72492 11844 72548
rect 11676 72380 11732 72436
rect 11900 69634 11956 69636
rect 11900 69582 11902 69634
rect 11902 69582 11954 69634
rect 11954 69582 11956 69634
rect 11900 69580 11956 69582
rect 11788 68572 11844 68628
rect 12572 75570 12628 75572
rect 12572 75518 12574 75570
rect 12574 75518 12626 75570
rect 12626 75518 12628 75570
rect 12572 75516 12628 75518
rect 13468 84364 13524 84420
rect 13244 83692 13300 83748
rect 13468 83298 13524 83300
rect 13468 83246 13470 83298
rect 13470 83246 13522 83298
rect 13522 83246 13524 83298
rect 13468 83244 13524 83246
rect 13468 82066 13524 82068
rect 13468 82014 13470 82066
rect 13470 82014 13522 82066
rect 13522 82014 13524 82066
rect 13468 82012 13524 82014
rect 13356 80668 13412 80724
rect 13468 80780 13524 80836
rect 13132 79436 13188 79492
rect 13132 78988 13188 79044
rect 13020 78204 13076 78260
rect 12236 74060 12292 74116
rect 12348 74620 12404 74676
rect 12236 73106 12292 73108
rect 12236 73054 12238 73106
rect 12238 73054 12290 73106
rect 12290 73054 12292 73106
rect 12236 73052 12292 73054
rect 12236 69410 12292 69412
rect 12236 69358 12238 69410
rect 12238 69358 12290 69410
rect 12290 69358 12292 69410
rect 12236 69356 12292 69358
rect 12460 70588 12516 70644
rect 12348 68684 12404 68740
rect 12908 76748 12964 76804
rect 12908 76578 12964 76580
rect 12908 76526 12910 76578
rect 12910 76526 12962 76578
rect 12962 76526 12964 76578
rect 12908 76524 12964 76526
rect 13468 77084 13524 77140
rect 13244 76466 13300 76468
rect 13244 76414 13246 76466
rect 13246 76414 13298 76466
rect 13298 76414 13300 76466
rect 13244 76412 13300 76414
rect 14140 89740 14196 89796
rect 13916 86492 13972 86548
rect 14028 88284 14084 88340
rect 13804 85932 13860 85988
rect 14476 97804 14532 97860
rect 14476 97522 14532 97524
rect 14476 97470 14478 97522
rect 14478 97470 14530 97522
rect 14530 97470 14532 97522
rect 14476 97468 14532 97470
rect 15148 106370 15204 106372
rect 15148 106318 15150 106370
rect 15150 106318 15202 106370
rect 15202 106318 15204 106370
rect 15148 106316 15204 106318
rect 15596 112812 15652 112868
rect 15820 111020 15876 111076
rect 16380 113260 16436 113316
rect 16380 113090 16436 113092
rect 16380 113038 16382 113090
rect 16382 113038 16434 113090
rect 16434 113038 16436 113090
rect 16380 113036 16436 113038
rect 16156 112588 16212 112644
rect 16716 112700 16772 112756
rect 15932 110572 15988 110628
rect 15820 110460 15876 110516
rect 15708 110124 15764 110180
rect 15932 110012 15988 110068
rect 15484 109676 15540 109732
rect 15372 108668 15428 108724
rect 16940 113372 16996 113428
rect 17500 113372 17556 113428
rect 17052 112588 17108 112644
rect 16828 111522 16884 111524
rect 16828 111470 16830 111522
rect 16830 111470 16882 111522
rect 16882 111470 16884 111522
rect 16828 111468 16884 111470
rect 16380 111356 16436 111412
rect 16268 110572 16324 110628
rect 16268 109788 16324 109844
rect 15372 108498 15428 108500
rect 15372 108446 15374 108498
rect 15374 108446 15426 108498
rect 15426 108446 15428 108498
rect 15372 108444 15428 108446
rect 16380 109394 16436 109396
rect 16380 109342 16382 109394
rect 16382 109342 16434 109394
rect 16434 109342 16436 109394
rect 16380 109340 16436 109342
rect 16156 108722 16212 108724
rect 16156 108670 16158 108722
rect 16158 108670 16210 108722
rect 16210 108670 16212 108722
rect 16156 108668 16212 108670
rect 15708 107996 15764 108052
rect 14924 105586 14980 105588
rect 14924 105534 14926 105586
rect 14926 105534 14978 105586
rect 14978 105534 14980 105586
rect 14924 105532 14980 105534
rect 15260 104018 15316 104020
rect 15260 103966 15262 104018
rect 15262 103966 15314 104018
rect 15314 103966 15316 104018
rect 15260 103964 15316 103966
rect 15372 103682 15428 103684
rect 15372 103630 15374 103682
rect 15374 103630 15426 103682
rect 15426 103630 15428 103682
rect 15372 103628 15428 103630
rect 14924 101554 14980 101556
rect 14924 101502 14926 101554
rect 14926 101502 14978 101554
rect 14978 101502 14980 101554
rect 14924 101500 14980 101502
rect 15820 104972 15876 105028
rect 15932 107548 15988 107604
rect 15596 103906 15652 103908
rect 15596 103854 15598 103906
rect 15598 103854 15650 103906
rect 15650 103854 15652 103906
rect 15596 103852 15652 103854
rect 15260 102284 15316 102340
rect 15260 101388 15316 101444
rect 14812 98028 14868 98084
rect 14924 101052 14980 101108
rect 14588 97132 14644 97188
rect 14924 97132 14980 97188
rect 14700 97020 14756 97076
rect 14476 93324 14532 93380
rect 14476 92930 14532 92932
rect 14476 92878 14478 92930
rect 14478 92878 14530 92930
rect 14530 92878 14532 92930
rect 14476 92876 14532 92878
rect 14364 91362 14420 91364
rect 14364 91310 14366 91362
rect 14366 91310 14418 91362
rect 14418 91310 14420 91362
rect 14364 91308 14420 91310
rect 14476 91196 14532 91252
rect 14364 90076 14420 90132
rect 14812 94892 14868 94948
rect 14700 94498 14756 94500
rect 14700 94446 14702 94498
rect 14702 94446 14754 94498
rect 14754 94446 14756 94498
rect 14700 94444 14756 94446
rect 14812 93042 14868 93044
rect 14812 92990 14814 93042
rect 14814 92990 14866 93042
rect 14866 92990 14868 93042
rect 14812 92988 14868 92990
rect 14588 90300 14644 90356
rect 14700 92652 14756 92708
rect 14476 88956 14532 89012
rect 14812 91532 14868 91588
rect 15036 96348 15092 96404
rect 16268 104412 16324 104468
rect 15932 103740 15988 103796
rect 15484 101500 15540 101556
rect 15484 98476 15540 98532
rect 15708 98700 15764 98756
rect 16044 98476 16100 98532
rect 16156 98306 16212 98308
rect 16156 98254 16158 98306
rect 16158 98254 16210 98306
rect 16210 98254 16212 98306
rect 16156 98252 16212 98254
rect 16380 97916 16436 97972
rect 15932 97468 15988 97524
rect 16380 97468 16436 97524
rect 15372 96124 15428 96180
rect 15484 96348 15540 96404
rect 15260 95900 15316 95956
rect 15148 93714 15204 93716
rect 15148 93662 15150 93714
rect 15150 93662 15202 93714
rect 15202 93662 15204 93714
rect 15148 93660 15204 93662
rect 15036 92988 15092 93044
rect 15036 92540 15092 92596
rect 15148 91922 15204 91924
rect 15148 91870 15150 91922
rect 15150 91870 15202 91922
rect 15202 91870 15204 91922
rect 15148 91868 15204 91870
rect 15260 91308 15316 91364
rect 14812 88396 14868 88452
rect 15148 90300 15204 90356
rect 14252 86156 14308 86212
rect 14364 87052 14420 87108
rect 14140 85820 14196 85876
rect 14252 85932 14308 85988
rect 13804 85596 13860 85652
rect 14028 85484 14084 85540
rect 13916 84252 13972 84308
rect 13916 84028 13972 84084
rect 13692 81116 13748 81172
rect 14028 82684 14084 82740
rect 15036 89794 15092 89796
rect 15036 89742 15038 89794
rect 15038 89742 15090 89794
rect 15090 89742 15092 89794
rect 15036 89740 15092 89742
rect 14924 88172 14980 88228
rect 14700 87442 14756 87444
rect 14700 87390 14702 87442
rect 14702 87390 14754 87442
rect 14754 87390 14756 87442
rect 14700 87388 14756 87390
rect 14364 85708 14420 85764
rect 14700 86492 14756 86548
rect 14700 85932 14756 85988
rect 14588 85762 14644 85764
rect 14588 85710 14590 85762
rect 14590 85710 14642 85762
rect 14642 85710 14644 85762
rect 14588 85708 14644 85710
rect 15036 87612 15092 87668
rect 15708 96626 15764 96628
rect 15708 96574 15710 96626
rect 15710 96574 15762 96626
rect 15762 96574 15764 96626
rect 15708 96572 15764 96574
rect 15932 96236 15988 96292
rect 15708 95900 15764 95956
rect 15820 94386 15876 94388
rect 15820 94334 15822 94386
rect 15822 94334 15874 94386
rect 15874 94334 15876 94386
rect 15820 94332 15876 94334
rect 15484 93548 15540 93604
rect 15484 93324 15540 93380
rect 15596 92258 15652 92260
rect 15596 92206 15598 92258
rect 15598 92206 15650 92258
rect 15650 92206 15652 92258
rect 15596 92204 15652 92206
rect 15484 90636 15540 90692
rect 15372 87500 15428 87556
rect 14924 87276 14980 87332
rect 15484 87388 15540 87444
rect 15148 85986 15204 85988
rect 15148 85934 15150 85986
rect 15150 85934 15202 85986
rect 15202 85934 15204 85986
rect 15148 85932 15204 85934
rect 15372 85708 15428 85764
rect 14924 85090 14980 85092
rect 14924 85038 14926 85090
rect 14926 85038 14978 85090
rect 14978 85038 14980 85090
rect 14924 85036 14980 85038
rect 15148 84924 15204 84980
rect 15036 84418 15092 84420
rect 15036 84366 15038 84418
rect 15038 84366 15090 84418
rect 15090 84366 15092 84418
rect 15036 84364 15092 84366
rect 14924 84140 14980 84196
rect 15036 83916 15092 83972
rect 14476 83410 14532 83412
rect 14476 83358 14478 83410
rect 14478 83358 14530 83410
rect 14530 83358 14532 83410
rect 14476 83356 14532 83358
rect 14812 83356 14868 83412
rect 14588 83132 14644 83188
rect 14476 82908 14532 82964
rect 14476 82460 14532 82516
rect 14028 82236 14084 82292
rect 14028 81676 14084 81732
rect 13916 81340 13972 81396
rect 13692 78092 13748 78148
rect 12796 73442 12852 73444
rect 12796 73390 12798 73442
rect 12798 73390 12850 73442
rect 12850 73390 12852 73442
rect 12796 73388 12852 73390
rect 12796 72770 12852 72772
rect 12796 72718 12798 72770
rect 12798 72718 12850 72770
rect 12850 72718 12852 72770
rect 12796 72716 12852 72718
rect 13132 74898 13188 74900
rect 13132 74846 13134 74898
rect 13134 74846 13186 74898
rect 13186 74846 13188 74898
rect 13132 74844 13188 74846
rect 13020 74620 13076 74676
rect 13244 73276 13300 73332
rect 13020 70588 13076 70644
rect 12012 68012 12068 68068
rect 12348 68012 12404 68068
rect 12124 67954 12180 67956
rect 12124 67902 12126 67954
rect 12126 67902 12178 67954
rect 12178 67902 12180 67954
rect 12124 67900 12180 67902
rect 11788 63868 11844 63924
rect 11900 63362 11956 63364
rect 11900 63310 11902 63362
rect 11902 63310 11954 63362
rect 11954 63310 11956 63362
rect 11900 63308 11956 63310
rect 11676 62412 11732 62468
rect 11900 62860 11956 62916
rect 12348 61628 12404 61684
rect 12348 61180 12404 61236
rect 12460 60844 12516 60900
rect 11564 58604 11620 58660
rect 12236 56812 12292 56868
rect 11452 56364 11508 56420
rect 11676 56028 11732 56084
rect 11340 49308 11396 49364
rect 11452 51772 11508 51828
rect 11452 50652 11508 50708
rect 11228 48188 11284 48244
rect 11340 48524 11396 48580
rect 11564 51212 11620 51268
rect 12348 56028 12404 56084
rect 12236 52892 12292 52948
rect 11788 52332 11844 52388
rect 12236 52556 12292 52612
rect 11900 51324 11956 51380
rect 11788 50482 11844 50484
rect 11788 50430 11790 50482
rect 11790 50430 11842 50482
rect 11842 50430 11844 50482
rect 11788 50428 11844 50430
rect 12012 50428 12068 50484
rect 11676 48412 11732 48468
rect 11788 49420 11844 49476
rect 11228 47068 11284 47124
rect 11116 46620 11172 46676
rect 11452 48130 11508 48132
rect 11452 48078 11454 48130
rect 11454 48078 11506 48130
rect 11506 48078 11508 48130
rect 11452 48076 11508 48078
rect 11676 48130 11732 48132
rect 11676 48078 11678 48130
rect 11678 48078 11730 48130
rect 11730 48078 11732 48130
rect 11676 48076 11732 48078
rect 11228 45836 11284 45892
rect 11228 45388 11284 45444
rect 10892 44546 10948 44548
rect 10892 44494 10894 44546
rect 10894 44494 10946 44546
rect 10946 44494 10948 44546
rect 10892 44492 10948 44494
rect 10220 43820 10276 43876
rect 10332 43932 10388 43988
rect 11004 43932 11060 43988
rect 10892 43036 10948 43092
rect 9996 41074 10052 41076
rect 9996 41022 9998 41074
rect 9998 41022 10050 41074
rect 10050 41022 10052 41074
rect 9996 41020 10052 41022
rect 9884 39058 9940 39060
rect 9884 39006 9886 39058
rect 9886 39006 9938 39058
rect 9938 39006 9940 39058
rect 9884 39004 9940 39006
rect 9884 38274 9940 38276
rect 9884 38222 9886 38274
rect 9886 38222 9938 38274
rect 9938 38222 9940 38274
rect 9884 38220 9940 38222
rect 10556 41916 10612 41972
rect 10332 40572 10388 40628
rect 10220 40460 10276 40516
rect 11004 41410 11060 41412
rect 11004 41358 11006 41410
rect 11006 41358 11058 41410
rect 11058 41358 11060 41410
rect 11004 41356 11060 41358
rect 10668 40796 10724 40852
rect 10780 41186 10836 41188
rect 10780 41134 10782 41186
rect 10782 41134 10834 41186
rect 10834 41134 10836 41186
rect 10780 41132 10836 41134
rect 10108 40348 10164 40404
rect 10108 40124 10164 40180
rect 10220 39900 10276 39956
rect 10108 39116 10164 39172
rect 10220 38108 10276 38164
rect 9996 37100 10052 37156
rect 10444 39452 10500 39508
rect 9772 36540 9828 36596
rect 9324 30044 9380 30100
rect 9436 35420 9492 35476
rect 8652 28588 8708 28644
rect 8988 28700 9044 28756
rect 8316 27692 8372 27748
rect 8316 26290 8372 26292
rect 8316 26238 8318 26290
rect 8318 26238 8370 26290
rect 8370 26238 8372 26290
rect 8316 26236 8372 26238
rect 7756 23324 7812 23380
rect 8316 25116 8372 25172
rect 7532 20524 7588 20580
rect 8876 26796 8932 26852
rect 9100 28252 9156 28308
rect 9212 27580 9268 27636
rect 9100 27244 9156 27300
rect 9212 27074 9268 27076
rect 9212 27022 9214 27074
rect 9214 27022 9266 27074
rect 9266 27022 9268 27074
rect 9212 27020 9268 27022
rect 9100 26290 9156 26292
rect 9100 26238 9102 26290
rect 9102 26238 9154 26290
rect 9154 26238 9156 26290
rect 9100 26236 9156 26238
rect 8988 25564 9044 25620
rect 9100 25506 9156 25508
rect 9100 25454 9102 25506
rect 9102 25454 9154 25506
rect 9154 25454 9156 25506
rect 9100 25452 9156 25454
rect 8652 25116 8708 25172
rect 9324 24668 9380 24724
rect 8988 24610 9044 24612
rect 8988 24558 8990 24610
rect 8990 24558 9042 24610
rect 9042 24558 9044 24610
rect 8988 24556 9044 24558
rect 6860 19404 6916 19460
rect 6636 19122 6692 19124
rect 6636 19070 6638 19122
rect 6638 19070 6690 19122
rect 6690 19070 6692 19122
rect 6636 19068 6692 19070
rect 6636 17948 6692 18004
rect 7084 18508 7140 18564
rect 6748 17724 6804 17780
rect 6524 16268 6580 16324
rect 6636 17276 6692 17332
rect 6636 17052 6692 17108
rect 6412 11564 6468 11620
rect 6860 17612 6916 17668
rect 6972 17106 7028 17108
rect 6972 17054 6974 17106
rect 6974 17054 7026 17106
rect 7026 17054 7028 17106
rect 6972 17052 7028 17054
rect 7084 16322 7140 16324
rect 7084 16270 7086 16322
rect 7086 16270 7138 16322
rect 7138 16270 7140 16322
rect 7084 16268 7140 16270
rect 6300 11228 6356 11284
rect 6748 15036 6804 15092
rect 7532 19516 7588 19572
rect 7756 22092 7812 22148
rect 7868 21474 7924 21476
rect 7868 21422 7870 21474
rect 7870 21422 7922 21474
rect 7922 21422 7924 21474
rect 7868 21420 7924 21422
rect 7756 19404 7812 19460
rect 7868 21196 7924 21252
rect 7980 19516 8036 19572
rect 8092 20188 8148 20244
rect 7868 18284 7924 18340
rect 7868 17612 7924 17668
rect 7980 16716 8036 16772
rect 8204 19964 8260 20020
rect 8204 19458 8260 19460
rect 8204 19406 8206 19458
rect 8206 19406 8258 19458
rect 8258 19406 8260 19458
rect 8204 19404 8260 19406
rect 8540 20076 8596 20132
rect 8764 20076 8820 20132
rect 8652 19906 8708 19908
rect 8652 19854 8654 19906
rect 8654 19854 8706 19906
rect 8706 19854 8708 19906
rect 8652 19852 8708 19854
rect 8988 23212 9044 23268
rect 9324 22204 9380 22260
rect 9212 21084 9268 21140
rect 8988 19404 9044 19460
rect 8876 18844 8932 18900
rect 8988 18450 9044 18452
rect 8988 18398 8990 18450
rect 8990 18398 9042 18450
rect 9042 18398 9044 18450
rect 8988 18396 9044 18398
rect 9100 17666 9156 17668
rect 9100 17614 9102 17666
rect 9102 17614 9154 17666
rect 9154 17614 9156 17666
rect 9100 17612 9156 17614
rect 9660 35308 9716 35364
rect 9548 34860 9604 34916
rect 9772 34636 9828 34692
rect 9996 36652 10052 36708
rect 10556 39116 10612 39172
rect 10668 40460 10724 40516
rect 10556 37660 10612 37716
rect 10780 40348 10836 40404
rect 10892 41020 10948 41076
rect 11340 45052 11396 45108
rect 11452 43708 11508 43764
rect 11452 42754 11508 42756
rect 11452 42702 11454 42754
rect 11454 42702 11506 42754
rect 11506 42702 11508 42754
rect 11452 42700 11508 42702
rect 11340 42588 11396 42644
rect 11340 40572 11396 40628
rect 11228 40460 11284 40516
rect 10780 38892 10836 38948
rect 11900 48242 11956 48244
rect 11900 48190 11902 48242
rect 11902 48190 11954 48242
rect 11954 48190 11956 48242
rect 11900 48188 11956 48190
rect 12236 48524 12292 48580
rect 12348 48860 12404 48916
rect 12236 48188 12292 48244
rect 12012 46508 12068 46564
rect 12236 47458 12292 47460
rect 12236 47406 12238 47458
rect 12238 47406 12290 47458
rect 12290 47406 12292 47458
rect 12236 47404 12292 47406
rect 12572 50594 12628 50596
rect 12572 50542 12574 50594
rect 12574 50542 12626 50594
rect 12626 50542 12628 50594
rect 12572 50540 12628 50542
rect 12796 68572 12852 68628
rect 12908 68402 12964 68404
rect 12908 68350 12910 68402
rect 12910 68350 12962 68402
rect 12962 68350 12964 68402
rect 12908 68348 12964 68350
rect 12796 67900 12852 67956
rect 12908 67676 12964 67732
rect 13132 69356 13188 69412
rect 13580 75964 13636 76020
rect 13468 74060 13524 74116
rect 14028 75964 14084 76020
rect 14476 82124 14532 82180
rect 14252 81954 14308 81956
rect 14252 81902 14254 81954
rect 14254 81902 14306 81954
rect 14306 81902 14308 81954
rect 14252 81900 14308 81902
rect 14476 81676 14532 81732
rect 14924 82684 14980 82740
rect 15036 82236 15092 82292
rect 14924 81788 14980 81844
rect 14812 81676 14868 81732
rect 14588 81452 14644 81508
rect 14700 81340 14756 81396
rect 14588 81170 14644 81172
rect 14588 81118 14590 81170
rect 14590 81118 14642 81170
rect 14642 81118 14644 81170
rect 14588 81116 14644 81118
rect 17388 112306 17444 112308
rect 17388 112254 17390 112306
rect 17390 112254 17442 112306
rect 17442 112254 17444 112306
rect 17388 112252 17444 112254
rect 17052 110796 17108 110852
rect 17612 112140 17668 112196
rect 16828 108556 16884 108612
rect 16828 107826 16884 107828
rect 16828 107774 16830 107826
rect 16830 107774 16882 107826
rect 16882 107774 16884 107826
rect 16828 107772 16884 107774
rect 16828 107042 16884 107044
rect 16828 106990 16830 107042
rect 16830 106990 16882 107042
rect 16882 106990 16884 107042
rect 16828 106988 16884 106990
rect 16716 106258 16772 106260
rect 16716 106206 16718 106258
rect 16718 106206 16770 106258
rect 16770 106206 16772 106258
rect 16716 106204 16772 106206
rect 16604 105196 16660 105252
rect 16604 103068 16660 103124
rect 16716 104412 16772 104468
rect 16604 102898 16660 102900
rect 16604 102846 16606 102898
rect 16606 102846 16658 102898
rect 16658 102846 16660 102898
rect 16604 102844 16660 102846
rect 16828 104076 16884 104132
rect 17612 110012 17668 110068
rect 17500 109452 17556 109508
rect 17388 109116 17444 109172
rect 17164 105196 17220 105252
rect 17276 108892 17332 108948
rect 17276 103180 17332 103236
rect 17388 108556 17444 108612
rect 17052 103122 17108 103124
rect 17052 103070 17054 103122
rect 17054 103070 17106 103122
rect 17106 103070 17108 103122
rect 17052 103068 17108 103070
rect 16940 100604 16996 100660
rect 17276 102060 17332 102116
rect 17500 107100 17556 107156
rect 17948 111858 18004 111860
rect 17948 111806 17950 111858
rect 17950 111806 18002 111858
rect 18002 111806 18004 111858
rect 17948 111804 18004 111806
rect 17948 110962 18004 110964
rect 17948 110910 17950 110962
rect 17950 110910 18002 110962
rect 18002 110910 18004 110962
rect 17948 110908 18004 110910
rect 17836 110012 17892 110068
rect 17724 109340 17780 109396
rect 17948 108892 18004 108948
rect 17724 108332 17780 108388
rect 17612 106428 17668 106484
rect 17948 106652 18004 106708
rect 17836 103516 17892 103572
rect 17948 105644 18004 105700
rect 17724 102844 17780 102900
rect 17388 101948 17444 102004
rect 17276 100770 17332 100772
rect 17276 100718 17278 100770
rect 17278 100718 17330 100770
rect 17330 100718 17332 100770
rect 17276 100716 17332 100718
rect 17276 100492 17332 100548
rect 16716 97020 16772 97076
rect 16828 97468 16884 97524
rect 16492 96348 16548 96404
rect 16492 96124 16548 96180
rect 15932 93324 15988 93380
rect 15932 91980 15988 92036
rect 16044 92092 16100 92148
rect 15932 91196 15988 91252
rect 15708 90972 15764 91028
rect 15708 85932 15764 85988
rect 15820 90636 15876 90692
rect 15596 84700 15652 84756
rect 15148 81228 15204 81284
rect 14364 79602 14420 79604
rect 14364 79550 14366 79602
rect 14366 79550 14418 79602
rect 14418 79550 14420 79602
rect 14364 79548 14420 79550
rect 14252 78876 14308 78932
rect 14812 80668 14868 80724
rect 15036 80668 15092 80724
rect 14700 80220 14756 80276
rect 15148 80556 15204 80612
rect 14924 80108 14980 80164
rect 15484 81676 15540 81732
rect 15484 81228 15540 81284
rect 15484 80892 15540 80948
rect 16268 92652 16324 92708
rect 16380 93772 16436 93828
rect 16156 91308 16212 91364
rect 16268 92316 16324 92372
rect 16044 90188 16100 90244
rect 16044 85932 16100 85988
rect 16044 85484 16100 85540
rect 16044 85090 16100 85092
rect 16044 85038 16046 85090
rect 16046 85038 16098 85090
rect 16098 85038 16100 85090
rect 16044 85036 16100 85038
rect 16828 95788 16884 95844
rect 17164 97580 17220 97636
rect 17052 96178 17108 96180
rect 17052 96126 17054 96178
rect 17054 96126 17106 96178
rect 17106 96126 17108 96178
rect 17052 96124 17108 96126
rect 17164 94108 17220 94164
rect 16604 92428 16660 92484
rect 16492 92316 16548 92372
rect 16492 90188 16548 90244
rect 17052 93714 17108 93716
rect 17052 93662 17054 93714
rect 17054 93662 17106 93714
rect 17106 93662 17108 93714
rect 17052 93660 17108 93662
rect 17052 92930 17108 92932
rect 17052 92878 17054 92930
rect 17054 92878 17106 92930
rect 17106 92878 17108 92930
rect 17052 92876 17108 92878
rect 17052 92146 17108 92148
rect 17052 92094 17054 92146
rect 17054 92094 17106 92146
rect 17106 92094 17108 92146
rect 17052 92092 17108 92094
rect 17164 91980 17220 92036
rect 16716 90972 16772 91028
rect 16828 91084 16884 91140
rect 16716 90354 16772 90356
rect 16716 90302 16718 90354
rect 16718 90302 16770 90354
rect 16770 90302 16772 90354
rect 16716 90300 16772 90302
rect 16604 88844 16660 88900
rect 16716 87500 16772 87556
rect 16380 85820 16436 85876
rect 16492 87388 16548 87444
rect 16156 84924 16212 84980
rect 15932 84306 15988 84308
rect 15932 84254 15934 84306
rect 15934 84254 15986 84306
rect 15986 84254 15988 84306
rect 15932 84252 15988 84254
rect 16044 84194 16100 84196
rect 16044 84142 16046 84194
rect 16046 84142 16098 84194
rect 16098 84142 16100 84194
rect 16044 84140 16100 84142
rect 16156 84028 16212 84084
rect 16044 83522 16100 83524
rect 16044 83470 16046 83522
rect 16046 83470 16098 83522
rect 16098 83470 16100 83522
rect 16044 83468 16100 83470
rect 16044 82908 16100 82964
rect 15932 82460 15988 82516
rect 15708 82066 15764 82068
rect 15708 82014 15710 82066
rect 15710 82014 15762 82066
rect 15762 82014 15764 82066
rect 15708 82012 15764 82014
rect 15708 81282 15764 81284
rect 15708 81230 15710 81282
rect 15710 81230 15762 81282
rect 15762 81230 15764 81282
rect 15708 81228 15764 81230
rect 15148 79548 15204 79604
rect 15596 79602 15652 79604
rect 15596 79550 15598 79602
rect 15598 79550 15650 79602
rect 15650 79550 15652 79602
rect 15596 79548 15652 79550
rect 14924 79100 14980 79156
rect 14588 78316 14644 78372
rect 14812 78316 14868 78372
rect 15148 78652 15204 78708
rect 15484 78034 15540 78036
rect 15484 77982 15486 78034
rect 15486 77982 15538 78034
rect 15538 77982 15540 78034
rect 15484 77980 15540 77982
rect 13804 74786 13860 74788
rect 13804 74734 13806 74786
rect 13806 74734 13858 74786
rect 13858 74734 13860 74786
rect 13804 74732 13860 74734
rect 13692 74172 13748 74228
rect 13692 73330 13748 73332
rect 13692 73278 13694 73330
rect 13694 73278 13746 73330
rect 13746 73278 13748 73330
rect 13692 73276 13748 73278
rect 13804 73106 13860 73108
rect 13804 73054 13806 73106
rect 13806 73054 13858 73106
rect 13858 73054 13860 73106
rect 13804 73052 13860 73054
rect 13580 72828 13636 72884
rect 13804 72604 13860 72660
rect 13356 72268 13412 72324
rect 13916 72268 13972 72324
rect 14252 72716 14308 72772
rect 14252 71538 14308 71540
rect 14252 71486 14254 71538
rect 14254 71486 14306 71538
rect 14306 71486 14308 71538
rect 14252 71484 14308 71486
rect 14812 74732 14868 74788
rect 14476 74114 14532 74116
rect 14476 74062 14478 74114
rect 14478 74062 14530 74114
rect 14530 74062 14532 74114
rect 14476 74060 14532 74062
rect 14588 72940 14644 72996
rect 14476 71932 14532 71988
rect 13244 67676 13300 67732
rect 13356 68796 13412 68852
rect 13020 65602 13076 65604
rect 13020 65550 13022 65602
rect 13022 65550 13074 65602
rect 13074 65550 13076 65602
rect 13020 65548 13076 65550
rect 13580 68348 13636 68404
rect 14364 70476 14420 70532
rect 13804 66834 13860 66836
rect 13804 66782 13806 66834
rect 13806 66782 13858 66834
rect 13858 66782 13860 66834
rect 13804 66780 13860 66782
rect 13468 65660 13524 65716
rect 13580 65772 13636 65828
rect 13692 65100 13748 65156
rect 13132 63980 13188 64036
rect 13580 64316 13636 64372
rect 12908 63308 12964 63364
rect 13468 63308 13524 63364
rect 12908 62860 12964 62916
rect 13468 62748 13524 62804
rect 13020 61570 13076 61572
rect 13020 61518 13022 61570
rect 13022 61518 13074 61570
rect 13074 61518 13076 61570
rect 13020 61516 13076 61518
rect 13132 61292 13188 61348
rect 13132 60620 13188 60676
rect 15484 76860 15540 76916
rect 15036 73330 15092 73332
rect 15036 73278 15038 73330
rect 15038 73278 15090 73330
rect 15090 73278 15092 73330
rect 15036 73276 15092 73278
rect 14924 72940 14980 72996
rect 14476 69356 14532 69412
rect 14476 69020 14532 69076
rect 14588 68796 14644 68852
rect 14140 68684 14196 68740
rect 14140 67842 14196 67844
rect 14140 67790 14142 67842
rect 14142 67790 14194 67842
rect 14194 67790 14196 67842
rect 14140 67788 14196 67790
rect 14140 67340 14196 67396
rect 13916 66108 13972 66164
rect 13916 65772 13972 65828
rect 14924 72604 14980 72660
rect 14812 71090 14868 71092
rect 14812 71038 14814 71090
rect 14814 71038 14866 71090
rect 14866 71038 14868 71090
rect 14812 71036 14868 71038
rect 14252 65548 14308 65604
rect 14812 68460 14868 68516
rect 14252 64034 14308 64036
rect 14252 63982 14254 64034
rect 14254 63982 14306 64034
rect 14306 63982 14308 64034
rect 14252 63980 14308 63982
rect 14924 67564 14980 67620
rect 15260 71596 15316 71652
rect 14700 67116 14756 67172
rect 14924 67058 14980 67060
rect 14924 67006 14926 67058
rect 14926 67006 14978 67058
rect 14978 67006 14980 67058
rect 14924 67004 14980 67006
rect 15372 70476 15428 70532
rect 15260 68626 15316 68628
rect 15260 68574 15262 68626
rect 15262 68574 15314 68626
rect 15314 68574 15316 68626
rect 15260 68572 15316 68574
rect 15260 67900 15316 67956
rect 15260 67228 15316 67284
rect 15148 66834 15204 66836
rect 15148 66782 15150 66834
rect 15150 66782 15202 66834
rect 15202 66782 15204 66834
rect 15148 66780 15204 66782
rect 15036 66556 15092 66612
rect 14476 63308 14532 63364
rect 13916 63138 13972 63140
rect 13916 63086 13918 63138
rect 13918 63086 13970 63138
rect 13970 63086 13972 63138
rect 13916 63084 13972 63086
rect 14252 62466 14308 62468
rect 14252 62414 14254 62466
rect 14254 62414 14306 62466
rect 14306 62414 14308 62466
rect 14252 62412 14308 62414
rect 15820 80556 15876 80612
rect 15932 81452 15988 81508
rect 16156 81452 16212 81508
rect 16604 85762 16660 85764
rect 16604 85710 16606 85762
rect 16606 85710 16658 85762
rect 16658 85710 16660 85762
rect 16604 85708 16660 85710
rect 16604 85484 16660 85540
rect 16604 84252 16660 84308
rect 16828 85932 16884 85988
rect 16940 89740 16996 89796
rect 17388 98924 17444 98980
rect 17612 102450 17668 102452
rect 17612 102398 17614 102450
rect 17614 102398 17666 102450
rect 17666 102398 17668 102450
rect 17612 102396 17668 102398
rect 17836 100716 17892 100772
rect 17724 99874 17780 99876
rect 17724 99822 17726 99874
rect 17726 99822 17778 99874
rect 17778 99822 17780 99874
rect 17724 99820 17780 99822
rect 17612 99708 17668 99764
rect 18508 113932 18564 113988
rect 18844 113932 18900 113988
rect 18620 113708 18676 113764
rect 19180 113596 19236 113652
rect 18284 111580 18340 111636
rect 18284 111132 18340 111188
rect 18284 109788 18340 109844
rect 18172 108108 18228 108164
rect 19068 113260 19124 113316
rect 18956 112700 19012 112756
rect 19516 113484 19572 113540
rect 19628 113708 19684 113764
rect 19516 113148 19572 113204
rect 19516 112812 19572 112868
rect 19068 110850 19124 110852
rect 19068 110798 19070 110850
rect 19070 110798 19122 110850
rect 19122 110798 19124 110850
rect 19068 110796 19124 110798
rect 18396 106764 18452 106820
rect 18508 109788 18564 109844
rect 18620 109394 18676 109396
rect 18620 109342 18622 109394
rect 18622 109342 18674 109394
rect 18674 109342 18676 109394
rect 18620 109340 18676 109342
rect 18732 106652 18788 106708
rect 18620 106428 18676 106484
rect 18508 106204 18564 106260
rect 18956 110124 19012 110180
rect 18956 109340 19012 109396
rect 19292 110178 19348 110180
rect 19292 110126 19294 110178
rect 19294 110126 19346 110178
rect 19346 110126 19348 110178
rect 19292 110124 19348 110126
rect 19516 111132 19572 111188
rect 19852 114268 19908 114324
rect 19852 112812 19908 112868
rect 20188 113260 20244 113316
rect 20412 113260 20468 113316
rect 20524 114380 20580 114436
rect 19740 112476 19796 112532
rect 19964 112588 20020 112644
rect 19852 111916 19908 111972
rect 18172 104466 18228 104468
rect 18172 104414 18174 104466
rect 18174 104414 18226 104466
rect 18226 104414 18228 104466
rect 18172 104412 18228 104414
rect 19180 108892 19236 108948
rect 19068 105586 19124 105588
rect 19068 105534 19070 105586
rect 19070 105534 19122 105586
rect 19122 105534 19124 105586
rect 19068 105532 19124 105534
rect 19068 105196 19124 105252
rect 18956 104018 19012 104020
rect 18956 103966 18958 104018
rect 18958 103966 19010 104018
rect 19010 103966 19012 104018
rect 18956 103964 19012 103966
rect 18844 101724 18900 101780
rect 18508 101052 18564 101108
rect 19404 109116 19460 109172
rect 19404 105586 19460 105588
rect 19404 105534 19406 105586
rect 19406 105534 19458 105586
rect 19458 105534 19460 105586
rect 19404 105532 19460 105534
rect 19740 110572 19796 110628
rect 19628 109004 19684 109060
rect 20300 112476 20356 112532
rect 20076 110908 20132 110964
rect 19964 110402 20020 110404
rect 19964 110350 19966 110402
rect 19966 110350 20018 110402
rect 20018 110350 20020 110402
rect 19964 110348 20020 110350
rect 19964 109452 20020 109508
rect 19740 108892 19796 108948
rect 19852 106428 19908 106484
rect 19516 104412 19572 104468
rect 19628 103964 19684 104020
rect 19516 102898 19572 102900
rect 19516 102846 19518 102898
rect 19518 102846 19570 102898
rect 19570 102846 19572 102898
rect 19516 102844 19572 102846
rect 18060 100492 18116 100548
rect 18956 99426 19012 99428
rect 18956 99374 18958 99426
rect 18958 99374 19010 99426
rect 19010 99374 19012 99426
rect 18956 99372 19012 99374
rect 19292 99314 19348 99316
rect 19292 99262 19294 99314
rect 19294 99262 19346 99314
rect 19346 99262 19348 99314
rect 19292 99260 19348 99262
rect 18844 99148 18900 99204
rect 18844 98530 18900 98532
rect 18844 98478 18846 98530
rect 18846 98478 18898 98530
rect 18898 98478 18900 98530
rect 18844 98476 18900 98478
rect 18172 98418 18228 98420
rect 18172 98366 18174 98418
rect 18174 98366 18226 98418
rect 18226 98366 18228 98418
rect 18172 98364 18228 98366
rect 18620 98364 18676 98420
rect 18284 98140 18340 98196
rect 18060 97916 18116 97972
rect 17500 94444 17556 94500
rect 18284 97580 18340 97636
rect 18396 97692 18452 97748
rect 19292 98418 19348 98420
rect 19292 98366 19294 98418
rect 19294 98366 19346 98418
rect 19346 98366 19348 98418
rect 19292 98364 19348 98366
rect 19516 99148 19572 99204
rect 18732 97468 18788 97524
rect 18284 96460 18340 96516
rect 17724 96012 17780 96068
rect 17836 96124 17892 96180
rect 17724 93996 17780 94052
rect 18060 96012 18116 96068
rect 17836 93884 17892 93940
rect 17948 95676 18004 95732
rect 17836 93714 17892 93716
rect 17836 93662 17838 93714
rect 17838 93662 17890 93714
rect 17890 93662 17892 93714
rect 17836 93660 17892 93662
rect 17724 92876 17780 92932
rect 17500 92540 17556 92596
rect 17836 92316 17892 92372
rect 17948 92092 18004 92148
rect 17724 91474 17780 91476
rect 17724 91422 17726 91474
rect 17726 91422 17778 91474
rect 17778 91422 17780 91474
rect 17724 91420 17780 91422
rect 18172 94722 18228 94724
rect 18172 94670 18174 94722
rect 18174 94670 18226 94722
rect 18226 94670 18228 94722
rect 18172 94668 18228 94670
rect 18172 94444 18228 94500
rect 18396 95900 18452 95956
rect 18396 93996 18452 94052
rect 18172 91362 18228 91364
rect 18172 91310 18174 91362
rect 18174 91310 18226 91362
rect 18226 91310 18228 91362
rect 18172 91308 18228 91310
rect 17948 91196 18004 91252
rect 17724 91084 17780 91140
rect 17500 90188 17556 90244
rect 17724 90188 17780 90244
rect 17276 89292 17332 89348
rect 17164 85874 17220 85876
rect 17164 85822 17166 85874
rect 17166 85822 17218 85874
rect 17218 85822 17220 85874
rect 17164 85820 17220 85822
rect 17164 85372 17220 85428
rect 16828 84812 16884 84868
rect 16716 84028 16772 84084
rect 16940 84476 16996 84532
rect 15820 78540 15876 78596
rect 15820 78092 15876 78148
rect 16044 78764 16100 78820
rect 15932 77922 15988 77924
rect 15932 77870 15934 77922
rect 15934 77870 15986 77922
rect 15986 77870 15988 77922
rect 15932 77868 15988 77870
rect 16156 78652 16212 78708
rect 16156 75516 16212 75572
rect 16044 74844 16100 74900
rect 15932 73276 15988 73332
rect 15820 72156 15876 72212
rect 15708 71596 15764 71652
rect 15596 71538 15652 71540
rect 15596 71486 15598 71538
rect 15598 71486 15650 71538
rect 15650 71486 15652 71538
rect 15596 71484 15652 71486
rect 15708 71260 15764 71316
rect 16604 82460 16660 82516
rect 16380 78988 16436 79044
rect 17052 83522 17108 83524
rect 17052 83470 17054 83522
rect 17054 83470 17106 83522
rect 17106 83470 17108 83522
rect 17052 83468 17108 83470
rect 16940 82796 16996 82852
rect 16716 79548 16772 79604
rect 16604 79490 16660 79492
rect 16604 79438 16606 79490
rect 16606 79438 16658 79490
rect 16658 79438 16660 79490
rect 16604 79436 16660 79438
rect 16492 76860 16548 76916
rect 17052 78818 17108 78820
rect 17052 78766 17054 78818
rect 17054 78766 17106 78818
rect 17106 78766 17108 78818
rect 17052 78764 17108 78766
rect 16268 75068 16324 75124
rect 16828 77980 16884 78036
rect 16380 74396 16436 74452
rect 16268 68514 16324 68516
rect 16268 68462 16270 68514
rect 16270 68462 16322 68514
rect 16322 68462 16324 68514
rect 16268 68460 16324 68462
rect 16156 67954 16212 67956
rect 16156 67902 16158 67954
rect 16158 67902 16210 67954
rect 16210 67902 16212 67954
rect 16156 67900 16212 67902
rect 16044 67340 16100 67396
rect 16156 67676 16212 67732
rect 15932 67116 15988 67172
rect 15484 67004 15540 67060
rect 16156 65660 16212 65716
rect 16268 66668 16324 66724
rect 15820 65602 15876 65604
rect 15820 65550 15822 65602
rect 15822 65550 15874 65602
rect 15874 65550 15876 65602
rect 15820 65548 15876 65550
rect 15484 63756 15540 63812
rect 15260 63138 15316 63140
rect 15260 63086 15262 63138
rect 15262 63086 15314 63138
rect 15314 63086 15316 63138
rect 15260 63084 15316 63086
rect 15148 62412 15204 62468
rect 15036 62188 15092 62244
rect 15260 62130 15316 62132
rect 15260 62078 15262 62130
rect 15262 62078 15314 62130
rect 15314 62078 15316 62130
rect 15260 62076 15316 62078
rect 13804 61068 13860 61124
rect 13580 60172 13636 60228
rect 13692 59164 13748 59220
rect 13580 57538 13636 57540
rect 13580 57486 13582 57538
rect 13582 57486 13634 57538
rect 13634 57486 13636 57538
rect 13580 57484 13636 57486
rect 13132 56866 13188 56868
rect 13132 56814 13134 56866
rect 13134 56814 13186 56866
rect 13186 56814 13188 56866
rect 13132 56812 13188 56814
rect 13132 52220 13188 52276
rect 12796 50706 12852 50708
rect 12796 50654 12798 50706
rect 12798 50654 12850 50706
rect 12850 50654 12852 50706
rect 12796 50652 12852 50654
rect 12684 49420 12740 49476
rect 12796 50316 12852 50372
rect 12684 49250 12740 49252
rect 12684 49198 12686 49250
rect 12686 49198 12738 49250
rect 12738 49198 12740 49250
rect 12684 49196 12740 49198
rect 12460 46956 12516 47012
rect 11900 43148 11956 43204
rect 12012 42476 12068 42532
rect 11900 42364 11956 42420
rect 11900 42082 11956 42084
rect 11900 42030 11902 42082
rect 11902 42030 11954 42082
rect 11954 42030 11956 42082
rect 11900 42028 11956 42030
rect 11788 41916 11844 41972
rect 11676 39900 11732 39956
rect 11788 40236 11844 40292
rect 11676 39452 11732 39508
rect 11228 39004 11284 39060
rect 11564 38892 11620 38948
rect 10668 37042 10724 37044
rect 10668 36990 10670 37042
rect 10670 36990 10722 37042
rect 10722 36990 10724 37042
rect 10668 36988 10724 36990
rect 10444 36876 10500 36932
rect 10780 36764 10836 36820
rect 10332 36482 10388 36484
rect 10332 36430 10334 36482
rect 10334 36430 10386 36482
rect 10386 36430 10388 36482
rect 10332 36428 10388 36430
rect 10220 35420 10276 35476
rect 9884 34076 9940 34132
rect 9996 34300 10052 34356
rect 9660 33404 9716 33460
rect 9996 33740 10052 33796
rect 9548 31612 9604 31668
rect 10108 33292 10164 33348
rect 9884 32786 9940 32788
rect 9884 32734 9886 32786
rect 9886 32734 9938 32786
rect 9938 32734 9940 32786
rect 9884 32732 9940 32734
rect 9884 31948 9940 32004
rect 9772 30268 9828 30324
rect 9996 31612 10052 31668
rect 9884 28754 9940 28756
rect 9884 28702 9886 28754
rect 9886 28702 9938 28754
rect 9938 28702 9940 28754
rect 9884 28700 9940 28702
rect 9772 28252 9828 28308
rect 9772 27244 9828 27300
rect 9884 27186 9940 27188
rect 9884 27134 9886 27186
rect 9886 27134 9938 27186
rect 9938 27134 9940 27186
rect 9884 27132 9940 27134
rect 9548 26290 9604 26292
rect 9548 26238 9550 26290
rect 9550 26238 9602 26290
rect 9602 26238 9604 26290
rect 9548 26236 9604 26238
rect 9884 26236 9940 26292
rect 9772 26066 9828 26068
rect 9772 26014 9774 26066
rect 9774 26014 9826 26066
rect 9826 26014 9828 26066
rect 9772 26012 9828 26014
rect 9660 25900 9716 25956
rect 9436 20748 9492 20804
rect 9548 25116 9604 25172
rect 9548 24220 9604 24276
rect 9548 20300 9604 20356
rect 9436 20076 9492 20132
rect 9660 20076 9716 20132
rect 9660 19794 9716 19796
rect 9660 19742 9662 19794
rect 9662 19742 9714 19794
rect 9714 19742 9716 19794
rect 9660 19740 9716 19742
rect 9660 18956 9716 19012
rect 8204 16770 8260 16772
rect 8204 16718 8206 16770
rect 8206 16718 8258 16770
rect 8258 16718 8260 16770
rect 8204 16716 8260 16718
rect 7868 15260 7924 15316
rect 7756 13916 7812 13972
rect 8092 15090 8148 15092
rect 8092 15038 8094 15090
rect 8094 15038 8146 15090
rect 8146 15038 8148 15090
rect 8092 15036 8148 15038
rect 7980 14588 8036 14644
rect 7532 13692 7588 13748
rect 7868 13692 7924 13748
rect 6748 13634 6804 13636
rect 6748 13582 6750 13634
rect 6750 13582 6802 13634
rect 6802 13582 6804 13634
rect 6748 13580 6804 13582
rect 6972 13244 7028 13300
rect 6748 12962 6804 12964
rect 6748 12910 6750 12962
rect 6750 12910 6802 12962
rect 6802 12910 6804 12962
rect 6748 12908 6804 12910
rect 6748 11954 6804 11956
rect 6748 11902 6750 11954
rect 6750 11902 6802 11954
rect 6802 11902 6804 11954
rect 6748 11900 6804 11902
rect 6636 11564 6692 11620
rect 6524 11340 6580 11396
rect 6076 9100 6132 9156
rect 6188 9996 6244 10052
rect 5964 9042 6020 9044
rect 5964 8990 5966 9042
rect 5966 8990 6018 9042
rect 6018 8990 6020 9042
rect 5964 8988 6020 8990
rect 5964 8204 6020 8260
rect 6076 7532 6132 7588
rect 4464 5514 4520 5516
rect 4464 5462 4466 5514
rect 4466 5462 4518 5514
rect 4518 5462 4520 5514
rect 4464 5460 4520 5462
rect 4568 5514 4624 5516
rect 4568 5462 4570 5514
rect 4570 5462 4622 5514
rect 4622 5462 4624 5514
rect 4568 5460 4624 5462
rect 4672 5514 4728 5516
rect 4672 5462 4674 5514
rect 4674 5462 4726 5514
rect 4726 5462 4728 5514
rect 4672 5460 4728 5462
rect 4956 6188 5012 6244
rect 5068 5906 5124 5908
rect 5068 5854 5070 5906
rect 5070 5854 5122 5906
rect 5122 5854 5124 5906
rect 5068 5852 5124 5854
rect 4844 5068 4900 5124
rect 5964 6972 6020 7028
rect 5852 6860 5908 6916
rect 5740 6748 5796 6804
rect 5292 5292 5348 5348
rect 6076 5852 6132 5908
rect 5852 5180 5908 5236
rect 6076 5628 6132 5684
rect 5404 4226 5460 4228
rect 5404 4174 5406 4226
rect 5406 4174 5458 4226
rect 5458 4174 5460 4226
rect 5404 4172 5460 4174
rect 4464 3946 4520 3948
rect 4464 3894 4466 3946
rect 4466 3894 4518 3946
rect 4518 3894 4520 3946
rect 4464 3892 4520 3894
rect 4568 3946 4624 3948
rect 4568 3894 4570 3946
rect 4570 3894 4622 3946
rect 4622 3894 4624 3946
rect 4568 3892 4624 3894
rect 4672 3946 4728 3948
rect 4672 3894 4674 3946
rect 4674 3894 4726 3946
rect 4726 3894 4728 3946
rect 4672 3892 4728 3894
rect 4956 3948 5012 4004
rect 5404 3778 5460 3780
rect 5404 3726 5406 3778
rect 5406 3726 5458 3778
rect 5458 3726 5460 3778
rect 5404 3724 5460 3726
rect 5740 4114 5796 4116
rect 5740 4062 5742 4114
rect 5742 4062 5794 4114
rect 5794 4062 5796 4114
rect 5740 4060 5796 4062
rect 6076 3836 6132 3892
rect 6636 10108 6692 10164
rect 7196 12908 7252 12964
rect 8092 12962 8148 12964
rect 8092 12910 8094 12962
rect 8094 12910 8146 12962
rect 8146 12910 8148 12962
rect 8092 12908 8148 12910
rect 7308 11618 7364 11620
rect 7308 11566 7310 11618
rect 7310 11566 7362 11618
rect 7362 11566 7364 11618
rect 7308 11564 7364 11566
rect 7756 11506 7812 11508
rect 7756 11454 7758 11506
rect 7758 11454 7810 11506
rect 7810 11454 7812 11506
rect 7756 11452 7812 11454
rect 7308 10780 7364 10836
rect 7084 10668 7140 10724
rect 6412 7644 6468 7700
rect 6300 3724 6356 3780
rect 6412 5516 6468 5572
rect 6636 8092 6692 8148
rect 6748 7644 6804 7700
rect 6636 7420 6692 7476
rect 6524 4172 6580 4228
rect 6636 6524 6692 6580
rect 6076 3276 6132 3332
rect 3804 3162 3860 3164
rect 3804 3110 3806 3162
rect 3806 3110 3858 3162
rect 3858 3110 3860 3162
rect 3804 3108 3860 3110
rect 3908 3162 3964 3164
rect 3908 3110 3910 3162
rect 3910 3110 3962 3162
rect 3962 3110 3964 3162
rect 3908 3108 3964 3110
rect 4012 3162 4068 3164
rect 4012 3110 4014 3162
rect 4014 3110 4066 3162
rect 4066 3110 4068 3162
rect 4012 3108 4068 3110
rect 4172 3052 4228 3108
rect 3836 2770 3892 2772
rect 3836 2718 3838 2770
rect 3838 2718 3890 2770
rect 3890 2718 3892 2770
rect 3836 2716 3892 2718
rect 5740 2658 5796 2660
rect 5740 2606 5742 2658
rect 5742 2606 5794 2658
rect 5794 2606 5796 2658
rect 5740 2604 5796 2606
rect 4464 2378 4520 2380
rect 4464 2326 4466 2378
rect 4466 2326 4518 2378
rect 4518 2326 4520 2378
rect 4464 2324 4520 2326
rect 4568 2378 4624 2380
rect 4568 2326 4570 2378
rect 4570 2326 4622 2378
rect 4622 2326 4624 2378
rect 4568 2324 4624 2326
rect 4672 2378 4728 2380
rect 4672 2326 4674 2378
rect 4674 2326 4726 2378
rect 4726 2326 4728 2378
rect 5292 2380 5348 2436
rect 5628 2380 5684 2436
rect 4672 2324 4728 2326
rect 4956 2210 5012 2212
rect 4956 2158 4958 2210
rect 4958 2158 5010 2210
rect 5010 2158 5012 2210
rect 4956 2156 5012 2158
rect 6748 5234 6804 5236
rect 6748 5182 6750 5234
rect 6750 5182 6802 5234
rect 6802 5182 6804 5234
rect 6748 5180 6804 5182
rect 6972 6972 7028 7028
rect 7644 10556 7700 10612
rect 7980 10386 8036 10388
rect 7980 10334 7982 10386
rect 7982 10334 8034 10386
rect 8034 10334 8036 10386
rect 7980 10332 8036 10334
rect 7532 10220 7588 10276
rect 7420 8818 7476 8820
rect 7420 8766 7422 8818
rect 7422 8766 7474 8818
rect 7474 8766 7476 8818
rect 7420 8764 7476 8766
rect 7308 8370 7364 8372
rect 7308 8318 7310 8370
rect 7310 8318 7362 8370
rect 7362 8318 7364 8370
rect 7308 8316 7364 8318
rect 7420 7420 7476 7476
rect 6972 6748 7028 6804
rect 6972 5906 7028 5908
rect 6972 5854 6974 5906
rect 6974 5854 7026 5906
rect 7026 5854 7028 5906
rect 6972 5852 7028 5854
rect 7084 5346 7140 5348
rect 7084 5294 7086 5346
rect 7086 5294 7138 5346
rect 7138 5294 7140 5346
rect 7084 5292 7140 5294
rect 6972 4060 7028 4116
rect 7308 6802 7364 6804
rect 7308 6750 7310 6802
rect 7310 6750 7362 6802
rect 7362 6750 7364 6802
rect 7308 6748 7364 6750
rect 7308 5180 7364 5236
rect 7196 3276 7252 3332
rect 5628 2044 5684 2100
rect 3836 1820 3892 1876
rect 6412 2380 6468 2436
rect 3804 1594 3860 1596
rect 3804 1542 3806 1594
rect 3806 1542 3858 1594
rect 3858 1542 3860 1594
rect 3804 1540 3860 1542
rect 3908 1594 3964 1596
rect 3908 1542 3910 1594
rect 3910 1542 3962 1594
rect 3962 1542 3964 1594
rect 3908 1540 3964 1542
rect 4012 1594 4068 1596
rect 4012 1542 4014 1594
rect 4014 1542 4066 1594
rect 4066 1542 4068 1594
rect 4012 1540 4068 1542
rect 5628 1260 5684 1316
rect 4172 1148 4228 1204
rect 4844 1090 4900 1092
rect 4844 1038 4846 1090
rect 4846 1038 4898 1090
rect 4898 1038 4900 1090
rect 4844 1036 4900 1038
rect 4464 810 4520 812
rect 4464 758 4466 810
rect 4466 758 4518 810
rect 4518 758 4520 810
rect 4464 756 4520 758
rect 4568 810 4624 812
rect 4568 758 4570 810
rect 4570 758 4622 810
rect 4622 758 4624 810
rect 4568 756 4624 758
rect 4672 810 4728 812
rect 4672 758 4674 810
rect 4674 758 4726 810
rect 4726 758 4728 810
rect 4672 756 4728 758
rect 5180 700 5236 756
rect 5628 924 5684 980
rect 1596 252 1652 308
rect 5404 364 5460 420
rect 5852 812 5908 868
rect 6076 1596 6132 1652
rect 6300 1484 6356 1540
rect 6524 1596 6580 1652
rect 6748 1596 6804 1652
rect 7868 8930 7924 8932
rect 7868 8878 7870 8930
rect 7870 8878 7922 8930
rect 7922 8878 7924 8930
rect 7868 8876 7924 8878
rect 8988 16098 9044 16100
rect 8988 16046 8990 16098
rect 8990 16046 9042 16098
rect 9042 16046 9044 16098
rect 8988 16044 9044 16046
rect 9212 17052 9268 17108
rect 8764 15314 8820 15316
rect 8764 15262 8766 15314
rect 8766 15262 8818 15314
rect 8818 15262 8820 15314
rect 8764 15260 8820 15262
rect 8316 15148 8372 15204
rect 8428 14812 8484 14868
rect 9324 15708 9380 15764
rect 9436 15202 9492 15204
rect 9436 15150 9438 15202
rect 9438 15150 9490 15202
rect 9490 15150 9492 15202
rect 9436 15148 9492 15150
rect 8988 14700 9044 14756
rect 8652 13746 8708 13748
rect 8652 13694 8654 13746
rect 8654 13694 8706 13746
rect 8706 13694 8708 13746
rect 8652 13692 8708 13694
rect 8540 13580 8596 13636
rect 8428 12796 8484 12852
rect 8428 12178 8484 12180
rect 8428 12126 8430 12178
rect 8430 12126 8482 12178
rect 8482 12126 8484 12178
rect 8428 12124 8484 12126
rect 8204 11004 8260 11060
rect 8428 10556 8484 10612
rect 8316 9772 8372 9828
rect 8204 9602 8260 9604
rect 8204 9550 8206 9602
rect 8206 9550 8258 9602
rect 8258 9550 8260 9602
rect 8204 9548 8260 9550
rect 7644 8370 7700 8372
rect 7644 8318 7646 8370
rect 7646 8318 7698 8370
rect 7698 8318 7700 8370
rect 7644 8316 7700 8318
rect 7644 7425 7646 7476
rect 7646 7425 7698 7476
rect 7698 7425 7700 7476
rect 7644 7420 7700 7425
rect 7644 5740 7700 5796
rect 8092 8428 8148 8484
rect 7980 7980 8036 8036
rect 7980 6690 8036 6692
rect 7980 6638 7982 6690
rect 7982 6638 8034 6690
rect 8034 6638 8036 6690
rect 7980 6636 8036 6638
rect 8204 8258 8260 8260
rect 8204 8206 8206 8258
rect 8206 8206 8258 8258
rect 8258 8206 8260 8258
rect 8204 8204 8260 8206
rect 7868 6412 7924 6468
rect 7868 5906 7924 5908
rect 7868 5854 7870 5906
rect 7870 5854 7922 5906
rect 7922 5854 7924 5906
rect 7868 5852 7924 5854
rect 8092 5292 8148 5348
rect 7868 5068 7924 5124
rect 8876 13468 8932 13524
rect 8876 13186 8932 13188
rect 8876 13134 8878 13186
rect 8878 13134 8930 13186
rect 8930 13134 8932 13186
rect 8876 13132 8932 13134
rect 9100 14140 9156 14196
rect 9324 15036 9380 15092
rect 9660 15148 9716 15204
rect 8764 11900 8820 11956
rect 8988 11954 9044 11956
rect 8988 11902 8990 11954
rect 8990 11902 9042 11954
rect 9042 11902 9044 11954
rect 8988 11900 9044 11902
rect 9212 12124 9268 12180
rect 9548 14028 9604 14084
rect 9436 12908 9492 12964
rect 9436 11788 9492 11844
rect 8764 11228 8820 11284
rect 8764 10668 8820 10724
rect 8428 8316 8484 8372
rect 8652 8652 8708 8708
rect 8876 9938 8932 9940
rect 8876 9886 8878 9938
rect 8878 9886 8930 9938
rect 8930 9886 8932 9938
rect 8876 9884 8932 9886
rect 9100 9996 9156 10052
rect 8764 8540 8820 8596
rect 8652 7980 8708 8036
rect 8428 6748 8484 6804
rect 8316 6636 8372 6692
rect 8316 5852 8372 5908
rect 8316 4956 8372 5012
rect 8316 3388 8372 3444
rect 7756 2770 7812 2772
rect 7756 2718 7758 2770
rect 7758 2718 7810 2770
rect 7810 2718 7812 2770
rect 7756 2716 7812 2718
rect 7532 2492 7588 2548
rect 7644 2098 7700 2100
rect 7644 2046 7646 2098
rect 7646 2046 7698 2098
rect 7698 2046 7700 2098
rect 7644 2044 7700 2046
rect 7980 2828 8036 2884
rect 8092 2716 8148 2772
rect 6972 1596 7028 1652
rect 7420 1596 7476 1652
rect 7196 252 7252 308
rect 7644 1596 7700 1652
rect 7868 1596 7924 1652
rect 8316 2268 8372 2324
rect 8428 2156 8484 2212
rect 9884 25564 9940 25620
rect 10668 35868 10724 35924
rect 10332 32732 10388 32788
rect 11004 36876 11060 36932
rect 11116 36316 11172 36372
rect 11676 37938 11732 37940
rect 11676 37886 11678 37938
rect 11678 37886 11730 37938
rect 11730 37886 11732 37938
rect 11676 37884 11732 37886
rect 11564 36764 11620 36820
rect 11340 36594 11396 36596
rect 11340 36542 11342 36594
rect 11342 36542 11394 36594
rect 11394 36542 11396 36594
rect 11340 36540 11396 36542
rect 11228 35868 11284 35924
rect 11564 36204 11620 36260
rect 11116 35084 11172 35140
rect 10780 34300 10836 34356
rect 10780 34130 10836 34132
rect 10780 34078 10782 34130
rect 10782 34078 10834 34130
rect 10834 34078 10836 34130
rect 10780 34076 10836 34078
rect 11116 34524 11172 34580
rect 11340 35308 11396 35364
rect 11564 35308 11620 35364
rect 11788 35308 11844 35364
rect 11228 33628 11284 33684
rect 10780 32732 10836 32788
rect 10780 32284 10836 32340
rect 11004 32620 11060 32676
rect 11004 32284 11060 32340
rect 11116 32508 11172 32564
rect 10444 30994 10500 30996
rect 10444 30942 10446 30994
rect 10446 30942 10498 30994
rect 10498 30942 10500 30994
rect 10444 30940 10500 30942
rect 10108 28700 10164 28756
rect 10220 28588 10276 28644
rect 10444 30268 10500 30324
rect 10668 30716 10724 30772
rect 10556 29426 10612 29428
rect 10556 29374 10558 29426
rect 10558 29374 10610 29426
rect 10610 29374 10612 29426
rect 10556 29372 10612 29374
rect 10332 28028 10388 28084
rect 10332 27580 10388 27636
rect 10556 27858 10612 27860
rect 10556 27806 10558 27858
rect 10558 27806 10610 27858
rect 10610 27806 10612 27858
rect 10556 27804 10612 27806
rect 10444 27020 10500 27076
rect 11004 31948 11060 32004
rect 11004 30716 11060 30772
rect 10780 30380 10836 30436
rect 11004 29314 11060 29316
rect 11004 29262 11006 29314
rect 11006 29262 11058 29314
rect 11058 29262 11060 29314
rect 11004 29260 11060 29262
rect 11452 32732 11508 32788
rect 11228 31612 11284 31668
rect 11340 32284 11396 32340
rect 11340 29986 11396 29988
rect 11340 29934 11342 29986
rect 11342 29934 11394 29986
rect 11394 29934 11396 29986
rect 11340 29932 11396 29934
rect 11340 29484 11396 29540
rect 12348 45612 12404 45668
rect 12348 42924 12404 42980
rect 12348 42140 12404 42196
rect 12572 48524 12628 48580
rect 12684 47404 12740 47460
rect 14252 60620 14308 60676
rect 14028 58546 14084 58548
rect 14028 58494 14030 58546
rect 14030 58494 14082 58546
rect 14082 58494 14084 58546
rect 14028 58492 14084 58494
rect 13916 58380 13972 58436
rect 15036 61404 15092 61460
rect 14812 61010 14868 61012
rect 14812 60958 14814 61010
rect 14814 60958 14866 61010
rect 14866 60958 14868 61010
rect 14812 60956 14868 60958
rect 14812 60732 14868 60788
rect 14812 59724 14868 59780
rect 14700 59218 14756 59220
rect 14700 59166 14702 59218
rect 14702 59166 14754 59218
rect 14754 59166 14756 59218
rect 14700 59164 14756 59166
rect 14588 58828 14644 58884
rect 14028 58156 14084 58212
rect 14252 57426 14308 57428
rect 14252 57374 14254 57426
rect 14254 57374 14306 57426
rect 14306 57374 14308 57426
rect 14252 57372 14308 57374
rect 13692 52780 13748 52836
rect 14140 56588 14196 56644
rect 14140 54684 14196 54740
rect 14140 54348 14196 54404
rect 14028 53618 14084 53620
rect 14028 53566 14030 53618
rect 14030 53566 14082 53618
rect 14082 53566 14084 53618
rect 14028 53564 14084 53566
rect 14028 52556 14084 52612
rect 13244 50988 13300 51044
rect 13580 50652 13636 50708
rect 14476 56194 14532 56196
rect 14476 56142 14478 56194
rect 14478 56142 14530 56194
rect 14530 56142 14532 56194
rect 14476 56140 14532 56142
rect 14588 55020 14644 55076
rect 14476 52780 14532 52836
rect 14476 52556 14532 52612
rect 14588 51996 14644 52052
rect 14588 50876 14644 50932
rect 13692 50540 13748 50596
rect 13804 50764 13860 50820
rect 12908 48860 12964 48916
rect 12908 48636 12964 48692
rect 13020 48130 13076 48132
rect 13020 48078 13022 48130
rect 13022 48078 13074 48130
rect 13074 48078 13076 48130
rect 13020 48076 13076 48078
rect 13580 48242 13636 48244
rect 13580 48190 13582 48242
rect 13582 48190 13634 48242
rect 13634 48190 13636 48242
rect 13580 48188 13636 48190
rect 13356 46956 13412 47012
rect 14028 46284 14084 46340
rect 13468 45218 13524 45220
rect 13468 45166 13470 45218
rect 13470 45166 13522 45218
rect 13522 45166 13524 45218
rect 13468 45164 13524 45166
rect 13020 43596 13076 43652
rect 12684 42924 12740 42980
rect 12908 42700 12964 42756
rect 12572 40236 12628 40292
rect 12684 41132 12740 41188
rect 12684 39564 12740 39620
rect 13020 41186 13076 41188
rect 13020 41134 13022 41186
rect 13022 41134 13074 41186
rect 13074 41134 13076 41186
rect 13020 41132 13076 41134
rect 13020 40514 13076 40516
rect 13020 40462 13022 40514
rect 13022 40462 13074 40514
rect 13074 40462 13076 40514
rect 13020 40460 13076 40462
rect 12012 36428 12068 36484
rect 12124 38274 12180 38276
rect 12124 38222 12126 38274
rect 12126 38222 12178 38274
rect 12178 38222 12180 38274
rect 12124 38220 12180 38222
rect 12236 37772 12292 37828
rect 12236 37324 12292 37380
rect 12236 35810 12292 35812
rect 12236 35758 12238 35810
rect 12238 35758 12290 35810
rect 12290 35758 12292 35810
rect 12236 35756 12292 35758
rect 12348 35644 12404 35700
rect 12124 34524 12180 34580
rect 11676 32060 11732 32116
rect 11564 31948 11620 32004
rect 11900 34130 11956 34132
rect 11900 34078 11902 34130
rect 11902 34078 11954 34130
rect 11954 34078 11956 34130
rect 11900 34076 11956 34078
rect 11788 31836 11844 31892
rect 11900 31724 11956 31780
rect 12124 31500 12180 31556
rect 12572 37324 12628 37380
rect 11564 31388 11620 31444
rect 11564 30940 11620 30996
rect 11676 30828 11732 30884
rect 11452 29372 11508 29428
rect 11340 28476 11396 28532
rect 10892 27804 10948 27860
rect 10108 24892 10164 24948
rect 10220 26572 10276 26628
rect 10892 27074 10948 27076
rect 10892 27022 10894 27074
rect 10894 27022 10946 27074
rect 10946 27022 10948 27074
rect 10892 27020 10948 27022
rect 11228 28028 11284 28084
rect 12124 28588 12180 28644
rect 11564 28028 11620 28084
rect 11228 26572 11284 26628
rect 11452 27468 11508 27524
rect 11900 27804 11956 27860
rect 10556 25340 10612 25396
rect 10220 22988 10276 23044
rect 9996 22428 10052 22484
rect 10108 21980 10164 22036
rect 9996 21084 10052 21140
rect 9884 20300 9940 20356
rect 10108 20018 10164 20020
rect 10108 19966 10110 20018
rect 10110 19966 10162 20018
rect 10162 19966 10164 20018
rect 10108 19964 10164 19966
rect 9996 19346 10052 19348
rect 9996 19294 9998 19346
rect 9998 19294 10050 19346
rect 10050 19294 10052 19346
rect 9996 19292 10052 19294
rect 10220 19292 10276 19348
rect 9884 18956 9940 19012
rect 10444 23826 10500 23828
rect 10444 23774 10446 23826
rect 10446 23774 10498 23826
rect 10498 23774 10500 23826
rect 10444 23772 10500 23774
rect 10444 22092 10500 22148
rect 10892 24892 10948 24948
rect 10668 23100 10724 23156
rect 10780 24556 10836 24612
rect 10556 20076 10612 20132
rect 10556 18956 10612 19012
rect 10668 18620 10724 18676
rect 10332 18508 10388 18564
rect 9996 16882 10052 16884
rect 9996 16830 9998 16882
rect 9998 16830 10050 16882
rect 10050 16830 10052 16882
rect 9996 16828 10052 16830
rect 9884 15932 9940 15988
rect 10108 15820 10164 15876
rect 10668 15874 10724 15876
rect 10668 15822 10670 15874
rect 10670 15822 10722 15874
rect 10722 15822 10724 15874
rect 10668 15820 10724 15822
rect 10668 15314 10724 15316
rect 10668 15262 10670 15314
rect 10670 15262 10722 15314
rect 10722 15262 10724 15314
rect 10668 15260 10724 15262
rect 9884 14530 9940 14532
rect 9884 14478 9886 14530
rect 9886 14478 9938 14530
rect 9938 14478 9940 14530
rect 9884 14476 9940 14478
rect 9772 13692 9828 13748
rect 9996 13468 10052 13524
rect 9884 11452 9940 11508
rect 9436 10668 9492 10724
rect 9324 9996 9380 10052
rect 9324 9100 9380 9156
rect 9660 10610 9716 10612
rect 9660 10558 9662 10610
rect 9662 10558 9714 10610
rect 9714 10558 9716 10610
rect 9660 10556 9716 10558
rect 9436 8540 9492 8596
rect 9212 7756 9268 7812
rect 9324 8204 9380 8260
rect 9100 7420 9156 7476
rect 8652 6748 8708 6804
rect 8652 4226 8708 4228
rect 8652 4174 8654 4226
rect 8654 4174 8706 4226
rect 8706 4174 8708 4226
rect 8652 4172 8708 4174
rect 8652 2770 8708 2772
rect 8652 2718 8654 2770
rect 8654 2718 8706 2770
rect 8706 2718 8708 2770
rect 8652 2716 8708 2718
rect 8540 1932 8596 1988
rect 8876 6076 8932 6132
rect 9100 5794 9156 5796
rect 9100 5742 9102 5794
rect 9102 5742 9154 5794
rect 9154 5742 9156 5794
rect 9100 5740 9156 5742
rect 9100 5404 9156 5460
rect 9100 4620 9156 4676
rect 9436 6860 9492 6916
rect 9548 7532 9604 7588
rect 9772 9826 9828 9828
rect 9772 9774 9774 9826
rect 9774 9774 9826 9826
rect 9826 9774 9828 9826
rect 9772 9772 9828 9774
rect 9772 8316 9828 8372
rect 9772 7980 9828 8036
rect 9772 7474 9828 7476
rect 9772 7422 9774 7474
rect 9774 7422 9826 7474
rect 9826 7422 9828 7474
rect 9772 7420 9828 7422
rect 9772 6524 9828 6580
rect 9324 4620 9380 4676
rect 9548 5404 9604 5460
rect 9212 4508 9268 4564
rect 9660 5516 9716 5572
rect 9548 5068 9604 5124
rect 9548 4060 9604 4116
rect 8988 3052 9044 3108
rect 9100 3724 9156 3780
rect 8316 1596 8372 1652
rect 8540 1596 8596 1652
rect 9324 3276 9380 3332
rect 9212 2940 9268 2996
rect 9436 3164 9492 3220
rect 9212 2716 9268 2772
rect 9772 4732 9828 4788
rect 9996 10556 10052 10612
rect 9996 9772 10052 9828
rect 10108 9436 10164 9492
rect 9996 8370 10052 8372
rect 9996 8318 9998 8370
rect 9998 8318 10050 8370
rect 10050 8318 10052 8370
rect 9996 8316 10052 8318
rect 10444 14700 10500 14756
rect 10444 13916 10500 13972
rect 10332 13468 10388 13524
rect 10332 12850 10388 12852
rect 10332 12798 10334 12850
rect 10334 12798 10386 12850
rect 10386 12798 10388 12850
rect 10332 12796 10388 12798
rect 10668 13580 10724 13636
rect 10556 11676 10612 11732
rect 10444 11564 10500 11620
rect 10444 11394 10500 11396
rect 10444 11342 10446 11394
rect 10446 11342 10498 11394
rect 10498 11342 10500 11394
rect 10444 11340 10500 11342
rect 10332 10332 10388 10388
rect 11004 23154 11060 23156
rect 11004 23102 11006 23154
rect 11006 23102 11058 23154
rect 11058 23102 11060 23154
rect 11004 23100 11060 23102
rect 11228 20802 11284 20804
rect 11228 20750 11230 20802
rect 11230 20750 11282 20802
rect 11282 20750 11284 20802
rect 11228 20748 11284 20750
rect 11228 19292 11284 19348
rect 11116 19234 11172 19236
rect 11116 19182 11118 19234
rect 11118 19182 11170 19234
rect 11170 19182 11172 19234
rect 11116 19180 11172 19182
rect 10892 14812 10948 14868
rect 11676 27132 11732 27188
rect 11564 26236 11620 26292
rect 11564 25452 11620 25508
rect 11900 26290 11956 26292
rect 11900 26238 11902 26290
rect 11902 26238 11954 26290
rect 11954 26238 11956 26290
rect 11900 26236 11956 26238
rect 12124 26348 12180 26404
rect 11900 25788 11956 25844
rect 11564 22540 11620 22596
rect 11676 22146 11732 22148
rect 11676 22094 11678 22146
rect 11678 22094 11730 22146
rect 11730 22094 11732 22146
rect 11676 22092 11732 22094
rect 11676 20188 11732 20244
rect 11228 17948 11284 18004
rect 11340 18956 11396 19012
rect 11564 17836 11620 17892
rect 11676 18284 11732 18340
rect 11452 17724 11508 17780
rect 11340 17276 11396 17332
rect 11116 16658 11172 16660
rect 11116 16606 11118 16658
rect 11118 16606 11170 16658
rect 11170 16606 11172 16658
rect 11116 16604 11172 16606
rect 11228 16210 11284 16212
rect 11228 16158 11230 16210
rect 11230 16158 11282 16210
rect 11282 16158 11284 16210
rect 11228 16156 11284 16158
rect 11004 14588 11060 14644
rect 11116 15596 11172 15652
rect 10780 13244 10836 13300
rect 10668 10108 10724 10164
rect 10892 12796 10948 12852
rect 10892 12066 10948 12068
rect 10892 12014 10894 12066
rect 10894 12014 10946 12066
rect 10946 12014 10948 12066
rect 10892 12012 10948 12014
rect 10780 11788 10836 11844
rect 10444 9436 10500 9492
rect 10668 9100 10724 9156
rect 10220 8428 10276 8484
rect 11564 17276 11620 17332
rect 11564 16210 11620 16212
rect 11564 16158 11566 16210
rect 11566 16158 11618 16210
rect 11618 16158 11620 16210
rect 11564 16156 11620 16158
rect 11564 15932 11620 15988
rect 11340 14364 11396 14420
rect 11228 13692 11284 13748
rect 11228 12236 11284 12292
rect 11004 11004 11060 11060
rect 11004 10780 11060 10836
rect 10892 10498 10948 10500
rect 10892 10446 10894 10498
rect 10894 10446 10946 10498
rect 10946 10446 10948 10498
rect 10892 10444 10948 10446
rect 10780 8316 10836 8372
rect 11228 11564 11284 11620
rect 11004 8988 11060 9044
rect 11004 8428 11060 8484
rect 11116 8540 11172 8596
rect 10220 7644 10276 7700
rect 10108 6690 10164 6692
rect 10108 6638 10110 6690
rect 10110 6638 10162 6690
rect 10162 6638 10164 6690
rect 10108 6636 10164 6638
rect 9996 6524 10052 6580
rect 10556 7586 10612 7588
rect 10556 7534 10558 7586
rect 10558 7534 10610 7586
rect 10610 7534 10612 7586
rect 10556 7532 10612 7534
rect 10780 7084 10836 7140
rect 10332 5964 10388 6020
rect 9996 5516 10052 5572
rect 8652 1148 8708 1204
rect 8764 1596 8820 1652
rect 8988 1372 9044 1428
rect 10556 5682 10612 5684
rect 10556 5630 10558 5682
rect 10558 5630 10610 5682
rect 10610 5630 10612 5682
rect 10556 5628 10612 5630
rect 10668 5404 10724 5460
rect 11004 7756 11060 7812
rect 11004 7532 11060 7588
rect 11564 10780 11620 10836
rect 11564 10610 11620 10612
rect 11564 10558 11566 10610
rect 11566 10558 11618 10610
rect 11618 10558 11620 10610
rect 11564 10556 11620 10558
rect 11340 8540 11396 8596
rect 11004 7250 11060 7252
rect 11004 7198 11006 7250
rect 11006 7198 11058 7250
rect 11058 7198 11060 7250
rect 11004 7196 11060 7198
rect 11564 7868 11620 7924
rect 11452 6860 11508 6916
rect 12124 24108 12180 24164
rect 12236 25116 12292 25172
rect 11900 23996 11956 24052
rect 12012 23042 12068 23044
rect 12012 22990 12014 23042
rect 12014 22990 12066 23042
rect 12066 22990 12068 23042
rect 12012 22988 12068 22990
rect 11900 19404 11956 19460
rect 12012 22428 12068 22484
rect 11900 19234 11956 19236
rect 11900 19182 11902 19234
rect 11902 19182 11954 19234
rect 11954 19182 11956 19234
rect 11900 19180 11956 19182
rect 11900 18508 11956 18564
rect 12012 18450 12068 18452
rect 12012 18398 12014 18450
rect 12014 18398 12066 18450
rect 12066 18398 12068 18450
rect 12012 18396 12068 18398
rect 12124 20524 12180 20580
rect 11900 16268 11956 16324
rect 12012 16044 12068 16100
rect 11788 15820 11844 15876
rect 11788 15372 11844 15428
rect 11900 14924 11956 14980
rect 11900 14252 11956 14308
rect 12460 35026 12516 35028
rect 12460 34974 12462 35026
rect 12462 34974 12514 35026
rect 12514 34974 12516 35026
rect 12460 34972 12516 34974
rect 12460 34748 12516 34804
rect 12684 36540 12740 36596
rect 12908 34802 12964 34804
rect 12908 34750 12910 34802
rect 12910 34750 12962 34802
rect 12962 34750 12964 34802
rect 12908 34748 12964 34750
rect 12796 33906 12852 33908
rect 12796 33854 12798 33906
rect 12798 33854 12850 33906
rect 12850 33854 12852 33906
rect 12796 33852 12852 33854
rect 13244 38780 13300 38836
rect 13468 42028 13524 42084
rect 13468 40290 13524 40292
rect 13468 40238 13470 40290
rect 13470 40238 13522 40290
rect 13522 40238 13524 40290
rect 13468 40236 13524 40238
rect 13468 39116 13524 39172
rect 14700 52780 14756 52836
rect 14924 59164 14980 59220
rect 15708 63026 15764 63028
rect 15708 62974 15710 63026
rect 15710 62974 15762 63026
rect 15762 62974 15764 63026
rect 15708 62972 15764 62974
rect 15932 63084 15988 63140
rect 15596 61570 15652 61572
rect 15596 61518 15598 61570
rect 15598 61518 15650 61570
rect 15650 61518 15652 61570
rect 15596 61516 15652 61518
rect 15596 60620 15652 60676
rect 15372 59164 15428 59220
rect 15372 57820 15428 57876
rect 14924 54514 14980 54516
rect 14924 54462 14926 54514
rect 14926 54462 14978 54514
rect 14978 54462 14980 54514
rect 14924 54460 14980 54462
rect 14924 53788 14980 53844
rect 14812 51378 14868 51380
rect 14812 51326 14814 51378
rect 14814 51326 14866 51378
rect 14866 51326 14868 51378
rect 14812 51324 14868 51326
rect 14924 50988 14980 51044
rect 15596 57426 15652 57428
rect 15596 57374 15598 57426
rect 15598 57374 15650 57426
rect 15650 57374 15652 57426
rect 15596 57372 15652 57374
rect 15260 55074 15316 55076
rect 15260 55022 15262 55074
rect 15262 55022 15314 55074
rect 15314 55022 15316 55074
rect 15260 55020 15316 55022
rect 14364 50652 14420 50708
rect 14476 49980 14532 50036
rect 14364 49196 14420 49252
rect 14812 50594 14868 50596
rect 14812 50542 14814 50594
rect 14814 50542 14866 50594
rect 14866 50542 14868 50594
rect 14812 50540 14868 50542
rect 15036 50540 15092 50596
rect 14588 48524 14644 48580
rect 14364 47740 14420 47796
rect 14364 46508 14420 46564
rect 14588 46284 14644 46340
rect 14252 44268 14308 44324
rect 14364 45164 14420 45220
rect 14364 44044 14420 44100
rect 14476 43538 14532 43540
rect 14476 43486 14478 43538
rect 14478 43486 14530 43538
rect 14530 43486 14532 43538
rect 14476 43484 14532 43486
rect 14028 43426 14084 43428
rect 14028 43374 14030 43426
rect 14030 43374 14082 43426
rect 14082 43374 14084 43426
rect 14028 43372 14084 43374
rect 13916 42476 13972 42532
rect 14588 42700 14644 42756
rect 14476 41916 14532 41972
rect 13804 40460 13860 40516
rect 14476 40460 14532 40516
rect 14812 49644 14868 49700
rect 15036 48524 15092 48580
rect 15596 53452 15652 53508
rect 15260 52892 15316 52948
rect 15372 52050 15428 52052
rect 15372 51998 15374 52050
rect 15374 51998 15426 52050
rect 15426 51998 15428 52050
rect 15372 51996 15428 51998
rect 15260 50876 15316 50932
rect 15932 61740 15988 61796
rect 15820 61516 15876 61572
rect 16268 62636 16324 62692
rect 16156 62076 16212 62132
rect 15932 61346 15988 61348
rect 15932 61294 15934 61346
rect 15934 61294 15986 61346
rect 15986 61294 15988 61346
rect 15932 61292 15988 61294
rect 15932 60674 15988 60676
rect 15932 60622 15934 60674
rect 15934 60622 15986 60674
rect 15986 60622 15988 60674
rect 15932 60620 15988 60622
rect 16156 53564 16212 53620
rect 15820 50428 15876 50484
rect 15260 50092 15316 50148
rect 15484 50204 15540 50260
rect 15148 49868 15204 49924
rect 15036 48300 15092 48356
rect 14924 48188 14980 48244
rect 14812 48018 14868 48020
rect 14812 47966 14814 48018
rect 14814 47966 14866 48018
rect 14866 47966 14868 48018
rect 14812 47964 14868 47966
rect 14924 47404 14980 47460
rect 14812 46396 14868 46452
rect 14812 43036 14868 43092
rect 14812 40908 14868 40964
rect 13916 39618 13972 39620
rect 13916 39566 13918 39618
rect 13918 39566 13970 39618
rect 13970 39566 13972 39618
rect 13916 39564 13972 39566
rect 13580 38332 13636 38388
rect 14028 38834 14084 38836
rect 14028 38782 14030 38834
rect 14030 38782 14082 38834
rect 14082 38782 14084 38834
rect 14028 38780 14084 38782
rect 14252 38332 14308 38388
rect 13916 37938 13972 37940
rect 13916 37886 13918 37938
rect 13918 37886 13970 37938
rect 13970 37886 13972 37938
rect 13916 37884 13972 37886
rect 14364 37884 14420 37940
rect 13580 36428 13636 36484
rect 14476 37212 14532 37268
rect 14364 36482 14420 36484
rect 14364 36430 14366 36482
rect 14366 36430 14418 36482
rect 14418 36430 14420 36482
rect 14364 36428 14420 36430
rect 14252 36092 14308 36148
rect 13244 34972 13300 35028
rect 13132 31554 13188 31556
rect 13132 31502 13134 31554
rect 13134 31502 13186 31554
rect 13186 31502 13188 31554
rect 13132 31500 13188 31502
rect 13356 32732 13412 32788
rect 12796 30828 12852 30884
rect 12460 30044 12516 30100
rect 13020 29372 13076 29428
rect 12684 27804 12740 27860
rect 12572 27020 12628 27076
rect 12684 26908 12740 26964
rect 12348 22428 12404 22484
rect 12460 26236 12516 26292
rect 12348 21980 12404 22036
rect 13468 29932 13524 29988
rect 13244 28642 13300 28644
rect 13244 28590 13246 28642
rect 13246 28590 13298 28642
rect 13298 28590 13300 28642
rect 13244 28588 13300 28590
rect 13020 27244 13076 27300
rect 12908 25788 12964 25844
rect 12908 25618 12964 25620
rect 12908 25566 12910 25618
rect 12910 25566 12962 25618
rect 12962 25566 12964 25618
rect 12908 25564 12964 25566
rect 12572 25228 12628 25284
rect 12684 24444 12740 24500
rect 12460 21420 12516 21476
rect 12572 24108 12628 24164
rect 12460 19740 12516 19796
rect 13020 24834 13076 24836
rect 13020 24782 13022 24834
rect 13022 24782 13074 24834
rect 13074 24782 13076 24834
rect 13020 24780 13076 24782
rect 12908 23996 12964 24052
rect 13916 35980 13972 36036
rect 13916 35138 13972 35140
rect 13916 35086 13918 35138
rect 13918 35086 13970 35138
rect 13970 35086 13972 35138
rect 13916 35084 13972 35086
rect 13804 34914 13860 34916
rect 13804 34862 13806 34914
rect 13806 34862 13858 34914
rect 13858 34862 13860 34914
rect 13804 34860 13860 34862
rect 14140 34076 14196 34132
rect 13692 33628 13748 33684
rect 14252 32508 14308 32564
rect 14028 32338 14084 32340
rect 14028 32286 14030 32338
rect 14030 32286 14082 32338
rect 14082 32286 14084 32338
rect 14028 32284 14084 32286
rect 14700 38722 14756 38724
rect 14700 38670 14702 38722
rect 14702 38670 14754 38722
rect 14754 38670 14756 38722
rect 14700 38668 14756 38670
rect 15372 49698 15428 49700
rect 15372 49646 15374 49698
rect 15374 49646 15426 49698
rect 15426 49646 15428 49698
rect 15372 49644 15428 49646
rect 15260 48914 15316 48916
rect 15260 48862 15262 48914
rect 15262 48862 15314 48914
rect 15314 48862 15316 48914
rect 15260 48860 15316 48862
rect 15260 45276 15316 45332
rect 15036 43484 15092 43540
rect 15036 43314 15092 43316
rect 15036 43262 15038 43314
rect 15038 43262 15090 43314
rect 15090 43262 15092 43314
rect 15036 43260 15092 43262
rect 15036 42924 15092 42980
rect 15484 43932 15540 43988
rect 14700 35980 14756 36036
rect 15036 37996 15092 38052
rect 15036 37266 15092 37268
rect 15036 37214 15038 37266
rect 15038 37214 15090 37266
rect 15090 37214 15092 37266
rect 15036 37212 15092 37214
rect 15036 35980 15092 36036
rect 14812 34972 14868 35028
rect 14924 34188 14980 34244
rect 14700 34130 14756 34132
rect 14700 34078 14702 34130
rect 14702 34078 14754 34130
rect 14754 34078 14756 34130
rect 14700 34076 14756 34078
rect 13692 31388 13748 31444
rect 13580 29372 13636 29428
rect 14252 30156 14308 30212
rect 14028 29372 14084 29428
rect 13804 28812 13860 28868
rect 13916 28754 13972 28756
rect 13916 28702 13918 28754
rect 13918 28702 13970 28754
rect 13970 28702 13972 28754
rect 13916 28700 13972 28702
rect 13580 27692 13636 27748
rect 13916 28252 13972 28308
rect 13356 24332 13412 24388
rect 12796 23436 12852 23492
rect 13244 23212 13300 23268
rect 13020 22652 13076 22708
rect 13132 22540 13188 22596
rect 13132 22092 13188 22148
rect 12796 21756 12852 21812
rect 13244 21868 13300 21924
rect 13468 22652 13524 22708
rect 13468 22092 13524 22148
rect 13916 26796 13972 26852
rect 14140 27356 14196 27412
rect 14364 29426 14420 29428
rect 14364 29374 14366 29426
rect 14366 29374 14418 29426
rect 14418 29374 14420 29426
rect 14364 29372 14420 29374
rect 14252 27244 14308 27300
rect 14364 28812 14420 28868
rect 14028 26236 14084 26292
rect 13916 25788 13972 25844
rect 14028 25676 14084 25732
rect 13580 21868 13636 21924
rect 12796 21196 12852 21252
rect 13468 21196 13524 21252
rect 12684 21084 12740 21140
rect 12348 19516 12404 19572
rect 12236 16098 12292 16100
rect 12236 16046 12238 16098
rect 12238 16046 12290 16098
rect 12290 16046 12292 16098
rect 12236 16044 12292 16046
rect 12572 19346 12628 19348
rect 12572 19294 12574 19346
rect 12574 19294 12626 19346
rect 12626 19294 12628 19346
rect 12572 19292 12628 19294
rect 12124 15372 12180 15428
rect 12460 18396 12516 18452
rect 12236 13634 12292 13636
rect 12236 13582 12238 13634
rect 12238 13582 12290 13634
rect 12290 13582 12292 13634
rect 12236 13580 12292 13582
rect 13132 20802 13188 20804
rect 13132 20750 13134 20802
rect 13134 20750 13186 20802
rect 13186 20750 13188 20802
rect 13132 20748 13188 20750
rect 13132 20018 13188 20020
rect 13132 19966 13134 20018
rect 13134 19966 13186 20018
rect 13186 19966 13188 20018
rect 13132 19964 13188 19966
rect 13244 19292 13300 19348
rect 13020 19068 13076 19124
rect 13020 18562 13076 18564
rect 13020 18510 13022 18562
rect 13022 18510 13074 18562
rect 13074 18510 13076 18562
rect 13020 18508 13076 18510
rect 12908 17106 12964 17108
rect 12908 17054 12910 17106
rect 12910 17054 12962 17106
rect 12962 17054 12964 17106
rect 12908 17052 12964 17054
rect 12908 16210 12964 16212
rect 12908 16158 12910 16210
rect 12910 16158 12962 16210
rect 12962 16158 12964 16210
rect 12908 16156 12964 16158
rect 12796 15820 12852 15876
rect 12460 15372 12516 15428
rect 12460 14924 12516 14980
rect 12572 15260 12628 15316
rect 12460 14754 12516 14756
rect 12460 14702 12462 14754
rect 12462 14702 12514 14754
rect 12514 14702 12516 14754
rect 12460 14700 12516 14702
rect 12348 13468 12404 13524
rect 12460 14140 12516 14196
rect 12012 12684 12068 12740
rect 11900 12572 11956 12628
rect 11900 12236 11956 12292
rect 12124 12178 12180 12180
rect 12124 12126 12126 12178
rect 12126 12126 12178 12178
rect 12178 12126 12180 12178
rect 12124 12124 12180 12126
rect 12012 11900 12068 11956
rect 11900 10892 11956 10948
rect 12012 11340 12068 11396
rect 11900 10332 11956 10388
rect 11788 9826 11844 9828
rect 11788 9774 11790 9826
rect 11790 9774 11842 9826
rect 11842 9774 11844 9826
rect 11788 9772 11844 9774
rect 12684 14476 12740 14532
rect 12348 11004 12404 11060
rect 11900 9548 11956 9604
rect 10892 6578 10948 6580
rect 10892 6526 10894 6578
rect 10894 6526 10946 6578
rect 10946 6526 10948 6578
rect 10892 6524 10948 6526
rect 10892 5404 10948 5460
rect 10108 2940 10164 2996
rect 9548 1708 9604 1764
rect 9660 1596 9716 1652
rect 9436 924 9492 980
rect 9548 364 9604 420
rect 10220 2044 10276 2100
rect 10556 4338 10612 4340
rect 10556 4286 10558 4338
rect 10558 4286 10610 4338
rect 10610 4286 10612 4338
rect 10556 4284 10612 4286
rect 11228 5122 11284 5124
rect 11228 5070 11230 5122
rect 11230 5070 11282 5122
rect 11282 5070 11284 5122
rect 11228 5068 11284 5070
rect 11228 4114 11284 4116
rect 11228 4062 11230 4114
rect 11230 4062 11282 4114
rect 11282 4062 11284 4114
rect 11228 4060 11284 4062
rect 10668 3948 10724 4004
rect 10556 2380 10612 2436
rect 10444 1932 10500 1988
rect 10108 1874 10164 1876
rect 10108 1822 10110 1874
rect 10110 1822 10162 1874
rect 10162 1822 10164 1874
rect 10108 1820 10164 1822
rect 10108 1596 10164 1652
rect 10332 1596 10388 1652
rect 10220 1036 10276 1092
rect 10892 3778 10948 3780
rect 10892 3726 10894 3778
rect 10894 3726 10946 3778
rect 10946 3726 10948 3778
rect 10892 3724 10948 3726
rect 11228 3500 11284 3556
rect 10892 3276 10948 3332
rect 12124 9772 12180 9828
rect 12236 10892 12292 10948
rect 12124 9042 12180 9044
rect 12124 8990 12126 9042
rect 12126 8990 12178 9042
rect 12178 8990 12180 9042
rect 12124 8988 12180 8990
rect 12124 8316 12180 8372
rect 12572 12850 12628 12852
rect 12572 12798 12574 12850
rect 12574 12798 12626 12850
rect 12626 12798 12628 12850
rect 12572 12796 12628 12798
rect 12460 10332 12516 10388
rect 12460 10108 12516 10164
rect 12908 15202 12964 15204
rect 12908 15150 12910 15202
rect 12910 15150 12962 15202
rect 12962 15150 12964 15202
rect 12908 15148 12964 15150
rect 12908 14924 12964 14980
rect 13020 13580 13076 13636
rect 13020 13244 13076 13300
rect 13020 13020 13076 13076
rect 12796 12236 12852 12292
rect 12796 10892 12852 10948
rect 12908 10556 12964 10612
rect 12572 9100 12628 9156
rect 12796 8204 12852 8260
rect 13020 8876 13076 8932
rect 13132 8818 13188 8820
rect 13132 8766 13134 8818
rect 13134 8766 13186 8818
rect 13186 8766 13188 8818
rect 13132 8764 13188 8766
rect 13020 8370 13076 8372
rect 13020 8318 13022 8370
rect 13022 8318 13074 8370
rect 13074 8318 13076 8370
rect 13020 8316 13076 8318
rect 12908 7980 12964 8036
rect 14252 25004 14308 25060
rect 14140 24780 14196 24836
rect 14140 23884 14196 23940
rect 14812 31836 14868 31892
rect 14924 32508 14980 32564
rect 14812 30210 14868 30212
rect 14812 30158 14814 30210
rect 14814 30158 14866 30210
rect 14866 30158 14868 30210
rect 14812 30156 14868 30158
rect 15372 41916 15428 41972
rect 15260 38780 15316 38836
rect 15484 38444 15540 38500
rect 15260 37042 15316 37044
rect 15260 36990 15262 37042
rect 15262 36990 15314 37042
rect 15314 36990 15316 37042
rect 15260 36988 15316 36990
rect 15260 33906 15316 33908
rect 15260 33854 15262 33906
rect 15262 33854 15314 33906
rect 15314 33854 15316 33906
rect 15260 33852 15316 33854
rect 15148 33068 15204 33124
rect 15148 32732 15204 32788
rect 15148 32396 15204 32452
rect 16156 49810 16212 49812
rect 16156 49758 16158 49810
rect 16158 49758 16210 49810
rect 16210 49758 16212 49810
rect 16156 49756 16212 49758
rect 16828 75068 16884 75124
rect 16716 74786 16772 74788
rect 16716 74734 16718 74786
rect 16718 74734 16770 74786
rect 16770 74734 16772 74786
rect 16716 74732 16772 74734
rect 16716 74338 16772 74340
rect 16716 74286 16718 74338
rect 16718 74286 16770 74338
rect 16770 74286 16772 74338
rect 16716 74284 16772 74286
rect 16604 74060 16660 74116
rect 16716 73276 16772 73332
rect 16828 71708 16884 71764
rect 17052 75068 17108 75124
rect 17052 74898 17108 74900
rect 17052 74846 17054 74898
rect 17054 74846 17106 74898
rect 17106 74846 17108 74898
rect 17052 74844 17108 74846
rect 17052 74620 17108 74676
rect 16940 71372 16996 71428
rect 17052 74060 17108 74116
rect 16828 70476 16884 70532
rect 16940 69410 16996 69412
rect 16940 69358 16942 69410
rect 16942 69358 16994 69410
rect 16994 69358 16996 69410
rect 16940 69356 16996 69358
rect 16828 68012 16884 68068
rect 16716 67676 16772 67732
rect 17388 88898 17444 88900
rect 17388 88846 17390 88898
rect 17390 88846 17442 88898
rect 17442 88846 17444 88898
rect 17388 88844 17444 88846
rect 17500 88732 17556 88788
rect 17500 87388 17556 87444
rect 17388 86828 17444 86884
rect 17388 85314 17444 85316
rect 17388 85262 17390 85314
rect 17390 85262 17442 85314
rect 17442 85262 17444 85314
rect 17388 85260 17444 85262
rect 17276 84476 17332 84532
rect 17276 78988 17332 79044
rect 17500 83916 17556 83972
rect 17836 85932 17892 85988
rect 18060 89292 18116 89348
rect 18172 90300 18228 90356
rect 18284 88732 18340 88788
rect 18508 92764 18564 92820
rect 18508 92540 18564 92596
rect 18956 96178 19012 96180
rect 18956 96126 18958 96178
rect 18958 96126 19010 96178
rect 19010 96126 19012 96178
rect 18956 96124 19012 96126
rect 18956 95452 19012 95508
rect 18844 94444 18900 94500
rect 18732 92706 18788 92708
rect 18732 92654 18734 92706
rect 18734 92654 18786 92706
rect 18786 92654 18788 92706
rect 18732 92652 18788 92654
rect 18620 91532 18676 91588
rect 18732 91084 18788 91140
rect 18844 91308 18900 91364
rect 18508 88786 18564 88788
rect 18508 88734 18510 88786
rect 18510 88734 18562 88786
rect 18562 88734 18564 88786
rect 18508 88732 18564 88734
rect 18396 88338 18452 88340
rect 18396 88286 18398 88338
rect 18398 88286 18450 88338
rect 18450 88286 18452 88338
rect 18396 88284 18452 88286
rect 18060 87612 18116 87668
rect 17724 84252 17780 84308
rect 17836 84028 17892 84084
rect 18060 84306 18116 84308
rect 18060 84254 18062 84306
rect 18062 84254 18114 84306
rect 18114 84254 18116 84306
rect 18060 84252 18116 84254
rect 17612 79100 17668 79156
rect 18060 82796 18116 82852
rect 17500 78988 17556 79044
rect 17836 79602 17892 79604
rect 17836 79550 17838 79602
rect 17838 79550 17890 79602
rect 17890 79550 17892 79602
rect 17836 79548 17892 79550
rect 17612 78764 17668 78820
rect 17388 77362 17444 77364
rect 17388 77310 17390 77362
rect 17390 77310 17442 77362
rect 17442 77310 17444 77362
rect 17388 77308 17444 77310
rect 17276 76300 17332 76356
rect 17612 77308 17668 77364
rect 17388 75516 17444 75572
rect 17500 75906 17556 75908
rect 17500 75854 17502 75906
rect 17502 75854 17554 75906
rect 17554 75854 17556 75906
rect 17500 75852 17556 75854
rect 17724 76524 17780 76580
rect 17948 76412 18004 76468
rect 17836 75068 17892 75124
rect 17724 74674 17780 74676
rect 17724 74622 17726 74674
rect 17726 74622 17778 74674
rect 17778 74622 17780 74674
rect 17724 74620 17780 74622
rect 17388 74060 17444 74116
rect 17388 72770 17444 72772
rect 17388 72718 17390 72770
rect 17390 72718 17442 72770
rect 17442 72718 17444 72770
rect 17388 72716 17444 72718
rect 17276 70028 17332 70084
rect 17276 69522 17332 69524
rect 17276 69470 17278 69522
rect 17278 69470 17330 69522
rect 17330 69470 17332 69522
rect 17276 69468 17332 69470
rect 17276 68908 17332 68964
rect 17164 67172 17220 67228
rect 17164 66892 17220 66948
rect 16828 63756 16884 63812
rect 16828 63084 16884 63140
rect 16940 65548 16996 65604
rect 17388 66668 17444 66724
rect 17724 74060 17780 74116
rect 17612 74002 17668 74004
rect 17612 73950 17614 74002
rect 17614 73950 17666 74002
rect 17666 73950 17668 74002
rect 17612 73948 17668 73950
rect 17612 72156 17668 72212
rect 17724 70194 17780 70196
rect 17724 70142 17726 70194
rect 17726 70142 17778 70194
rect 17778 70142 17780 70194
rect 17724 70140 17780 70142
rect 17612 68796 17668 68852
rect 17612 67452 17668 67508
rect 16828 62636 16884 62692
rect 16940 62076 16996 62132
rect 16716 61346 16772 61348
rect 16716 61294 16718 61346
rect 16718 61294 16770 61346
rect 16770 61294 16772 61346
rect 16716 61292 16772 61294
rect 16604 60172 16660 60228
rect 17836 67954 17892 67956
rect 17836 67902 17838 67954
rect 17838 67902 17890 67954
rect 17890 67902 17892 67954
rect 17836 67900 17892 67902
rect 17836 66220 17892 66276
rect 17388 63868 17444 63924
rect 17388 63532 17444 63588
rect 17276 62354 17332 62356
rect 17276 62302 17278 62354
rect 17278 62302 17330 62354
rect 17330 62302 17332 62354
rect 17276 62300 17332 62302
rect 17500 63362 17556 63364
rect 17500 63310 17502 63362
rect 17502 63310 17554 63362
rect 17554 63310 17556 63362
rect 17500 63308 17556 63310
rect 17500 63084 17556 63140
rect 17276 61852 17332 61908
rect 17164 61628 17220 61684
rect 17052 61570 17108 61572
rect 17052 61518 17054 61570
rect 17054 61518 17106 61570
rect 17106 61518 17108 61570
rect 17052 61516 17108 61518
rect 17164 60956 17220 61012
rect 17388 61180 17444 61236
rect 16604 60002 16660 60004
rect 16604 59950 16606 60002
rect 16606 59950 16658 60002
rect 16658 59950 16660 60002
rect 16604 59948 16660 59950
rect 16828 59218 16884 59220
rect 16828 59166 16830 59218
rect 16830 59166 16882 59218
rect 16882 59166 16884 59218
rect 16828 59164 16884 59166
rect 16492 58828 16548 58884
rect 16716 59052 16772 59108
rect 17724 63698 17780 63700
rect 17724 63646 17726 63698
rect 17726 63646 17778 63698
rect 17778 63646 17780 63698
rect 17724 63644 17780 63646
rect 18732 90636 18788 90692
rect 18844 90578 18900 90580
rect 18844 90526 18846 90578
rect 18846 90526 18898 90578
rect 18898 90526 18900 90578
rect 18844 90524 18900 90526
rect 18732 88956 18788 89012
rect 18844 87218 18900 87220
rect 18844 87166 18846 87218
rect 18846 87166 18898 87218
rect 18898 87166 18900 87218
rect 18844 87164 18900 87166
rect 18956 86604 19012 86660
rect 19516 97020 19572 97076
rect 19516 95954 19572 95956
rect 19516 95902 19518 95954
rect 19518 95902 19570 95954
rect 19570 95902 19572 95954
rect 19516 95900 19572 95902
rect 19628 94668 19684 94724
rect 20076 107548 20132 107604
rect 20636 112588 20692 112644
rect 20748 112700 20804 112756
rect 20412 111020 20468 111076
rect 20524 111580 20580 111636
rect 20076 105084 20132 105140
rect 20636 111468 20692 111524
rect 20860 111132 20916 111188
rect 20636 109228 20692 109284
rect 19964 103794 20020 103796
rect 19964 103742 19966 103794
rect 19966 103742 20018 103794
rect 20018 103742 20020 103794
rect 19964 103740 20020 103742
rect 19852 98812 19908 98868
rect 19964 99148 20020 99204
rect 19852 98194 19908 98196
rect 19852 98142 19854 98194
rect 19854 98142 19906 98194
rect 19906 98142 19908 98194
rect 19852 98140 19908 98142
rect 19964 96290 20020 96292
rect 19964 96238 19966 96290
rect 19966 96238 20018 96290
rect 20018 96238 20020 96290
rect 19964 96236 20020 96238
rect 20300 98812 20356 98868
rect 19852 95228 19908 95284
rect 19292 94274 19348 94276
rect 19292 94222 19294 94274
rect 19294 94222 19346 94274
rect 19346 94222 19348 94274
rect 19292 94220 19348 94222
rect 19180 93490 19236 93492
rect 19180 93438 19182 93490
rect 19182 93438 19234 93490
rect 19234 93438 19236 93490
rect 19180 93436 19236 93438
rect 19516 93490 19572 93492
rect 19516 93438 19518 93490
rect 19518 93438 19570 93490
rect 19570 93438 19572 93490
rect 19516 93436 19572 93438
rect 19404 92652 19460 92708
rect 19292 92428 19348 92484
rect 19292 91644 19348 91700
rect 19180 90860 19236 90916
rect 19516 91922 19572 91924
rect 19516 91870 19518 91922
rect 19518 91870 19570 91922
rect 19570 91870 19572 91922
rect 19516 91868 19572 91870
rect 19516 91644 19572 91700
rect 19740 93100 19796 93156
rect 19964 94444 20020 94500
rect 20076 94668 20132 94724
rect 19852 92540 19908 92596
rect 19740 91362 19796 91364
rect 19740 91310 19742 91362
rect 19742 91310 19794 91362
rect 19794 91310 19796 91362
rect 19740 91308 19796 91310
rect 20188 94498 20244 94500
rect 20188 94446 20190 94498
rect 20190 94446 20242 94498
rect 20242 94446 20244 94498
rect 20188 94444 20244 94446
rect 20188 94220 20244 94276
rect 20188 91420 20244 91476
rect 19292 87948 19348 88004
rect 19180 85932 19236 85988
rect 18620 84812 18676 84868
rect 18508 82514 18564 82516
rect 18508 82462 18510 82514
rect 18510 82462 18562 82514
rect 18562 82462 18564 82514
rect 18508 82460 18564 82462
rect 18172 82236 18228 82292
rect 18396 81340 18452 81396
rect 18172 78818 18228 78820
rect 18172 78766 18174 78818
rect 18174 78766 18226 78818
rect 18226 78766 18228 78818
rect 18172 78764 18228 78766
rect 18844 80780 18900 80836
rect 18732 79548 18788 79604
rect 18172 76972 18228 77028
rect 18508 77026 18564 77028
rect 18508 76974 18510 77026
rect 18510 76974 18562 77026
rect 18562 76974 18564 77026
rect 18508 76972 18564 76974
rect 18396 76412 18452 76468
rect 18732 78204 18788 78260
rect 18732 77810 18788 77812
rect 18732 77758 18734 77810
rect 18734 77758 18786 77810
rect 18786 77758 18788 77810
rect 18732 77756 18788 77758
rect 18060 75852 18116 75908
rect 18732 75068 18788 75124
rect 18844 76300 18900 76356
rect 18396 74172 18452 74228
rect 18620 74060 18676 74116
rect 18060 73500 18116 73556
rect 18172 73948 18228 74004
rect 18396 73554 18452 73556
rect 18396 73502 18398 73554
rect 18398 73502 18450 73554
rect 18450 73502 18452 73554
rect 18396 73500 18452 73502
rect 19068 84476 19124 84532
rect 19068 84140 19124 84196
rect 19628 88002 19684 88004
rect 19628 87950 19630 88002
rect 19630 87950 19682 88002
rect 19682 87950 19684 88002
rect 19628 87948 19684 87950
rect 19628 87052 19684 87108
rect 20076 90748 20132 90804
rect 19852 87052 19908 87108
rect 19852 86770 19908 86772
rect 19852 86718 19854 86770
rect 19854 86718 19906 86770
rect 19906 86718 19908 86770
rect 19852 86716 19908 86718
rect 19404 85932 19460 85988
rect 19404 85762 19460 85764
rect 19404 85710 19406 85762
rect 19406 85710 19458 85762
rect 19458 85710 19460 85762
rect 19404 85708 19460 85710
rect 20188 87052 20244 87108
rect 19628 85260 19684 85316
rect 19740 85090 19796 85092
rect 19740 85038 19742 85090
rect 19742 85038 19794 85090
rect 19794 85038 19796 85090
rect 19740 85036 19796 85038
rect 19964 85036 20020 85092
rect 19404 84700 19460 84756
rect 19852 84812 19908 84868
rect 19292 84364 19348 84420
rect 19628 84588 19684 84644
rect 19740 84364 19796 84420
rect 19292 84028 19348 84084
rect 19516 83244 19572 83300
rect 19404 81954 19460 81956
rect 19404 81902 19406 81954
rect 19406 81902 19458 81954
rect 19458 81902 19460 81954
rect 19404 81900 19460 81902
rect 19292 81228 19348 81284
rect 18284 71762 18340 71764
rect 18284 71710 18286 71762
rect 18286 71710 18338 71762
rect 18338 71710 18340 71762
rect 18284 71708 18340 71710
rect 18172 70082 18228 70084
rect 18172 70030 18174 70082
rect 18174 70030 18226 70082
rect 18226 70030 18228 70082
rect 18172 70028 18228 70030
rect 18284 68908 18340 68964
rect 18060 68012 18116 68068
rect 18172 68796 18228 68852
rect 18396 68236 18452 68292
rect 18172 67452 18228 67508
rect 18284 67116 18340 67172
rect 18172 67004 18228 67060
rect 18172 65548 18228 65604
rect 18508 66444 18564 66500
rect 18508 66274 18564 66276
rect 18508 66222 18510 66274
rect 18510 66222 18562 66274
rect 18562 66222 18564 66274
rect 18508 66220 18564 66222
rect 17724 61852 17780 61908
rect 18508 65996 18564 66052
rect 17612 61794 17668 61796
rect 17612 61742 17614 61794
rect 17614 61742 17666 61794
rect 17666 61742 17668 61794
rect 17612 61740 17668 61742
rect 17612 61068 17668 61124
rect 17948 61852 18004 61908
rect 18396 63308 18452 63364
rect 18172 61682 18228 61684
rect 18172 61630 18174 61682
rect 18174 61630 18226 61682
rect 18226 61630 18228 61682
rect 18172 61628 18228 61630
rect 17724 60956 17780 61012
rect 17836 60844 17892 60900
rect 17500 60060 17556 60116
rect 17724 60284 17780 60340
rect 17052 58658 17108 58660
rect 17052 58606 17054 58658
rect 17054 58606 17106 58658
rect 17106 58606 17108 58658
rect 17052 58604 17108 58606
rect 16716 57148 16772 57204
rect 17948 60284 18004 60340
rect 17948 58604 18004 58660
rect 16380 54460 16436 54516
rect 17164 54514 17220 54516
rect 17164 54462 17166 54514
rect 17166 54462 17218 54514
rect 17218 54462 17220 54514
rect 17164 54460 17220 54462
rect 17164 53676 17220 53732
rect 16492 53340 16548 53396
rect 16828 52722 16884 52724
rect 16828 52670 16830 52722
rect 16830 52670 16882 52722
rect 16882 52670 16884 52722
rect 16828 52668 16884 52670
rect 16828 52444 16884 52500
rect 17052 52274 17108 52276
rect 17052 52222 17054 52274
rect 17054 52222 17106 52274
rect 17106 52222 17108 52274
rect 17052 52220 17108 52222
rect 16380 50204 16436 50260
rect 16268 49644 16324 49700
rect 16156 49532 16212 49588
rect 15932 47458 15988 47460
rect 15932 47406 15934 47458
rect 15934 47406 15986 47458
rect 15986 47406 15988 47458
rect 15932 47404 15988 47406
rect 16044 46060 16100 46116
rect 16044 43148 16100 43204
rect 15708 42754 15764 42756
rect 15708 42702 15710 42754
rect 15710 42702 15762 42754
rect 15762 42702 15764 42754
rect 15708 42700 15764 42702
rect 15820 41468 15876 41524
rect 15820 40348 15876 40404
rect 16380 49586 16436 49588
rect 16380 49534 16382 49586
rect 16382 49534 16434 49586
rect 16434 49534 16436 49586
rect 16380 49532 16436 49534
rect 16604 48524 16660 48580
rect 16940 48300 16996 48356
rect 16604 47852 16660 47908
rect 16828 48188 16884 48244
rect 16604 47292 16660 47348
rect 16380 46562 16436 46564
rect 16380 46510 16382 46562
rect 16382 46510 16434 46562
rect 16434 46510 16436 46562
rect 16380 46508 16436 46510
rect 16268 41804 16324 41860
rect 16380 45948 16436 46004
rect 16604 45948 16660 46004
rect 16604 45500 16660 45556
rect 16604 42924 16660 42980
rect 16492 41916 16548 41972
rect 16268 40460 16324 40516
rect 15932 40236 15988 40292
rect 15708 38834 15764 38836
rect 15708 38782 15710 38834
rect 15710 38782 15762 38834
rect 15762 38782 15764 38834
rect 15708 38780 15764 38782
rect 16044 38444 16100 38500
rect 17276 51154 17332 51156
rect 17276 51102 17278 51154
rect 17278 51102 17330 51154
rect 17330 51102 17332 51154
rect 17276 51100 17332 51102
rect 17948 51548 18004 51604
rect 17948 50652 18004 50708
rect 17948 50428 18004 50484
rect 17388 48860 17444 48916
rect 17500 47516 17556 47572
rect 17052 47458 17108 47460
rect 17052 47406 17054 47458
rect 17054 47406 17106 47458
rect 17106 47406 17108 47458
rect 17052 47404 17108 47406
rect 16828 41916 16884 41972
rect 17276 46284 17332 46340
rect 17164 43538 17220 43540
rect 17164 43486 17166 43538
rect 17166 43486 17218 43538
rect 17218 43486 17220 43538
rect 17164 43484 17220 43486
rect 17836 49084 17892 49140
rect 17948 48524 18004 48580
rect 17836 46114 17892 46116
rect 17836 46062 17838 46114
rect 17838 46062 17890 46114
rect 17890 46062 17892 46114
rect 17836 46060 17892 46062
rect 18172 60674 18228 60676
rect 18172 60622 18174 60674
rect 18174 60622 18226 60674
rect 18226 60622 18228 60674
rect 18172 60620 18228 60622
rect 18732 69804 18788 69860
rect 18844 69468 18900 69524
rect 18956 70476 19012 70532
rect 18956 68908 19012 68964
rect 19628 77868 19684 77924
rect 19404 76748 19460 76804
rect 19516 76466 19572 76468
rect 19516 76414 19518 76466
rect 19518 76414 19570 76466
rect 19570 76414 19572 76466
rect 19516 76412 19572 76414
rect 19740 75068 19796 75124
rect 19740 74114 19796 74116
rect 19740 74062 19742 74114
rect 19742 74062 19794 74114
rect 19794 74062 19796 74114
rect 19740 74060 19796 74062
rect 19292 71932 19348 71988
rect 19180 70140 19236 70196
rect 19628 71820 19684 71876
rect 18844 68124 18900 68180
rect 18844 67676 18900 67732
rect 19068 68514 19124 68516
rect 19068 68462 19070 68514
rect 19070 68462 19122 68514
rect 19122 68462 19124 68514
rect 19068 68460 19124 68462
rect 19292 69132 19348 69188
rect 18732 65996 18788 66052
rect 19180 68012 19236 68068
rect 18844 67004 18900 67060
rect 18732 65100 18788 65156
rect 18956 66444 19012 66500
rect 19516 69522 19572 69524
rect 19516 69470 19518 69522
rect 19518 69470 19570 69522
rect 19570 69470 19572 69522
rect 19516 69468 19572 69470
rect 20076 84700 20132 84756
rect 19964 82066 20020 82068
rect 19964 82014 19966 82066
rect 19966 82014 20018 82066
rect 20018 82014 20020 82066
rect 19964 82012 20020 82014
rect 19964 80780 20020 80836
rect 19964 79548 20020 79604
rect 20076 79212 20132 79268
rect 19964 77250 20020 77252
rect 19964 77198 19966 77250
rect 19966 77198 20018 77250
rect 20018 77198 20020 77250
rect 19964 77196 20020 77198
rect 21084 111916 21140 111972
rect 21196 113260 21252 113316
rect 21532 113484 21588 113540
rect 21756 113372 21812 113428
rect 21868 114044 21924 114100
rect 21308 112812 21364 112868
rect 21084 111020 21140 111076
rect 20860 108780 20916 108836
rect 20860 104130 20916 104132
rect 20860 104078 20862 104130
rect 20862 104078 20914 104130
rect 20914 104078 20916 104130
rect 20860 104076 20916 104078
rect 21308 110962 21364 110964
rect 21308 110910 21310 110962
rect 21310 110910 21362 110962
rect 21362 110910 21364 110962
rect 21308 110908 21364 110910
rect 21084 100940 21140 100996
rect 20972 100268 21028 100324
rect 21756 112700 21812 112756
rect 21980 112924 22036 112980
rect 22428 114044 22484 114100
rect 22316 113820 22372 113876
rect 22876 114492 22932 114548
rect 22988 114604 23044 114660
rect 22652 113820 22708 113876
rect 23324 114380 23380 114436
rect 21532 112028 21588 112084
rect 21532 111858 21588 111860
rect 21532 111806 21534 111858
rect 21534 111806 21586 111858
rect 21586 111806 21588 111858
rect 21532 111804 21588 111806
rect 22204 112700 22260 112756
rect 21868 111970 21924 111972
rect 21868 111918 21870 111970
rect 21870 111918 21922 111970
rect 21922 111918 21924 111970
rect 21868 111916 21924 111918
rect 22204 111858 22260 111860
rect 22204 111806 22206 111858
rect 22206 111806 22258 111858
rect 22258 111806 22260 111858
rect 22204 111804 22260 111806
rect 22204 111468 22260 111524
rect 21756 111020 21812 111076
rect 21980 111132 22036 111188
rect 22092 110796 22148 110852
rect 21644 110460 21700 110516
rect 21532 110236 21588 110292
rect 22316 110908 22372 110964
rect 22316 110012 22372 110068
rect 21756 106204 21812 106260
rect 22204 109900 22260 109956
rect 21420 105420 21476 105476
rect 21868 104300 21924 104356
rect 21196 98812 21252 98868
rect 22876 113260 22932 113316
rect 22652 112140 22708 112196
rect 22764 112028 22820 112084
rect 22428 107324 22484 107380
rect 22652 110572 22708 110628
rect 22652 110402 22708 110404
rect 22652 110350 22654 110402
rect 22654 110350 22706 110402
rect 22706 110350 22708 110402
rect 22652 110348 22708 110350
rect 22652 106092 22708 106148
rect 21756 96684 21812 96740
rect 20972 95900 21028 95956
rect 20412 90748 20468 90804
rect 20524 94892 20580 94948
rect 20636 90524 20692 90580
rect 20860 92988 20916 93044
rect 20860 92764 20916 92820
rect 20860 90748 20916 90804
rect 21084 93884 21140 93940
rect 21868 96626 21924 96628
rect 21868 96574 21870 96626
rect 21870 96574 21922 96626
rect 21922 96574 21924 96626
rect 21868 96572 21924 96574
rect 21756 95954 21812 95956
rect 21756 95902 21758 95954
rect 21758 95902 21810 95954
rect 21810 95902 21812 95954
rect 21756 95900 21812 95902
rect 21084 92146 21140 92148
rect 21084 92094 21086 92146
rect 21086 92094 21138 92146
rect 21138 92094 21140 92146
rect 21084 92092 21140 92094
rect 21308 92092 21364 92148
rect 21644 92876 21700 92932
rect 21644 92652 21700 92708
rect 20972 90636 21028 90692
rect 21196 90636 21252 90692
rect 20636 89404 20692 89460
rect 20524 87500 20580 87556
rect 20636 89180 20692 89236
rect 20524 87164 20580 87220
rect 20412 85314 20468 85316
rect 20412 85262 20414 85314
rect 20414 85262 20466 85314
rect 20466 85262 20468 85314
rect 20412 85260 20468 85262
rect 21196 88226 21252 88228
rect 21196 88174 21198 88226
rect 21198 88174 21250 88226
rect 21250 88174 21252 88226
rect 21196 88172 21252 88174
rect 21532 92316 21588 92372
rect 21868 92204 21924 92260
rect 21756 92092 21812 92148
rect 22204 96796 22260 96852
rect 22316 96684 22372 96740
rect 22092 94444 22148 94500
rect 22204 94220 22260 94276
rect 22988 110908 23044 110964
rect 22876 104860 22932 104916
rect 23996 114716 24052 114772
rect 23772 114268 23828 114324
rect 24220 114156 24276 114212
rect 24668 114604 24724 114660
rect 24444 113932 24500 113988
rect 24464 113706 24520 113708
rect 24464 113654 24466 113706
rect 24466 113654 24518 113706
rect 24518 113654 24520 113706
rect 24464 113652 24520 113654
rect 24568 113706 24624 113708
rect 24568 113654 24570 113706
rect 24570 113654 24622 113706
rect 24622 113654 24624 113706
rect 24568 113652 24624 113654
rect 24672 113706 24728 113708
rect 24672 113654 24674 113706
rect 24674 113654 24726 113706
rect 24726 113654 24728 113706
rect 24672 113652 24728 113654
rect 24556 113538 24612 113540
rect 24556 113486 24558 113538
rect 24558 113486 24610 113538
rect 24610 113486 24612 113538
rect 24556 113484 24612 113486
rect 23548 113148 23604 113204
rect 23436 113036 23492 113092
rect 23324 112924 23380 112980
rect 23212 111356 23268 111412
rect 23324 111244 23380 111300
rect 23324 110572 23380 110628
rect 23212 109340 23268 109396
rect 23100 106316 23156 106372
rect 24668 113372 24724 113428
rect 23804 112922 23860 112924
rect 23804 112870 23806 112922
rect 23806 112870 23858 112922
rect 23858 112870 23860 112922
rect 23804 112868 23860 112870
rect 23908 112922 23964 112924
rect 23908 112870 23910 112922
rect 23910 112870 23962 112922
rect 23962 112870 23964 112922
rect 23908 112868 23964 112870
rect 24012 112922 24068 112924
rect 24012 112870 24014 112922
rect 24014 112870 24066 112922
rect 24066 112870 24068 112922
rect 24012 112868 24068 112870
rect 23660 112364 23716 112420
rect 23996 112700 24052 112756
rect 24220 112700 24276 112756
rect 24332 112812 24388 112868
rect 23660 111580 23716 111636
rect 23996 111468 24052 111524
rect 24220 112252 24276 112308
rect 23804 111354 23860 111356
rect 23804 111302 23806 111354
rect 23806 111302 23858 111354
rect 23858 111302 23860 111354
rect 23804 111300 23860 111302
rect 23908 111354 23964 111356
rect 23908 111302 23910 111354
rect 23910 111302 23962 111354
rect 23962 111302 23964 111354
rect 23908 111300 23964 111302
rect 24012 111354 24068 111356
rect 24012 111302 24014 111354
rect 24014 111302 24066 111354
rect 24066 111302 24068 111354
rect 24012 111300 24068 111302
rect 23884 111132 23940 111188
rect 23660 111020 23716 111076
rect 23548 110348 23604 110404
rect 23996 110962 24052 110964
rect 23996 110910 23998 110962
rect 23998 110910 24050 110962
rect 24050 110910 24052 110962
rect 23996 110908 24052 110910
rect 23804 109786 23860 109788
rect 23804 109734 23806 109786
rect 23806 109734 23858 109786
rect 23858 109734 23860 109786
rect 23804 109732 23860 109734
rect 23908 109786 23964 109788
rect 23908 109734 23910 109786
rect 23910 109734 23962 109786
rect 23962 109734 23964 109786
rect 23908 109732 23964 109734
rect 24012 109786 24068 109788
rect 24012 109734 24014 109786
rect 24014 109734 24066 109786
rect 24066 109734 24068 109786
rect 24012 109732 24068 109734
rect 23660 108332 23716 108388
rect 23804 108218 23860 108220
rect 23804 108166 23806 108218
rect 23806 108166 23858 108218
rect 23858 108166 23860 108218
rect 23804 108164 23860 108166
rect 23908 108218 23964 108220
rect 23908 108166 23910 108218
rect 23910 108166 23962 108218
rect 23962 108166 23964 108218
rect 23908 108164 23964 108166
rect 24012 108218 24068 108220
rect 24012 108166 24014 108218
rect 24014 108166 24066 108218
rect 24066 108166 24068 108218
rect 24012 108164 24068 108166
rect 23804 106650 23860 106652
rect 23804 106598 23806 106650
rect 23806 106598 23858 106650
rect 23858 106598 23860 106650
rect 23804 106596 23860 106598
rect 23908 106650 23964 106652
rect 23908 106598 23910 106650
rect 23910 106598 23962 106650
rect 23962 106598 23964 106650
rect 23908 106596 23964 106598
rect 24012 106650 24068 106652
rect 24012 106598 24014 106650
rect 24014 106598 24066 106650
rect 24066 106598 24068 106650
rect 24012 106596 24068 106598
rect 22988 97692 23044 97748
rect 24780 113314 24836 113316
rect 24780 113262 24782 113314
rect 24782 113262 24834 113314
rect 24834 113262 24836 113314
rect 24780 113260 24836 113262
rect 25116 113036 25172 113092
rect 24892 112476 24948 112532
rect 24892 112252 24948 112308
rect 24464 112138 24520 112140
rect 24464 112086 24466 112138
rect 24466 112086 24518 112138
rect 24518 112086 24520 112138
rect 24464 112084 24520 112086
rect 24568 112138 24624 112140
rect 24568 112086 24570 112138
rect 24570 112086 24622 112138
rect 24622 112086 24624 112138
rect 24568 112084 24624 112086
rect 24672 112138 24728 112140
rect 24672 112086 24674 112138
rect 24674 112086 24726 112138
rect 24726 112086 24728 112138
rect 24672 112084 24728 112086
rect 24668 111692 24724 111748
rect 25116 111916 25172 111972
rect 24780 110796 24836 110852
rect 24892 111356 24948 111412
rect 24556 110684 24612 110740
rect 24464 110570 24520 110572
rect 24464 110518 24466 110570
rect 24466 110518 24518 110570
rect 24518 110518 24520 110570
rect 24464 110516 24520 110518
rect 24568 110570 24624 110572
rect 24568 110518 24570 110570
rect 24570 110518 24622 110570
rect 24622 110518 24624 110570
rect 24568 110516 24624 110518
rect 24672 110570 24728 110572
rect 24672 110518 24674 110570
rect 24674 110518 24726 110570
rect 24726 110518 24728 110570
rect 24672 110516 24728 110518
rect 25004 111132 25060 111188
rect 25116 111020 25172 111076
rect 25452 114044 25508 114100
rect 25564 112700 25620 112756
rect 25676 113820 25732 113876
rect 25340 112588 25396 112644
rect 25788 113596 25844 113652
rect 28476 114716 28532 114772
rect 26012 113484 26068 113540
rect 26124 114492 26180 114548
rect 26796 114380 26852 114436
rect 28364 114268 28420 114324
rect 27692 113932 27748 113988
rect 25340 112028 25396 112084
rect 25564 111858 25620 111860
rect 25564 111806 25566 111858
rect 25566 111806 25618 111858
rect 25618 111806 25620 111858
rect 25564 111804 25620 111806
rect 25676 111244 25732 111300
rect 25564 111020 25620 111076
rect 25340 110572 25396 110628
rect 24668 110178 24724 110180
rect 24668 110126 24670 110178
rect 24670 110126 24722 110178
rect 24722 110126 24724 110178
rect 24668 110124 24724 110126
rect 24464 109002 24520 109004
rect 24464 108950 24466 109002
rect 24466 108950 24518 109002
rect 24518 108950 24520 109002
rect 24464 108948 24520 108950
rect 24568 109002 24624 109004
rect 24568 108950 24570 109002
rect 24570 108950 24622 109002
rect 24622 108950 24624 109002
rect 24568 108948 24624 108950
rect 24672 109002 24728 109004
rect 24672 108950 24674 109002
rect 24674 108950 24726 109002
rect 24726 108950 24728 109002
rect 24672 108948 24728 108950
rect 25228 110290 25284 110292
rect 25228 110238 25230 110290
rect 25230 110238 25282 110290
rect 25282 110238 25284 110290
rect 25228 110236 25284 110238
rect 25340 110012 25396 110068
rect 25228 109004 25284 109060
rect 25116 108498 25172 108500
rect 25116 108446 25118 108498
rect 25118 108446 25170 108498
rect 25170 108446 25172 108498
rect 25116 108444 25172 108446
rect 25116 107938 25172 107940
rect 25116 107886 25118 107938
rect 25118 107886 25170 107938
rect 25170 107886 25172 107938
rect 25116 107884 25172 107886
rect 24464 107434 24520 107436
rect 24464 107382 24466 107434
rect 24466 107382 24518 107434
rect 24518 107382 24520 107434
rect 24464 107380 24520 107382
rect 24568 107434 24624 107436
rect 24568 107382 24570 107434
rect 24570 107382 24622 107434
rect 24622 107382 24624 107434
rect 24568 107380 24624 107382
rect 24672 107434 24728 107436
rect 24672 107382 24674 107434
rect 24674 107382 24726 107434
rect 24726 107382 24728 107434
rect 24672 107380 24728 107382
rect 25116 106876 25172 106932
rect 24220 105756 24276 105812
rect 24464 105866 24520 105868
rect 24464 105814 24466 105866
rect 24466 105814 24518 105866
rect 24518 105814 24520 105866
rect 24464 105812 24520 105814
rect 24568 105866 24624 105868
rect 24568 105814 24570 105866
rect 24570 105814 24622 105866
rect 24622 105814 24624 105866
rect 24568 105812 24624 105814
rect 24672 105866 24728 105868
rect 24672 105814 24674 105866
rect 24674 105814 24726 105866
rect 24726 105814 24728 105866
rect 24672 105812 24728 105814
rect 23804 105082 23860 105084
rect 23804 105030 23806 105082
rect 23806 105030 23858 105082
rect 23858 105030 23860 105082
rect 23804 105028 23860 105030
rect 23908 105082 23964 105084
rect 23908 105030 23910 105082
rect 23910 105030 23962 105082
rect 23962 105030 23964 105082
rect 23908 105028 23964 105030
rect 24012 105082 24068 105084
rect 24012 105030 24014 105082
rect 24014 105030 24066 105082
rect 24066 105030 24068 105082
rect 24012 105028 24068 105030
rect 24464 104298 24520 104300
rect 24464 104246 24466 104298
rect 24466 104246 24518 104298
rect 24518 104246 24520 104298
rect 24464 104244 24520 104246
rect 24568 104298 24624 104300
rect 24568 104246 24570 104298
rect 24570 104246 24622 104298
rect 24622 104246 24624 104298
rect 24568 104244 24624 104246
rect 24672 104298 24728 104300
rect 24672 104246 24674 104298
rect 24674 104246 24726 104298
rect 24726 104246 24728 104298
rect 24672 104244 24728 104246
rect 23804 103514 23860 103516
rect 23804 103462 23806 103514
rect 23806 103462 23858 103514
rect 23858 103462 23860 103514
rect 23804 103460 23860 103462
rect 23908 103514 23964 103516
rect 23908 103462 23910 103514
rect 23910 103462 23962 103514
rect 23962 103462 23964 103514
rect 23908 103460 23964 103462
rect 24012 103514 24068 103516
rect 24012 103462 24014 103514
rect 24014 103462 24066 103514
rect 24066 103462 24068 103514
rect 24012 103460 24068 103462
rect 24464 102730 24520 102732
rect 24464 102678 24466 102730
rect 24466 102678 24518 102730
rect 24518 102678 24520 102730
rect 24464 102676 24520 102678
rect 24568 102730 24624 102732
rect 24568 102678 24570 102730
rect 24570 102678 24622 102730
rect 24622 102678 24624 102730
rect 24568 102676 24624 102678
rect 24672 102730 24728 102732
rect 24672 102678 24674 102730
rect 24674 102678 24726 102730
rect 24726 102678 24728 102730
rect 24672 102676 24728 102678
rect 23804 101946 23860 101948
rect 23804 101894 23806 101946
rect 23806 101894 23858 101946
rect 23858 101894 23860 101946
rect 23804 101892 23860 101894
rect 23908 101946 23964 101948
rect 23908 101894 23910 101946
rect 23910 101894 23962 101946
rect 23962 101894 23964 101946
rect 23908 101892 23964 101894
rect 24012 101946 24068 101948
rect 24012 101894 24014 101946
rect 24014 101894 24066 101946
rect 24066 101894 24068 101946
rect 24012 101892 24068 101894
rect 24464 101162 24520 101164
rect 24464 101110 24466 101162
rect 24466 101110 24518 101162
rect 24518 101110 24520 101162
rect 24464 101108 24520 101110
rect 24568 101162 24624 101164
rect 24568 101110 24570 101162
rect 24570 101110 24622 101162
rect 24622 101110 24624 101162
rect 24568 101108 24624 101110
rect 24672 101162 24728 101164
rect 24672 101110 24674 101162
rect 24674 101110 24726 101162
rect 24726 101110 24728 101162
rect 24672 101108 24728 101110
rect 23804 100378 23860 100380
rect 23804 100326 23806 100378
rect 23806 100326 23858 100378
rect 23858 100326 23860 100378
rect 23804 100324 23860 100326
rect 23908 100378 23964 100380
rect 23908 100326 23910 100378
rect 23910 100326 23962 100378
rect 23962 100326 23964 100378
rect 23908 100324 23964 100326
rect 24012 100378 24068 100380
rect 24012 100326 24014 100378
rect 24014 100326 24066 100378
rect 24066 100326 24068 100378
rect 24012 100324 24068 100326
rect 24464 99594 24520 99596
rect 24464 99542 24466 99594
rect 24466 99542 24518 99594
rect 24518 99542 24520 99594
rect 24464 99540 24520 99542
rect 24568 99594 24624 99596
rect 24568 99542 24570 99594
rect 24570 99542 24622 99594
rect 24622 99542 24624 99594
rect 24568 99540 24624 99542
rect 24672 99594 24728 99596
rect 24672 99542 24674 99594
rect 24674 99542 24726 99594
rect 24726 99542 24728 99594
rect 24672 99540 24728 99542
rect 23804 98810 23860 98812
rect 23804 98758 23806 98810
rect 23806 98758 23858 98810
rect 23858 98758 23860 98810
rect 23804 98756 23860 98758
rect 23908 98810 23964 98812
rect 23908 98758 23910 98810
rect 23910 98758 23962 98810
rect 23962 98758 23964 98810
rect 23908 98756 23964 98758
rect 24012 98810 24068 98812
rect 24012 98758 24014 98810
rect 24014 98758 24066 98810
rect 24066 98758 24068 98810
rect 24012 98756 24068 98758
rect 24464 98026 24520 98028
rect 24464 97974 24466 98026
rect 24466 97974 24518 98026
rect 24518 97974 24520 98026
rect 24464 97972 24520 97974
rect 24568 98026 24624 98028
rect 24568 97974 24570 98026
rect 24570 97974 24622 98026
rect 24622 97974 24624 98026
rect 24568 97972 24624 97974
rect 24672 98026 24728 98028
rect 24672 97974 24674 98026
rect 24674 97974 24726 98026
rect 24726 97974 24728 98026
rect 24672 97972 24728 97974
rect 22428 94220 22484 94276
rect 21980 91644 22036 91700
rect 21532 90860 21588 90916
rect 21532 90636 21588 90692
rect 21420 88172 21476 88228
rect 21308 87276 21364 87332
rect 20748 87218 20804 87220
rect 20748 87166 20750 87218
rect 20750 87166 20802 87218
rect 20802 87166 20804 87218
rect 20748 87164 20804 87166
rect 20860 86380 20916 86436
rect 20860 86156 20916 86212
rect 20748 85762 20804 85764
rect 20748 85710 20750 85762
rect 20750 85710 20802 85762
rect 20802 85710 20804 85762
rect 20748 85708 20804 85710
rect 21308 85708 21364 85764
rect 20972 85036 21028 85092
rect 21084 84252 21140 84308
rect 21196 84924 21252 84980
rect 20412 81900 20468 81956
rect 20524 82124 20580 82180
rect 20300 80556 20356 80612
rect 20188 78876 20244 78932
rect 21196 82124 21252 82180
rect 21196 81900 21252 81956
rect 20860 81282 20916 81284
rect 20860 81230 20862 81282
rect 20862 81230 20914 81282
rect 20914 81230 20916 81282
rect 20860 81228 20916 81230
rect 21196 81116 21252 81172
rect 21532 85820 21588 85876
rect 21420 84924 21476 84980
rect 21308 81004 21364 81060
rect 21420 84700 21476 84756
rect 22092 91084 22148 91140
rect 21868 90860 21924 90916
rect 21756 90748 21812 90804
rect 21756 87276 21812 87332
rect 22204 90860 22260 90916
rect 22316 92876 22372 92932
rect 22764 94220 22820 94276
rect 22652 92146 22708 92148
rect 22652 92094 22654 92146
rect 22654 92094 22706 92146
rect 22706 92094 22708 92146
rect 22652 92092 22708 92094
rect 22764 91138 22820 91140
rect 22764 91086 22766 91138
rect 22766 91086 22818 91138
rect 22818 91086 22820 91138
rect 22764 91084 22820 91086
rect 22204 90524 22260 90580
rect 21980 88956 22036 89012
rect 21868 86828 21924 86884
rect 21868 86156 21924 86212
rect 21644 84700 21700 84756
rect 21644 84476 21700 84532
rect 21532 81004 21588 81060
rect 20524 78764 20580 78820
rect 20300 78540 20356 78596
rect 20188 77644 20244 77700
rect 20188 75404 20244 75460
rect 20188 74060 20244 74116
rect 20076 72546 20132 72548
rect 20076 72494 20078 72546
rect 20078 72494 20130 72546
rect 20130 72494 20132 72546
rect 20076 72492 20132 72494
rect 19964 71986 20020 71988
rect 19964 71934 19966 71986
rect 19966 71934 20018 71986
rect 20018 71934 20020 71986
rect 19964 71932 20020 71934
rect 19852 70476 19908 70532
rect 20748 79548 20804 79604
rect 20972 79602 21028 79604
rect 20972 79550 20974 79602
rect 20974 79550 21026 79602
rect 21026 79550 21028 79602
rect 20972 79548 21028 79550
rect 21084 78540 21140 78596
rect 20412 77308 20468 77364
rect 21420 80610 21476 80612
rect 21420 80558 21422 80610
rect 21422 80558 21474 80610
rect 21474 80558 21476 80610
rect 21420 80556 21476 80558
rect 20748 77532 20804 77588
rect 20748 77308 20804 77364
rect 20636 77250 20692 77252
rect 20636 77198 20638 77250
rect 20638 77198 20690 77250
rect 20690 77198 20692 77250
rect 20636 77196 20692 77198
rect 20524 76300 20580 76356
rect 20412 75794 20468 75796
rect 20412 75742 20414 75794
rect 20414 75742 20466 75794
rect 20466 75742 20468 75794
rect 20412 75740 20468 75742
rect 20748 76242 20804 76244
rect 20748 76190 20750 76242
rect 20750 76190 20802 76242
rect 20802 76190 20804 76242
rect 20748 76188 20804 76190
rect 20524 74956 20580 75012
rect 20188 70140 20244 70196
rect 20076 69970 20132 69972
rect 20076 69918 20078 69970
rect 20078 69918 20130 69970
rect 20130 69918 20132 69970
rect 20076 69916 20132 69918
rect 19404 67788 19460 67844
rect 19292 67116 19348 67172
rect 19964 68738 20020 68740
rect 19964 68686 19966 68738
rect 19966 68686 20018 68738
rect 20018 68686 20020 68738
rect 19964 68684 20020 68686
rect 20076 68626 20132 68628
rect 20076 68574 20078 68626
rect 20078 68574 20130 68626
rect 20130 68574 20132 68626
rect 20076 68572 20132 68574
rect 20188 68236 20244 68292
rect 19964 67452 20020 67508
rect 19740 67340 19796 67396
rect 19628 67228 19684 67284
rect 19068 65996 19124 66052
rect 18732 63810 18788 63812
rect 18732 63758 18734 63810
rect 18734 63758 18786 63810
rect 18786 63758 18788 63810
rect 18732 63756 18788 63758
rect 18508 60732 18564 60788
rect 18732 61404 18788 61460
rect 18732 60620 18788 60676
rect 18284 59836 18340 59892
rect 18732 59948 18788 60004
rect 18732 59500 18788 59556
rect 19068 64818 19124 64820
rect 19068 64766 19070 64818
rect 19070 64766 19122 64818
rect 19122 64766 19124 64818
rect 19068 64764 19124 64766
rect 19180 63644 19236 63700
rect 18956 62188 19012 62244
rect 19068 62076 19124 62132
rect 19068 61740 19124 61796
rect 19068 61068 19124 61124
rect 18956 60002 19012 60004
rect 18956 59950 18958 60002
rect 18958 59950 19010 60002
rect 19010 59950 19012 60002
rect 18956 59948 19012 59950
rect 18956 59330 19012 59332
rect 18956 59278 18958 59330
rect 18958 59278 19010 59330
rect 19010 59278 19012 59330
rect 18956 59276 19012 59278
rect 19292 60786 19348 60788
rect 19292 60734 19294 60786
rect 19294 60734 19346 60786
rect 19346 60734 19348 60786
rect 19292 60732 19348 60734
rect 19292 60172 19348 60228
rect 19180 59500 19236 59556
rect 18732 54796 18788 54852
rect 18172 54124 18228 54180
rect 18396 50482 18452 50484
rect 18396 50430 18398 50482
rect 18398 50430 18450 50482
rect 18450 50430 18452 50482
rect 18396 50428 18452 50430
rect 18060 45052 18116 45108
rect 17612 43596 17668 43652
rect 17836 43372 17892 43428
rect 18172 43932 18228 43988
rect 18396 50092 18452 50148
rect 18956 48188 19012 48244
rect 18620 46844 18676 46900
rect 18732 47458 18788 47460
rect 18732 47406 18734 47458
rect 18734 47406 18786 47458
rect 18786 47406 18788 47458
rect 18732 47404 18788 47406
rect 17612 41916 17668 41972
rect 17052 40908 17108 40964
rect 16716 40460 16772 40516
rect 17164 40460 17220 40516
rect 16940 40402 16996 40404
rect 16940 40350 16942 40402
rect 16942 40350 16994 40402
rect 16994 40350 16996 40402
rect 16940 40348 16996 40350
rect 16156 37324 16212 37380
rect 16268 38332 16324 38388
rect 15932 35474 15988 35476
rect 15932 35422 15934 35474
rect 15934 35422 15986 35474
rect 15986 35422 15988 35474
rect 15932 35420 15988 35422
rect 16044 35308 16100 35364
rect 15932 35084 15988 35140
rect 15708 33404 15764 33460
rect 15148 31218 15204 31220
rect 15148 31166 15150 31218
rect 15150 31166 15202 31218
rect 15202 31166 15204 31218
rect 15148 31164 15204 31166
rect 15036 30268 15092 30324
rect 14700 28588 14756 28644
rect 14700 26908 14756 26964
rect 14476 26290 14532 26292
rect 14476 26238 14478 26290
rect 14478 26238 14530 26290
rect 14530 26238 14532 26290
rect 14476 26236 14532 26238
rect 14476 24668 14532 24724
rect 14924 28812 14980 28868
rect 15372 31666 15428 31668
rect 15372 31614 15374 31666
rect 15374 31614 15426 31666
rect 15426 31614 15428 31666
rect 15372 31612 15428 31614
rect 15260 27580 15316 27636
rect 15596 32284 15652 32340
rect 15148 27186 15204 27188
rect 15148 27134 15150 27186
rect 15150 27134 15202 27186
rect 15202 27134 15204 27186
rect 15148 27132 15204 27134
rect 15260 27074 15316 27076
rect 15260 27022 15262 27074
rect 15262 27022 15314 27074
rect 15314 27022 15316 27074
rect 15260 27020 15316 27022
rect 15036 26066 15092 26068
rect 15036 26014 15038 26066
rect 15038 26014 15090 26066
rect 15090 26014 15092 26066
rect 15036 26012 15092 26014
rect 14924 25788 14980 25844
rect 14924 25506 14980 25508
rect 14924 25454 14926 25506
rect 14926 25454 14978 25506
rect 14978 25454 14980 25506
rect 14924 25452 14980 25454
rect 14924 25228 14980 25284
rect 14364 23324 14420 23380
rect 13916 23100 13972 23156
rect 13916 22764 13972 22820
rect 14588 23154 14644 23156
rect 14588 23102 14590 23154
rect 14590 23102 14642 23154
rect 14642 23102 14644 23154
rect 14588 23100 14644 23102
rect 14364 23042 14420 23044
rect 14364 22990 14366 23042
rect 14366 22990 14418 23042
rect 14418 22990 14420 23042
rect 14364 22988 14420 22990
rect 13804 21756 13860 21812
rect 14140 21532 14196 21588
rect 13804 21196 13860 21252
rect 13916 21084 13972 21140
rect 13692 19906 13748 19908
rect 13692 19854 13694 19906
rect 13694 19854 13746 19906
rect 13746 19854 13748 19906
rect 13692 19852 13748 19854
rect 13580 19404 13636 19460
rect 13580 19234 13636 19236
rect 13580 19182 13582 19234
rect 13582 19182 13634 19234
rect 13634 19182 13636 19234
rect 13580 19180 13636 19182
rect 13468 18338 13524 18340
rect 13468 18286 13470 18338
rect 13470 18286 13522 18338
rect 13522 18286 13524 18338
rect 13468 18284 13524 18286
rect 14364 22092 14420 22148
rect 14812 24050 14868 24052
rect 14812 23998 14814 24050
rect 14814 23998 14866 24050
rect 14866 23998 14868 24050
rect 14812 23996 14868 23998
rect 14924 23436 14980 23492
rect 15260 26236 15316 26292
rect 15708 31500 15764 31556
rect 16380 35698 16436 35700
rect 16380 35646 16382 35698
rect 16382 35646 16434 35698
rect 16434 35646 16436 35698
rect 16380 35644 16436 35646
rect 16716 37212 16772 37268
rect 16940 35980 16996 36036
rect 17388 40236 17444 40292
rect 17276 37266 17332 37268
rect 17276 37214 17278 37266
rect 17278 37214 17330 37266
rect 17330 37214 17332 37266
rect 17276 37212 17332 37214
rect 17052 35756 17108 35812
rect 17276 35980 17332 36036
rect 16828 35644 16884 35700
rect 17164 35698 17220 35700
rect 17164 35646 17166 35698
rect 17166 35646 17218 35698
rect 17218 35646 17220 35698
rect 17164 35644 17220 35646
rect 16828 35420 16884 35476
rect 16604 34748 16660 34804
rect 16828 34690 16884 34692
rect 16828 34638 16830 34690
rect 16830 34638 16882 34690
rect 16882 34638 16884 34690
rect 16828 34636 16884 34638
rect 16716 34412 16772 34468
rect 16828 34242 16884 34244
rect 16828 34190 16830 34242
rect 16830 34190 16882 34242
rect 16882 34190 16884 34242
rect 16828 34188 16884 34190
rect 16492 34076 16548 34132
rect 16828 33234 16884 33236
rect 16828 33182 16830 33234
rect 16830 33182 16882 33234
rect 16882 33182 16884 33234
rect 16828 33180 16884 33182
rect 16716 33068 16772 33124
rect 17500 39900 17556 39956
rect 17500 38668 17556 38724
rect 17500 36764 17556 36820
rect 17836 41916 17892 41972
rect 17836 37996 17892 38052
rect 18620 43372 18676 43428
rect 18172 40402 18228 40404
rect 18172 40350 18174 40402
rect 18174 40350 18226 40402
rect 18226 40350 18228 40402
rect 18172 40348 18228 40350
rect 18844 43932 18900 43988
rect 18732 41916 18788 41972
rect 18844 40796 18900 40852
rect 19964 66444 20020 66500
rect 19628 63980 19684 64036
rect 19628 62860 19684 62916
rect 20636 73388 20692 73444
rect 20412 67900 20468 67956
rect 21196 77532 21252 77588
rect 21420 77308 21476 77364
rect 21980 85596 22036 85652
rect 22092 84306 22148 84308
rect 22092 84254 22094 84306
rect 22094 84254 22146 84306
rect 22146 84254 22148 84306
rect 22092 84252 22148 84254
rect 21980 81228 22036 81284
rect 21868 80668 21924 80724
rect 21980 80444 22036 80500
rect 21084 76188 21140 76244
rect 21084 74060 21140 74116
rect 20972 73106 21028 73108
rect 20972 73054 20974 73106
rect 20974 73054 21026 73106
rect 21026 73054 21028 73106
rect 20972 73052 21028 73054
rect 20860 72546 20916 72548
rect 20860 72494 20862 72546
rect 20862 72494 20914 72546
rect 20914 72494 20916 72546
rect 20860 72492 20916 72494
rect 20412 67004 20468 67060
rect 20860 71596 20916 71652
rect 20636 70028 20692 70084
rect 20636 68348 20692 68404
rect 20748 68012 20804 68068
rect 20636 67900 20692 67956
rect 20076 63532 20132 63588
rect 20748 67842 20804 67844
rect 20748 67790 20750 67842
rect 20750 67790 20802 67842
rect 20802 67790 20804 67842
rect 20748 67788 20804 67790
rect 20748 67116 20804 67172
rect 19852 62860 19908 62916
rect 19404 58546 19460 58548
rect 19404 58494 19406 58546
rect 19406 58494 19458 58546
rect 19458 58494 19460 58546
rect 19404 58492 19460 58494
rect 19292 53788 19348 53844
rect 19516 57260 19572 57316
rect 19292 51996 19348 52052
rect 19516 49980 19572 50036
rect 19404 47740 19460 47796
rect 19740 49138 19796 49140
rect 19740 49086 19742 49138
rect 19742 49086 19794 49138
rect 19794 49086 19796 49138
rect 19740 49084 19796 49086
rect 19740 47292 19796 47348
rect 19516 44492 19572 44548
rect 19964 62636 20020 62692
rect 20748 63756 20804 63812
rect 20188 62188 20244 62244
rect 20188 59500 20244 59556
rect 19964 59276 20020 59332
rect 20636 61964 20692 62020
rect 20524 61628 20580 61684
rect 20636 61740 20692 61796
rect 20412 60844 20468 60900
rect 20300 53900 20356 53956
rect 20412 60620 20468 60676
rect 20300 51884 20356 51940
rect 20188 48972 20244 49028
rect 20188 46956 20244 47012
rect 20076 45836 20132 45892
rect 19740 45164 19796 45220
rect 19404 44210 19460 44212
rect 19404 44158 19406 44210
rect 19406 44158 19458 44210
rect 19458 44158 19460 44210
rect 19404 44156 19460 44158
rect 19852 44546 19908 44548
rect 19852 44494 19854 44546
rect 19854 44494 19906 44546
rect 19906 44494 19908 44546
rect 19852 44492 19908 44494
rect 19740 44044 19796 44100
rect 19292 41858 19348 41860
rect 19292 41806 19294 41858
rect 19294 41806 19346 41858
rect 19346 41806 19348 41858
rect 19292 41804 19348 41806
rect 20188 42700 20244 42756
rect 19740 42028 19796 42084
rect 19628 41804 19684 41860
rect 18956 40460 19012 40516
rect 18620 40236 18676 40292
rect 18060 37548 18116 37604
rect 18396 38220 18452 38276
rect 18396 37884 18452 37940
rect 17948 37212 18004 37268
rect 18060 36764 18116 36820
rect 17948 36706 18004 36708
rect 17948 36654 17950 36706
rect 17950 36654 18002 36706
rect 18002 36654 18004 36706
rect 17948 36652 18004 36654
rect 17724 35868 17780 35924
rect 17612 35756 17668 35812
rect 17388 35196 17444 35252
rect 17500 35420 17556 35476
rect 17276 34914 17332 34916
rect 17276 34862 17278 34914
rect 17278 34862 17330 34914
rect 17330 34862 17332 34914
rect 17276 34860 17332 34862
rect 17164 34076 17220 34132
rect 16380 32508 16436 32564
rect 16604 32562 16660 32564
rect 16604 32510 16606 32562
rect 16606 32510 16658 32562
rect 16658 32510 16660 32562
rect 16604 32508 16660 32510
rect 15932 31612 15988 31668
rect 16156 31778 16212 31780
rect 16156 31726 16158 31778
rect 16158 31726 16210 31778
rect 16210 31726 16212 31778
rect 16156 31724 16212 31726
rect 16044 31276 16100 31332
rect 16156 31388 16212 31444
rect 16044 30882 16100 30884
rect 16044 30830 16046 30882
rect 16046 30830 16098 30882
rect 16098 30830 16100 30882
rect 16044 30828 16100 30830
rect 15932 30716 15988 30772
rect 16380 30716 16436 30772
rect 16268 30434 16324 30436
rect 16268 30382 16270 30434
rect 16270 30382 16322 30434
rect 16322 30382 16324 30434
rect 16268 30380 16324 30382
rect 16044 30322 16100 30324
rect 16044 30270 16046 30322
rect 16046 30270 16098 30322
rect 16098 30270 16100 30322
rect 16044 30268 16100 30270
rect 15708 28812 15764 28868
rect 15708 26908 15764 26964
rect 15820 26236 15876 26292
rect 15820 26012 15876 26068
rect 15596 25788 15652 25844
rect 15484 25564 15540 25620
rect 15708 25506 15764 25508
rect 15708 25454 15710 25506
rect 15710 25454 15762 25506
rect 15762 25454 15764 25506
rect 15708 25452 15764 25454
rect 16156 28364 16212 28420
rect 16156 27580 16212 27636
rect 16156 26796 16212 26852
rect 16268 27020 16324 27076
rect 16604 30380 16660 30436
rect 17836 35756 17892 35812
rect 17724 35084 17780 35140
rect 17948 35308 18004 35364
rect 17836 35026 17892 35028
rect 17836 34974 17838 35026
rect 17838 34974 17890 35026
rect 17890 34974 17892 35026
rect 17836 34972 17892 34974
rect 17612 34130 17668 34132
rect 17612 34078 17614 34130
rect 17614 34078 17666 34130
rect 17666 34078 17668 34130
rect 17612 34076 17668 34078
rect 17836 34076 17892 34132
rect 18060 34748 18116 34804
rect 18284 35980 18340 36036
rect 18172 34076 18228 34132
rect 16828 29538 16884 29540
rect 16828 29486 16830 29538
rect 16830 29486 16882 29538
rect 16882 29486 16884 29538
rect 16828 29484 16884 29486
rect 17276 32562 17332 32564
rect 17276 32510 17278 32562
rect 17278 32510 17330 32562
rect 17330 32510 17332 32562
rect 17276 32508 17332 32510
rect 17724 33292 17780 33348
rect 17500 33180 17556 33236
rect 17500 32844 17556 32900
rect 17052 31778 17108 31780
rect 17052 31726 17054 31778
rect 17054 31726 17106 31778
rect 17106 31726 17108 31778
rect 17052 31724 17108 31726
rect 17052 31554 17108 31556
rect 17052 31502 17054 31554
rect 17054 31502 17106 31554
rect 17106 31502 17108 31554
rect 17052 31500 17108 31502
rect 17164 31106 17220 31108
rect 17164 31054 17166 31106
rect 17166 31054 17218 31106
rect 17218 31054 17220 31106
rect 17164 31052 17220 31054
rect 16940 29372 16996 29428
rect 17052 30994 17108 30996
rect 17052 30942 17054 30994
rect 17054 30942 17106 30994
rect 17106 30942 17108 30994
rect 17052 30940 17108 30942
rect 17724 33068 17780 33124
rect 17052 30322 17108 30324
rect 17052 30270 17054 30322
rect 17054 30270 17106 30322
rect 17106 30270 17108 30322
rect 17052 30268 17108 30270
rect 17276 30210 17332 30212
rect 17276 30158 17278 30210
rect 17278 30158 17330 30210
rect 17330 30158 17332 30210
rect 17276 30156 17332 30158
rect 17276 29932 17332 29988
rect 17052 27244 17108 27300
rect 16940 27186 16996 27188
rect 16940 27134 16942 27186
rect 16942 27134 16994 27186
rect 16994 27134 16996 27186
rect 16940 27132 16996 27134
rect 16828 27074 16884 27076
rect 16828 27022 16830 27074
rect 16830 27022 16882 27074
rect 16882 27022 16884 27074
rect 16828 27020 16884 27022
rect 16716 26684 16772 26740
rect 16380 26236 16436 26292
rect 17164 26290 17220 26292
rect 17164 26238 17166 26290
rect 17166 26238 17218 26290
rect 17218 26238 17220 26290
rect 17164 26236 17220 26238
rect 16604 26066 16660 26068
rect 16604 26014 16606 26066
rect 16606 26014 16658 26066
rect 16658 26014 16660 26066
rect 16604 26012 16660 26014
rect 15932 25228 15988 25284
rect 15372 23996 15428 24052
rect 17388 29596 17444 29652
rect 17500 30940 17556 30996
rect 17388 29372 17444 29428
rect 18060 33628 18116 33684
rect 18060 33180 18116 33236
rect 18396 35756 18452 35812
rect 18284 33628 18340 33684
rect 18396 35532 18452 35588
rect 18284 33458 18340 33460
rect 18284 33406 18286 33458
rect 18286 33406 18338 33458
rect 18338 33406 18340 33458
rect 18284 33404 18340 33406
rect 18172 32562 18228 32564
rect 18172 32510 18174 32562
rect 18174 32510 18226 32562
rect 18226 32510 18228 32562
rect 18172 32508 18228 32510
rect 17948 31724 18004 31780
rect 17612 29986 17668 29988
rect 17612 29934 17614 29986
rect 17614 29934 17666 29986
rect 17666 29934 17668 29986
rect 17612 29932 17668 29934
rect 17612 29426 17668 29428
rect 17612 29374 17614 29426
rect 17614 29374 17666 29426
rect 17666 29374 17668 29426
rect 17612 29372 17668 29374
rect 17388 27916 17444 27972
rect 17612 28700 17668 28756
rect 17836 30434 17892 30436
rect 17836 30382 17838 30434
rect 17838 30382 17890 30434
rect 17890 30382 17892 30434
rect 17836 30380 17892 30382
rect 17836 30210 17892 30212
rect 17836 30158 17838 30210
rect 17838 30158 17890 30210
rect 17890 30158 17892 30210
rect 17836 30156 17892 30158
rect 19404 40236 19460 40292
rect 19964 40348 20020 40404
rect 19180 36540 19236 36596
rect 18732 35308 18788 35364
rect 18620 34972 18676 35028
rect 18732 35084 18788 35140
rect 19404 37772 19460 37828
rect 19404 36258 19460 36260
rect 19404 36206 19406 36258
rect 19406 36206 19458 36258
rect 19458 36206 19460 36258
rect 19404 36204 19460 36206
rect 19292 35980 19348 36036
rect 19180 35644 19236 35700
rect 19068 34860 19124 34916
rect 18956 34636 19012 34692
rect 18844 34130 18900 34132
rect 18844 34078 18846 34130
rect 18846 34078 18898 34130
rect 18898 34078 18900 34130
rect 18844 34076 18900 34078
rect 18732 33740 18788 33796
rect 18508 33346 18564 33348
rect 18508 33294 18510 33346
rect 18510 33294 18562 33346
rect 18562 33294 18564 33346
rect 18508 33292 18564 33294
rect 18732 33068 18788 33124
rect 19068 34524 19124 34580
rect 19404 34972 19460 35028
rect 19068 33570 19124 33572
rect 19068 33518 19070 33570
rect 19070 33518 19122 33570
rect 19122 33518 19124 33570
rect 19068 33516 19124 33518
rect 19292 33516 19348 33572
rect 19180 33068 19236 33124
rect 18956 32956 19012 33012
rect 19852 38050 19908 38052
rect 19852 37998 19854 38050
rect 19854 37998 19906 38050
rect 19906 37998 19908 38050
rect 19852 37996 19908 37998
rect 19740 37100 19796 37156
rect 19628 36594 19684 36596
rect 19628 36542 19630 36594
rect 19630 36542 19682 36594
rect 19682 36542 19684 36594
rect 19628 36540 19684 36542
rect 20188 38332 20244 38388
rect 20636 59276 20692 59332
rect 21084 71762 21140 71764
rect 21084 71710 21086 71762
rect 21086 71710 21138 71762
rect 21138 71710 21140 71762
rect 21084 71708 21140 71710
rect 21532 76748 21588 76804
rect 21420 76412 21476 76468
rect 21308 76300 21364 76356
rect 22652 90354 22708 90356
rect 22652 90302 22654 90354
rect 22654 90302 22706 90354
rect 22706 90302 22708 90354
rect 22652 90300 22708 90302
rect 22876 89180 22932 89236
rect 23804 97242 23860 97244
rect 23804 97190 23806 97242
rect 23806 97190 23858 97242
rect 23858 97190 23860 97242
rect 23804 97188 23860 97190
rect 23908 97242 23964 97244
rect 23908 97190 23910 97242
rect 23910 97190 23962 97242
rect 23962 97190 23964 97242
rect 23908 97188 23964 97190
rect 24012 97242 24068 97244
rect 24012 97190 24014 97242
rect 24014 97190 24066 97242
rect 24066 97190 24068 97242
rect 24012 97188 24068 97190
rect 24464 96458 24520 96460
rect 24464 96406 24466 96458
rect 24466 96406 24518 96458
rect 24518 96406 24520 96458
rect 24464 96404 24520 96406
rect 24568 96458 24624 96460
rect 24568 96406 24570 96458
rect 24570 96406 24622 96458
rect 24622 96406 24624 96458
rect 24568 96404 24624 96406
rect 24672 96458 24728 96460
rect 24672 96406 24674 96458
rect 24674 96406 24726 96458
rect 24726 96406 24728 96458
rect 24672 96404 24728 96406
rect 23804 95674 23860 95676
rect 23804 95622 23806 95674
rect 23806 95622 23858 95674
rect 23858 95622 23860 95674
rect 23804 95620 23860 95622
rect 23908 95674 23964 95676
rect 23908 95622 23910 95674
rect 23910 95622 23962 95674
rect 23962 95622 23964 95674
rect 23908 95620 23964 95622
rect 24012 95674 24068 95676
rect 24012 95622 24014 95674
rect 24014 95622 24066 95674
rect 24066 95622 24068 95674
rect 24012 95620 24068 95622
rect 23324 95004 23380 95060
rect 24892 95004 24948 95060
rect 23772 94780 23828 94836
rect 24464 94890 24520 94892
rect 24464 94838 24466 94890
rect 24466 94838 24518 94890
rect 24518 94838 24520 94890
rect 24464 94836 24520 94838
rect 24568 94890 24624 94892
rect 24568 94838 24570 94890
rect 24570 94838 24622 94890
rect 24622 94838 24624 94890
rect 24568 94836 24624 94838
rect 24672 94890 24728 94892
rect 24672 94838 24674 94890
rect 24674 94838 24726 94890
rect 24726 94838 24728 94890
rect 24672 94836 24728 94838
rect 23660 94722 23716 94724
rect 23660 94670 23662 94722
rect 23662 94670 23714 94722
rect 23714 94670 23716 94722
rect 23660 94668 23716 94670
rect 23324 94610 23380 94612
rect 23324 94558 23326 94610
rect 23326 94558 23378 94610
rect 23378 94558 23380 94610
rect 23324 94556 23380 94558
rect 23804 94106 23860 94108
rect 23804 94054 23806 94106
rect 23806 94054 23858 94106
rect 23858 94054 23860 94106
rect 23804 94052 23860 94054
rect 23908 94106 23964 94108
rect 23908 94054 23910 94106
rect 23910 94054 23962 94106
rect 23962 94054 23964 94106
rect 23908 94052 23964 94054
rect 24012 94106 24068 94108
rect 24012 94054 24014 94106
rect 24014 94054 24066 94106
rect 24066 94054 24068 94106
rect 24012 94052 24068 94054
rect 24464 93322 24520 93324
rect 24464 93270 24466 93322
rect 24466 93270 24518 93322
rect 24518 93270 24520 93322
rect 24464 93268 24520 93270
rect 24568 93322 24624 93324
rect 24568 93270 24570 93322
rect 24570 93270 24622 93322
rect 24622 93270 24624 93322
rect 24568 93268 24624 93270
rect 24672 93322 24728 93324
rect 24672 93270 24674 93322
rect 24674 93270 24726 93322
rect 24726 93270 24728 93322
rect 24672 93268 24728 93270
rect 24668 93042 24724 93044
rect 24668 92990 24670 93042
rect 24670 92990 24722 93042
rect 24722 92990 24724 93042
rect 24668 92988 24724 92990
rect 23804 92538 23860 92540
rect 23804 92486 23806 92538
rect 23806 92486 23858 92538
rect 23858 92486 23860 92538
rect 23804 92484 23860 92486
rect 23908 92538 23964 92540
rect 23908 92486 23910 92538
rect 23910 92486 23962 92538
rect 23962 92486 23964 92538
rect 23908 92484 23964 92486
rect 24012 92538 24068 92540
rect 24012 92486 24014 92538
rect 24014 92486 24066 92538
rect 24066 92486 24068 92538
rect 24012 92484 24068 92486
rect 23804 90970 23860 90972
rect 23804 90918 23806 90970
rect 23806 90918 23858 90970
rect 23858 90918 23860 90970
rect 23804 90916 23860 90918
rect 23908 90970 23964 90972
rect 23908 90918 23910 90970
rect 23910 90918 23962 90970
rect 23962 90918 23964 90970
rect 23908 90916 23964 90918
rect 24012 90970 24068 90972
rect 24012 90918 24014 90970
rect 24014 90918 24066 90970
rect 24066 90918 24068 90970
rect 24012 90916 24068 90918
rect 23804 89402 23860 89404
rect 23804 89350 23806 89402
rect 23806 89350 23858 89402
rect 23858 89350 23860 89402
rect 23804 89348 23860 89350
rect 23908 89402 23964 89404
rect 23908 89350 23910 89402
rect 23910 89350 23962 89402
rect 23962 89350 23964 89402
rect 23908 89348 23964 89350
rect 24012 89402 24068 89404
rect 24012 89350 24014 89402
rect 24014 89350 24066 89402
rect 24066 89350 24068 89402
rect 24012 89348 24068 89350
rect 22316 87612 22372 87668
rect 22652 86604 22708 86660
rect 22540 86156 22596 86212
rect 22540 85820 22596 85876
rect 22540 85090 22596 85092
rect 22540 85038 22542 85090
rect 22542 85038 22594 85090
rect 22594 85038 22596 85090
rect 22540 85036 22596 85038
rect 22428 82572 22484 82628
rect 22876 87442 22932 87444
rect 22876 87390 22878 87442
rect 22878 87390 22930 87442
rect 22930 87390 22932 87442
rect 22876 87388 22932 87390
rect 23804 87834 23860 87836
rect 23804 87782 23806 87834
rect 23806 87782 23858 87834
rect 23858 87782 23860 87834
rect 23804 87780 23860 87782
rect 23908 87834 23964 87836
rect 23908 87782 23910 87834
rect 23910 87782 23962 87834
rect 23962 87782 23964 87834
rect 23908 87780 23964 87782
rect 24012 87834 24068 87836
rect 24012 87782 24014 87834
rect 24014 87782 24066 87834
rect 24066 87782 24068 87834
rect 24012 87780 24068 87782
rect 23884 87500 23940 87556
rect 23212 87388 23268 87444
rect 23548 86940 23604 86996
rect 23436 86770 23492 86772
rect 23436 86718 23438 86770
rect 23438 86718 23490 86770
rect 23490 86718 23492 86770
rect 23436 86716 23492 86718
rect 22876 86044 22932 86100
rect 22988 85932 23044 85988
rect 22764 85820 22820 85876
rect 23324 86098 23380 86100
rect 23324 86046 23326 86098
rect 23326 86046 23378 86098
rect 23378 86046 23380 86098
rect 23324 86044 23380 86046
rect 23548 86044 23604 86100
rect 23436 85932 23492 85988
rect 23548 85874 23604 85876
rect 23548 85822 23550 85874
rect 23550 85822 23602 85874
rect 23602 85822 23604 85874
rect 23548 85820 23604 85822
rect 23996 86380 24052 86436
rect 23804 86266 23860 86268
rect 23804 86214 23806 86266
rect 23806 86214 23858 86266
rect 23858 86214 23860 86266
rect 23804 86212 23860 86214
rect 23908 86266 23964 86268
rect 23908 86214 23910 86266
rect 23910 86214 23962 86266
rect 23962 86214 23964 86266
rect 23908 86212 23964 86214
rect 24012 86266 24068 86268
rect 24012 86214 24014 86266
rect 24014 86214 24066 86266
rect 24066 86214 24068 86266
rect 24012 86212 24068 86214
rect 24108 85762 24164 85764
rect 24108 85710 24110 85762
rect 24110 85710 24162 85762
rect 24162 85710 24164 85762
rect 24108 85708 24164 85710
rect 23884 85650 23940 85652
rect 23884 85598 23886 85650
rect 23886 85598 23938 85650
rect 23938 85598 23940 85650
rect 23884 85596 23940 85598
rect 23100 85314 23156 85316
rect 23100 85262 23102 85314
rect 23102 85262 23154 85314
rect 23154 85262 23156 85314
rect 23100 85260 23156 85262
rect 23548 85314 23604 85316
rect 23548 85262 23550 85314
rect 23550 85262 23602 85314
rect 23602 85262 23604 85314
rect 23548 85260 23604 85262
rect 23884 85202 23940 85204
rect 23884 85150 23886 85202
rect 23886 85150 23938 85202
rect 23938 85150 23940 85202
rect 23884 85148 23940 85150
rect 22540 82012 22596 82068
rect 23436 85036 23492 85092
rect 22876 82626 22932 82628
rect 22876 82574 22878 82626
rect 22878 82574 22930 82626
rect 22930 82574 22932 82626
rect 22876 82572 22932 82574
rect 22428 80946 22484 80948
rect 22428 80894 22430 80946
rect 22430 80894 22482 80946
rect 22482 80894 22484 80946
rect 22428 80892 22484 80894
rect 22204 80780 22260 80836
rect 22092 79772 22148 79828
rect 22204 80108 22260 80164
rect 22092 78876 22148 78932
rect 22092 77420 22148 77476
rect 21868 76354 21924 76356
rect 21868 76302 21870 76354
rect 21870 76302 21922 76354
rect 21922 76302 21924 76354
rect 21868 76300 21924 76302
rect 21420 74114 21476 74116
rect 21420 74062 21422 74114
rect 21422 74062 21474 74114
rect 21474 74062 21476 74114
rect 21420 74060 21476 74062
rect 21756 75794 21812 75796
rect 21756 75742 21758 75794
rect 21758 75742 21810 75794
rect 21810 75742 21812 75794
rect 21756 75740 21812 75742
rect 22428 79772 22484 79828
rect 22316 79602 22372 79604
rect 22316 79550 22318 79602
rect 22318 79550 22370 79602
rect 22370 79550 22372 79602
rect 22316 79548 22372 79550
rect 22316 78818 22372 78820
rect 22316 78766 22318 78818
rect 22318 78766 22370 78818
rect 22370 78766 22372 78818
rect 22316 78764 22372 78766
rect 22316 76466 22372 76468
rect 22316 76414 22318 76466
rect 22318 76414 22370 76466
rect 22370 76414 22372 76466
rect 22316 76412 22372 76414
rect 22428 74284 22484 74340
rect 21308 72604 21364 72660
rect 21532 73052 21588 73108
rect 21196 71596 21252 71652
rect 21196 71372 21252 71428
rect 21084 69356 21140 69412
rect 21420 71650 21476 71652
rect 21420 71598 21422 71650
rect 21422 71598 21474 71650
rect 21474 71598 21476 71650
rect 21420 71596 21476 71598
rect 20972 68796 21028 68852
rect 21084 68908 21140 68964
rect 21308 68908 21364 68964
rect 20972 68236 21028 68292
rect 21420 68348 21476 68404
rect 21308 67900 21364 67956
rect 21196 67564 21252 67620
rect 21084 67170 21140 67172
rect 21084 67118 21086 67170
rect 21086 67118 21138 67170
rect 21138 67118 21140 67170
rect 21084 67116 21140 67118
rect 21196 67228 21252 67284
rect 20972 66444 21028 66500
rect 20972 64034 21028 64036
rect 20972 63982 20974 64034
rect 20974 63982 21026 64034
rect 21026 63982 21028 64034
rect 20972 63980 21028 63982
rect 20972 63756 21028 63812
rect 21644 69916 21700 69972
rect 21756 69804 21812 69860
rect 21756 68796 21812 68852
rect 21868 68012 21924 68068
rect 21308 65100 21364 65156
rect 21868 67452 21924 67508
rect 21084 62524 21140 62580
rect 21308 63420 21364 63476
rect 21420 63084 21476 63140
rect 21420 62636 21476 62692
rect 20972 61068 21028 61124
rect 21196 62076 21252 62132
rect 20972 60786 21028 60788
rect 20972 60734 20974 60786
rect 20974 60734 21026 60786
rect 21026 60734 21028 60786
rect 20972 60732 21028 60734
rect 20860 58492 20916 58548
rect 21644 62412 21700 62468
rect 21756 62524 21812 62580
rect 21644 62242 21700 62244
rect 21644 62190 21646 62242
rect 21646 62190 21698 62242
rect 21698 62190 21700 62242
rect 21644 62188 21700 62190
rect 22652 80780 22708 80836
rect 23212 81842 23268 81844
rect 23212 81790 23214 81842
rect 23214 81790 23266 81842
rect 23266 81790 23268 81842
rect 23212 81788 23268 81790
rect 22764 80444 22820 80500
rect 22876 80668 22932 80724
rect 23804 84698 23860 84700
rect 23804 84646 23806 84698
rect 23806 84646 23858 84698
rect 23858 84646 23860 84698
rect 23804 84644 23860 84646
rect 23908 84698 23964 84700
rect 23908 84646 23910 84698
rect 23910 84646 23962 84698
rect 23962 84646 23964 84698
rect 23908 84644 23964 84646
rect 24012 84698 24068 84700
rect 24012 84646 24014 84698
rect 24014 84646 24066 84698
rect 24066 84646 24068 84698
rect 24012 84644 24068 84646
rect 22876 78876 22932 78932
rect 23660 84028 23716 84084
rect 23804 83130 23860 83132
rect 23804 83078 23806 83130
rect 23806 83078 23858 83130
rect 23858 83078 23860 83130
rect 23804 83076 23860 83078
rect 23908 83130 23964 83132
rect 23908 83078 23910 83130
rect 23910 83078 23962 83130
rect 23962 83078 23964 83130
rect 23908 83076 23964 83078
rect 24012 83130 24068 83132
rect 24012 83078 24014 83130
rect 24014 83078 24066 83130
rect 24066 83078 24068 83130
rect 24012 83076 24068 83078
rect 23804 81562 23860 81564
rect 23804 81510 23806 81562
rect 23806 81510 23858 81562
rect 23858 81510 23860 81562
rect 23804 81508 23860 81510
rect 23908 81562 23964 81564
rect 23908 81510 23910 81562
rect 23910 81510 23962 81562
rect 23962 81510 23964 81562
rect 23908 81508 23964 81510
rect 24012 81562 24068 81564
rect 24012 81510 24014 81562
rect 24014 81510 24066 81562
rect 24066 81510 24068 81562
rect 24012 81508 24068 81510
rect 23548 80386 23604 80388
rect 23548 80334 23550 80386
rect 23550 80334 23602 80386
rect 23602 80334 23604 80386
rect 23548 80332 23604 80334
rect 23804 79994 23860 79996
rect 23804 79942 23806 79994
rect 23806 79942 23858 79994
rect 23858 79942 23860 79994
rect 23804 79940 23860 79942
rect 23908 79994 23964 79996
rect 23908 79942 23910 79994
rect 23910 79942 23962 79994
rect 23962 79942 23964 79994
rect 23908 79940 23964 79942
rect 24012 79994 24068 79996
rect 24012 79942 24014 79994
rect 24014 79942 24066 79994
rect 24066 79942 24068 79994
rect 24012 79940 24068 79942
rect 23772 79602 23828 79604
rect 23772 79550 23774 79602
rect 23774 79550 23826 79602
rect 23826 79550 23828 79602
rect 23772 79548 23828 79550
rect 23804 78426 23860 78428
rect 23804 78374 23806 78426
rect 23806 78374 23858 78426
rect 23858 78374 23860 78426
rect 23804 78372 23860 78374
rect 23908 78426 23964 78428
rect 23908 78374 23910 78426
rect 23910 78374 23962 78426
rect 23962 78374 23964 78426
rect 23908 78372 23964 78374
rect 24012 78426 24068 78428
rect 24012 78374 24014 78426
rect 24014 78374 24066 78426
rect 24066 78374 24068 78426
rect 24012 78372 24068 78374
rect 23804 76858 23860 76860
rect 23804 76806 23806 76858
rect 23806 76806 23858 76858
rect 23858 76806 23860 76858
rect 23804 76804 23860 76806
rect 23908 76858 23964 76860
rect 23908 76806 23910 76858
rect 23910 76806 23962 76858
rect 23962 76806 23964 76858
rect 23908 76804 23964 76806
rect 24012 76858 24068 76860
rect 24012 76806 24014 76858
rect 24014 76806 24066 76858
rect 24066 76806 24068 76858
rect 24012 76804 24068 76806
rect 22988 75404 23044 75460
rect 22652 73276 22708 73332
rect 23324 74620 23380 74676
rect 22988 74338 23044 74340
rect 22988 74286 22990 74338
rect 22990 74286 23042 74338
rect 23042 74286 23044 74338
rect 22988 74284 23044 74286
rect 23436 74060 23492 74116
rect 22988 71820 23044 71876
rect 22428 69804 22484 69860
rect 22652 68348 22708 68404
rect 22428 68236 22484 68292
rect 22652 67340 22708 67396
rect 22092 63138 22148 63140
rect 22092 63086 22094 63138
rect 22094 63086 22146 63138
rect 22146 63086 22148 63138
rect 22092 63084 22148 63086
rect 21644 61964 21700 62020
rect 21756 60732 21812 60788
rect 21196 57148 21252 57204
rect 20972 51772 21028 51828
rect 20860 45612 20916 45668
rect 20412 44380 20468 44436
rect 20524 44492 20580 44548
rect 20412 41356 20468 41412
rect 20636 41970 20692 41972
rect 20636 41918 20638 41970
rect 20638 41918 20690 41970
rect 20690 41918 20692 41970
rect 20636 41916 20692 41918
rect 20636 40684 20692 40740
rect 20972 41970 21028 41972
rect 20972 41918 20974 41970
rect 20974 41918 21026 41970
rect 21026 41918 21028 41970
rect 20972 41916 21028 41918
rect 21868 60620 21924 60676
rect 21868 59948 21924 60004
rect 21644 59500 21700 59556
rect 21308 56028 21364 56084
rect 21420 53730 21476 53732
rect 21420 53678 21422 53730
rect 21422 53678 21474 53730
rect 21474 53678 21476 53730
rect 21420 53676 21476 53678
rect 21308 45666 21364 45668
rect 21308 45614 21310 45666
rect 21310 45614 21362 45666
rect 21362 45614 21364 45666
rect 21308 45612 21364 45614
rect 21532 43484 21588 43540
rect 22876 69410 22932 69412
rect 22876 69358 22878 69410
rect 22878 69358 22930 69410
rect 22930 69358 22932 69410
rect 22876 69356 22932 69358
rect 23100 68684 23156 68740
rect 22876 67676 22932 67732
rect 23212 68460 23268 68516
rect 23804 75290 23860 75292
rect 23804 75238 23806 75290
rect 23806 75238 23858 75290
rect 23858 75238 23860 75290
rect 23804 75236 23860 75238
rect 23908 75290 23964 75292
rect 23908 75238 23910 75290
rect 23910 75238 23962 75290
rect 23962 75238 23964 75290
rect 23908 75236 23964 75238
rect 24012 75290 24068 75292
rect 24012 75238 24014 75290
rect 24014 75238 24066 75290
rect 24066 75238 24068 75290
rect 24012 75236 24068 75238
rect 23804 73722 23860 73724
rect 23804 73670 23806 73722
rect 23806 73670 23858 73722
rect 23858 73670 23860 73722
rect 23804 73668 23860 73670
rect 23908 73722 23964 73724
rect 23908 73670 23910 73722
rect 23910 73670 23962 73722
rect 23962 73670 23964 73722
rect 23908 73668 23964 73670
rect 24012 73722 24068 73724
rect 24012 73670 24014 73722
rect 24014 73670 24066 73722
rect 24066 73670 24068 73722
rect 24012 73668 24068 73670
rect 23436 68460 23492 68516
rect 23804 72154 23860 72156
rect 23804 72102 23806 72154
rect 23806 72102 23858 72154
rect 23858 72102 23860 72154
rect 23804 72100 23860 72102
rect 23908 72154 23964 72156
rect 23908 72102 23910 72154
rect 23910 72102 23962 72154
rect 23962 72102 23964 72154
rect 23908 72100 23964 72102
rect 24012 72154 24068 72156
rect 24012 72102 24014 72154
rect 24014 72102 24066 72154
rect 24066 72102 24068 72154
rect 24012 72100 24068 72102
rect 23804 70586 23860 70588
rect 23804 70534 23806 70586
rect 23806 70534 23858 70586
rect 23858 70534 23860 70586
rect 23804 70532 23860 70534
rect 23908 70586 23964 70588
rect 23908 70534 23910 70586
rect 23910 70534 23962 70586
rect 23962 70534 23964 70586
rect 23908 70532 23964 70534
rect 24012 70586 24068 70588
rect 24012 70534 24014 70586
rect 24014 70534 24066 70586
rect 24066 70534 24068 70586
rect 24012 70532 24068 70534
rect 24464 91754 24520 91756
rect 24464 91702 24466 91754
rect 24466 91702 24518 91754
rect 24518 91702 24520 91754
rect 24464 91700 24520 91702
rect 24568 91754 24624 91756
rect 24568 91702 24570 91754
rect 24570 91702 24622 91754
rect 24622 91702 24624 91754
rect 24568 91700 24624 91702
rect 24672 91754 24728 91756
rect 24672 91702 24674 91754
rect 24674 91702 24726 91754
rect 24726 91702 24728 91754
rect 24672 91700 24728 91702
rect 24464 90186 24520 90188
rect 24464 90134 24466 90186
rect 24466 90134 24518 90186
rect 24518 90134 24520 90186
rect 24464 90132 24520 90134
rect 24568 90186 24624 90188
rect 24568 90134 24570 90186
rect 24570 90134 24622 90186
rect 24622 90134 24624 90186
rect 24568 90132 24624 90134
rect 24672 90186 24728 90188
rect 24672 90134 24674 90186
rect 24674 90134 24726 90186
rect 24726 90134 24728 90186
rect 24672 90132 24728 90134
rect 24332 88956 24388 89012
rect 24892 88732 24948 88788
rect 24464 88618 24520 88620
rect 24464 88566 24466 88618
rect 24466 88566 24518 88618
rect 24518 88566 24520 88618
rect 24464 88564 24520 88566
rect 24568 88618 24624 88620
rect 24568 88566 24570 88618
rect 24570 88566 24622 88618
rect 24622 88566 24624 88618
rect 24568 88564 24624 88566
rect 24672 88618 24728 88620
rect 24672 88566 24674 88618
rect 24674 88566 24726 88618
rect 24726 88566 24728 88618
rect 24672 88564 24728 88566
rect 24464 87050 24520 87052
rect 24464 86998 24466 87050
rect 24466 86998 24518 87050
rect 24518 86998 24520 87050
rect 24464 86996 24520 86998
rect 24568 87050 24624 87052
rect 24568 86998 24570 87050
rect 24570 86998 24622 87050
rect 24622 86998 24624 87050
rect 24568 86996 24624 86998
rect 24672 87050 24728 87052
rect 24672 86998 24674 87050
rect 24674 86998 24726 87050
rect 24726 86998 24728 87050
rect 24672 86996 24728 86998
rect 24444 85762 24500 85764
rect 24444 85710 24446 85762
rect 24446 85710 24498 85762
rect 24498 85710 24500 85762
rect 24444 85708 24500 85710
rect 24464 85482 24520 85484
rect 24464 85430 24466 85482
rect 24466 85430 24518 85482
rect 24518 85430 24520 85482
rect 24464 85428 24520 85430
rect 24568 85482 24624 85484
rect 24568 85430 24570 85482
rect 24570 85430 24622 85482
rect 24622 85430 24624 85482
rect 24568 85428 24624 85430
rect 24672 85482 24728 85484
rect 24672 85430 24674 85482
rect 24674 85430 24726 85482
rect 24726 85430 24728 85482
rect 24672 85428 24728 85430
rect 24332 85260 24388 85316
rect 24464 83914 24520 83916
rect 24464 83862 24466 83914
rect 24466 83862 24518 83914
rect 24518 83862 24520 83914
rect 24464 83860 24520 83862
rect 24568 83914 24624 83916
rect 24568 83862 24570 83914
rect 24570 83862 24622 83914
rect 24622 83862 24624 83914
rect 24568 83860 24624 83862
rect 24672 83914 24728 83916
rect 24672 83862 24674 83914
rect 24674 83862 24726 83914
rect 24726 83862 24728 83914
rect 24672 83860 24728 83862
rect 24464 82346 24520 82348
rect 24464 82294 24466 82346
rect 24466 82294 24518 82346
rect 24518 82294 24520 82346
rect 24464 82292 24520 82294
rect 24568 82346 24624 82348
rect 24568 82294 24570 82346
rect 24570 82294 24622 82346
rect 24622 82294 24624 82346
rect 24568 82292 24624 82294
rect 24672 82346 24728 82348
rect 24672 82294 24674 82346
rect 24674 82294 24726 82346
rect 24726 82294 24728 82346
rect 24672 82292 24728 82294
rect 24464 80778 24520 80780
rect 24464 80726 24466 80778
rect 24466 80726 24518 80778
rect 24518 80726 24520 80778
rect 24464 80724 24520 80726
rect 24568 80778 24624 80780
rect 24568 80726 24570 80778
rect 24570 80726 24622 80778
rect 24622 80726 24624 80778
rect 24568 80724 24624 80726
rect 24672 80778 24728 80780
rect 24672 80726 24674 80778
rect 24674 80726 24726 80778
rect 24726 80726 24728 80778
rect 24672 80724 24728 80726
rect 24464 79210 24520 79212
rect 24464 79158 24466 79210
rect 24466 79158 24518 79210
rect 24518 79158 24520 79210
rect 24464 79156 24520 79158
rect 24568 79210 24624 79212
rect 24568 79158 24570 79210
rect 24570 79158 24622 79210
rect 24622 79158 24624 79210
rect 24568 79156 24624 79158
rect 24672 79210 24728 79212
rect 24672 79158 24674 79210
rect 24674 79158 24726 79210
rect 24726 79158 24728 79210
rect 24672 79156 24728 79158
rect 24464 77642 24520 77644
rect 24464 77590 24466 77642
rect 24466 77590 24518 77642
rect 24518 77590 24520 77642
rect 24464 77588 24520 77590
rect 24568 77642 24624 77644
rect 24568 77590 24570 77642
rect 24570 77590 24622 77642
rect 24622 77590 24624 77642
rect 24568 77588 24624 77590
rect 24672 77642 24728 77644
rect 24672 77590 24674 77642
rect 24674 77590 24726 77642
rect 24726 77590 24728 77642
rect 24672 77588 24728 77590
rect 24464 76074 24520 76076
rect 24464 76022 24466 76074
rect 24466 76022 24518 76074
rect 24518 76022 24520 76074
rect 24464 76020 24520 76022
rect 24568 76074 24624 76076
rect 24568 76022 24570 76074
rect 24570 76022 24622 76074
rect 24622 76022 24624 76074
rect 24568 76020 24624 76022
rect 24672 76074 24728 76076
rect 24672 76022 24674 76074
rect 24674 76022 24726 76074
rect 24726 76022 24728 76074
rect 24672 76020 24728 76022
rect 24464 74506 24520 74508
rect 24464 74454 24466 74506
rect 24466 74454 24518 74506
rect 24518 74454 24520 74506
rect 24464 74452 24520 74454
rect 24568 74506 24624 74508
rect 24568 74454 24570 74506
rect 24570 74454 24622 74506
rect 24622 74454 24624 74506
rect 24568 74452 24624 74454
rect 24672 74506 24728 74508
rect 24672 74454 24674 74506
rect 24674 74454 24726 74506
rect 24726 74454 24728 74506
rect 24672 74452 24728 74454
rect 24464 72938 24520 72940
rect 24464 72886 24466 72938
rect 24466 72886 24518 72938
rect 24518 72886 24520 72938
rect 24464 72884 24520 72886
rect 24568 72938 24624 72940
rect 24568 72886 24570 72938
rect 24570 72886 24622 72938
rect 24622 72886 24624 72938
rect 24568 72884 24624 72886
rect 24672 72938 24728 72940
rect 24672 72886 24674 72938
rect 24674 72886 24726 72938
rect 24726 72886 24728 72938
rect 24672 72884 24728 72886
rect 24464 71370 24520 71372
rect 24464 71318 24466 71370
rect 24466 71318 24518 71370
rect 24518 71318 24520 71370
rect 24464 71316 24520 71318
rect 24568 71370 24624 71372
rect 24568 71318 24570 71370
rect 24570 71318 24622 71370
rect 24622 71318 24624 71370
rect 24568 71316 24624 71318
rect 24672 71370 24728 71372
rect 24672 71318 24674 71370
rect 24674 71318 24726 71370
rect 24726 71318 24728 71370
rect 24672 71316 24728 71318
rect 24464 69802 24520 69804
rect 24464 69750 24466 69802
rect 24466 69750 24518 69802
rect 24518 69750 24520 69802
rect 24464 69748 24520 69750
rect 24568 69802 24624 69804
rect 24568 69750 24570 69802
rect 24570 69750 24622 69802
rect 24622 69750 24624 69802
rect 24568 69748 24624 69750
rect 24672 69802 24728 69804
rect 24672 69750 24674 69802
rect 24674 69750 24726 69802
rect 24726 69750 24728 69802
rect 24672 69748 24728 69750
rect 23804 69018 23860 69020
rect 23804 68966 23806 69018
rect 23806 68966 23858 69018
rect 23858 68966 23860 69018
rect 23804 68964 23860 68966
rect 23908 69018 23964 69020
rect 23908 68966 23910 69018
rect 23910 68966 23962 69018
rect 23962 68966 23964 69018
rect 23908 68964 23964 68966
rect 24012 69018 24068 69020
rect 24012 68966 24014 69018
rect 24014 68966 24066 69018
rect 24066 68966 24068 69018
rect 24012 68964 24068 68966
rect 24220 68908 24276 68964
rect 24332 68796 24388 68852
rect 24668 68626 24724 68628
rect 24668 68574 24670 68626
rect 24670 68574 24722 68626
rect 24722 68574 24724 68626
rect 24668 68572 24724 68574
rect 24444 68348 24500 68404
rect 24464 68234 24520 68236
rect 24464 68182 24466 68234
rect 24466 68182 24518 68234
rect 24518 68182 24520 68234
rect 24464 68180 24520 68182
rect 24568 68234 24624 68236
rect 24568 68182 24570 68234
rect 24570 68182 24622 68234
rect 24622 68182 24624 68234
rect 24568 68180 24624 68182
rect 24672 68234 24728 68236
rect 24672 68182 24674 68234
rect 24674 68182 24726 68234
rect 24726 68182 24728 68234
rect 24672 68180 24728 68182
rect 23660 67452 23716 67508
rect 23804 67450 23860 67452
rect 23804 67398 23806 67450
rect 23806 67398 23858 67450
rect 23858 67398 23860 67450
rect 23804 67396 23860 67398
rect 23908 67450 23964 67452
rect 23908 67398 23910 67450
rect 23910 67398 23962 67450
rect 23962 67398 23964 67450
rect 23908 67396 23964 67398
rect 24012 67450 24068 67452
rect 24012 67398 24014 67450
rect 24014 67398 24066 67450
rect 24066 67398 24068 67450
rect 24012 67396 24068 67398
rect 23436 67228 23492 67284
rect 24464 66666 24520 66668
rect 24464 66614 24466 66666
rect 24466 66614 24518 66666
rect 24518 66614 24520 66666
rect 24464 66612 24520 66614
rect 24568 66666 24624 66668
rect 24568 66614 24570 66666
rect 24570 66614 24622 66666
rect 24622 66614 24624 66666
rect 24568 66612 24624 66614
rect 24672 66666 24728 66668
rect 24672 66614 24674 66666
rect 24674 66614 24726 66666
rect 24726 66614 24728 66666
rect 24672 66612 24728 66614
rect 23804 65882 23860 65884
rect 23804 65830 23806 65882
rect 23806 65830 23858 65882
rect 23858 65830 23860 65882
rect 23804 65828 23860 65830
rect 23908 65882 23964 65884
rect 23908 65830 23910 65882
rect 23910 65830 23962 65882
rect 23962 65830 23964 65882
rect 23908 65828 23964 65830
rect 24012 65882 24068 65884
rect 24012 65830 24014 65882
rect 24014 65830 24066 65882
rect 24066 65830 24068 65882
rect 24012 65828 24068 65830
rect 24464 65098 24520 65100
rect 24464 65046 24466 65098
rect 24466 65046 24518 65098
rect 24518 65046 24520 65098
rect 24464 65044 24520 65046
rect 24568 65098 24624 65100
rect 24568 65046 24570 65098
rect 24570 65046 24622 65098
rect 24622 65046 24624 65098
rect 24568 65044 24624 65046
rect 24672 65098 24728 65100
rect 24672 65046 24674 65098
rect 24674 65046 24726 65098
rect 24726 65046 24728 65098
rect 24672 65044 24728 65046
rect 23804 64314 23860 64316
rect 23804 64262 23806 64314
rect 23806 64262 23858 64314
rect 23858 64262 23860 64314
rect 23804 64260 23860 64262
rect 23908 64314 23964 64316
rect 23908 64262 23910 64314
rect 23910 64262 23962 64314
rect 23962 64262 23964 64314
rect 23908 64260 23964 64262
rect 24012 64314 24068 64316
rect 24012 64262 24014 64314
rect 24014 64262 24066 64314
rect 24066 64262 24068 64314
rect 24012 64260 24068 64262
rect 24464 63530 24520 63532
rect 24464 63478 24466 63530
rect 24466 63478 24518 63530
rect 24518 63478 24520 63530
rect 24464 63476 24520 63478
rect 24568 63530 24624 63532
rect 24568 63478 24570 63530
rect 24570 63478 24622 63530
rect 24622 63478 24624 63530
rect 24568 63476 24624 63478
rect 24672 63530 24728 63532
rect 24672 63478 24674 63530
rect 24674 63478 24726 63530
rect 24726 63478 24728 63530
rect 24672 63476 24728 63478
rect 23804 62746 23860 62748
rect 23804 62694 23806 62746
rect 23806 62694 23858 62746
rect 23858 62694 23860 62746
rect 23804 62692 23860 62694
rect 23908 62746 23964 62748
rect 23908 62694 23910 62746
rect 23910 62694 23962 62746
rect 23962 62694 23964 62746
rect 23908 62692 23964 62694
rect 24012 62746 24068 62748
rect 24012 62694 24014 62746
rect 24014 62694 24066 62746
rect 24066 62694 24068 62746
rect 24012 62692 24068 62694
rect 23772 62354 23828 62356
rect 23772 62302 23774 62354
rect 23774 62302 23826 62354
rect 23826 62302 23828 62354
rect 23772 62300 23828 62302
rect 22764 61180 22820 61236
rect 22204 60732 22260 60788
rect 22428 60844 22484 60900
rect 22204 59890 22260 59892
rect 22204 59838 22206 59890
rect 22206 59838 22258 59890
rect 22258 59838 22260 59890
rect 22204 59836 22260 59838
rect 22092 59276 22148 59332
rect 21756 53676 21812 53732
rect 21868 44828 21924 44884
rect 20860 41580 20916 41636
rect 21084 41186 21140 41188
rect 21084 41134 21086 41186
rect 21086 41134 21138 41186
rect 21138 41134 21140 41186
rect 21084 41132 21140 41134
rect 20972 40402 21028 40404
rect 20972 40350 20974 40402
rect 20974 40350 21026 40402
rect 21026 40350 21028 40402
rect 20972 40348 21028 40350
rect 20860 40236 20916 40292
rect 20860 39004 20916 39060
rect 19964 36092 20020 36148
rect 19740 35586 19796 35588
rect 19740 35534 19742 35586
rect 19742 35534 19794 35586
rect 19794 35534 19796 35586
rect 19740 35532 19796 35534
rect 19852 34300 19908 34356
rect 19628 33852 19684 33908
rect 19740 33628 19796 33684
rect 19516 33346 19572 33348
rect 19516 33294 19518 33346
rect 19518 33294 19570 33346
rect 19570 33294 19572 33346
rect 19516 33292 19572 33294
rect 20188 35308 20244 35364
rect 20188 35084 20244 35140
rect 19852 33234 19908 33236
rect 19852 33182 19854 33234
rect 19854 33182 19906 33234
rect 19906 33182 19908 33234
rect 19852 33180 19908 33182
rect 18172 31388 18228 31444
rect 18060 30156 18116 30212
rect 18508 31218 18564 31220
rect 18508 31166 18510 31218
rect 18510 31166 18562 31218
rect 18562 31166 18564 31218
rect 18508 31164 18564 31166
rect 18620 31052 18676 31108
rect 18396 30098 18452 30100
rect 18396 30046 18398 30098
rect 18398 30046 18450 30098
rect 18450 30046 18452 30098
rect 18396 30044 18452 30046
rect 18284 29932 18340 29988
rect 16380 25228 16436 25284
rect 16268 25116 16324 25172
rect 16156 24892 16212 24948
rect 14812 23100 14868 23156
rect 15260 23436 15316 23492
rect 15484 23154 15540 23156
rect 15484 23102 15486 23154
rect 15486 23102 15538 23154
rect 15538 23102 15540 23154
rect 15484 23100 15540 23102
rect 15036 22988 15092 23044
rect 14924 22594 14980 22596
rect 14924 22542 14926 22594
rect 14926 22542 14978 22594
rect 14978 22542 14980 22594
rect 14924 22540 14980 22542
rect 14812 22092 14868 22148
rect 14364 21532 14420 21588
rect 14812 21868 14868 21924
rect 14140 21084 14196 21140
rect 13916 20802 13972 20804
rect 13916 20750 13918 20802
rect 13918 20750 13970 20802
rect 13970 20750 13972 20802
rect 13916 20748 13972 20750
rect 14476 20412 14532 20468
rect 14700 21532 14756 21588
rect 14812 20972 14868 21028
rect 15596 22764 15652 22820
rect 15708 22540 15764 22596
rect 15372 22204 15428 22260
rect 15820 21644 15876 21700
rect 15708 20860 15764 20916
rect 16044 20860 16100 20916
rect 17388 25506 17444 25508
rect 17388 25454 17390 25506
rect 17390 25454 17442 25506
rect 17442 25454 17444 25506
rect 17388 25452 17444 25454
rect 17164 24892 17220 24948
rect 17276 24722 17332 24724
rect 17276 24670 17278 24722
rect 17278 24670 17330 24722
rect 17330 24670 17332 24722
rect 17276 24668 17332 24670
rect 16716 24610 16772 24612
rect 16716 24558 16718 24610
rect 16718 24558 16770 24610
rect 16770 24558 16772 24610
rect 16716 24556 16772 24558
rect 17724 26236 17780 26292
rect 17724 24668 17780 24724
rect 16380 22204 16436 22260
rect 17164 23660 17220 23716
rect 16940 22428 16996 22484
rect 17052 23100 17108 23156
rect 16828 22204 16884 22260
rect 15708 20636 15764 20692
rect 15260 19964 15316 20020
rect 13916 18732 13972 18788
rect 14588 18732 14644 18788
rect 14476 18508 14532 18564
rect 15148 18956 15204 19012
rect 15260 18732 15316 18788
rect 15148 18508 15204 18564
rect 15596 20578 15652 20580
rect 15596 20526 15598 20578
rect 15598 20526 15650 20578
rect 15650 20526 15652 20578
rect 15596 20524 15652 20526
rect 15372 18508 15428 18564
rect 15484 19852 15540 19908
rect 14700 17612 14756 17668
rect 14924 17778 14980 17780
rect 14924 17726 14926 17778
rect 14926 17726 14978 17778
rect 14978 17726 14980 17778
rect 14924 17724 14980 17726
rect 14924 17052 14980 17108
rect 15036 17164 15092 17220
rect 14028 16098 14084 16100
rect 14028 16046 14030 16098
rect 14030 16046 14082 16098
rect 14082 16046 14084 16098
rect 14028 16044 14084 16046
rect 13916 15260 13972 15316
rect 14028 15372 14084 15428
rect 14140 15148 14196 15204
rect 13468 14700 13524 14756
rect 13580 14476 13636 14532
rect 13356 13132 13412 13188
rect 13468 13356 13524 13412
rect 13468 12796 13524 12852
rect 14028 14812 14084 14868
rect 13916 14754 13972 14756
rect 13916 14702 13918 14754
rect 13918 14702 13970 14754
rect 13970 14702 13972 14754
rect 13916 14700 13972 14702
rect 13916 13916 13972 13972
rect 13804 13468 13860 13524
rect 13804 13244 13860 13300
rect 13916 12908 13972 12964
rect 14364 16604 14420 16660
rect 14140 13186 14196 13188
rect 14140 13134 14142 13186
rect 14142 13134 14194 13186
rect 14194 13134 14196 13186
rect 14140 13132 14196 13134
rect 14028 12066 14084 12068
rect 14028 12014 14030 12066
rect 14030 12014 14082 12066
rect 14082 12014 14084 12066
rect 14028 12012 14084 12014
rect 13916 11506 13972 11508
rect 13916 11454 13918 11506
rect 13918 11454 13970 11506
rect 13970 11454 13972 11506
rect 13916 11452 13972 11454
rect 13468 10556 13524 10612
rect 13356 8204 13412 8260
rect 11564 4620 11620 4676
rect 11564 4338 11620 4340
rect 11564 4286 11566 4338
rect 11566 4286 11618 4338
rect 11618 4286 11620 4338
rect 11564 4284 11620 4286
rect 11452 3507 11454 3556
rect 11454 3507 11506 3556
rect 11506 3507 11508 3556
rect 11452 3500 11508 3507
rect 11340 2940 11396 2996
rect 11900 5628 11956 5684
rect 12236 7196 12292 7252
rect 12460 6690 12516 6692
rect 12460 6638 12462 6690
rect 12462 6638 12514 6690
rect 12514 6638 12516 6690
rect 12460 6636 12516 6638
rect 12908 6412 12964 6468
rect 12236 5234 12292 5236
rect 12236 5182 12238 5234
rect 12238 5182 12290 5234
rect 12290 5182 12292 5234
rect 12236 5180 12292 5182
rect 12236 4338 12292 4340
rect 12236 4286 12238 4338
rect 12238 4286 12290 4338
rect 12290 4286 12292 4338
rect 12236 4284 12292 4286
rect 12908 5068 12964 5124
rect 12684 3724 12740 3780
rect 11004 924 11060 980
rect 10780 588 10836 644
rect 10556 476 10612 532
rect 11788 3500 11844 3556
rect 11676 2604 11732 2660
rect 11564 2546 11620 2548
rect 11564 2494 11566 2546
rect 11566 2494 11618 2546
rect 11618 2494 11620 2546
rect 11564 2492 11620 2494
rect 11788 2492 11844 2548
rect 11788 2156 11844 2212
rect 11116 252 11172 308
rect 11228 1596 11284 1652
rect 11452 1596 11508 1652
rect 11564 1260 11620 1316
rect 11676 1484 11732 1540
rect 11900 1596 11956 1652
rect 12012 1372 12068 1428
rect 12124 1596 12180 1652
rect 13356 7420 13412 7476
rect 13244 7362 13300 7364
rect 13244 7310 13246 7362
rect 13246 7310 13298 7362
rect 13298 7310 13300 7362
rect 13244 7308 13300 7310
rect 13244 5292 13300 5348
rect 13580 9884 13636 9940
rect 13692 9436 13748 9492
rect 13580 9154 13636 9156
rect 13580 9102 13582 9154
rect 13582 9102 13634 9154
rect 13634 9102 13636 9154
rect 13580 9100 13636 9102
rect 13580 7980 13636 8036
rect 13916 10892 13972 10948
rect 14140 10892 14196 10948
rect 14476 15596 14532 15652
rect 15596 19740 15652 19796
rect 16044 20636 16100 20692
rect 16044 19906 16100 19908
rect 16044 19854 16046 19906
rect 16046 19854 16098 19906
rect 16098 19854 16100 19906
rect 16044 19852 16100 19854
rect 15932 19346 15988 19348
rect 15932 19294 15934 19346
rect 15934 19294 15986 19346
rect 15986 19294 15988 19346
rect 15932 19292 15988 19294
rect 15596 18956 15652 19012
rect 15596 18338 15652 18340
rect 15596 18286 15598 18338
rect 15598 18286 15650 18338
rect 15650 18286 15652 18338
rect 15596 18284 15652 18286
rect 15484 15148 15540 15204
rect 15596 18060 15652 18116
rect 17724 23548 17780 23604
rect 17500 23154 17556 23156
rect 17500 23102 17502 23154
rect 17502 23102 17554 23154
rect 17554 23102 17556 23154
rect 17500 23100 17556 23102
rect 17276 22204 17332 22260
rect 16604 21196 16660 21252
rect 16492 20972 16548 21028
rect 16156 18172 16212 18228
rect 15932 15314 15988 15316
rect 15932 15262 15934 15314
rect 15934 15262 15986 15314
rect 15986 15262 15988 15314
rect 15932 15260 15988 15262
rect 15372 14700 15428 14756
rect 14812 14364 14868 14420
rect 15036 14364 15092 14420
rect 14588 14028 14644 14084
rect 15036 14028 15092 14084
rect 14700 13692 14756 13748
rect 14588 13580 14644 13636
rect 14364 10556 14420 10612
rect 14252 10332 14308 10388
rect 15708 12460 15764 12516
rect 15708 11340 15764 11396
rect 14700 11004 14756 11060
rect 14028 9826 14084 9828
rect 14028 9774 14030 9826
rect 14030 9774 14082 9826
rect 14082 9774 14084 9826
rect 14028 9772 14084 9774
rect 14924 10780 14980 10836
rect 13916 9042 13972 9044
rect 13916 8990 13918 9042
rect 13918 8990 13970 9042
rect 13970 8990 13972 9042
rect 13916 8988 13972 8990
rect 13804 7868 13860 7924
rect 13580 7532 13636 7588
rect 13692 7420 13748 7476
rect 13580 6972 13636 7028
rect 13916 7250 13972 7252
rect 13916 7198 13918 7250
rect 13918 7198 13970 7250
rect 13970 7198 13972 7250
rect 13916 7196 13972 7198
rect 13580 6524 13636 6580
rect 13580 6300 13636 6356
rect 13356 5068 13412 5124
rect 13468 5404 13524 5460
rect 13356 4338 13412 4340
rect 13356 4286 13358 4338
rect 13358 4286 13410 4338
rect 13410 4286 13412 4338
rect 13356 4284 13412 4286
rect 12908 2156 12964 2212
rect 12796 2098 12852 2100
rect 12796 2046 12798 2098
rect 12798 2046 12850 2098
rect 12850 2046 12852 2098
rect 12796 2044 12852 2046
rect 12348 1986 12404 1988
rect 12348 1934 12350 1986
rect 12350 1934 12402 1986
rect 12402 1934 12404 1986
rect 12348 1932 12404 1934
rect 12236 588 12292 644
rect 12348 1596 12404 1652
rect 12572 1596 12628 1652
rect 12796 1596 12852 1652
rect 12684 1036 12740 1092
rect 13020 1596 13076 1652
rect 13356 3388 13412 3444
rect 13244 2940 13300 2996
rect 14588 9212 14644 9268
rect 14700 9436 14756 9492
rect 14476 9100 14532 9156
rect 14364 9042 14420 9044
rect 14364 8990 14366 9042
rect 14366 8990 14418 9042
rect 14418 8990 14420 9042
rect 14364 8988 14420 8990
rect 14588 8930 14644 8932
rect 14588 8878 14590 8930
rect 14590 8878 14642 8930
rect 14642 8878 14644 8930
rect 14588 8876 14644 8878
rect 14588 8258 14644 8260
rect 14588 8206 14590 8258
rect 14590 8206 14642 8258
rect 14642 8206 14644 8258
rect 14588 8204 14644 8206
rect 14364 6690 14420 6692
rect 14364 6638 14366 6690
rect 14366 6638 14418 6690
rect 14418 6638 14420 6690
rect 14364 6636 14420 6638
rect 14476 6412 14532 6468
rect 15708 11116 15764 11172
rect 15708 10108 15764 10164
rect 15260 9660 15316 9716
rect 15484 8764 15540 8820
rect 15148 6748 15204 6804
rect 14700 6300 14756 6356
rect 14812 6412 14868 6468
rect 13580 5292 13636 5348
rect 14028 5292 14084 5348
rect 13916 5068 13972 5124
rect 13580 4508 13636 4564
rect 13692 3554 13748 3556
rect 13692 3502 13694 3554
rect 13694 3502 13746 3554
rect 13746 3502 13748 3554
rect 13692 3500 13748 3502
rect 13692 2940 13748 2996
rect 13244 1932 13300 1988
rect 13132 1148 13188 1204
rect 13244 1596 13300 1652
rect 13132 252 13188 308
rect 14028 2940 14084 2996
rect 14252 5122 14308 5124
rect 14252 5070 14254 5122
rect 14254 5070 14306 5122
rect 14306 5070 14308 5122
rect 14252 5068 14308 5070
rect 14140 2716 14196 2772
rect 14028 2658 14084 2660
rect 14028 2606 14030 2658
rect 14030 2606 14082 2658
rect 14082 2606 14084 2658
rect 14028 2604 14084 2606
rect 13916 1260 13972 1316
rect 14028 252 14084 308
rect 14140 2492 14196 2548
rect 14700 5628 14756 5684
rect 14476 3948 14532 4004
rect 14588 3554 14644 3556
rect 14588 3502 14590 3554
rect 14590 3502 14642 3554
rect 14642 3502 14644 3554
rect 14588 3500 14644 3502
rect 15372 7474 15428 7476
rect 15372 7422 15374 7474
rect 15374 7422 15426 7474
rect 15426 7422 15428 7474
rect 15372 7420 15428 7422
rect 14924 5516 14980 5572
rect 15148 4844 15204 4900
rect 15148 3388 15204 3444
rect 14700 2604 14756 2660
rect 14364 1986 14420 1988
rect 14364 1934 14366 1986
rect 14366 1934 14418 1986
rect 14418 1934 14420 1986
rect 14364 1932 14420 1934
rect 14700 1596 14756 1652
rect 14812 1202 14868 1204
rect 14812 1150 14814 1202
rect 14814 1150 14866 1202
rect 14866 1150 14868 1202
rect 14812 1148 14868 1150
rect 15596 7868 15652 7924
rect 15596 5906 15652 5908
rect 15596 5854 15598 5906
rect 15598 5854 15650 5906
rect 15650 5854 15652 5906
rect 15596 5852 15652 5854
rect 16044 13356 16100 13412
rect 16044 10220 16100 10276
rect 16268 15202 16324 15204
rect 16268 15150 16270 15202
rect 16270 15150 16322 15202
rect 16322 15150 16324 15202
rect 16268 15148 16324 15150
rect 16380 12124 16436 12180
rect 15932 6524 15988 6580
rect 15484 5516 15540 5572
rect 15372 5346 15428 5348
rect 15372 5294 15374 5346
rect 15374 5294 15426 5346
rect 15426 5294 15428 5346
rect 15372 5292 15428 5294
rect 15708 5292 15764 5348
rect 15372 5068 15428 5124
rect 15036 2828 15092 2884
rect 15260 2268 15316 2324
rect 14812 924 14868 980
rect 15036 978 15092 980
rect 15036 926 15038 978
rect 15038 926 15090 978
rect 15090 926 15092 978
rect 15036 924 15092 926
rect 14588 700 14644 756
rect 15036 700 15092 756
rect 14812 364 14868 420
rect 15596 4562 15652 4564
rect 15596 4510 15598 4562
rect 15598 4510 15650 4562
rect 15650 4510 15652 4562
rect 15596 4508 15652 4510
rect 15372 1708 15428 1764
rect 15932 5180 15988 5236
rect 15708 2770 15764 2772
rect 15708 2718 15710 2770
rect 15710 2718 15762 2770
rect 15762 2718 15764 2770
rect 15708 2716 15764 2718
rect 16268 7980 16324 8036
rect 16156 6636 16212 6692
rect 16268 4508 16324 4564
rect 17052 20748 17108 20804
rect 16940 19740 16996 19796
rect 17388 21756 17444 21812
rect 17164 19292 17220 19348
rect 17388 19180 17444 19236
rect 16940 18396 16996 18452
rect 16716 17836 16772 17892
rect 17612 22540 17668 22596
rect 17612 22258 17668 22260
rect 17612 22206 17614 22258
rect 17614 22206 17666 22258
rect 17666 22206 17668 22258
rect 17612 22204 17668 22206
rect 17948 26850 18004 26852
rect 17948 26798 17950 26850
rect 17950 26798 18002 26850
rect 18002 26798 18004 26850
rect 17948 26796 18004 26798
rect 19068 31890 19124 31892
rect 19068 31838 19070 31890
rect 19070 31838 19122 31890
rect 19122 31838 19124 31890
rect 19068 31836 19124 31838
rect 19292 31778 19348 31780
rect 19292 31726 19294 31778
rect 19294 31726 19346 31778
rect 19346 31726 19348 31778
rect 19292 31724 19348 31726
rect 19852 32508 19908 32564
rect 19740 32396 19796 32452
rect 19404 31500 19460 31556
rect 18844 31388 18900 31444
rect 19628 31666 19684 31668
rect 19628 31614 19630 31666
rect 19630 31614 19682 31666
rect 19682 31614 19684 31666
rect 19628 31612 19684 31614
rect 18844 30770 18900 30772
rect 18844 30718 18846 30770
rect 18846 30718 18898 30770
rect 18898 30718 18900 30770
rect 18844 30716 18900 30718
rect 18844 30492 18900 30548
rect 18732 29484 18788 29540
rect 18620 28866 18676 28868
rect 18620 28814 18622 28866
rect 18622 28814 18674 28866
rect 18674 28814 18676 28866
rect 18620 28812 18676 28814
rect 18396 28588 18452 28644
rect 18508 28476 18564 28532
rect 19068 30044 19124 30100
rect 18844 29426 18900 29428
rect 18844 29374 18846 29426
rect 18846 29374 18898 29426
rect 18898 29374 18900 29426
rect 18844 29372 18900 29374
rect 19068 28530 19124 28532
rect 19068 28478 19070 28530
rect 19070 28478 19122 28530
rect 19122 28478 19124 28530
rect 19068 28476 19124 28478
rect 19180 28028 19236 28084
rect 18732 27746 18788 27748
rect 18732 27694 18734 27746
rect 18734 27694 18786 27746
rect 18786 27694 18788 27746
rect 18732 27692 18788 27694
rect 18732 27468 18788 27524
rect 18620 27298 18676 27300
rect 18620 27246 18622 27298
rect 18622 27246 18674 27298
rect 18674 27246 18676 27298
rect 18620 27244 18676 27246
rect 19292 27580 19348 27636
rect 19628 30044 19684 30100
rect 19516 29932 19572 29988
rect 19516 29372 19572 29428
rect 20076 33122 20132 33124
rect 20076 33070 20078 33122
rect 20078 33070 20130 33122
rect 20130 33070 20132 33122
rect 20076 33068 20132 33070
rect 20076 30994 20132 30996
rect 20076 30942 20078 30994
rect 20078 30942 20130 30994
rect 20130 30942 20132 30994
rect 20076 30940 20132 30942
rect 20076 30492 20132 30548
rect 19852 28812 19908 28868
rect 19964 29986 20020 29988
rect 19964 29934 19966 29986
rect 19966 29934 20018 29986
rect 20018 29934 20020 29986
rect 19964 29932 20020 29934
rect 20076 28588 20132 28644
rect 19516 28028 19572 28084
rect 20076 28418 20132 28420
rect 20076 28366 20078 28418
rect 20078 28366 20130 28418
rect 20130 28366 20132 28418
rect 20076 28364 20132 28366
rect 19292 27244 19348 27300
rect 19964 28082 20020 28084
rect 19964 28030 19966 28082
rect 19966 28030 20018 28082
rect 20018 28030 20020 28082
rect 19964 28028 20020 28030
rect 19852 27692 19908 27748
rect 18844 27020 18900 27076
rect 19180 27020 19236 27076
rect 18060 26012 18116 26068
rect 17948 25730 18004 25732
rect 17948 25678 17950 25730
rect 17950 25678 18002 25730
rect 18002 25678 18004 25730
rect 17948 25676 18004 25678
rect 17836 21532 17892 21588
rect 17948 24556 18004 24612
rect 17612 20860 17668 20916
rect 17724 19404 17780 19460
rect 17724 19180 17780 19236
rect 18060 24332 18116 24388
rect 18172 23660 18228 23716
rect 18284 26348 18340 26404
rect 18060 22988 18116 23044
rect 19068 26796 19124 26852
rect 18732 26460 18788 26516
rect 18620 25340 18676 25396
rect 18396 23884 18452 23940
rect 18396 23154 18452 23156
rect 18396 23102 18398 23154
rect 18398 23102 18450 23154
rect 18450 23102 18452 23154
rect 18396 23100 18452 23102
rect 18060 22316 18116 22372
rect 18396 22204 18452 22260
rect 18172 21532 18228 21588
rect 17948 19852 18004 19908
rect 18060 20524 18116 20580
rect 17948 19068 18004 19124
rect 17836 18172 17892 18228
rect 17052 15596 17108 15652
rect 17388 15484 17444 15540
rect 17500 14530 17556 14532
rect 17500 14478 17502 14530
rect 17502 14478 17554 14530
rect 17554 14478 17556 14530
rect 17500 14476 17556 14478
rect 16604 13468 16660 13524
rect 16828 13692 16884 13748
rect 16940 13634 16996 13636
rect 16940 13582 16942 13634
rect 16942 13582 16994 13634
rect 16994 13582 16996 13634
rect 16940 13580 16996 13582
rect 17276 13580 17332 13636
rect 16716 13356 16772 13412
rect 16716 12178 16772 12180
rect 16716 12126 16718 12178
rect 16718 12126 16770 12178
rect 16770 12126 16772 12178
rect 16716 12124 16772 12126
rect 16828 12572 16884 12628
rect 16716 10050 16772 10052
rect 16716 9998 16718 10050
rect 16718 9998 16770 10050
rect 16770 9998 16772 10050
rect 16716 9996 16772 9998
rect 17052 12348 17108 12404
rect 17164 11676 17220 11732
rect 16828 8988 16884 9044
rect 17948 16604 18004 16660
rect 17724 15596 17780 15652
rect 17724 13692 17780 13748
rect 17836 13468 17892 13524
rect 17948 15372 18004 15428
rect 17612 11788 17668 11844
rect 17724 12684 17780 12740
rect 17388 11564 17444 11620
rect 16940 9772 16996 9828
rect 16828 8034 16884 8036
rect 16828 7982 16830 8034
rect 16830 7982 16882 8034
rect 16882 7982 16884 8034
rect 16828 7980 16884 7982
rect 16940 7756 16996 7812
rect 16604 6524 16660 6580
rect 16828 5516 16884 5572
rect 16940 6300 16996 6356
rect 16492 5068 16548 5124
rect 16268 4338 16324 4340
rect 16268 4286 16270 4338
rect 16270 4286 16322 4338
rect 16322 4286 16324 4338
rect 16268 4284 16324 4286
rect 17276 9154 17332 9156
rect 17276 9102 17278 9154
rect 17278 9102 17330 9154
rect 17330 9102 17332 9154
rect 17276 9100 17332 9102
rect 17388 8876 17444 8932
rect 17388 8428 17444 8484
rect 18060 15932 18116 15988
rect 18060 15314 18116 15316
rect 18060 15262 18062 15314
rect 18062 15262 18114 15314
rect 18114 15262 18116 15314
rect 18060 15260 18116 15262
rect 18396 21586 18452 21588
rect 18396 21534 18398 21586
rect 18398 21534 18450 21586
rect 18450 21534 18452 21586
rect 18396 21532 18452 21534
rect 18396 19852 18452 19908
rect 18620 19852 18676 19908
rect 18284 19404 18340 19460
rect 18508 19458 18564 19460
rect 18508 19406 18510 19458
rect 18510 19406 18562 19458
rect 18562 19406 18564 19458
rect 18508 19404 18564 19406
rect 18508 17948 18564 18004
rect 18284 17388 18340 17444
rect 18620 17778 18676 17780
rect 18620 17726 18622 17778
rect 18622 17726 18674 17778
rect 18674 17726 18676 17778
rect 18620 17724 18676 17726
rect 18508 16828 18564 16884
rect 18172 15708 18228 15764
rect 18956 25228 19012 25284
rect 18844 23042 18900 23044
rect 18844 22990 18846 23042
rect 18846 22990 18898 23042
rect 18898 22990 18900 23042
rect 18844 22988 18900 22990
rect 18844 22092 18900 22148
rect 19516 26908 19572 26964
rect 20076 27244 20132 27300
rect 19516 25228 19572 25284
rect 19404 23212 19460 23268
rect 19180 21532 19236 21588
rect 19292 21196 19348 21252
rect 19180 19852 19236 19908
rect 19068 19516 19124 19572
rect 18956 17836 19012 17892
rect 18844 16716 18900 16772
rect 18396 14476 18452 14532
rect 18284 13804 18340 13860
rect 18284 12796 18340 12852
rect 17948 11676 18004 11732
rect 18732 14812 18788 14868
rect 18956 15820 19012 15876
rect 19180 18844 19236 18900
rect 18732 14530 18788 14532
rect 18732 14478 18734 14530
rect 18734 14478 18786 14530
rect 18786 14478 18788 14530
rect 18732 14476 18788 14478
rect 18732 13468 18788 13524
rect 18732 12908 18788 12964
rect 18620 12012 18676 12068
rect 18508 10332 18564 10388
rect 18396 9884 18452 9940
rect 18060 9826 18116 9828
rect 18060 9774 18062 9826
rect 18062 9774 18114 9826
rect 18114 9774 18116 9826
rect 18060 9772 18116 9774
rect 17724 7980 17780 8036
rect 17500 7084 17556 7140
rect 17948 8370 18004 8372
rect 17948 8318 17950 8370
rect 17950 8318 18002 8370
rect 18002 8318 18004 8370
rect 17948 8316 18004 8318
rect 18396 8092 18452 8148
rect 18508 8652 18564 8708
rect 17836 7196 17892 7252
rect 18060 6748 18116 6804
rect 17612 6524 17668 6580
rect 18284 6524 18340 6580
rect 17052 4956 17108 5012
rect 17164 4508 17220 4564
rect 16828 3554 16884 3556
rect 16828 3502 16830 3554
rect 16830 3502 16882 3554
rect 16882 3502 16884 3554
rect 16828 3500 16884 3502
rect 15708 2210 15764 2212
rect 15708 2158 15710 2210
rect 15710 2158 15762 2210
rect 15762 2158 15764 2210
rect 15708 2156 15764 2158
rect 16044 2098 16100 2100
rect 16044 2046 16046 2098
rect 16046 2046 16098 2098
rect 16098 2046 16100 2098
rect 16044 2044 16100 2046
rect 16716 3052 16772 3108
rect 16604 2940 16660 2996
rect 16716 2828 16772 2884
rect 17052 2828 17108 2884
rect 16940 2492 16996 2548
rect 15708 812 15764 868
rect 15596 476 15652 532
rect 15708 588 15764 644
rect 16156 812 16212 868
rect 17836 5404 17892 5460
rect 17724 5068 17780 5124
rect 17500 2156 17556 2212
rect 17612 2940 17668 2996
rect 17164 2098 17220 2100
rect 17164 2046 17166 2098
rect 17166 2046 17218 2098
rect 17218 2046 17220 2098
rect 17164 2044 17220 2046
rect 17836 1820 17892 1876
rect 17500 1036 17556 1092
rect 18284 5068 18340 5124
rect 18284 4338 18340 4340
rect 18284 4286 18286 4338
rect 18286 4286 18338 4338
rect 18338 4286 18340 4338
rect 18284 4284 18340 4286
rect 18396 3612 18452 3668
rect 18956 12908 19012 12964
rect 19068 14812 19124 14868
rect 18844 9154 18900 9156
rect 18844 9102 18846 9154
rect 18846 9102 18898 9154
rect 18898 9102 18900 9154
rect 18844 9100 18900 9102
rect 18956 8652 19012 8708
rect 19180 13132 19236 13188
rect 19180 11618 19236 11620
rect 19180 11566 19182 11618
rect 19182 11566 19234 11618
rect 19234 11566 19236 11618
rect 19180 11564 19236 11566
rect 19068 8316 19124 8372
rect 19180 9436 19236 9492
rect 19180 8988 19236 9044
rect 18732 7644 18788 7700
rect 18844 7420 18900 7476
rect 18956 7308 19012 7364
rect 19068 6636 19124 6692
rect 19180 6524 19236 6580
rect 19516 21868 19572 21924
rect 19628 21084 19684 21140
rect 20524 36316 20580 36372
rect 20300 32508 20356 32564
rect 20524 35308 20580 35364
rect 21084 38108 21140 38164
rect 20748 35868 20804 35924
rect 20748 35420 20804 35476
rect 20860 35196 20916 35252
rect 20972 35810 21028 35812
rect 20972 35758 20974 35810
rect 20974 35758 21026 35810
rect 21026 35758 21028 35810
rect 20972 35756 21028 35758
rect 21308 41916 21364 41972
rect 21532 41916 21588 41972
rect 21644 41858 21700 41860
rect 21644 41806 21646 41858
rect 21646 41806 21698 41858
rect 21698 41806 21700 41858
rect 21644 41804 21700 41806
rect 21420 41468 21476 41524
rect 21756 41692 21812 41748
rect 21308 40684 21364 40740
rect 21532 40796 21588 40852
rect 21644 40460 21700 40516
rect 21308 40236 21364 40292
rect 22204 44492 22260 44548
rect 22092 43538 22148 43540
rect 22092 43486 22094 43538
rect 22094 43486 22146 43538
rect 22146 43486 22148 43538
rect 22092 43484 22148 43486
rect 21420 38722 21476 38724
rect 21420 38670 21422 38722
rect 21422 38670 21474 38722
rect 21474 38670 21476 38722
rect 21420 38668 21476 38670
rect 21308 37884 21364 37940
rect 21308 37436 21364 37492
rect 21420 37042 21476 37044
rect 21420 36990 21422 37042
rect 21422 36990 21474 37042
rect 21474 36990 21476 37042
rect 21420 36988 21476 36990
rect 21308 36316 21364 36372
rect 21196 35084 21252 35140
rect 21196 34914 21252 34916
rect 21196 34862 21198 34914
rect 21198 34862 21250 34914
rect 21250 34862 21252 34914
rect 21196 34860 21252 34862
rect 21420 35698 21476 35700
rect 21420 35646 21422 35698
rect 21422 35646 21474 35698
rect 21474 35646 21476 35698
rect 21420 35644 21476 35646
rect 22092 41916 22148 41972
rect 22652 60620 22708 60676
rect 24464 61962 24520 61964
rect 24464 61910 24466 61962
rect 24466 61910 24518 61962
rect 24518 61910 24520 61962
rect 24464 61908 24520 61910
rect 24568 61962 24624 61964
rect 24568 61910 24570 61962
rect 24570 61910 24622 61962
rect 24622 61910 24624 61962
rect 24568 61908 24624 61910
rect 24672 61962 24728 61964
rect 24672 61910 24674 61962
rect 24674 61910 24726 61962
rect 24726 61910 24728 61962
rect 24672 61908 24728 61910
rect 23804 61178 23860 61180
rect 23804 61126 23806 61178
rect 23806 61126 23858 61178
rect 23858 61126 23860 61178
rect 23804 61124 23860 61126
rect 23908 61178 23964 61180
rect 23908 61126 23910 61178
rect 23910 61126 23962 61178
rect 23962 61126 23964 61178
rect 23908 61124 23964 61126
rect 24012 61178 24068 61180
rect 24012 61126 24014 61178
rect 24014 61126 24066 61178
rect 24066 61126 24068 61178
rect 24012 61124 24068 61126
rect 23660 60786 23716 60788
rect 23660 60734 23662 60786
rect 23662 60734 23714 60786
rect 23714 60734 23716 60786
rect 23660 60732 23716 60734
rect 24464 60394 24520 60396
rect 24464 60342 24466 60394
rect 24466 60342 24518 60394
rect 24518 60342 24520 60394
rect 24464 60340 24520 60342
rect 24568 60394 24624 60396
rect 24568 60342 24570 60394
rect 24570 60342 24622 60394
rect 24622 60342 24624 60394
rect 24568 60340 24624 60342
rect 24672 60394 24728 60396
rect 24672 60342 24674 60394
rect 24674 60342 24726 60394
rect 24726 60342 24728 60394
rect 24672 60340 24728 60342
rect 23804 59610 23860 59612
rect 23804 59558 23806 59610
rect 23806 59558 23858 59610
rect 23858 59558 23860 59610
rect 23804 59556 23860 59558
rect 23908 59610 23964 59612
rect 23908 59558 23910 59610
rect 23910 59558 23962 59610
rect 23962 59558 23964 59610
rect 23908 59556 23964 59558
rect 24012 59610 24068 59612
rect 24012 59558 24014 59610
rect 24014 59558 24066 59610
rect 24066 59558 24068 59610
rect 24012 59556 24068 59558
rect 24464 58826 24520 58828
rect 24464 58774 24466 58826
rect 24466 58774 24518 58826
rect 24518 58774 24520 58826
rect 24464 58772 24520 58774
rect 24568 58826 24624 58828
rect 24568 58774 24570 58826
rect 24570 58774 24622 58826
rect 24622 58774 24624 58826
rect 24568 58772 24624 58774
rect 24672 58826 24728 58828
rect 24672 58774 24674 58826
rect 24674 58774 24726 58826
rect 24726 58774 24728 58826
rect 24672 58772 24728 58774
rect 23804 58042 23860 58044
rect 23804 57990 23806 58042
rect 23806 57990 23858 58042
rect 23858 57990 23860 58042
rect 23804 57988 23860 57990
rect 23908 58042 23964 58044
rect 23908 57990 23910 58042
rect 23910 57990 23962 58042
rect 23962 57990 23964 58042
rect 23908 57988 23964 57990
rect 24012 58042 24068 58044
rect 24012 57990 24014 58042
rect 24014 57990 24066 58042
rect 24066 57990 24068 58042
rect 24012 57988 24068 57990
rect 23436 57820 23492 57876
rect 22652 47404 22708 47460
rect 23212 46450 23268 46452
rect 23212 46398 23214 46450
rect 23214 46398 23266 46450
rect 23266 46398 23268 46450
rect 23212 46396 23268 46398
rect 22764 46172 22820 46228
rect 22652 45836 22708 45892
rect 22428 40908 22484 40964
rect 22540 44492 22596 44548
rect 22092 40460 22148 40516
rect 23212 45164 23268 45220
rect 23100 44210 23156 44212
rect 23100 44158 23102 44210
rect 23102 44158 23154 44210
rect 23154 44158 23156 44210
rect 23100 44156 23156 44158
rect 22652 42028 22708 42084
rect 22876 41410 22932 41412
rect 22876 41358 22878 41410
rect 22878 41358 22930 41410
rect 22930 41358 22932 41410
rect 22876 41356 22932 41358
rect 22204 40684 22260 40740
rect 22988 40796 23044 40852
rect 21980 37884 22036 37940
rect 22204 38332 22260 38388
rect 21196 34300 21252 34356
rect 21084 33628 21140 33684
rect 20748 32844 20804 32900
rect 20300 30380 20356 30436
rect 20300 28812 20356 28868
rect 20300 27356 20356 27412
rect 20300 26236 20356 26292
rect 20300 25394 20356 25396
rect 20300 25342 20302 25394
rect 20302 25342 20354 25394
rect 20354 25342 20356 25394
rect 20300 25340 20356 25342
rect 19516 20914 19572 20916
rect 19516 20862 19518 20914
rect 19518 20862 19570 20914
rect 19570 20862 19572 20914
rect 19516 20860 19572 20862
rect 20524 31612 20580 31668
rect 20636 30716 20692 30772
rect 21084 32674 21140 32676
rect 21084 32622 21086 32674
rect 21086 32622 21138 32674
rect 21138 32622 21140 32674
rect 21084 32620 21140 32622
rect 20972 32562 21028 32564
rect 20972 32510 20974 32562
rect 20974 32510 21026 32562
rect 21026 32510 21028 32562
rect 20972 32508 21028 32510
rect 20860 31836 20916 31892
rect 21420 34188 21476 34244
rect 21980 35474 22036 35476
rect 21980 35422 21982 35474
rect 21982 35422 22034 35474
rect 22034 35422 22036 35474
rect 21980 35420 22036 35422
rect 21868 34972 21924 35028
rect 22092 34524 22148 34580
rect 21980 34076 22036 34132
rect 21868 33964 21924 34020
rect 21644 32956 21700 33012
rect 20972 30940 21028 30996
rect 20636 29426 20692 29428
rect 20636 29374 20638 29426
rect 20638 29374 20690 29426
rect 20690 29374 20692 29426
rect 20636 29372 20692 29374
rect 21420 30156 21476 30212
rect 21308 29484 21364 29540
rect 21644 29372 21700 29428
rect 21532 29314 21588 29316
rect 21532 29262 21534 29314
rect 21534 29262 21586 29314
rect 21586 29262 21588 29314
rect 21532 29260 21588 29262
rect 21308 29036 21364 29092
rect 20860 28530 20916 28532
rect 20860 28478 20862 28530
rect 20862 28478 20914 28530
rect 20914 28478 20916 28530
rect 20860 28476 20916 28478
rect 20636 28028 20692 28084
rect 20524 27356 20580 27412
rect 21084 27858 21140 27860
rect 21084 27806 21086 27858
rect 21086 27806 21138 27858
rect 21138 27806 21140 27858
rect 21084 27804 21140 27806
rect 21868 32396 21924 32452
rect 22428 37996 22484 38052
rect 22428 35644 22484 35700
rect 22540 34860 22596 34916
rect 22316 34188 22372 34244
rect 22764 37436 22820 37492
rect 22652 33628 22708 33684
rect 22764 33852 22820 33908
rect 22316 32338 22372 32340
rect 22316 32286 22318 32338
rect 22318 32286 22370 32338
rect 22370 32286 22372 32338
rect 22316 32284 22372 32286
rect 21868 30492 21924 30548
rect 22204 29426 22260 29428
rect 22204 29374 22206 29426
rect 22206 29374 22258 29426
rect 22258 29374 22260 29426
rect 22204 29372 22260 29374
rect 21084 27298 21140 27300
rect 21084 27246 21086 27298
rect 21086 27246 21138 27298
rect 21138 27246 21140 27298
rect 21084 27244 21140 27246
rect 20748 26796 20804 26852
rect 20748 26514 20804 26516
rect 20748 26462 20750 26514
rect 20750 26462 20802 26514
rect 20802 26462 20804 26514
rect 20748 26460 20804 26462
rect 20748 26124 20804 26180
rect 20860 24834 20916 24836
rect 20860 24782 20862 24834
rect 20862 24782 20914 24834
rect 20914 24782 20916 24834
rect 20860 24780 20916 24782
rect 20076 23436 20132 23492
rect 19852 21586 19908 21588
rect 19852 21534 19854 21586
rect 19854 21534 19906 21586
rect 19906 21534 19908 21586
rect 19852 21532 19908 21534
rect 19852 21308 19908 21364
rect 19852 21084 19908 21140
rect 19964 20300 20020 20356
rect 19852 19516 19908 19572
rect 19964 19458 20020 19460
rect 19964 19406 19966 19458
rect 19966 19406 20018 19458
rect 20018 19406 20020 19458
rect 19964 19404 20020 19406
rect 21308 26962 21364 26964
rect 21308 26910 21310 26962
rect 21310 26910 21362 26962
rect 21362 26910 21364 26962
rect 21308 26908 21364 26910
rect 20412 23826 20468 23828
rect 20412 23774 20414 23826
rect 20414 23774 20466 23826
rect 20466 23774 20468 23826
rect 20412 23772 20468 23774
rect 20300 23660 20356 23716
rect 20524 23436 20580 23492
rect 20524 22764 20580 22820
rect 20524 22092 20580 22148
rect 20188 17836 20244 17892
rect 19964 17778 20020 17780
rect 19964 17726 19966 17778
rect 19966 17726 20018 17778
rect 20018 17726 20020 17778
rect 19964 17724 20020 17726
rect 19852 16322 19908 16324
rect 19852 16270 19854 16322
rect 19854 16270 19906 16322
rect 19906 16270 19908 16322
rect 19852 16268 19908 16270
rect 19404 15986 19460 15988
rect 19404 15934 19406 15986
rect 19406 15934 19458 15986
rect 19458 15934 19460 15986
rect 19404 15932 19460 15934
rect 20188 17052 20244 17108
rect 20076 16828 20132 16884
rect 19740 14252 19796 14308
rect 19740 13244 19796 13300
rect 19404 11452 19460 11508
rect 19964 12962 20020 12964
rect 19964 12910 19966 12962
rect 19966 12910 20018 12962
rect 20018 12910 20020 12962
rect 19964 12908 20020 12910
rect 20748 21196 20804 21252
rect 20636 20300 20692 20356
rect 20860 19964 20916 20020
rect 21196 21868 21252 21924
rect 21420 21474 21476 21476
rect 21420 21422 21422 21474
rect 21422 21422 21474 21474
rect 21474 21422 21476 21474
rect 21420 21420 21476 21422
rect 21308 21084 21364 21140
rect 21868 28082 21924 28084
rect 21868 28030 21870 28082
rect 21870 28030 21922 28082
rect 21922 28030 21924 28082
rect 21868 28028 21924 28030
rect 21980 27970 22036 27972
rect 21980 27918 21982 27970
rect 21982 27918 22034 27970
rect 22034 27918 22036 27970
rect 21980 27916 22036 27918
rect 21756 26962 21812 26964
rect 21756 26910 21758 26962
rect 21758 26910 21810 26962
rect 21810 26910 21812 26962
rect 21756 26908 21812 26910
rect 22540 28028 22596 28084
rect 22428 27916 22484 27972
rect 21644 26460 21700 26516
rect 22204 26908 22260 26964
rect 23100 40348 23156 40404
rect 21868 25900 21924 25956
rect 21868 25506 21924 25508
rect 21868 25454 21870 25506
rect 21870 25454 21922 25506
rect 21922 25454 21924 25506
rect 21868 25452 21924 25454
rect 21644 24834 21700 24836
rect 21644 24782 21646 24834
rect 21646 24782 21698 24834
rect 21698 24782 21700 24834
rect 21644 24780 21700 24782
rect 21644 24220 21700 24276
rect 21756 23772 21812 23828
rect 21644 23548 21700 23604
rect 21532 20802 21588 20804
rect 21532 20750 21534 20802
rect 21534 20750 21586 20802
rect 21586 20750 21588 20802
rect 21532 20748 21588 20750
rect 21868 23324 21924 23380
rect 21868 23042 21924 23044
rect 21868 22990 21870 23042
rect 21870 22990 21922 23042
rect 21922 22990 21924 23042
rect 21868 22988 21924 22990
rect 22988 32284 23044 32340
rect 22316 26290 22372 26292
rect 22316 26238 22318 26290
rect 22318 26238 22370 26290
rect 22370 26238 22372 26290
rect 22316 26236 22372 26238
rect 22092 25452 22148 25508
rect 22540 25506 22596 25508
rect 22540 25454 22542 25506
rect 22542 25454 22594 25506
rect 22594 25454 22596 25506
rect 22540 25452 22596 25454
rect 22764 25228 22820 25284
rect 22092 21980 22148 22036
rect 20636 16716 20692 16772
rect 20412 14588 20468 14644
rect 20188 12012 20244 12068
rect 20300 13580 20356 13636
rect 20412 13468 20468 13524
rect 20412 12908 20468 12964
rect 19516 8370 19572 8372
rect 19516 8318 19518 8370
rect 19518 8318 19570 8370
rect 19570 8318 19572 8370
rect 19516 8316 19572 8318
rect 19404 7420 19460 7476
rect 19740 8204 19796 8260
rect 19740 6860 19796 6916
rect 19628 6636 19684 6692
rect 18844 5852 18900 5908
rect 18844 5628 18900 5684
rect 19068 5628 19124 5684
rect 18956 4844 19012 4900
rect 18844 3948 18900 4004
rect 18620 2940 18676 2996
rect 18620 2770 18676 2772
rect 18620 2718 18622 2770
rect 18622 2718 18674 2770
rect 18674 2718 18676 2770
rect 18620 2716 18676 2718
rect 18284 2604 18340 2660
rect 18172 2210 18228 2212
rect 18172 2158 18174 2210
rect 18174 2158 18226 2210
rect 18226 2158 18228 2210
rect 18172 2156 18228 2158
rect 16940 978 16996 980
rect 16940 926 16942 978
rect 16942 926 16994 978
rect 16994 926 16996 978
rect 16940 924 16996 926
rect 17276 924 17332 980
rect 17052 476 17108 532
rect 18620 2268 18676 2324
rect 18396 812 18452 868
rect 17948 588 18004 644
rect 17724 140 17780 196
rect 19404 5516 19460 5572
rect 19740 5404 19796 5460
rect 20076 8818 20132 8820
rect 20076 8766 20078 8818
rect 20078 8766 20130 8818
rect 20130 8766 20132 8818
rect 20076 8764 20132 8766
rect 19964 8204 20020 8260
rect 20076 7756 20132 7812
rect 20076 7084 20132 7140
rect 19964 6860 20020 6916
rect 20412 7532 20468 7588
rect 20524 10556 20580 10612
rect 20972 16492 21028 16548
rect 21644 17052 21700 17108
rect 21196 16492 21252 16548
rect 21196 16044 21252 16100
rect 20748 13634 20804 13636
rect 20748 13582 20750 13634
rect 20750 13582 20802 13634
rect 20802 13582 20804 13634
rect 20748 13580 20804 13582
rect 20748 13244 20804 13300
rect 21980 19404 22036 19460
rect 21532 14700 21588 14756
rect 21196 14476 21252 14532
rect 21532 14364 21588 14420
rect 21308 13468 21364 13524
rect 21196 13244 21252 13300
rect 21196 11228 21252 11284
rect 21196 10556 21252 10612
rect 20748 10498 20804 10500
rect 20748 10446 20750 10498
rect 20750 10446 20802 10498
rect 20802 10446 20804 10498
rect 20748 10444 20804 10446
rect 20636 10332 20692 10388
rect 21084 9660 21140 9716
rect 21308 9660 21364 9716
rect 20860 9042 20916 9044
rect 20860 8990 20862 9042
rect 20862 8990 20914 9042
rect 20914 8990 20916 9042
rect 20860 8988 20916 8990
rect 21196 8540 21252 8596
rect 21084 8092 21140 8148
rect 20748 7756 20804 7812
rect 20188 6524 20244 6580
rect 20300 6972 20356 7028
rect 20524 7308 20580 7364
rect 19964 5852 20020 5908
rect 19292 4338 19348 4340
rect 19292 4286 19294 4338
rect 19294 4286 19346 4338
rect 19346 4286 19348 4338
rect 19292 4284 19348 4286
rect 19404 3388 19460 3444
rect 19292 2546 19348 2548
rect 19292 2494 19294 2546
rect 19294 2494 19346 2546
rect 19346 2494 19348 2546
rect 19292 2492 19348 2494
rect 19852 4956 19908 5012
rect 19628 4396 19684 4452
rect 19964 4844 20020 4900
rect 20636 7084 20692 7140
rect 20524 6748 20580 6804
rect 20412 6578 20468 6580
rect 20412 6526 20414 6578
rect 20414 6526 20466 6578
rect 20466 6526 20468 6578
rect 20412 6524 20468 6526
rect 20412 5516 20468 5572
rect 20076 4620 20132 4676
rect 20300 4620 20356 4676
rect 19628 2940 19684 2996
rect 19852 2492 19908 2548
rect 20188 2380 20244 2436
rect 19852 1708 19908 1764
rect 19964 1820 20020 1876
rect 19292 1260 19348 1316
rect 19964 1260 20020 1316
rect 20412 4284 20468 4340
rect 20748 5516 20804 5572
rect 20524 3612 20580 3668
rect 20860 5404 20916 5460
rect 20748 3164 20804 3220
rect 20860 3052 20916 3108
rect 21756 14476 21812 14532
rect 21756 13634 21812 13636
rect 21756 13582 21758 13634
rect 21758 13582 21810 13634
rect 21810 13582 21812 13634
rect 21756 13580 21812 13582
rect 21532 9660 21588 9716
rect 21644 9996 21700 10052
rect 21644 8988 21700 9044
rect 21644 8764 21700 8820
rect 21420 8146 21476 8148
rect 21420 8094 21422 8146
rect 21422 8094 21474 8146
rect 21474 8094 21476 8146
rect 21420 8092 21476 8094
rect 21420 7532 21476 7588
rect 21420 6636 21476 6692
rect 22428 23154 22484 23156
rect 22428 23102 22430 23154
rect 22430 23102 22482 23154
rect 22482 23102 22484 23154
rect 22428 23100 22484 23102
rect 24464 57258 24520 57260
rect 24464 57206 24466 57258
rect 24466 57206 24518 57258
rect 24518 57206 24520 57258
rect 24464 57204 24520 57206
rect 24568 57258 24624 57260
rect 24568 57206 24570 57258
rect 24570 57206 24622 57258
rect 24622 57206 24624 57258
rect 24568 57204 24624 57206
rect 24672 57258 24728 57260
rect 24672 57206 24674 57258
rect 24674 57206 24726 57258
rect 24726 57206 24728 57258
rect 24672 57204 24728 57206
rect 23804 56474 23860 56476
rect 23804 56422 23806 56474
rect 23806 56422 23858 56474
rect 23858 56422 23860 56474
rect 23804 56420 23860 56422
rect 23908 56474 23964 56476
rect 23908 56422 23910 56474
rect 23910 56422 23962 56474
rect 23962 56422 23964 56474
rect 23908 56420 23964 56422
rect 24012 56474 24068 56476
rect 24012 56422 24014 56474
rect 24014 56422 24066 56474
rect 24066 56422 24068 56474
rect 24012 56420 24068 56422
rect 24464 55690 24520 55692
rect 24464 55638 24466 55690
rect 24466 55638 24518 55690
rect 24518 55638 24520 55690
rect 24464 55636 24520 55638
rect 24568 55690 24624 55692
rect 24568 55638 24570 55690
rect 24570 55638 24622 55690
rect 24622 55638 24624 55690
rect 24568 55636 24624 55638
rect 24672 55690 24728 55692
rect 24672 55638 24674 55690
rect 24674 55638 24726 55690
rect 24726 55638 24728 55690
rect 24672 55636 24728 55638
rect 23660 55132 23716 55188
rect 23548 47964 23604 48020
rect 24780 55186 24836 55188
rect 24780 55134 24782 55186
rect 24782 55134 24834 55186
rect 24834 55134 24836 55186
rect 24780 55132 24836 55134
rect 23804 54906 23860 54908
rect 23804 54854 23806 54906
rect 23806 54854 23858 54906
rect 23858 54854 23860 54906
rect 23804 54852 23860 54854
rect 23908 54906 23964 54908
rect 23908 54854 23910 54906
rect 23910 54854 23962 54906
rect 23962 54854 23964 54906
rect 23908 54852 23964 54854
rect 24012 54906 24068 54908
rect 24012 54854 24014 54906
rect 24014 54854 24066 54906
rect 24066 54854 24068 54906
rect 24012 54852 24068 54854
rect 24464 54122 24520 54124
rect 24464 54070 24466 54122
rect 24466 54070 24518 54122
rect 24518 54070 24520 54122
rect 24464 54068 24520 54070
rect 24568 54122 24624 54124
rect 24568 54070 24570 54122
rect 24570 54070 24622 54122
rect 24622 54070 24624 54122
rect 24568 54068 24624 54070
rect 24672 54122 24728 54124
rect 24672 54070 24674 54122
rect 24674 54070 24726 54122
rect 24726 54070 24728 54122
rect 24672 54068 24728 54070
rect 23804 53338 23860 53340
rect 23804 53286 23806 53338
rect 23806 53286 23858 53338
rect 23858 53286 23860 53338
rect 23804 53284 23860 53286
rect 23908 53338 23964 53340
rect 23908 53286 23910 53338
rect 23910 53286 23962 53338
rect 23962 53286 23964 53338
rect 23908 53284 23964 53286
rect 24012 53338 24068 53340
rect 24012 53286 24014 53338
rect 24014 53286 24066 53338
rect 24066 53286 24068 53338
rect 24012 53284 24068 53286
rect 24464 52554 24520 52556
rect 24464 52502 24466 52554
rect 24466 52502 24518 52554
rect 24518 52502 24520 52554
rect 24464 52500 24520 52502
rect 24568 52554 24624 52556
rect 24568 52502 24570 52554
rect 24570 52502 24622 52554
rect 24622 52502 24624 52554
rect 24568 52500 24624 52502
rect 24672 52554 24728 52556
rect 24672 52502 24674 52554
rect 24674 52502 24726 52554
rect 24726 52502 24728 52554
rect 24672 52500 24728 52502
rect 23804 51770 23860 51772
rect 23804 51718 23806 51770
rect 23806 51718 23858 51770
rect 23858 51718 23860 51770
rect 23804 51716 23860 51718
rect 23908 51770 23964 51772
rect 23908 51718 23910 51770
rect 23910 51718 23962 51770
rect 23962 51718 23964 51770
rect 23908 51716 23964 51718
rect 24012 51770 24068 51772
rect 24012 51718 24014 51770
rect 24014 51718 24066 51770
rect 24066 51718 24068 51770
rect 24012 51716 24068 51718
rect 24464 50986 24520 50988
rect 24464 50934 24466 50986
rect 24466 50934 24518 50986
rect 24518 50934 24520 50986
rect 24464 50932 24520 50934
rect 24568 50986 24624 50988
rect 24568 50934 24570 50986
rect 24570 50934 24622 50986
rect 24622 50934 24624 50986
rect 24568 50932 24624 50934
rect 24672 50986 24728 50988
rect 24672 50934 24674 50986
rect 24674 50934 24726 50986
rect 24726 50934 24728 50986
rect 24672 50932 24728 50934
rect 23804 50202 23860 50204
rect 23804 50150 23806 50202
rect 23806 50150 23858 50202
rect 23858 50150 23860 50202
rect 23804 50148 23860 50150
rect 23908 50202 23964 50204
rect 23908 50150 23910 50202
rect 23910 50150 23962 50202
rect 23962 50150 23964 50202
rect 23908 50148 23964 50150
rect 24012 50202 24068 50204
rect 24012 50150 24014 50202
rect 24014 50150 24066 50202
rect 24066 50150 24068 50202
rect 24012 50148 24068 50150
rect 24464 49418 24520 49420
rect 24464 49366 24466 49418
rect 24466 49366 24518 49418
rect 24518 49366 24520 49418
rect 24464 49364 24520 49366
rect 24568 49418 24624 49420
rect 24568 49366 24570 49418
rect 24570 49366 24622 49418
rect 24622 49366 24624 49418
rect 24568 49364 24624 49366
rect 24672 49418 24728 49420
rect 24672 49366 24674 49418
rect 24674 49366 24726 49418
rect 24726 49366 24728 49418
rect 24672 49364 24728 49366
rect 23804 48634 23860 48636
rect 23804 48582 23806 48634
rect 23806 48582 23858 48634
rect 23858 48582 23860 48634
rect 23804 48580 23860 48582
rect 23908 48634 23964 48636
rect 23908 48582 23910 48634
rect 23910 48582 23962 48634
rect 23962 48582 23964 48634
rect 23908 48580 23964 48582
rect 24012 48634 24068 48636
rect 24012 48582 24014 48634
rect 24014 48582 24066 48634
rect 24066 48582 24068 48634
rect 24012 48580 24068 48582
rect 24464 47850 24520 47852
rect 24464 47798 24466 47850
rect 24466 47798 24518 47850
rect 24518 47798 24520 47850
rect 24464 47796 24520 47798
rect 24568 47850 24624 47852
rect 24568 47798 24570 47850
rect 24570 47798 24622 47850
rect 24622 47798 24624 47850
rect 24568 47796 24624 47798
rect 24672 47850 24728 47852
rect 24672 47798 24674 47850
rect 24674 47798 24726 47850
rect 24726 47798 24728 47850
rect 24672 47796 24728 47798
rect 23804 47066 23860 47068
rect 23804 47014 23806 47066
rect 23806 47014 23858 47066
rect 23858 47014 23860 47066
rect 23804 47012 23860 47014
rect 23908 47066 23964 47068
rect 23908 47014 23910 47066
rect 23910 47014 23962 47066
rect 23962 47014 23964 47066
rect 23908 47012 23964 47014
rect 24012 47066 24068 47068
rect 24012 47014 24014 47066
rect 24014 47014 24066 47066
rect 24066 47014 24068 47066
rect 24012 47012 24068 47014
rect 24464 46282 24520 46284
rect 24464 46230 24466 46282
rect 24466 46230 24518 46282
rect 24518 46230 24520 46282
rect 24464 46228 24520 46230
rect 24568 46282 24624 46284
rect 24568 46230 24570 46282
rect 24570 46230 24622 46282
rect 24622 46230 24624 46282
rect 24568 46228 24624 46230
rect 24672 46282 24728 46284
rect 24672 46230 24674 46282
rect 24674 46230 24726 46282
rect 24726 46230 24728 46282
rect 24672 46228 24728 46230
rect 23804 45498 23860 45500
rect 23804 45446 23806 45498
rect 23806 45446 23858 45498
rect 23858 45446 23860 45498
rect 23804 45444 23860 45446
rect 23908 45498 23964 45500
rect 23908 45446 23910 45498
rect 23910 45446 23962 45498
rect 23962 45446 23964 45498
rect 23908 45444 23964 45446
rect 24012 45498 24068 45500
rect 24012 45446 24014 45498
rect 24014 45446 24066 45498
rect 24066 45446 24068 45498
rect 24012 45444 24068 45446
rect 25004 79548 25060 79604
rect 25004 62300 25060 62356
rect 25116 63868 25172 63924
rect 25116 57484 25172 57540
rect 24892 45276 24948 45332
rect 25004 53004 25060 53060
rect 24464 44714 24520 44716
rect 24464 44662 24466 44714
rect 24466 44662 24518 44714
rect 24518 44662 24520 44714
rect 24464 44660 24520 44662
rect 24568 44714 24624 44716
rect 24568 44662 24570 44714
rect 24570 44662 24622 44714
rect 24622 44662 24624 44714
rect 24568 44660 24624 44662
rect 24672 44714 24728 44716
rect 24672 44662 24674 44714
rect 24674 44662 24726 44714
rect 24726 44662 24728 44714
rect 24672 44660 24728 44662
rect 23804 43930 23860 43932
rect 23804 43878 23806 43930
rect 23806 43878 23858 43930
rect 23858 43878 23860 43930
rect 23804 43876 23860 43878
rect 23908 43930 23964 43932
rect 23908 43878 23910 43930
rect 23910 43878 23962 43930
rect 23962 43878 23964 43930
rect 23908 43876 23964 43878
rect 24012 43930 24068 43932
rect 24012 43878 24014 43930
rect 24014 43878 24066 43930
rect 24066 43878 24068 43930
rect 24012 43876 24068 43878
rect 24464 43146 24520 43148
rect 24464 43094 24466 43146
rect 24466 43094 24518 43146
rect 24518 43094 24520 43146
rect 24464 43092 24520 43094
rect 24568 43146 24624 43148
rect 24568 43094 24570 43146
rect 24570 43094 24622 43146
rect 24622 43094 24624 43146
rect 24568 43092 24624 43094
rect 24672 43146 24728 43148
rect 24672 43094 24674 43146
rect 24674 43094 24726 43146
rect 24726 43094 24728 43146
rect 24672 43092 24728 43094
rect 23804 42362 23860 42364
rect 23804 42310 23806 42362
rect 23806 42310 23858 42362
rect 23858 42310 23860 42362
rect 23804 42308 23860 42310
rect 23908 42362 23964 42364
rect 23908 42310 23910 42362
rect 23910 42310 23962 42362
rect 23962 42310 23964 42362
rect 23908 42308 23964 42310
rect 24012 42362 24068 42364
rect 24012 42310 24014 42362
rect 24014 42310 24066 42362
rect 24066 42310 24068 42362
rect 24012 42308 24068 42310
rect 23660 41580 23716 41636
rect 24464 41578 24520 41580
rect 24464 41526 24466 41578
rect 24466 41526 24518 41578
rect 24518 41526 24520 41578
rect 24464 41524 24520 41526
rect 24568 41578 24624 41580
rect 24568 41526 24570 41578
rect 24570 41526 24622 41578
rect 24622 41526 24624 41578
rect 24568 41524 24624 41526
rect 24672 41578 24728 41580
rect 24672 41526 24674 41578
rect 24674 41526 24726 41578
rect 24726 41526 24728 41578
rect 24672 41524 24728 41526
rect 23772 41132 23828 41188
rect 23804 40794 23860 40796
rect 23804 40742 23806 40794
rect 23806 40742 23858 40794
rect 23858 40742 23860 40794
rect 23804 40740 23860 40742
rect 23908 40794 23964 40796
rect 23908 40742 23910 40794
rect 23910 40742 23962 40794
rect 23962 40742 23964 40794
rect 23908 40740 23964 40742
rect 24012 40794 24068 40796
rect 24012 40742 24014 40794
rect 24014 40742 24066 40794
rect 24066 40742 24068 40794
rect 24012 40740 24068 40742
rect 23660 40402 23716 40404
rect 23660 40350 23662 40402
rect 23662 40350 23714 40402
rect 23714 40350 23716 40402
rect 23660 40348 23716 40350
rect 24464 40010 24520 40012
rect 24464 39958 24466 40010
rect 24466 39958 24518 40010
rect 24518 39958 24520 40010
rect 24464 39956 24520 39958
rect 24568 40010 24624 40012
rect 24568 39958 24570 40010
rect 24570 39958 24622 40010
rect 24622 39958 24624 40010
rect 24568 39956 24624 39958
rect 24672 40010 24728 40012
rect 24672 39958 24674 40010
rect 24674 39958 24726 40010
rect 24726 39958 24728 40010
rect 24672 39956 24728 39958
rect 23804 39226 23860 39228
rect 23804 39174 23806 39226
rect 23806 39174 23858 39226
rect 23858 39174 23860 39226
rect 23804 39172 23860 39174
rect 23908 39226 23964 39228
rect 23908 39174 23910 39226
rect 23910 39174 23962 39226
rect 23962 39174 23964 39226
rect 23908 39172 23964 39174
rect 24012 39226 24068 39228
rect 24012 39174 24014 39226
rect 24014 39174 24066 39226
rect 24066 39174 24068 39226
rect 24012 39172 24068 39174
rect 23212 31890 23268 31892
rect 23212 31838 23214 31890
rect 23214 31838 23266 31890
rect 23266 31838 23268 31890
rect 23212 31836 23268 31838
rect 23212 29036 23268 29092
rect 22764 22652 22820 22708
rect 22540 22316 22596 22372
rect 24464 38442 24520 38444
rect 24464 38390 24466 38442
rect 24466 38390 24518 38442
rect 24518 38390 24520 38442
rect 24464 38388 24520 38390
rect 24568 38442 24624 38444
rect 24568 38390 24570 38442
rect 24570 38390 24622 38442
rect 24622 38390 24624 38442
rect 24568 38388 24624 38390
rect 24672 38442 24728 38444
rect 24672 38390 24674 38442
rect 24674 38390 24726 38442
rect 24726 38390 24728 38442
rect 24672 38388 24728 38390
rect 24332 38220 24388 38276
rect 23804 37658 23860 37660
rect 23804 37606 23806 37658
rect 23806 37606 23858 37658
rect 23858 37606 23860 37658
rect 23804 37604 23860 37606
rect 23908 37658 23964 37660
rect 23908 37606 23910 37658
rect 23910 37606 23962 37658
rect 23962 37606 23964 37658
rect 23908 37604 23964 37606
rect 24012 37658 24068 37660
rect 24012 37606 24014 37658
rect 24014 37606 24066 37658
rect 24066 37606 24068 37658
rect 24012 37604 24068 37606
rect 23996 36594 24052 36596
rect 23996 36542 23998 36594
rect 23998 36542 24050 36594
rect 24050 36542 24052 36594
rect 23996 36540 24052 36542
rect 23804 36090 23860 36092
rect 23804 36038 23806 36090
rect 23806 36038 23858 36090
rect 23858 36038 23860 36090
rect 23804 36036 23860 36038
rect 23908 36090 23964 36092
rect 23908 36038 23910 36090
rect 23910 36038 23962 36090
rect 23962 36038 23964 36090
rect 23908 36036 23964 36038
rect 24012 36090 24068 36092
rect 24012 36038 24014 36090
rect 24014 36038 24066 36090
rect 24066 36038 24068 36090
rect 24012 36036 24068 36038
rect 23436 34860 23492 34916
rect 23804 34522 23860 34524
rect 23804 34470 23806 34522
rect 23806 34470 23858 34522
rect 23858 34470 23860 34522
rect 23804 34468 23860 34470
rect 23908 34522 23964 34524
rect 23908 34470 23910 34522
rect 23910 34470 23962 34522
rect 23962 34470 23964 34522
rect 23908 34468 23964 34470
rect 24012 34522 24068 34524
rect 24012 34470 24014 34522
rect 24014 34470 24066 34522
rect 24066 34470 24068 34522
rect 24012 34468 24068 34470
rect 23772 33404 23828 33460
rect 23804 32954 23860 32956
rect 23804 32902 23806 32954
rect 23806 32902 23858 32954
rect 23858 32902 23860 32954
rect 23804 32900 23860 32902
rect 23908 32954 23964 32956
rect 23908 32902 23910 32954
rect 23910 32902 23962 32954
rect 23962 32902 23964 32954
rect 23908 32900 23964 32902
rect 24012 32954 24068 32956
rect 24012 32902 24014 32954
rect 24014 32902 24066 32954
rect 24066 32902 24068 32954
rect 24012 32900 24068 32902
rect 23660 32732 23716 32788
rect 23804 31386 23860 31388
rect 23804 31334 23806 31386
rect 23806 31334 23858 31386
rect 23858 31334 23860 31386
rect 23804 31332 23860 31334
rect 23908 31386 23964 31388
rect 23908 31334 23910 31386
rect 23910 31334 23962 31386
rect 23962 31334 23964 31386
rect 23908 31332 23964 31334
rect 24012 31386 24068 31388
rect 24012 31334 24014 31386
rect 24014 31334 24066 31386
rect 24066 31334 24068 31386
rect 24012 31332 24068 31334
rect 23804 29818 23860 29820
rect 23804 29766 23806 29818
rect 23806 29766 23858 29818
rect 23858 29766 23860 29818
rect 23804 29764 23860 29766
rect 23908 29818 23964 29820
rect 23908 29766 23910 29818
rect 23910 29766 23962 29818
rect 23962 29766 23964 29818
rect 23908 29764 23964 29766
rect 24012 29818 24068 29820
rect 24012 29766 24014 29818
rect 24014 29766 24066 29818
rect 24066 29766 24068 29818
rect 24012 29764 24068 29766
rect 23804 28250 23860 28252
rect 23804 28198 23806 28250
rect 23806 28198 23858 28250
rect 23858 28198 23860 28250
rect 23804 28196 23860 28198
rect 23908 28250 23964 28252
rect 23908 28198 23910 28250
rect 23910 28198 23962 28250
rect 23962 28198 23964 28250
rect 23908 28196 23964 28198
rect 24012 28250 24068 28252
rect 24012 28198 24014 28250
rect 24014 28198 24066 28250
rect 24066 28198 24068 28250
rect 24012 28196 24068 28198
rect 23212 23548 23268 23604
rect 23804 26682 23860 26684
rect 23804 26630 23806 26682
rect 23806 26630 23858 26682
rect 23858 26630 23860 26682
rect 23804 26628 23860 26630
rect 23908 26682 23964 26684
rect 23908 26630 23910 26682
rect 23910 26630 23962 26682
rect 23962 26630 23964 26682
rect 23908 26628 23964 26630
rect 24012 26682 24068 26684
rect 24012 26630 24014 26682
rect 24014 26630 24066 26682
rect 24066 26630 24068 26682
rect 24012 26628 24068 26630
rect 23804 25114 23860 25116
rect 23804 25062 23806 25114
rect 23806 25062 23858 25114
rect 23858 25062 23860 25114
rect 23804 25060 23860 25062
rect 23908 25114 23964 25116
rect 23908 25062 23910 25114
rect 23910 25062 23962 25114
rect 23962 25062 23964 25114
rect 23908 25060 23964 25062
rect 24012 25114 24068 25116
rect 24012 25062 24014 25114
rect 24014 25062 24066 25114
rect 24066 25062 24068 25114
rect 24012 25060 24068 25062
rect 23804 23546 23860 23548
rect 23804 23494 23806 23546
rect 23806 23494 23858 23546
rect 23858 23494 23860 23546
rect 23804 23492 23860 23494
rect 23908 23546 23964 23548
rect 23908 23494 23910 23546
rect 23910 23494 23962 23546
rect 23962 23494 23964 23546
rect 23908 23492 23964 23494
rect 24012 23546 24068 23548
rect 24012 23494 24014 23546
rect 24014 23494 24066 23546
rect 24066 23494 24068 23546
rect 24012 23492 24068 23494
rect 23212 23154 23268 23156
rect 23212 23102 23214 23154
rect 23214 23102 23266 23154
rect 23266 23102 23268 23154
rect 23212 23100 23268 23102
rect 22988 22988 23044 23044
rect 23100 22876 23156 22932
rect 22540 21810 22596 21812
rect 22540 21758 22542 21810
rect 22542 21758 22594 21810
rect 22594 21758 22596 21810
rect 22540 21756 22596 21758
rect 23212 22764 23268 22820
rect 23436 23100 23492 23156
rect 23548 22652 23604 22708
rect 23324 21756 23380 21812
rect 22764 21532 22820 21588
rect 24108 22930 24164 22932
rect 24108 22878 24110 22930
rect 24110 22878 24162 22930
rect 24162 22878 24164 22930
rect 24108 22876 24164 22878
rect 23772 22258 23828 22260
rect 23772 22206 23774 22258
rect 23774 22206 23826 22258
rect 23826 22206 23828 22258
rect 23772 22204 23828 22206
rect 24220 22092 24276 22148
rect 23804 21978 23860 21980
rect 23804 21926 23806 21978
rect 23806 21926 23858 21978
rect 23858 21926 23860 21978
rect 23804 21924 23860 21926
rect 23908 21978 23964 21980
rect 23908 21926 23910 21978
rect 23910 21926 23962 21978
rect 23962 21926 23964 21978
rect 23908 21924 23964 21926
rect 24012 21978 24068 21980
rect 24012 21926 24014 21978
rect 24014 21926 24066 21978
rect 24066 21926 24068 21978
rect 24012 21924 24068 21926
rect 21868 12908 21924 12964
rect 21868 11788 21924 11844
rect 22204 14700 22260 14756
rect 22316 13916 22372 13972
rect 22092 13580 22148 13636
rect 22540 13074 22596 13076
rect 22540 13022 22542 13074
rect 22542 13022 22594 13074
rect 22594 13022 22596 13074
rect 22540 13020 22596 13022
rect 22428 12178 22484 12180
rect 22428 12126 22430 12178
rect 22430 12126 22482 12178
rect 22482 12126 22484 12178
rect 22428 12124 22484 12126
rect 21980 9324 22036 9380
rect 21868 9212 21924 9268
rect 21756 8540 21812 8596
rect 21868 8988 21924 9044
rect 21756 7980 21812 8036
rect 21756 6076 21812 6132
rect 22428 9996 22484 10052
rect 23212 19852 23268 19908
rect 23100 16098 23156 16100
rect 23100 16046 23102 16098
rect 23102 16046 23154 16098
rect 23154 16046 23156 16098
rect 23100 16044 23156 16046
rect 22988 12124 23044 12180
rect 22764 9324 22820 9380
rect 22428 9266 22484 9268
rect 22428 9214 22430 9266
rect 22430 9214 22482 9266
rect 22482 9214 22484 9266
rect 22428 9212 22484 9214
rect 22316 9100 22372 9156
rect 22092 6690 22148 6692
rect 22092 6638 22094 6690
rect 22094 6638 22146 6690
rect 22146 6638 22148 6690
rect 22092 6636 22148 6638
rect 22204 6412 22260 6468
rect 21532 4508 21588 4564
rect 21868 5852 21924 5908
rect 21196 4060 21252 4116
rect 21196 3836 21252 3892
rect 21420 4060 21476 4116
rect 20972 2716 21028 2772
rect 21084 3500 21140 3556
rect 20860 1932 20916 1988
rect 19740 364 19796 420
rect 19964 252 20020 308
rect 20636 252 20692 308
rect 20972 1708 21028 1764
rect 21420 2828 21476 2884
rect 21420 2492 21476 2548
rect 21868 4172 21924 4228
rect 21756 2716 21812 2772
rect 21532 1484 21588 1540
rect 21868 2156 21924 2212
rect 21756 1202 21812 1204
rect 21756 1150 21758 1202
rect 21758 1150 21810 1202
rect 21810 1150 21812 1202
rect 21756 1148 21812 1150
rect 22092 2210 22148 2212
rect 22092 2158 22094 2210
rect 22094 2158 22146 2210
rect 22146 2158 22148 2210
rect 22092 2156 22148 2158
rect 22316 5906 22372 5908
rect 22316 5854 22318 5906
rect 22318 5854 22370 5906
rect 22370 5854 22372 5906
rect 22316 5852 22372 5854
rect 22316 5404 22372 5460
rect 22428 5292 22484 5348
rect 22428 5122 22484 5124
rect 22428 5070 22430 5122
rect 22430 5070 22482 5122
rect 22482 5070 22484 5122
rect 22428 5068 22484 5070
rect 22876 7868 22932 7924
rect 22876 6972 22932 7028
rect 22988 6636 23044 6692
rect 22876 6524 22932 6580
rect 22988 6188 23044 6244
rect 22988 4956 23044 5012
rect 22764 4620 22820 4676
rect 22988 4732 23044 4788
rect 22428 4284 22484 4340
rect 22316 2770 22372 2772
rect 22316 2718 22318 2770
rect 22318 2718 22370 2770
rect 22370 2718 22372 2770
rect 22316 2716 22372 2718
rect 22316 476 22372 532
rect 22540 3836 22596 3892
rect 22876 3724 22932 3780
rect 22988 3164 23044 3220
rect 22876 2380 22932 2436
rect 22652 2156 22708 2212
rect 22540 1596 22596 1652
rect 22988 978 23044 980
rect 22988 926 22990 978
rect 22990 926 23042 978
rect 23042 926 23044 978
rect 22988 924 23044 926
rect 23804 20410 23860 20412
rect 23804 20358 23806 20410
rect 23806 20358 23858 20410
rect 23858 20358 23860 20410
rect 23804 20356 23860 20358
rect 23908 20410 23964 20412
rect 23908 20358 23910 20410
rect 23910 20358 23962 20410
rect 23962 20358 23964 20410
rect 23908 20356 23964 20358
rect 24012 20410 24068 20412
rect 24012 20358 24014 20410
rect 24014 20358 24066 20410
rect 24066 20358 24068 20410
rect 24012 20356 24068 20358
rect 23804 18842 23860 18844
rect 23804 18790 23806 18842
rect 23806 18790 23858 18842
rect 23858 18790 23860 18842
rect 23804 18788 23860 18790
rect 23908 18842 23964 18844
rect 23908 18790 23910 18842
rect 23910 18790 23962 18842
rect 23962 18790 23964 18842
rect 23908 18788 23964 18790
rect 24012 18842 24068 18844
rect 24012 18790 24014 18842
rect 24014 18790 24066 18842
rect 24066 18790 24068 18842
rect 24012 18788 24068 18790
rect 23436 15260 23492 15316
rect 23660 18620 23716 18676
rect 23804 17274 23860 17276
rect 23804 17222 23806 17274
rect 23806 17222 23858 17274
rect 23858 17222 23860 17274
rect 23804 17220 23860 17222
rect 23908 17274 23964 17276
rect 23908 17222 23910 17274
rect 23910 17222 23962 17274
rect 23962 17222 23964 17274
rect 23908 17220 23964 17222
rect 24012 17274 24068 17276
rect 24012 17222 24014 17274
rect 24014 17222 24066 17274
rect 24066 17222 24068 17274
rect 24012 17220 24068 17222
rect 23804 15706 23860 15708
rect 23804 15654 23806 15706
rect 23806 15654 23858 15706
rect 23858 15654 23860 15706
rect 23804 15652 23860 15654
rect 23908 15706 23964 15708
rect 23908 15654 23910 15706
rect 23910 15654 23962 15706
rect 23962 15654 23964 15706
rect 23908 15652 23964 15654
rect 24012 15706 24068 15708
rect 24012 15654 24014 15706
rect 24014 15654 24066 15706
rect 24066 15654 24068 15706
rect 24012 15652 24068 15654
rect 23804 14138 23860 14140
rect 23804 14086 23806 14138
rect 23806 14086 23858 14138
rect 23858 14086 23860 14138
rect 23804 14084 23860 14086
rect 23908 14138 23964 14140
rect 23908 14086 23910 14138
rect 23910 14086 23962 14138
rect 23962 14086 23964 14138
rect 23908 14084 23964 14086
rect 24012 14138 24068 14140
rect 24012 14086 24014 14138
rect 24014 14086 24066 14138
rect 24066 14086 24068 14138
rect 24012 14084 24068 14086
rect 23804 12570 23860 12572
rect 23804 12518 23806 12570
rect 23806 12518 23858 12570
rect 23858 12518 23860 12570
rect 23804 12516 23860 12518
rect 23908 12570 23964 12572
rect 23908 12518 23910 12570
rect 23910 12518 23962 12570
rect 23962 12518 23964 12570
rect 23908 12516 23964 12518
rect 24012 12570 24068 12572
rect 24012 12518 24014 12570
rect 24014 12518 24066 12570
rect 24066 12518 24068 12570
rect 24012 12516 24068 12518
rect 23212 6412 23268 6468
rect 23660 11340 23716 11396
rect 23804 11002 23860 11004
rect 23804 10950 23806 11002
rect 23806 10950 23858 11002
rect 23858 10950 23860 11002
rect 23804 10948 23860 10950
rect 23908 11002 23964 11004
rect 23908 10950 23910 11002
rect 23910 10950 23962 11002
rect 23962 10950 23964 11002
rect 23908 10948 23964 10950
rect 24012 11002 24068 11004
rect 24012 10950 24014 11002
rect 24014 10950 24066 11002
rect 24066 10950 24068 11002
rect 24012 10948 24068 10950
rect 23804 9434 23860 9436
rect 23804 9382 23806 9434
rect 23806 9382 23858 9434
rect 23858 9382 23860 9434
rect 23804 9380 23860 9382
rect 23908 9434 23964 9436
rect 23908 9382 23910 9434
rect 23910 9382 23962 9434
rect 23962 9382 23964 9434
rect 23908 9380 23964 9382
rect 24012 9434 24068 9436
rect 24012 9382 24014 9434
rect 24014 9382 24066 9434
rect 24066 9382 24068 9434
rect 24012 9380 24068 9382
rect 24108 8930 24164 8932
rect 24108 8878 24110 8930
rect 24110 8878 24162 8930
rect 24162 8878 24164 8930
rect 24108 8876 24164 8878
rect 23212 5964 23268 6020
rect 23324 5346 23380 5348
rect 23324 5294 23326 5346
rect 23326 5294 23378 5346
rect 23378 5294 23380 5346
rect 23324 5292 23380 5294
rect 23436 5068 23492 5124
rect 23548 8092 23604 8148
rect 23436 4620 23492 4676
rect 23212 2098 23268 2100
rect 23212 2046 23214 2098
rect 23214 2046 23266 2098
rect 23266 2046 23268 2098
rect 23212 2044 23268 2046
rect 23804 7866 23860 7868
rect 23660 7756 23716 7812
rect 23804 7814 23806 7866
rect 23806 7814 23858 7866
rect 23858 7814 23860 7866
rect 23804 7812 23860 7814
rect 23908 7866 23964 7868
rect 23908 7814 23910 7866
rect 23910 7814 23962 7866
rect 23962 7814 23964 7866
rect 23908 7812 23964 7814
rect 24012 7866 24068 7868
rect 24012 7814 24014 7866
rect 24014 7814 24066 7866
rect 24066 7814 24068 7866
rect 24012 7812 24068 7814
rect 23660 7532 23716 7588
rect 23804 6298 23860 6300
rect 23804 6246 23806 6298
rect 23806 6246 23858 6298
rect 23858 6246 23860 6298
rect 23804 6244 23860 6246
rect 23908 6298 23964 6300
rect 23908 6246 23910 6298
rect 23910 6246 23962 6298
rect 23962 6246 23964 6298
rect 23908 6244 23964 6246
rect 24012 6298 24068 6300
rect 24012 6246 24014 6298
rect 24014 6246 24066 6298
rect 24066 6246 24068 6298
rect 24012 6244 24068 6246
rect 24108 6076 24164 6132
rect 23996 5346 24052 5348
rect 23996 5294 23998 5346
rect 23998 5294 24050 5346
rect 24050 5294 24052 5346
rect 23996 5292 24052 5294
rect 23804 4730 23860 4732
rect 23804 4678 23806 4730
rect 23806 4678 23858 4730
rect 23858 4678 23860 4730
rect 23804 4676 23860 4678
rect 23908 4730 23964 4732
rect 23908 4678 23910 4730
rect 23910 4678 23962 4730
rect 23962 4678 23964 4730
rect 23908 4676 23964 4678
rect 24012 4730 24068 4732
rect 24012 4678 24014 4730
rect 24014 4678 24066 4730
rect 24066 4678 24068 4730
rect 24012 4676 24068 4678
rect 23660 4396 23716 4452
rect 23772 4284 23828 4340
rect 23548 3778 23604 3780
rect 23548 3726 23550 3778
rect 23550 3726 23602 3778
rect 23602 3726 23604 3778
rect 23548 3724 23604 3726
rect 24108 4226 24164 4228
rect 24108 4174 24110 4226
rect 24110 4174 24162 4226
rect 24162 4174 24164 4226
rect 24108 4172 24164 4174
rect 23772 3500 23828 3556
rect 23884 3276 23940 3332
rect 23804 3162 23860 3164
rect 23804 3110 23806 3162
rect 23806 3110 23858 3162
rect 23858 3110 23860 3162
rect 23804 3108 23860 3110
rect 23908 3162 23964 3164
rect 23908 3110 23910 3162
rect 23910 3110 23962 3162
rect 23962 3110 23964 3162
rect 23908 3108 23964 3110
rect 24012 3162 24068 3164
rect 24012 3110 24014 3162
rect 24014 3110 24066 3162
rect 24066 3110 24068 3162
rect 24012 3108 24068 3110
rect 23660 2940 23716 2996
rect 24108 2546 24164 2548
rect 24108 2494 24110 2546
rect 24110 2494 24162 2546
rect 24162 2494 24164 2546
rect 24108 2492 24164 2494
rect 23660 2380 23716 2436
rect 23804 1594 23860 1596
rect 23804 1542 23806 1594
rect 23806 1542 23858 1594
rect 23858 1542 23860 1594
rect 23804 1540 23860 1542
rect 23908 1594 23964 1596
rect 23908 1542 23910 1594
rect 23910 1542 23962 1594
rect 23962 1542 23964 1594
rect 23908 1540 23964 1542
rect 24012 1594 24068 1596
rect 24012 1542 24014 1594
rect 24014 1542 24066 1594
rect 24066 1542 24068 1594
rect 24012 1540 24068 1542
rect 23772 1372 23828 1428
rect 24464 36874 24520 36876
rect 24464 36822 24466 36874
rect 24466 36822 24518 36874
rect 24518 36822 24520 36874
rect 24464 36820 24520 36822
rect 24568 36874 24624 36876
rect 24568 36822 24570 36874
rect 24570 36822 24622 36874
rect 24622 36822 24624 36874
rect 24568 36820 24624 36822
rect 24672 36874 24728 36876
rect 24672 36822 24674 36874
rect 24674 36822 24726 36874
rect 24726 36822 24728 36874
rect 24672 36820 24728 36822
rect 24464 35306 24520 35308
rect 24464 35254 24466 35306
rect 24466 35254 24518 35306
rect 24518 35254 24520 35306
rect 24464 35252 24520 35254
rect 24568 35306 24624 35308
rect 24568 35254 24570 35306
rect 24570 35254 24622 35306
rect 24622 35254 24624 35306
rect 24568 35252 24624 35254
rect 24672 35306 24728 35308
rect 24672 35254 24674 35306
rect 24674 35254 24726 35306
rect 24726 35254 24728 35306
rect 24672 35252 24728 35254
rect 24780 35026 24836 35028
rect 24780 34974 24782 35026
rect 24782 34974 24834 35026
rect 24834 34974 24836 35026
rect 24780 34972 24836 34974
rect 24668 34914 24724 34916
rect 24668 34862 24670 34914
rect 24670 34862 24722 34914
rect 24722 34862 24724 34914
rect 24668 34860 24724 34862
rect 24668 34018 24724 34020
rect 24668 33966 24670 34018
rect 24670 33966 24722 34018
rect 24722 33966 24724 34018
rect 24668 33964 24724 33966
rect 24464 33738 24520 33740
rect 24464 33686 24466 33738
rect 24466 33686 24518 33738
rect 24518 33686 24520 33738
rect 24464 33684 24520 33686
rect 24568 33738 24624 33740
rect 24568 33686 24570 33738
rect 24570 33686 24622 33738
rect 24622 33686 24624 33738
rect 24568 33684 24624 33686
rect 24672 33738 24728 33740
rect 24672 33686 24674 33738
rect 24674 33686 24726 33738
rect 24726 33686 24728 33738
rect 24672 33684 24728 33686
rect 24464 32170 24520 32172
rect 24464 32118 24466 32170
rect 24466 32118 24518 32170
rect 24518 32118 24520 32170
rect 24464 32116 24520 32118
rect 24568 32170 24624 32172
rect 24568 32118 24570 32170
rect 24570 32118 24622 32170
rect 24622 32118 24624 32170
rect 24568 32116 24624 32118
rect 24672 32170 24728 32172
rect 24672 32118 24674 32170
rect 24674 32118 24726 32170
rect 24726 32118 24728 32170
rect 24672 32116 24728 32118
rect 24892 31836 24948 31892
rect 24464 30602 24520 30604
rect 24464 30550 24466 30602
rect 24466 30550 24518 30602
rect 24518 30550 24520 30602
rect 24464 30548 24520 30550
rect 24568 30602 24624 30604
rect 24568 30550 24570 30602
rect 24570 30550 24622 30602
rect 24622 30550 24624 30602
rect 24568 30548 24624 30550
rect 24672 30602 24728 30604
rect 24672 30550 24674 30602
rect 24674 30550 24726 30602
rect 24726 30550 24728 30602
rect 24672 30548 24728 30550
rect 24464 29034 24520 29036
rect 24464 28982 24466 29034
rect 24466 28982 24518 29034
rect 24518 28982 24520 29034
rect 24464 28980 24520 28982
rect 24568 29034 24624 29036
rect 24568 28982 24570 29034
rect 24570 28982 24622 29034
rect 24622 28982 24624 29034
rect 24568 28980 24624 28982
rect 24672 29034 24728 29036
rect 24672 28982 24674 29034
rect 24674 28982 24726 29034
rect 24726 28982 24728 29034
rect 24672 28980 24728 28982
rect 24464 27466 24520 27468
rect 24464 27414 24466 27466
rect 24466 27414 24518 27466
rect 24518 27414 24520 27466
rect 24464 27412 24520 27414
rect 24568 27466 24624 27468
rect 24568 27414 24570 27466
rect 24570 27414 24622 27466
rect 24622 27414 24624 27466
rect 24568 27412 24624 27414
rect 24672 27466 24728 27468
rect 24672 27414 24674 27466
rect 24674 27414 24726 27466
rect 24726 27414 24728 27466
rect 24672 27412 24728 27414
rect 24464 25898 24520 25900
rect 24464 25846 24466 25898
rect 24466 25846 24518 25898
rect 24518 25846 24520 25898
rect 24464 25844 24520 25846
rect 24568 25898 24624 25900
rect 24568 25846 24570 25898
rect 24570 25846 24622 25898
rect 24622 25846 24624 25898
rect 24568 25844 24624 25846
rect 24672 25898 24728 25900
rect 24672 25846 24674 25898
rect 24674 25846 24726 25898
rect 24726 25846 24728 25898
rect 24672 25844 24728 25846
rect 24464 24330 24520 24332
rect 24464 24278 24466 24330
rect 24466 24278 24518 24330
rect 24518 24278 24520 24330
rect 24464 24276 24520 24278
rect 24568 24330 24624 24332
rect 24568 24278 24570 24330
rect 24570 24278 24622 24330
rect 24622 24278 24624 24330
rect 24568 24276 24624 24278
rect 24672 24330 24728 24332
rect 24672 24278 24674 24330
rect 24674 24278 24726 24330
rect 24726 24278 24728 24330
rect 24672 24276 24728 24278
rect 24464 22762 24520 22764
rect 24464 22710 24466 22762
rect 24466 22710 24518 22762
rect 24518 22710 24520 22762
rect 24464 22708 24520 22710
rect 24568 22762 24624 22764
rect 24568 22710 24570 22762
rect 24570 22710 24622 22762
rect 24622 22710 24624 22762
rect 24568 22708 24624 22710
rect 24672 22762 24728 22764
rect 24672 22710 24674 22762
rect 24674 22710 24726 22762
rect 24726 22710 24728 22762
rect 24672 22708 24728 22710
rect 24464 21194 24520 21196
rect 24464 21142 24466 21194
rect 24466 21142 24518 21194
rect 24518 21142 24520 21194
rect 24464 21140 24520 21142
rect 24568 21194 24624 21196
rect 24568 21142 24570 21194
rect 24570 21142 24622 21194
rect 24622 21142 24624 21194
rect 24568 21140 24624 21142
rect 24672 21194 24728 21196
rect 24672 21142 24674 21194
rect 24674 21142 24726 21194
rect 24726 21142 24728 21194
rect 24672 21140 24728 21142
rect 24464 19626 24520 19628
rect 24464 19574 24466 19626
rect 24466 19574 24518 19626
rect 24518 19574 24520 19626
rect 24464 19572 24520 19574
rect 24568 19626 24624 19628
rect 24568 19574 24570 19626
rect 24570 19574 24622 19626
rect 24622 19574 24624 19626
rect 24568 19572 24624 19574
rect 24672 19626 24728 19628
rect 24672 19574 24674 19626
rect 24674 19574 24726 19626
rect 24726 19574 24728 19626
rect 24672 19572 24728 19574
rect 25004 18396 25060 18452
rect 24464 18058 24520 18060
rect 24464 18006 24466 18058
rect 24466 18006 24518 18058
rect 24518 18006 24520 18058
rect 24464 18004 24520 18006
rect 24568 18058 24624 18060
rect 24568 18006 24570 18058
rect 24570 18006 24622 18058
rect 24622 18006 24624 18058
rect 24568 18004 24624 18006
rect 24672 18058 24728 18060
rect 24672 18006 24674 18058
rect 24674 18006 24726 18058
rect 24726 18006 24728 18058
rect 24672 18004 24728 18006
rect 24892 16716 24948 16772
rect 24464 16490 24520 16492
rect 24464 16438 24466 16490
rect 24466 16438 24518 16490
rect 24518 16438 24520 16490
rect 24464 16436 24520 16438
rect 24568 16490 24624 16492
rect 24568 16438 24570 16490
rect 24570 16438 24622 16490
rect 24622 16438 24624 16490
rect 24568 16436 24624 16438
rect 24672 16490 24728 16492
rect 24672 16438 24674 16490
rect 24674 16438 24726 16490
rect 24726 16438 24728 16490
rect 24672 16436 24728 16438
rect 24464 14922 24520 14924
rect 24464 14870 24466 14922
rect 24466 14870 24518 14922
rect 24518 14870 24520 14922
rect 24464 14868 24520 14870
rect 24568 14922 24624 14924
rect 24568 14870 24570 14922
rect 24570 14870 24622 14922
rect 24622 14870 24624 14922
rect 24568 14868 24624 14870
rect 24672 14922 24728 14924
rect 24672 14870 24674 14922
rect 24674 14870 24726 14922
rect 24726 14870 24728 14922
rect 24672 14868 24728 14870
rect 26012 111746 26068 111748
rect 26012 111694 26014 111746
rect 26014 111694 26066 111746
rect 26066 111694 26068 111746
rect 26012 111692 26068 111694
rect 25900 110066 25956 110068
rect 25900 110014 25902 110066
rect 25902 110014 25954 110066
rect 25954 110014 25956 110066
rect 25900 110012 25956 110014
rect 26572 113260 26628 113316
rect 26460 112924 26516 112980
rect 27020 112812 27076 112868
rect 27132 113148 27188 113204
rect 26908 112364 26964 112420
rect 26796 111916 26852 111972
rect 26124 110796 26180 110852
rect 26460 111692 26516 111748
rect 26012 109900 26068 109956
rect 25676 96124 25732 96180
rect 25452 92706 25508 92708
rect 25452 92654 25454 92706
rect 25454 92654 25506 92706
rect 25506 92654 25508 92706
rect 25452 92652 25508 92654
rect 25452 35420 25508 35476
rect 25452 34130 25508 34132
rect 25452 34078 25454 34130
rect 25454 34078 25506 34130
rect 25506 34078 25508 34130
rect 25452 34076 25508 34078
rect 24892 14812 24948 14868
rect 24464 13354 24520 13356
rect 24464 13302 24466 13354
rect 24466 13302 24518 13354
rect 24518 13302 24520 13354
rect 24464 13300 24520 13302
rect 24568 13354 24624 13356
rect 24568 13302 24570 13354
rect 24570 13302 24622 13354
rect 24622 13302 24624 13354
rect 24568 13300 24624 13302
rect 24672 13354 24728 13356
rect 24672 13302 24674 13354
rect 24674 13302 24726 13354
rect 24726 13302 24728 13354
rect 24672 13300 24728 13302
rect 25116 12796 25172 12852
rect 24464 11786 24520 11788
rect 24464 11734 24466 11786
rect 24466 11734 24518 11786
rect 24518 11734 24520 11786
rect 24464 11732 24520 11734
rect 24568 11786 24624 11788
rect 24568 11734 24570 11786
rect 24570 11734 24622 11786
rect 24622 11734 24624 11786
rect 24568 11732 24624 11734
rect 24672 11786 24728 11788
rect 24672 11734 24674 11786
rect 24674 11734 24726 11786
rect 24726 11734 24728 11786
rect 24672 11732 24728 11734
rect 25004 10332 25060 10388
rect 24464 10218 24520 10220
rect 24464 10166 24466 10218
rect 24466 10166 24518 10218
rect 24518 10166 24520 10218
rect 24464 10164 24520 10166
rect 24568 10218 24624 10220
rect 24568 10166 24570 10218
rect 24570 10166 24622 10218
rect 24622 10166 24624 10218
rect 24568 10164 24624 10166
rect 24672 10218 24728 10220
rect 24672 10166 24674 10218
rect 24674 10166 24726 10218
rect 24726 10166 24728 10218
rect 24672 10164 24728 10166
rect 24556 9154 24612 9156
rect 24556 9102 24558 9154
rect 24558 9102 24610 9154
rect 24610 9102 24612 9154
rect 24556 9100 24612 9102
rect 24892 9100 24948 9156
rect 24464 8650 24520 8652
rect 24464 8598 24466 8650
rect 24466 8598 24518 8650
rect 24518 8598 24520 8650
rect 24464 8596 24520 8598
rect 24568 8650 24624 8652
rect 24568 8598 24570 8650
rect 24570 8598 24622 8650
rect 24622 8598 24624 8650
rect 24568 8596 24624 8598
rect 24672 8650 24728 8652
rect 24672 8598 24674 8650
rect 24674 8598 24726 8650
rect 24726 8598 24728 8650
rect 24672 8596 24728 8598
rect 24464 7082 24520 7084
rect 24464 7030 24466 7082
rect 24466 7030 24518 7082
rect 24518 7030 24520 7082
rect 24464 7028 24520 7030
rect 24568 7082 24624 7084
rect 24568 7030 24570 7082
rect 24570 7030 24622 7082
rect 24622 7030 24624 7082
rect 24568 7028 24624 7030
rect 24672 7082 24728 7084
rect 24672 7030 24674 7082
rect 24674 7030 24726 7082
rect 24726 7030 24728 7082
rect 24672 7028 24728 7030
rect 24556 5906 24612 5908
rect 24556 5854 24558 5906
rect 24558 5854 24610 5906
rect 24610 5854 24612 5906
rect 24556 5852 24612 5854
rect 24464 5514 24520 5516
rect 24464 5462 24466 5514
rect 24466 5462 24518 5514
rect 24518 5462 24520 5514
rect 24464 5460 24520 5462
rect 24568 5514 24624 5516
rect 24568 5462 24570 5514
rect 24570 5462 24622 5514
rect 24622 5462 24624 5514
rect 24568 5460 24624 5462
rect 24672 5514 24728 5516
rect 24672 5462 24674 5514
rect 24674 5462 24726 5514
rect 24726 5462 24728 5514
rect 24672 5460 24728 5462
rect 25788 92706 25844 92708
rect 25788 92654 25790 92706
rect 25790 92654 25842 92706
rect 25842 92654 25844 92706
rect 25788 92652 25844 92654
rect 26124 108498 26180 108500
rect 26124 108446 26126 108498
rect 26126 108446 26178 108498
rect 26178 108446 26180 108498
rect 26124 108444 26180 108446
rect 26796 111692 26852 111748
rect 26796 110572 26852 110628
rect 26572 110290 26628 110292
rect 26572 110238 26574 110290
rect 26574 110238 26626 110290
rect 26626 110238 26628 110290
rect 26572 110236 26628 110238
rect 26460 110012 26516 110068
rect 27580 113036 27636 113092
rect 27468 112418 27524 112420
rect 27468 112366 27470 112418
rect 27470 112366 27522 112418
rect 27522 112366 27524 112418
rect 27468 112364 27524 112366
rect 27468 112028 27524 112084
rect 27244 111970 27300 111972
rect 27244 111918 27246 111970
rect 27246 111918 27298 111970
rect 27298 111918 27300 111970
rect 27244 111916 27300 111918
rect 27244 110796 27300 110852
rect 28252 112588 28308 112644
rect 29148 114604 29204 114660
rect 29036 114156 29092 114212
rect 28476 111746 28532 111748
rect 28476 111694 28478 111746
rect 28478 111694 28530 111746
rect 28530 111694 28532 111746
rect 28476 111692 28532 111694
rect 28924 112476 28980 112532
rect 28812 112306 28868 112308
rect 28812 112254 28814 112306
rect 28814 112254 28866 112306
rect 28866 112254 28868 112306
rect 28812 112252 28868 112254
rect 29820 113538 29876 113540
rect 29820 113486 29822 113538
rect 29822 113486 29874 113538
rect 29874 113486 29876 113538
rect 29820 113484 29876 113486
rect 29260 113314 29316 113316
rect 29260 113262 29262 113314
rect 29262 113262 29314 113314
rect 29314 113262 29316 113314
rect 29260 113260 29316 113262
rect 29932 112924 29988 112980
rect 29820 112700 29876 112756
rect 29260 111858 29316 111860
rect 29260 111806 29262 111858
rect 29262 111806 29314 111858
rect 29314 111806 29316 111858
rect 29260 111804 29316 111806
rect 28588 111468 28644 111524
rect 27916 111356 27972 111412
rect 30044 112028 30100 112084
rect 30156 111916 30212 111972
rect 30604 111858 30660 111860
rect 30604 111806 30606 111858
rect 30606 111806 30658 111858
rect 30658 111806 30660 111858
rect 30604 111804 30660 111806
rect 29484 111244 29540 111300
rect 30268 111580 30324 111636
rect 29596 111132 29652 111188
rect 27804 111020 27860 111076
rect 27020 110402 27076 110404
rect 27020 110350 27022 110402
rect 27022 110350 27074 110402
rect 27074 110350 27076 110402
rect 27020 110348 27076 110350
rect 27356 110402 27412 110404
rect 27356 110350 27358 110402
rect 27358 110350 27410 110402
rect 27410 110350 27412 110402
rect 27356 110348 27412 110350
rect 27692 110290 27748 110292
rect 27692 110238 27694 110290
rect 27694 110238 27746 110290
rect 27746 110238 27748 110290
rect 27692 110236 27748 110238
rect 26908 109340 26964 109396
rect 27244 110124 27300 110180
rect 26348 108444 26404 108500
rect 26572 109004 26628 109060
rect 26236 106092 26292 106148
rect 26348 94220 26404 94276
rect 25900 87500 25956 87556
rect 26236 89068 26292 89124
rect 26460 82460 26516 82516
rect 26236 76524 26292 76580
rect 27020 109004 27076 109060
rect 27020 108780 27076 108836
rect 26572 79996 26628 80052
rect 26684 76524 26740 76580
rect 26012 39788 26068 39844
rect 25788 32844 25844 32900
rect 25676 9996 25732 10052
rect 25788 17612 25844 17668
rect 26012 30156 26068 30212
rect 25900 16268 25956 16324
rect 26572 76412 26628 76468
rect 26572 15932 26628 15988
rect 26460 15148 26516 15204
rect 27132 108444 27188 108500
rect 27132 89068 27188 89124
rect 26796 17612 26852 17668
rect 27020 17724 27076 17780
rect 26348 15036 26404 15092
rect 26236 14812 26292 14868
rect 25788 6972 25844 7028
rect 26012 14588 26068 14644
rect 25788 6748 25844 6804
rect 25340 5906 25396 5908
rect 25340 5854 25342 5906
rect 25342 5854 25394 5906
rect 25394 5854 25396 5906
rect 25340 5852 25396 5854
rect 25116 5404 25172 5460
rect 25116 4732 25172 4788
rect 25116 4284 25172 4340
rect 24668 4172 24724 4228
rect 25004 4172 25060 4228
rect 24464 3946 24520 3948
rect 24464 3894 24466 3946
rect 24466 3894 24518 3946
rect 24518 3894 24520 3946
rect 24464 3892 24520 3894
rect 24568 3946 24624 3948
rect 24568 3894 24570 3946
rect 24570 3894 24622 3946
rect 24622 3894 24624 3946
rect 24568 3892 24624 3894
rect 24672 3946 24728 3948
rect 24672 3894 24674 3946
rect 24674 3894 24726 3946
rect 24726 3894 24728 3946
rect 24672 3892 24728 3894
rect 24892 3778 24948 3780
rect 24892 3726 24894 3778
rect 24894 3726 24946 3778
rect 24946 3726 24948 3778
rect 24892 3724 24948 3726
rect 24556 2940 24612 2996
rect 25228 3724 25284 3780
rect 25004 2940 25060 2996
rect 25228 3164 25284 3220
rect 24464 2378 24520 2380
rect 24464 2326 24466 2378
rect 24466 2326 24518 2378
rect 24518 2326 24520 2378
rect 24464 2324 24520 2326
rect 24568 2378 24624 2380
rect 24568 2326 24570 2378
rect 24570 2326 24622 2378
rect 24622 2326 24624 2378
rect 24568 2324 24624 2326
rect 24672 2378 24728 2380
rect 24672 2326 24674 2378
rect 24674 2326 24726 2378
rect 24726 2326 24728 2378
rect 24672 2324 24728 2326
rect 24892 2268 24948 2324
rect 25116 1820 25172 1876
rect 25116 1596 25172 1652
rect 24332 1484 24388 1540
rect 23996 1148 24052 1204
rect 24892 1260 24948 1316
rect 24464 810 24520 812
rect 24464 758 24466 810
rect 24466 758 24518 810
rect 24518 758 24520 810
rect 24464 756 24520 758
rect 24568 810 24624 812
rect 24568 758 24570 810
rect 24570 758 24622 810
rect 24622 758 24624 810
rect 24568 756 24624 758
rect 24672 810 24728 812
rect 24672 758 24674 810
rect 24674 758 24726 810
rect 24726 758 24728 810
rect 24672 756 24728 758
rect 24444 588 24500 644
rect 24668 588 24724 644
rect 25564 4732 25620 4788
rect 25452 3948 25508 4004
rect 25900 3500 25956 3556
rect 26012 3164 26068 3220
rect 26124 9884 26180 9940
rect 26460 14812 26516 14868
rect 26572 14588 26628 14644
rect 26572 7308 26628 7364
rect 26460 4396 26516 4452
rect 26348 4226 26404 4228
rect 26348 4174 26350 4226
rect 26350 4174 26402 4226
rect 26402 4174 26404 4226
rect 26348 4172 26404 4174
rect 25452 2770 25508 2772
rect 25452 2718 25454 2770
rect 25454 2718 25506 2770
rect 25506 2718 25508 2770
rect 25452 2716 25508 2718
rect 25788 2546 25844 2548
rect 25788 2494 25790 2546
rect 25790 2494 25842 2546
rect 25842 2494 25844 2546
rect 25788 2492 25844 2494
rect 25788 2268 25844 2324
rect 25452 2156 25508 2212
rect 25564 812 25620 868
rect 26124 2770 26180 2772
rect 26124 2718 26126 2770
rect 26126 2718 26178 2770
rect 26178 2718 26180 2770
rect 26124 2716 26180 2718
rect 26572 4060 26628 4116
rect 26908 5794 26964 5796
rect 26908 5742 26910 5794
rect 26910 5742 26962 5794
rect 26962 5742 26964 5794
rect 26908 5740 26964 5742
rect 26684 3836 26740 3892
rect 26796 3554 26852 3556
rect 26796 3502 26798 3554
rect 26798 3502 26850 3554
rect 26850 3502 26852 3554
rect 26796 3500 26852 3502
rect 26348 2156 26404 2212
rect 26236 1874 26292 1876
rect 26236 1822 26238 1874
rect 26238 1822 26290 1874
rect 26290 1822 26292 1874
rect 26236 1820 26292 1822
rect 26012 1596 26068 1652
rect 26124 1090 26180 1092
rect 26124 1038 26126 1090
rect 26126 1038 26178 1090
rect 26178 1038 26180 1090
rect 26124 1036 26180 1038
rect 26796 2098 26852 2100
rect 26796 2046 26798 2098
rect 26798 2046 26850 2098
rect 26850 2046 26852 2098
rect 26796 2044 26852 2046
rect 28476 109004 28532 109060
rect 27356 108332 27412 108388
rect 27804 94332 27860 94388
rect 27692 55244 27748 55300
rect 27356 6860 27412 6916
rect 27692 38108 27748 38164
rect 28028 92652 28084 92708
rect 27916 90300 27972 90356
rect 28028 35084 28084 35140
rect 28140 85596 28196 85652
rect 28252 56252 28308 56308
rect 28364 55298 28420 55300
rect 28364 55246 28366 55298
rect 28366 55246 28418 55298
rect 28418 55246 28420 55298
rect 28364 55244 28420 55246
rect 28140 27916 28196 27972
rect 28252 40908 28308 40964
rect 27916 19404 27972 19460
rect 28028 26796 28084 26852
rect 27804 17836 27860 17892
rect 27692 6524 27748 6580
rect 27804 15148 27860 15204
rect 27244 5068 27300 5124
rect 27468 6412 27524 6468
rect 27356 4844 27412 4900
rect 27132 1932 27188 1988
rect 27244 1148 27300 1204
rect 28028 11564 28084 11620
rect 28364 24668 28420 24724
rect 28252 9212 28308 9268
rect 30604 110738 30660 110740
rect 30604 110686 30606 110738
rect 30606 110686 30658 110738
rect 30658 110686 30660 110738
rect 30604 110684 30660 110686
rect 29484 109452 29540 109508
rect 30604 109564 30660 109620
rect 30380 108668 30436 108724
rect 30604 108444 30660 108500
rect 30604 107324 30660 107380
rect 30604 106204 30660 106260
rect 29596 105980 29652 106036
rect 30268 105586 30324 105588
rect 30268 105534 30270 105586
rect 30270 105534 30322 105586
rect 30322 105534 30324 105586
rect 30268 105532 30324 105534
rect 30604 105084 30660 105140
rect 30268 104076 30324 104132
rect 30604 103964 30660 104020
rect 30268 102898 30324 102900
rect 30268 102846 30270 102898
rect 30270 102846 30322 102898
rect 30322 102846 30324 102898
rect 30268 102844 30324 102846
rect 30604 102898 30660 102900
rect 30604 102846 30606 102898
rect 30606 102846 30658 102898
rect 30658 102846 30660 102898
rect 30604 102844 30660 102846
rect 30268 102450 30324 102452
rect 30268 102398 30270 102450
rect 30270 102398 30322 102450
rect 30322 102398 30324 102450
rect 30268 102396 30324 102398
rect 30604 101724 30660 101780
rect 29484 100770 29540 100772
rect 29484 100718 29486 100770
rect 29486 100718 29538 100770
rect 29538 100718 29540 100770
rect 29484 100716 29540 100718
rect 30604 100604 30660 100660
rect 30268 99762 30324 99764
rect 30268 99710 30270 99762
rect 30270 99710 30322 99762
rect 30322 99710 30324 99762
rect 30268 99708 30324 99710
rect 30604 99484 30660 99540
rect 30268 99314 30324 99316
rect 30268 99262 30270 99314
rect 30270 99262 30322 99314
rect 30322 99262 30324 99314
rect 30268 99260 30324 99262
rect 29372 99036 29428 99092
rect 29260 98924 29316 98980
rect 30604 98364 30660 98420
rect 30604 97244 30660 97300
rect 29484 96796 29540 96852
rect 29484 96572 29540 96628
rect 30604 96124 30660 96180
rect 30380 95228 30436 95284
rect 30268 94668 30324 94724
rect 30604 95058 30660 95060
rect 30604 95006 30606 95058
rect 30606 95006 30658 95058
rect 30658 95006 30660 95058
rect 30604 95004 30660 95006
rect 30604 93884 30660 93940
rect 30268 93436 30324 93492
rect 30604 92764 30660 92820
rect 30268 91922 30324 91924
rect 30268 91870 30270 91922
rect 30270 91870 30322 91922
rect 30322 91870 30324 91922
rect 30268 91868 30324 91870
rect 30604 91644 30660 91700
rect 30604 90524 30660 90580
rect 30268 90412 30324 90468
rect 30268 89906 30324 89908
rect 30268 89854 30270 89906
rect 30270 89854 30322 89906
rect 30322 89854 30324 89906
rect 30268 89852 30324 89854
rect 30604 89404 30660 89460
rect 30604 88284 30660 88340
rect 30268 87442 30324 87444
rect 30268 87390 30270 87442
rect 30270 87390 30322 87442
rect 30322 87390 30324 87442
rect 30268 87388 30324 87390
rect 30604 87218 30660 87220
rect 30604 87166 30606 87218
rect 30606 87166 30658 87218
rect 30658 87166 30660 87218
rect 30604 87164 30660 87166
rect 30604 86044 30660 86100
rect 30268 85708 30324 85764
rect 30268 85202 30324 85204
rect 30268 85150 30270 85202
rect 30270 85150 30322 85202
rect 30322 85150 30324 85202
rect 30268 85148 30324 85150
rect 30604 84924 30660 84980
rect 30268 84082 30324 84084
rect 30268 84030 30270 84082
rect 30270 84030 30322 84082
rect 30322 84030 30324 84082
rect 30268 84028 30324 84030
rect 30604 83804 30660 83860
rect 30604 82684 30660 82740
rect 30268 82572 30324 82628
rect 29484 81954 29540 81956
rect 29484 81902 29486 81954
rect 29486 81902 29538 81954
rect 29538 81902 29540 81954
rect 29484 81900 29540 81902
rect 30604 81564 30660 81620
rect 30604 80444 30660 80500
rect 29484 79660 29540 79716
rect 30604 79378 30660 79380
rect 30604 79326 30606 79378
rect 30606 79326 30658 79378
rect 30658 79326 30660 79378
rect 30604 79324 30660 79326
rect 29484 78876 29540 78932
rect 29484 77922 29540 77924
rect 29484 77870 29486 77922
rect 29486 77870 29538 77922
rect 29538 77870 29540 77922
rect 29484 77868 29540 77870
rect 30604 78204 30660 78260
rect 29372 77756 29428 77812
rect 30268 74674 30324 74676
rect 30268 74622 30270 74674
rect 30270 74622 30322 74674
rect 30322 74622 30324 74674
rect 30268 74620 30324 74622
rect 30604 74674 30660 74676
rect 30604 74622 30606 74674
rect 30606 74622 30658 74674
rect 30658 74622 30660 74674
rect 30604 74620 30660 74622
rect 30268 74114 30324 74116
rect 30268 74062 30270 74114
rect 30270 74062 30322 74114
rect 30322 74062 30324 74114
rect 30268 74060 30324 74062
rect 30604 73500 30660 73556
rect 30604 72380 30660 72436
rect 29484 70978 29540 70980
rect 29484 70926 29486 70978
rect 29486 70926 29538 70978
rect 29538 70926 29540 70978
rect 29484 70924 29540 70926
rect 28700 68348 28756 68404
rect 29484 68402 29540 68404
rect 29484 68350 29486 68402
rect 29486 68350 29538 68402
rect 29538 68350 29540 68402
rect 29484 68348 29540 68350
rect 28700 58156 28756 58212
rect 28812 63084 28868 63140
rect 29484 63138 29540 63140
rect 29484 63086 29486 63138
rect 29486 63086 29538 63138
rect 29538 63086 29540 63138
rect 29484 63084 29540 63086
rect 29596 60172 29652 60228
rect 30604 71260 30660 71316
rect 30604 70140 30660 70196
rect 30604 69020 30660 69076
rect 30604 67900 30660 67956
rect 30268 66444 30324 66500
rect 30380 64764 30436 64820
rect 30604 66834 30660 66836
rect 30604 66782 30606 66834
rect 30606 66782 30658 66834
rect 30658 66782 30660 66834
rect 30604 66780 30660 66782
rect 30604 65660 30660 65716
rect 30604 64540 30660 64596
rect 30492 63868 30548 63924
rect 30604 63420 30660 63476
rect 30604 62300 30660 62356
rect 30604 61180 30660 61236
rect 29708 59724 29764 59780
rect 30604 60060 30660 60116
rect 29484 59388 29540 59444
rect 29484 57708 29540 57764
rect 30604 58994 30660 58996
rect 30604 58942 30606 58994
rect 30606 58942 30658 58994
rect 30658 58942 30660 58994
rect 30604 58940 30660 58942
rect 29260 56588 29316 56644
rect 30604 57820 30660 57876
rect 30268 56028 30324 56084
rect 30604 56700 30660 56756
rect 30604 55580 30660 55636
rect 29932 53676 29988 53732
rect 29484 51884 29540 51940
rect 29372 50652 29428 50708
rect 30604 54460 30660 54516
rect 30156 53452 30212 53508
rect 30604 53340 30660 53396
rect 30380 52668 30436 52724
rect 30268 52220 30324 52276
rect 30604 52220 30660 52276
rect 30268 51154 30324 51156
rect 30268 51102 30270 51154
rect 30270 51102 30322 51154
rect 30322 51102 30324 51154
rect 30268 51100 30324 51102
rect 30604 51154 30660 51156
rect 30604 51102 30606 51154
rect 30606 51102 30658 51154
rect 30658 51102 30660 51154
rect 30604 51100 30660 51102
rect 30604 49980 30660 50036
rect 30380 49084 30436 49140
rect 30492 49644 30548 49700
rect 30044 48300 30100 48356
rect 30268 48188 30324 48244
rect 28812 48076 28868 48132
rect 30268 48018 30324 48020
rect 30268 47966 30270 48018
rect 30270 47966 30322 48018
rect 30322 47966 30324 48018
rect 30268 47964 30324 47966
rect 30268 47458 30324 47460
rect 30268 47406 30270 47458
rect 30270 47406 30322 47458
rect 30322 47406 30324 47458
rect 30268 47404 30324 47406
rect 29708 45276 29764 45332
rect 29484 44882 29540 44884
rect 29484 44830 29486 44882
rect 29486 44830 29538 44882
rect 29538 44830 29540 44882
rect 29484 44828 29540 44830
rect 29484 40460 29540 40516
rect 29484 39452 29540 39508
rect 29484 37996 29540 38052
rect 29596 36652 29652 36708
rect 30380 42812 30436 42868
rect 30268 36540 30324 36596
rect 29596 32620 29652 32676
rect 29372 30716 29428 30772
rect 29148 29148 29204 29204
rect 29596 27858 29652 27860
rect 29596 27806 29598 27858
rect 29598 27806 29650 27858
rect 29650 27806 29652 27858
rect 29596 27804 29652 27806
rect 29708 27746 29764 27748
rect 29708 27694 29710 27746
rect 29710 27694 29762 27746
rect 29762 27694 29764 27746
rect 29708 27692 29764 27694
rect 30268 35138 30324 35140
rect 30268 35086 30270 35138
rect 30270 35086 30322 35138
rect 30322 35086 30324 35138
rect 30268 35084 30324 35086
rect 30268 34300 30324 34356
rect 30604 48860 30660 48916
rect 30604 47740 30660 47796
rect 30604 46620 30660 46676
rect 30604 45500 30660 45556
rect 30604 44380 30660 44436
rect 30604 43314 30660 43316
rect 30604 43262 30606 43314
rect 30606 43262 30658 43314
rect 30658 43262 30660 43314
rect 30604 43260 30660 43262
rect 30604 42140 30660 42196
rect 30604 41020 30660 41076
rect 30604 39900 30660 39956
rect 31276 37772 31332 37828
rect 30604 35196 30660 35252
rect 30604 34300 30660 34356
rect 30380 32844 30436 32900
rect 30156 30828 30212 30884
rect 30268 30210 30324 30212
rect 30268 30158 30270 30210
rect 30270 30158 30322 30210
rect 30322 30158 30324 30210
rect 30268 30156 30324 30158
rect 30268 28754 30324 28756
rect 30268 28702 30270 28754
rect 30270 28702 30322 28754
rect 30322 28702 30324 28754
rect 30268 28700 30324 28702
rect 30268 27916 30324 27972
rect 30268 25730 30324 25732
rect 30268 25678 30270 25730
rect 30270 25678 30322 25730
rect 30322 25678 30324 25730
rect 30268 25676 30324 25678
rect 30716 33404 30772 33460
rect 30604 32508 30660 32564
rect 30604 31612 30660 31668
rect 30604 30770 30660 30772
rect 30604 30718 30606 30770
rect 30606 30718 30658 30770
rect 30658 30718 30660 30770
rect 30604 30716 30660 30718
rect 30604 29820 30660 29876
rect 30604 28924 30660 28980
rect 30604 28028 30660 28084
rect 30716 27132 30772 27188
rect 30604 26236 30660 26292
rect 30604 25340 30660 25396
rect 29484 25004 29540 25060
rect 30268 24722 30324 24724
rect 30268 24670 30270 24722
rect 30270 24670 30322 24722
rect 30322 24670 30324 24722
rect 30268 24668 30324 24670
rect 30268 24050 30324 24052
rect 30268 23998 30270 24050
rect 30270 23998 30322 24050
rect 30322 23998 30324 24050
rect 30268 23996 30324 23998
rect 30268 23324 30324 23380
rect 30268 22594 30324 22596
rect 30268 22542 30270 22594
rect 30270 22542 30322 22594
rect 30322 22542 30324 22594
rect 30268 22540 30324 22542
rect 30268 20802 30324 20804
rect 30268 20750 30270 20802
rect 30270 20750 30322 20802
rect 30322 20750 30324 20802
rect 30268 20748 30324 20750
rect 30156 20636 30212 20692
rect 30268 19458 30324 19460
rect 30268 19406 30270 19458
rect 30270 19406 30322 19458
rect 30322 19406 30324 19458
rect 30268 19404 30324 19406
rect 30268 18450 30324 18452
rect 30268 18398 30270 18450
rect 30270 18398 30322 18450
rect 30322 18398 30324 18450
rect 30268 18396 30324 18398
rect 30268 17890 30324 17892
rect 30268 17838 30270 17890
rect 30270 17838 30322 17890
rect 30322 17838 30324 17890
rect 30268 17836 30324 17838
rect 30268 16658 30324 16660
rect 30268 16606 30270 16658
rect 30270 16606 30322 16658
rect 30322 16606 30324 16658
rect 30268 16604 30324 16606
rect 30268 16322 30324 16324
rect 30268 16270 30270 16322
rect 30270 16270 30322 16322
rect 30322 16270 30324 16322
rect 30268 16268 30324 16270
rect 30492 25004 30548 25060
rect 30268 14754 30324 14756
rect 30268 14702 30270 14754
rect 30270 14702 30322 14754
rect 30322 14702 30324 14754
rect 30268 14700 30324 14702
rect 30268 13186 30324 13188
rect 30268 13134 30270 13186
rect 30270 13134 30322 13186
rect 30322 13134 30324 13186
rect 30268 13132 30324 13134
rect 30604 24498 30660 24500
rect 30604 24446 30606 24498
rect 30606 24446 30658 24498
rect 30658 24446 30660 24498
rect 30604 24444 30660 24446
rect 30604 23548 30660 23604
rect 30604 22652 30660 22708
rect 30604 21756 30660 21812
rect 30716 20860 30772 20916
rect 30604 19964 30660 20020
rect 30604 19068 30660 19124
rect 30604 18226 30660 18228
rect 30604 18174 30606 18226
rect 30606 18174 30658 18226
rect 30658 18174 30660 18226
rect 30604 18172 30660 18174
rect 30604 17276 30660 17332
rect 30604 16380 30660 16436
rect 30604 15484 30660 15540
rect 30716 14588 30772 14644
rect 30604 13692 30660 13748
rect 30604 12796 30660 12852
rect 30604 11954 30660 11956
rect 30604 11902 30606 11954
rect 30606 11902 30658 11954
rect 30658 11902 30660 11954
rect 30604 11900 30660 11902
rect 30268 11618 30324 11620
rect 30268 11566 30270 11618
rect 30270 11566 30322 11618
rect 30322 11566 30324 11618
rect 30268 11564 30324 11566
rect 30604 11004 30660 11060
rect 28140 1708 28196 1764
rect 31500 27692 31556 27748
rect 31388 15260 31444 15316
rect 31500 10108 31556 10164
rect 31388 8316 31444 8372
rect 31276 7420 31332 7476
rect 29260 5628 29316 5684
rect 28476 3276 28532 3332
rect 28364 1596 28420 1652
rect 28588 1372 28644 1428
rect 27692 1260 27748 1316
rect 28028 1202 28084 1204
rect 28028 1150 28030 1202
rect 28030 1150 28082 1202
rect 28082 1150 28084 1202
rect 28028 1148 28084 1150
rect 28364 1090 28420 1092
rect 28364 1038 28366 1090
rect 28366 1038 28418 1090
rect 28418 1038 28420 1090
rect 28364 1036 28420 1038
rect 27468 476 27524 532
rect 29036 252 29092 308
rect 26796 140 26852 196
rect 26460 28 26516 84
<< metal3 >>
rect 9874 114716 9884 114772
rect 9940 114716 23044 114772
rect 23986 114716 23996 114772
rect 24052 114716 28476 114772
rect 28532 114716 28542 114772
rect 0 114660 112 114688
rect 22988 114660 23044 114716
rect 0 114604 6636 114660
rect 6692 114604 6702 114660
rect 22978 114604 22988 114660
rect 23044 114604 23054 114660
rect 24658 114604 24668 114660
rect 24724 114604 29148 114660
rect 29204 114604 29214 114660
rect 0 114576 112 114604
rect 4274 114492 4284 114548
rect 4340 114492 12460 114548
rect 12516 114492 12526 114548
rect 22866 114492 22876 114548
rect 22932 114492 26124 114548
rect 26180 114492 26190 114548
rect 9090 114380 9100 114436
rect 9156 114380 10556 114436
rect 10612 114380 10622 114436
rect 11890 114380 11900 114436
rect 11956 114380 20524 114436
rect 20580 114380 20590 114436
rect 23314 114380 23324 114436
rect 23380 114380 26796 114436
rect 26852 114380 26862 114436
rect 8978 114268 8988 114324
rect 9044 114268 19852 114324
rect 19908 114268 19918 114324
rect 23762 114268 23772 114324
rect 23828 114268 28364 114324
rect 28420 114268 28430 114324
rect 0 114212 112 114240
rect 0 114156 140 114212
rect 196 114156 206 114212
rect 4834 114156 4844 114212
rect 4900 114156 10220 114212
rect 10276 114156 10286 114212
rect 12114 114156 12124 114212
rect 12180 114156 15372 114212
rect 15428 114156 15438 114212
rect 24210 114156 24220 114212
rect 24276 114156 29036 114212
rect 29092 114156 29102 114212
rect 0 114128 112 114156
rect 9202 114044 9212 114100
rect 9268 114044 21868 114100
rect 21924 114044 21934 114100
rect 22418 114044 22428 114100
rect 22484 114044 25452 114100
rect 25508 114044 25518 114100
rect 1922 113932 1932 113988
rect 1988 113932 6300 113988
rect 6356 113932 6366 113988
rect 9650 113932 9660 113988
rect 9716 113932 18508 113988
rect 18564 113932 18574 113988
rect 18834 113932 18844 113988
rect 18900 113932 19964 113988
rect 20020 113932 20030 113988
rect 24434 113932 24444 113988
rect 24500 113932 27692 113988
rect 27748 113932 27758 113988
rect 5366 113820 5404 113876
rect 5460 113820 5470 113876
rect 5842 113820 5852 113876
rect 5908 113820 11900 113876
rect 11956 113820 11966 113876
rect 12338 113820 12348 113876
rect 12404 113820 22316 113876
rect 22372 113820 22382 113876
rect 22642 113820 22652 113876
rect 22708 113820 25676 113876
rect 25732 113820 25742 113876
rect 0 113764 112 113792
rect 0 113708 812 113764
rect 868 113708 878 113764
rect 8530 113708 8540 113764
rect 8596 113708 11900 113764
rect 11956 113708 11966 113764
rect 18610 113708 18620 113764
rect 18676 113708 19628 113764
rect 19684 113708 19694 113764
rect 0 113680 112 113708
rect 4454 113652 4464 113708
rect 4520 113652 4568 113708
rect 4624 113652 4672 113708
rect 4728 113652 4738 113708
rect 24454 113652 24464 113708
rect 24520 113652 24568 113708
rect 24624 113652 24672 113708
rect 24728 113652 24738 113708
rect 5170 113596 5180 113652
rect 5236 113596 10332 113652
rect 10388 113596 10398 113652
rect 12562 113596 12572 113652
rect 12628 113596 19180 113652
rect 19236 113596 19246 113652
rect 25778 113596 25788 113652
rect 25844 113596 27356 113652
rect 27412 113596 27422 113652
rect 1474 113484 1484 113540
rect 1540 113484 8092 113540
rect 8148 113484 8158 113540
rect 13010 113484 13020 113540
rect 13076 113484 14700 113540
rect 14756 113484 14766 113540
rect 14998 113484 15036 113540
rect 15092 113484 15102 113540
rect 19478 113484 19516 113540
rect 19572 113484 19582 113540
rect 21522 113484 21532 113540
rect 21588 113484 24556 113540
rect 24612 113484 24622 113540
rect 26002 113484 26012 113540
rect 26068 113484 29820 113540
rect 29876 113484 29886 113540
rect 1036 113372 3164 113428
rect 3220 113372 3230 113428
rect 5282 113372 5292 113428
rect 5348 113372 5516 113428
rect 5572 113372 5582 113428
rect 5842 113372 5852 113428
rect 5908 113372 8764 113428
rect 8820 113372 8830 113428
rect 9874 113372 9884 113428
rect 9940 113372 11564 113428
rect 11620 113372 11630 113428
rect 13654 113372 13692 113428
rect 13748 113372 13758 113428
rect 14102 113372 14140 113428
rect 14196 113372 14206 113428
rect 14550 113372 14588 113428
rect 14644 113372 14654 113428
rect 16930 113372 16940 113428
rect 16996 113372 17500 113428
rect 17556 113372 17566 113428
rect 21746 113372 21756 113428
rect 21812 113372 24668 113428
rect 24724 113372 24734 113428
rect 0 113316 112 113344
rect 1036 113316 1092 113372
rect 0 113260 1092 113316
rect 1250 113260 1260 113316
rect 1316 113260 3388 113316
rect 3444 113260 3454 113316
rect 6066 113260 6076 113316
rect 6132 113260 7308 113316
rect 7364 113260 7374 113316
rect 7522 113260 7532 113316
rect 7588 113260 15148 113316
rect 15204 113260 15214 113316
rect 15362 113260 15372 113316
rect 15428 113260 16380 113316
rect 16436 113260 16446 113316
rect 19058 113260 19068 113316
rect 19124 113260 20188 113316
rect 20244 113260 20254 113316
rect 20402 113260 20412 113316
rect 20468 113260 21196 113316
rect 21252 113260 21262 113316
rect 22866 113260 22876 113316
rect 22932 113260 24780 113316
rect 24836 113260 24846 113316
rect 26562 113260 26572 113316
rect 26628 113260 29260 113316
rect 29316 113260 29326 113316
rect 0 113232 112 113260
rect 1474 113148 1484 113204
rect 1540 113148 7084 113204
rect 7140 113148 7150 113204
rect 7308 113148 13524 113204
rect 14578 113148 14588 113204
rect 14644 113148 19516 113204
rect 19572 113148 19582 113204
rect 23538 113148 23548 113204
rect 23604 113148 27132 113204
rect 27188 113148 27198 113204
rect 7308 113092 7364 113148
rect 13468 113092 13524 113148
rect 6626 113036 6636 113092
rect 6692 113036 7364 113092
rect 7970 113036 7980 113092
rect 8036 113036 9324 113092
rect 9380 113036 9390 113092
rect 10210 113036 10220 113092
rect 10276 113036 10668 113092
rect 10724 113036 10734 113092
rect 12226 113036 12236 113092
rect 12292 113036 13244 113092
rect 13300 113036 13310 113092
rect 13468 113036 16380 113092
rect 16436 113036 16446 113092
rect 23426 113036 23436 113092
rect 23492 113036 24948 113092
rect 25106 113036 25116 113092
rect 25172 113036 27580 113092
rect 27636 113036 27646 113092
rect 24892 112980 24948 113036
rect 31584 112980 31696 113008
rect 4946 112924 4956 112980
rect 5012 112924 7420 112980
rect 7476 112924 7486 112980
rect 9314 112924 9324 112980
rect 9380 112924 11676 112980
rect 11732 112924 12012 112980
rect 12068 112924 12078 112980
rect 12786 112924 12796 112980
rect 12852 112924 21364 112980
rect 21970 112924 21980 112980
rect 22036 112924 23324 112980
rect 23380 112924 23390 112980
rect 24892 112924 26460 112980
rect 26516 112924 26526 112980
rect 29922 112924 29932 112980
rect 29988 112924 31696 112980
rect 0 112868 112 112896
rect 3794 112868 3804 112924
rect 3860 112868 3908 112924
rect 3964 112868 4012 112924
rect 4068 112868 4078 112924
rect 21308 112868 21364 112924
rect 23794 112868 23804 112924
rect 23860 112868 23908 112924
rect 23964 112868 24012 112924
rect 24068 112868 24078 112924
rect 31584 112896 31696 112924
rect 0 112812 3388 112868
rect 6066 112812 6076 112868
rect 6132 112812 15596 112868
rect 15652 112812 15662 112868
rect 19506 112812 19516 112868
rect 19572 112812 19852 112868
rect 19908 112812 19918 112868
rect 21298 112812 21308 112868
rect 21364 112812 21374 112868
rect 24322 112812 24332 112868
rect 24388 112812 27020 112868
rect 27076 112812 27086 112868
rect 0 112784 112 112812
rect 3332 112756 3388 112812
rect 3332 112700 5180 112756
rect 5236 112700 5246 112756
rect 5404 112700 7532 112756
rect 7588 112700 7598 112756
rect 8082 112700 8092 112756
rect 8148 112700 11676 112756
rect 11732 112700 11742 112756
rect 12674 112700 12684 112756
rect 12740 112700 14140 112756
rect 14196 112700 14476 112756
rect 14532 112700 16716 112756
rect 16772 112700 18956 112756
rect 19012 112700 20748 112756
rect 20804 112700 21756 112756
rect 21812 112700 21822 112756
rect 22194 112700 22204 112756
rect 22260 112700 23996 112756
rect 24052 112700 24062 112756
rect 24210 112700 24220 112756
rect 24276 112700 24286 112756
rect 25554 112700 25564 112756
rect 25620 112700 29820 112756
rect 29876 112700 29886 112756
rect 5404 112644 5460 112700
rect 4946 112588 4956 112644
rect 5012 112588 5460 112644
rect 5730 112588 5740 112644
rect 5796 112588 7196 112644
rect 7252 112588 7262 112644
rect 10098 112588 10108 112644
rect 10164 112588 12124 112644
rect 12180 112588 12190 112644
rect 14326 112588 14364 112644
rect 14420 112588 14430 112644
rect 14774 112588 14812 112644
rect 14868 112588 14878 112644
rect 15138 112588 15148 112644
rect 15204 112588 15260 112644
rect 15316 112588 15326 112644
rect 16034 112588 16044 112644
rect 16100 112588 16156 112644
rect 16212 112588 16222 112644
rect 17014 112588 17052 112644
rect 17108 112588 17118 112644
rect 19954 112588 19964 112644
rect 20020 112588 20636 112644
rect 20692 112588 20702 112644
rect 5506 112476 5516 112532
rect 5572 112476 6300 112532
rect 6356 112476 6366 112532
rect 6822 112476 6860 112532
rect 6916 112476 10220 112532
rect 10276 112476 10286 112532
rect 10630 112476 10668 112532
rect 10724 112476 10734 112532
rect 10892 112476 11116 112532
rect 11172 112476 11182 112532
rect 11890 112476 11900 112532
rect 11956 112476 19572 112532
rect 19730 112476 19740 112532
rect 19796 112476 20300 112532
rect 20356 112476 20366 112532
rect 0 112420 112 112448
rect 10892 112420 10948 112476
rect 19516 112420 19572 112476
rect 0 112364 1092 112420
rect 4834 112364 4844 112420
rect 4900 112364 10948 112420
rect 11218 112364 11228 112420
rect 11284 112364 11340 112420
rect 11396 112364 11564 112420
rect 11620 112364 11630 112420
rect 11890 112364 11900 112420
rect 11956 112364 18900 112420
rect 19516 112364 23660 112420
rect 23716 112364 23726 112420
rect 0 112336 112 112364
rect 1036 112196 1092 112364
rect 1782 112252 1820 112308
rect 1876 112252 1886 112308
rect 5030 112252 5068 112308
rect 5124 112252 5134 112308
rect 5730 112252 5740 112308
rect 5796 112252 6412 112308
rect 6468 112252 6478 112308
rect 7942 112252 7980 112308
rect 8036 112252 8046 112308
rect 8530 112252 8540 112308
rect 8596 112252 9100 112308
rect 9156 112252 9166 112308
rect 10556 112252 14700 112308
rect 14756 112252 16156 112308
rect 16212 112252 16222 112308
rect 17350 112252 17388 112308
rect 17444 112252 17454 112308
rect 10556 112196 10612 112252
rect 18844 112196 18900 112364
rect 24220 112308 24276 112700
rect 25330 112588 25340 112644
rect 25396 112588 28252 112644
rect 28308 112588 28318 112644
rect 24882 112476 24892 112532
rect 24948 112476 28924 112532
rect 28980 112476 28990 112532
rect 26898 112364 26908 112420
rect 26964 112364 27468 112420
rect 27524 112364 27534 112420
rect 24210 112252 24220 112308
rect 24276 112252 24286 112308
rect 24882 112252 24892 112308
rect 24948 112252 28812 112308
rect 28868 112252 28878 112308
rect 1036 112140 1708 112196
rect 1764 112140 1774 112196
rect 6626 112140 6636 112196
rect 6692 112140 10612 112196
rect 10770 112140 10780 112196
rect 10836 112140 12684 112196
rect 12740 112140 12750 112196
rect 12908 112140 17612 112196
rect 17668 112140 17678 112196
rect 18844 112140 22652 112196
rect 22708 112140 22718 112196
rect 4454 112084 4464 112140
rect 4520 112084 4568 112140
rect 4624 112084 4672 112140
rect 4728 112084 4738 112140
rect 12908 112084 12964 112140
rect 24454 112084 24464 112140
rect 24520 112084 24568 112140
rect 24624 112084 24672 112140
rect 24728 112084 24738 112140
rect 8866 112028 8876 112084
rect 8932 112028 9660 112084
rect 9716 112028 9726 112084
rect 11890 112028 11900 112084
rect 11956 112028 12236 112084
rect 12292 112028 12302 112084
rect 12450 112028 12460 112084
rect 12516 112028 12964 112084
rect 13458 112028 13468 112084
rect 13524 112028 15260 112084
rect 15316 112028 15326 112084
rect 16146 112028 16156 112084
rect 16212 112028 20132 112084
rect 21522 112028 21532 112084
rect 21588 112028 22764 112084
rect 22820 112028 22830 112084
rect 25302 112028 25340 112084
rect 25396 112028 25406 112084
rect 27458 112028 27468 112084
rect 27524 112028 30044 112084
rect 30100 112028 30110 112084
rect 0 111972 112 112000
rect 0 111916 588 111972
rect 644 111916 654 111972
rect 4386 111916 4396 111972
rect 4452 111916 10724 111972
rect 10882 111916 10892 111972
rect 10948 111916 19852 111972
rect 19908 111916 19918 111972
rect 0 111888 112 111916
rect 10668 111860 10724 111916
rect 802 111804 812 111860
rect 868 111804 1596 111860
rect 1652 111804 1662 111860
rect 5058 111804 5068 111860
rect 5124 111804 7644 111860
rect 7700 111804 7710 111860
rect 9426 111804 9436 111860
rect 9492 111804 10332 111860
rect 10388 111804 10398 111860
rect 10668 111804 13132 111860
rect 13188 111804 13198 111860
rect 13682 111804 13692 111860
rect 13748 111804 14924 111860
rect 14980 111804 15148 111860
rect 17910 111804 17948 111860
rect 18004 111804 18014 111860
rect 15092 111748 15148 111804
rect 20076 111748 20132 112028
rect 21074 111916 21084 111972
rect 21140 111916 21868 111972
rect 21924 111916 21934 111972
rect 25106 111916 25116 111972
rect 25172 111916 26796 111972
rect 26852 111916 26862 111972
rect 27234 111916 27244 111972
rect 27300 111916 30156 111972
rect 30212 111916 30222 111972
rect 31584 111860 31696 111888
rect 21522 111804 21532 111860
rect 21588 111804 21644 111860
rect 21700 111804 21710 111860
rect 22166 111804 22204 111860
rect 22260 111804 22270 111860
rect 25554 111804 25564 111860
rect 25620 111804 29260 111860
rect 29316 111804 29326 111860
rect 30594 111804 30604 111860
rect 30660 111804 31696 111860
rect 31584 111776 31696 111804
rect 3490 111692 3500 111748
rect 3556 111692 7084 111748
rect 7140 111692 7150 111748
rect 7746 111692 7756 111748
rect 7812 111692 10220 111748
rect 10276 111692 10286 111748
rect 10518 111692 10556 111748
rect 10612 111692 10622 111748
rect 10892 111692 14980 111748
rect 15092 111692 18564 111748
rect 20076 111692 24668 111748
rect 24724 111692 24734 111748
rect 26002 111692 26012 111748
rect 26068 111692 26460 111748
rect 26516 111692 26526 111748
rect 26786 111692 26796 111748
rect 26852 111692 28476 111748
rect 28532 111692 28542 111748
rect 10892 111636 10948 111692
rect 14924 111636 14980 111692
rect 18508 111636 18564 111692
rect 1250 111580 1260 111636
rect 1316 111580 2716 111636
rect 2772 111580 3500 111636
rect 3556 111580 8428 111636
rect 8484 111580 8494 111636
rect 8754 111580 8764 111636
rect 8820 111580 10948 111636
rect 11190 111580 11228 111636
rect 11284 111580 11294 111636
rect 11442 111580 11452 111636
rect 11508 111580 13692 111636
rect 13748 111580 13758 111636
rect 14438 111580 14476 111636
rect 14532 111580 14542 111636
rect 14914 111580 14924 111636
rect 14980 111580 14990 111636
rect 16604 111580 18284 111636
rect 18340 111580 18350 111636
rect 18508 111580 20524 111636
rect 20580 111580 20590 111636
rect 23650 111580 23660 111636
rect 23716 111580 30268 111636
rect 30324 111580 30334 111636
rect 0 111524 112 111552
rect 16604 111524 16660 111580
rect 0 111468 1484 111524
rect 1540 111468 1550 111524
rect 3154 111468 3164 111524
rect 3220 111468 4900 111524
rect 7970 111468 7980 111524
rect 8036 111468 16660 111524
rect 16790 111468 16828 111524
rect 16884 111468 16894 111524
rect 17714 111468 17724 111524
rect 17780 111468 20636 111524
rect 20692 111468 20702 111524
rect 22194 111468 22204 111524
rect 22260 111468 23996 111524
rect 24052 111468 24062 111524
rect 24220 111468 28588 111524
rect 28644 111468 28654 111524
rect 0 111440 112 111468
rect 3794 111300 3804 111356
rect 3860 111300 3908 111356
rect 3964 111300 4012 111356
rect 4068 111300 4078 111356
rect 4844 111300 4900 111468
rect 5394 111356 5404 111412
rect 5460 111356 8988 111412
rect 9044 111356 9054 111412
rect 10882 111356 10892 111412
rect 10948 111356 13244 111412
rect 13300 111356 13310 111412
rect 13458 111356 13468 111412
rect 13524 111356 15036 111412
rect 15092 111356 15102 111412
rect 16370 111356 16380 111412
rect 16436 111356 23212 111412
rect 23268 111356 23278 111412
rect 23794 111300 23804 111356
rect 23860 111300 23908 111356
rect 23964 111300 24012 111356
rect 24068 111300 24078 111356
rect 4844 111244 14028 111300
rect 14084 111244 18004 111300
rect 4274 111132 4284 111188
rect 4340 111132 6412 111188
rect 6468 111132 6478 111188
rect 7074 111132 7084 111188
rect 7140 111132 11452 111188
rect 11508 111132 11518 111188
rect 12226 111132 12236 111188
rect 12292 111132 17724 111188
rect 17780 111132 17790 111188
rect 0 111076 112 111104
rect 17948 111076 18004 111244
rect 19516 111244 23324 111300
rect 23380 111244 23390 111300
rect 19516 111188 19572 111244
rect 24220 111188 24276 111468
rect 24882 111356 24892 111412
rect 24948 111356 27916 111412
rect 27972 111356 27982 111412
rect 25666 111244 25676 111300
rect 25732 111244 29484 111300
rect 29540 111244 29550 111300
rect 18274 111132 18284 111188
rect 18340 111132 19516 111188
rect 19572 111132 19582 111188
rect 20850 111132 20860 111188
rect 20916 111132 21980 111188
rect 22036 111132 22046 111188
rect 23874 111132 23884 111188
rect 23940 111132 24276 111188
rect 24994 111132 25004 111188
rect 25060 111132 29596 111188
rect 29652 111132 29662 111188
rect 0 111020 3500 111076
rect 3556 111020 3566 111076
rect 3714 111020 3724 111076
rect 3780 111020 4844 111076
rect 4900 111020 4910 111076
rect 5292 111020 7532 111076
rect 7588 111020 7598 111076
rect 10658 111020 10668 111076
rect 10724 111020 12908 111076
rect 12964 111020 12974 111076
rect 14252 111020 15820 111076
rect 15876 111020 15886 111076
rect 17948 111020 18228 111076
rect 20402 111020 20412 111076
rect 20468 111020 21084 111076
rect 21140 111020 21150 111076
rect 21746 111020 21756 111076
rect 21812 111020 23548 111076
rect 23650 111020 23660 111076
rect 23716 111020 25116 111076
rect 25172 111020 25182 111076
rect 25554 111020 25564 111076
rect 25620 111020 27804 111076
rect 27860 111020 27870 111076
rect 0 110992 112 111020
rect 5292 110964 5348 111020
rect 14252 110964 14308 111020
rect 18172 110964 18228 111020
rect 23492 110964 23548 111020
rect 578 110908 588 110964
rect 644 110908 1596 110964
rect 1652 110908 1662 110964
rect 2818 110908 2828 110964
rect 2884 110908 5348 110964
rect 5478 110908 5516 110964
rect 5572 110908 5582 110964
rect 6850 110908 6860 110964
rect 6916 110908 7980 110964
rect 8036 110908 8046 110964
rect 10546 110908 10556 110964
rect 10612 110908 11116 110964
rect 11172 110908 11182 110964
rect 11554 110908 11564 110964
rect 11620 110908 12796 110964
rect 12852 110908 12862 110964
rect 13468 110908 13580 110964
rect 13636 110908 14252 110964
rect 14308 110908 14318 110964
rect 14578 110908 14588 110964
rect 14644 110908 15148 110964
rect 15204 110908 15214 110964
rect 17826 110908 17836 110964
rect 17892 110908 17948 110964
rect 18004 110908 18014 110964
rect 18172 110908 18620 110964
rect 18676 110908 18686 110964
rect 20066 110908 20076 110964
rect 20132 110908 21308 110964
rect 21364 110908 21374 110964
rect 22278 110908 22316 110964
rect 22372 110908 22382 110964
rect 22978 110908 22988 110964
rect 23044 110908 23212 110964
rect 23268 110908 23278 110964
rect 23492 110908 23996 110964
rect 24052 110908 24062 110964
rect 13468 110852 13524 110908
rect 1474 110796 1484 110852
rect 1540 110796 6748 110852
rect 6804 110796 6814 110852
rect 13356 110796 13524 110852
rect 13682 110796 13692 110852
rect 13748 110796 17052 110852
rect 17108 110796 17118 110852
rect 19058 110796 19068 110852
rect 19124 110796 19134 110852
rect 22082 110796 22092 110852
rect 22148 110796 24780 110852
rect 24836 110796 24846 110852
rect 26114 110796 26124 110852
rect 26180 110796 27020 110852
rect 27076 110796 27086 110852
rect 27234 110796 27244 110852
rect 27300 110796 27310 110852
rect 13356 110740 13412 110796
rect 19068 110740 19124 110796
rect 4050 110684 4060 110740
rect 4116 110684 4844 110740
rect 4900 110684 4910 110740
rect 10882 110684 10892 110740
rect 10948 110684 11676 110740
rect 11732 110684 13020 110740
rect 13076 110684 13412 110740
rect 13570 110684 13580 110740
rect 13636 110684 13916 110740
rect 13972 110684 13982 110740
rect 14466 110684 14476 110740
rect 14532 110684 19124 110740
rect 24546 110684 24556 110740
rect 24612 110684 26908 110740
rect 26964 110684 26974 110740
rect 0 110628 112 110656
rect 27244 110628 27300 110796
rect 31584 110740 31696 110768
rect 30594 110684 30604 110740
rect 30660 110684 31696 110740
rect 31584 110656 31696 110684
rect 0 110572 3220 110628
rect 5394 110572 5404 110628
rect 5460 110572 9156 110628
rect 11330 110572 11340 110628
rect 11396 110572 14588 110628
rect 14644 110572 14654 110628
rect 15810 110572 15820 110628
rect 15876 110572 15932 110628
rect 15988 110572 15998 110628
rect 16258 110572 16268 110628
rect 16324 110572 19740 110628
rect 19796 110572 19806 110628
rect 22642 110572 22652 110628
rect 22708 110572 23324 110628
rect 23380 110572 23390 110628
rect 25302 110572 25340 110628
rect 25396 110572 25406 110628
rect 26786 110572 26796 110628
rect 26852 110572 27300 110628
rect 0 110544 112 110572
rect 3164 110292 3220 110572
rect 4454 110516 4464 110572
rect 4520 110516 4568 110572
rect 4624 110516 4672 110572
rect 4728 110516 4738 110572
rect 9100 110516 9156 110572
rect 24454 110516 24464 110572
rect 24520 110516 24568 110572
rect 24624 110516 24672 110572
rect 24728 110516 24738 110572
rect 3938 110460 3948 110516
rect 4004 110460 4284 110516
rect 4340 110460 4350 110516
rect 6150 110460 6188 110516
rect 6244 110460 6254 110516
rect 6402 110460 6412 110516
rect 6468 110460 6636 110516
rect 6692 110460 8876 110516
rect 8932 110460 8942 110516
rect 9100 110460 11564 110516
rect 11620 110460 12460 110516
rect 12516 110460 12526 110516
rect 13878 110460 13916 110516
rect 13972 110460 13982 110516
rect 15810 110460 15820 110516
rect 15876 110460 21644 110516
rect 21700 110460 21710 110516
rect 3378 110348 3388 110404
rect 3444 110348 9996 110404
rect 10052 110348 10062 110404
rect 12226 110348 12236 110404
rect 12292 110348 19964 110404
rect 20020 110348 20030 110404
rect 22642 110348 22652 110404
rect 22708 110348 23548 110404
rect 23604 110348 23614 110404
rect 27010 110348 27020 110404
rect 27076 110348 27132 110404
rect 27188 110348 27198 110404
rect 27346 110348 27356 110404
rect 27412 110348 27450 110404
rect 3164 110236 4228 110292
rect 4386 110236 4396 110292
rect 4452 110236 4956 110292
rect 5012 110236 5022 110292
rect 5180 110236 5628 110292
rect 5684 110236 5694 110292
rect 9202 110236 9212 110292
rect 9268 110236 21532 110292
rect 21588 110236 21598 110292
rect 25190 110236 25228 110292
rect 25284 110236 25294 110292
rect 26562 110236 26572 110292
rect 26628 110236 27692 110292
rect 27748 110236 27758 110292
rect 0 110180 112 110208
rect 4172 110180 4228 110236
rect 5180 110180 5236 110236
rect 0 110124 3948 110180
rect 4004 110124 4014 110180
rect 4172 110124 5236 110180
rect 5404 110124 6412 110180
rect 6468 110124 6478 110180
rect 10294 110124 10332 110180
rect 10388 110124 10398 110180
rect 13234 110124 13244 110180
rect 13300 110124 14252 110180
rect 14308 110124 14756 110180
rect 14914 110124 14924 110180
rect 14980 110124 15708 110180
rect 15764 110124 15774 110180
rect 18946 110124 18956 110180
rect 19012 110124 19292 110180
rect 19348 110124 19358 110180
rect 24658 110124 24668 110180
rect 24724 110124 27244 110180
rect 27300 110124 27310 110180
rect 0 110096 112 110124
rect 5404 110068 5460 110124
rect 14700 110068 14756 110124
rect 3052 110012 5460 110068
rect 5618 110012 5628 110068
rect 5684 110012 10276 110068
rect 12870 110012 12908 110068
rect 12964 110012 12974 110068
rect 13990 110012 14028 110068
rect 14084 110012 14094 110068
rect 14700 110012 15932 110068
rect 15988 110012 15998 110068
rect 17602 110012 17612 110068
rect 17668 110012 17836 110068
rect 17892 110012 22316 110068
rect 22372 110012 22382 110068
rect 25330 110012 25340 110068
rect 25396 110012 25900 110068
rect 25956 110012 26460 110068
rect 26516 110012 26526 110068
rect 3052 109844 3108 110012
rect 10220 109956 10276 110012
rect 3266 109900 3276 109956
rect 3332 109900 5292 109956
rect 5348 109900 5358 109956
rect 5730 109900 5740 109956
rect 5796 109900 6636 109956
rect 6692 109900 6702 109956
rect 10210 109900 10220 109956
rect 10276 109900 10286 109956
rect 11218 109900 11228 109956
rect 11284 109900 14252 109956
rect 14308 109900 14318 109956
rect 22194 109900 22204 109956
rect 22260 109900 26012 109956
rect 26068 109900 26078 109956
rect 3052 109788 3220 109844
rect 4274 109788 4284 109844
rect 4340 109788 5404 109844
rect 5460 109788 5470 109844
rect 5618 109788 5628 109844
rect 5684 109788 16268 109844
rect 16324 109788 16334 109844
rect 18274 109788 18284 109844
rect 18340 109788 18508 109844
rect 18564 109788 18574 109844
rect 0 109732 112 109760
rect 0 109676 1820 109732
rect 1876 109676 2940 109732
rect 2996 109676 3006 109732
rect 0 109648 112 109676
rect 3164 109620 3220 109788
rect 3794 109732 3804 109788
rect 3860 109732 3908 109788
rect 3964 109732 4012 109788
rect 4068 109732 4078 109788
rect 23794 109732 23804 109788
rect 23860 109732 23908 109788
rect 23964 109732 24012 109788
rect 24068 109732 24078 109788
rect 4834 109676 4844 109732
rect 4900 109676 7980 109732
rect 8036 109676 8046 109732
rect 12898 109676 12908 109732
rect 12964 109676 15484 109732
rect 15540 109676 15550 109732
rect 31584 109620 31696 109648
rect 924 109564 3220 109620
rect 3378 109564 3388 109620
rect 3444 109564 4620 109620
rect 4676 109564 4686 109620
rect 5394 109564 5404 109620
rect 5460 109564 13244 109620
rect 13300 109564 13310 109620
rect 14914 109564 14924 109620
rect 14980 109564 15036 109620
rect 15092 109564 15102 109620
rect 30594 109564 30604 109620
rect 30660 109564 31696 109620
rect 0 109284 112 109312
rect 924 109284 980 109564
rect 31584 109536 31696 109564
rect 1138 109452 1148 109508
rect 1204 109452 5404 109508
rect 5460 109452 5470 109508
rect 7970 109452 7980 109508
rect 8036 109452 12852 109508
rect 13010 109452 13020 109508
rect 13076 109452 13468 109508
rect 13524 109452 13580 109508
rect 13636 109452 13646 109508
rect 15810 109452 15820 109508
rect 15876 109452 17500 109508
rect 17556 109452 17566 109508
rect 18610 109452 18620 109508
rect 18676 109452 19964 109508
rect 20020 109452 29484 109508
rect 29540 109452 29550 109508
rect 12796 109396 12852 109452
rect 3490 109340 3500 109396
rect 3556 109340 3612 109396
rect 3668 109340 3678 109396
rect 3826 109340 3836 109396
rect 3892 109340 4956 109396
rect 5012 109340 7084 109396
rect 7140 109340 7150 109396
rect 8054 109340 8092 109396
rect 8148 109340 8158 109396
rect 9874 109340 9884 109396
rect 9940 109340 9996 109396
rect 10052 109340 10062 109396
rect 12796 109340 13916 109396
rect 13972 109340 14476 109396
rect 14532 109340 14542 109396
rect 16370 109340 16380 109396
rect 16436 109340 17724 109396
rect 17780 109340 17790 109396
rect 18610 109340 18620 109396
rect 18676 109340 18956 109396
rect 19012 109340 19022 109396
rect 23202 109340 23212 109396
rect 23268 109340 26908 109396
rect 26964 109340 26974 109396
rect 0 109228 980 109284
rect 1586 109228 1596 109284
rect 1652 109228 3220 109284
rect 3714 109228 3724 109284
rect 3780 109228 4172 109284
rect 4228 109228 4238 109284
rect 4834 109228 4844 109284
rect 4900 109228 4910 109284
rect 5730 109228 5740 109284
rect 5796 109228 5852 109284
rect 5908 109228 5918 109284
rect 8642 109228 8652 109284
rect 8708 109228 12124 109284
rect 12180 109228 12190 109284
rect 20626 109228 20636 109284
rect 20692 109228 23044 109284
rect 0 109200 112 109228
rect 3164 109172 3220 109228
rect 4844 109172 4900 109228
rect 22988 109172 23044 109228
rect 3164 109116 4900 109172
rect 5282 109116 5292 109172
rect 5348 109116 8316 109172
rect 8372 109116 8382 109172
rect 9510 109116 9548 109172
rect 9604 109116 9614 109172
rect 10210 109116 10220 109172
rect 10276 109116 10780 109172
rect 10836 109116 10846 109172
rect 11666 109116 11676 109172
rect 11732 109116 17388 109172
rect 17444 109116 17454 109172
rect 19366 109116 19404 109172
rect 19460 109116 19470 109172
rect 22988 109116 28028 109172
rect 28084 109116 28094 109172
rect 10780 109060 10836 109116
rect 2258 109004 2268 109060
rect 2324 109004 2604 109060
rect 2660 109004 2670 109060
rect 3490 109004 3500 109060
rect 3556 109004 4172 109060
rect 4228 109004 4238 109060
rect 5058 109004 5068 109060
rect 5124 109004 10444 109060
rect 10500 109004 10510 109060
rect 10780 109004 12908 109060
rect 12964 109004 12974 109060
rect 13234 109004 13244 109060
rect 13300 109004 19628 109060
rect 19684 109004 19694 109060
rect 25218 109004 25228 109060
rect 25284 109004 25340 109060
rect 25396 109004 26572 109060
rect 26628 109004 26638 109060
rect 27010 109004 27020 109060
rect 27076 109004 27132 109060
rect 27188 109004 28476 109060
rect 28532 109004 28542 109060
rect 4454 108948 4464 109004
rect 4520 108948 4568 109004
rect 4624 108948 4672 109004
rect 4728 108948 4738 109004
rect 24454 108948 24464 109004
rect 24520 108948 24568 109004
rect 24624 108948 24672 109004
rect 24728 108948 24738 109004
rect 3938 108892 3948 108948
rect 4004 108892 4284 108948
rect 4340 108892 4350 108948
rect 4834 108892 4844 108948
rect 4900 108892 8596 108948
rect 8978 108892 8988 108948
rect 9044 108892 9548 108948
rect 9604 108892 9614 108948
rect 10546 108892 10556 108948
rect 10612 108892 13468 108948
rect 13524 108892 13534 108948
rect 15222 108892 15260 108948
rect 15316 108892 15326 108948
rect 17266 108892 17276 108948
rect 17332 108892 17948 108948
rect 18004 108892 18014 108948
rect 19170 108892 19180 108948
rect 19236 108892 19740 108948
rect 19796 108892 19806 108948
rect 0 108836 112 108864
rect 0 108780 1764 108836
rect 4050 108780 4060 108836
rect 4116 108780 5068 108836
rect 5124 108780 5134 108836
rect 5404 108780 7084 108836
rect 7140 108780 7150 108836
rect 0 108752 112 108780
rect 1708 108500 1764 108780
rect 3266 108556 3276 108612
rect 3332 108556 3388 108724
rect 3444 108668 3454 108724
rect 3602 108668 3612 108724
rect 3668 108668 4844 108724
rect 4900 108668 4910 108724
rect 5404 108612 5460 108780
rect 8540 108724 8596 108892
rect 9202 108780 9212 108836
rect 9268 108780 20860 108836
rect 20916 108780 20926 108836
rect 26898 108780 26908 108836
rect 26964 108780 27020 108836
rect 27076 108780 27086 108836
rect 6738 108668 6748 108724
rect 6804 108668 8092 108724
rect 8148 108668 8158 108724
rect 8502 108668 8540 108724
rect 8596 108668 9380 108724
rect 9986 108668 9996 108724
rect 10052 108668 15372 108724
rect 15428 108668 15438 108724
rect 16146 108668 16156 108724
rect 16212 108668 30380 108724
rect 30436 108668 30446 108724
rect 4284 108556 5460 108612
rect 5618 108556 5628 108612
rect 5684 108556 6860 108612
rect 6916 108556 6926 108612
rect 8838 108556 8876 108612
rect 8932 108556 8942 108612
rect 4284 108500 4340 108556
rect 9324 108500 9380 108668
rect 9538 108556 9548 108612
rect 9604 108556 9884 108612
rect 9940 108556 9950 108612
rect 13906 108556 13916 108612
rect 13972 108556 13982 108612
rect 16818 108556 16828 108612
rect 16884 108556 17388 108612
rect 17444 108556 17454 108612
rect 19394 108556 19404 108612
rect 19460 108556 26236 108612
rect 26292 108556 26302 108612
rect 13916 108500 13972 108556
rect 31584 108500 31696 108528
rect 1708 108444 4340 108500
rect 4610 108444 4620 108500
rect 4676 108444 4956 108500
rect 5012 108444 7196 108500
rect 7252 108444 7262 108500
rect 7858 108444 7868 108500
rect 7924 108444 9100 108500
rect 9156 108444 9166 108500
rect 9324 108444 13972 108500
rect 15250 108444 15260 108500
rect 15316 108444 15372 108500
rect 15428 108444 15438 108500
rect 23426 108444 23436 108500
rect 23492 108444 25116 108500
rect 25172 108444 25182 108500
rect 26114 108444 26124 108500
rect 26180 108444 26348 108500
rect 26404 108444 27132 108500
rect 27188 108444 27198 108500
rect 30594 108444 30604 108500
rect 30660 108444 31696 108500
rect 31584 108416 31696 108444
rect 0 108388 112 108416
rect 0 108332 476 108388
rect 532 108332 542 108388
rect 0 108304 112 108332
rect 3266 108220 3276 108276
rect 3332 108220 3388 108388
rect 3444 108332 3454 108388
rect 3612 108332 10668 108388
rect 10724 108332 10734 108388
rect 10892 108332 11564 108388
rect 11620 108332 17724 108388
rect 17780 108332 17790 108388
rect 23650 108332 23660 108388
rect 23716 108332 27356 108388
rect 27412 108332 27422 108388
rect 3612 108164 3668 108332
rect 10892 108276 10948 108332
rect 4722 108220 4732 108276
rect 4788 108220 6076 108276
rect 6132 108220 6142 108276
rect 10434 108220 10444 108276
rect 10500 108220 10948 108276
rect 13570 108220 13580 108276
rect 13636 108220 15148 108276
rect 3794 108164 3804 108220
rect 3860 108164 3908 108220
rect 3964 108164 4012 108220
rect 4068 108164 4078 108220
rect 15092 108164 15148 108220
rect 23794 108164 23804 108220
rect 23860 108164 23908 108220
rect 23964 108164 24012 108220
rect 24068 108164 24078 108220
rect 3332 108108 3668 108164
rect 6290 108108 6300 108164
rect 6356 108108 7756 108164
rect 7812 108108 7822 108164
rect 9314 108108 9324 108164
rect 9380 108108 14028 108164
rect 14084 108108 14094 108164
rect 15092 108108 18172 108164
rect 18228 108108 18238 108164
rect 3332 108052 3388 108108
rect 1250 107996 1260 108052
rect 1316 107996 1326 108052
rect 2930 107996 2940 108052
rect 2996 107996 3388 108052
rect 3490 107996 3500 108052
rect 3556 107996 15708 108052
rect 15764 107996 15774 108052
rect 0 107940 112 107968
rect 1260 107940 1316 107996
rect 0 107884 868 107940
rect 1260 107884 5516 107940
rect 5572 107884 5740 107940
rect 5796 107884 5806 107940
rect 6262 107884 6300 107940
rect 6356 107884 6366 107940
rect 9846 107884 9884 107940
rect 9940 107884 9950 107940
rect 13906 107884 13916 107940
rect 13972 107884 14028 107940
rect 14084 107884 14094 107940
rect 25106 107884 25116 107940
rect 25172 107884 25228 107940
rect 25284 107884 25294 107940
rect 0 107856 112 107884
rect 812 107828 868 107884
rect 812 107772 1708 107828
rect 1764 107772 1774 107828
rect 3266 107772 3276 107828
rect 3332 107772 3500 107828
rect 3556 107772 3566 107828
rect 5170 107772 5180 107828
rect 5236 107772 5292 107828
rect 5348 107772 5358 107828
rect 9286 107772 9324 107828
rect 9380 107772 9390 107828
rect 9762 107772 9772 107828
rect 9828 107772 9996 107828
rect 10052 107772 10062 107828
rect 10658 107772 10668 107828
rect 10724 107772 11004 107828
rect 11060 107772 11340 107828
rect 11396 107772 11406 107828
rect 13430 107772 13468 107828
rect 13524 107772 13534 107828
rect 13906 107772 13916 107828
rect 13972 107772 14140 107828
rect 14196 107772 14206 107828
rect 14578 107772 14588 107828
rect 14644 107772 16828 107828
rect 16884 107772 16894 107828
rect 2258 107660 2268 107716
rect 2324 107660 7084 107716
rect 7140 107660 7150 107716
rect 7858 107660 7868 107716
rect 7924 107660 10444 107716
rect 10500 107660 10510 107716
rect 13682 107660 13692 107716
rect 13748 107660 15036 107716
rect 15092 107660 15102 107716
rect 4274 107548 4284 107604
rect 4340 107548 4396 107604
rect 4452 107548 4462 107604
rect 6402 107548 6412 107604
rect 6468 107548 7308 107604
rect 7364 107548 7374 107604
rect 8754 107548 8764 107604
rect 8820 107548 11340 107604
rect 11396 107548 12012 107604
rect 12068 107548 12078 107604
rect 12786 107548 12796 107604
rect 12852 107548 13804 107604
rect 13860 107548 13870 107604
rect 14018 107548 14028 107604
rect 14084 107548 14700 107604
rect 14756 107548 14812 107604
rect 14868 107548 14878 107604
rect 15026 107548 15036 107604
rect 15092 107548 15932 107604
rect 15988 107548 15998 107604
rect 20066 107548 20076 107604
rect 20132 107548 26796 107604
rect 26852 107548 26862 107604
rect 0 107492 112 107520
rect 0 107436 4340 107492
rect 6066 107436 6076 107492
rect 6132 107436 13356 107492
rect 13412 107436 13422 107492
rect 14018 107436 14028 107492
rect 14084 107436 14364 107492
rect 14420 107436 14430 107492
rect 14690 107436 14700 107492
rect 14756 107436 14812 107492
rect 14868 107436 14878 107492
rect 0 107408 112 107436
rect 1586 107324 1596 107380
rect 1652 107324 3612 107380
rect 3668 107324 3678 107380
rect 4284 107268 4340 107436
rect 4454 107380 4464 107436
rect 4520 107380 4568 107436
rect 4624 107380 4672 107436
rect 4728 107380 4738 107436
rect 24454 107380 24464 107436
rect 24520 107380 24568 107436
rect 24624 107380 24672 107436
rect 24728 107380 24738 107436
rect 31584 107380 31696 107408
rect 5170 107324 5180 107380
rect 5236 107324 11788 107380
rect 11844 107324 11854 107380
rect 13122 107324 13132 107380
rect 13188 107324 22428 107380
rect 22484 107324 22494 107380
rect 30594 107324 30604 107380
rect 30660 107324 31696 107380
rect 31584 107296 31696 107324
rect 4284 107212 12684 107268
rect 12740 107212 15148 107268
rect 15092 107156 15148 107212
rect 3490 107100 3500 107156
rect 3556 107100 5404 107156
rect 5460 107100 5470 107156
rect 7298 107100 7308 107156
rect 7364 107100 11340 107156
rect 11396 107100 11406 107156
rect 15092 107100 17500 107156
rect 17556 107100 17566 107156
rect 0 107044 112 107072
rect 0 106988 2380 107044
rect 2436 106988 2446 107044
rect 3266 106988 3276 107044
rect 3332 106988 3612 107044
rect 3668 106988 3678 107044
rect 4722 106988 4732 107044
rect 4788 106988 16828 107044
rect 16884 106988 16894 107044
rect 0 106960 112 106988
rect 2370 106876 2380 106932
rect 2436 106876 4620 106932
rect 4676 106876 4686 106932
rect 7298 106876 7308 106932
rect 7364 106876 7756 106932
rect 7812 106876 7822 106932
rect 8278 106876 8316 106932
rect 8372 106876 8382 106932
rect 8754 106876 8764 106932
rect 8820 106876 8876 106932
rect 8932 106876 8942 106932
rect 9510 106876 9548 106932
rect 9604 106876 9614 106932
rect 10742 106876 10780 106932
rect 10836 106876 10846 106932
rect 14550 106876 14588 106932
rect 14644 106876 14654 106932
rect 21298 106876 21308 106932
rect 21364 106876 25116 106932
rect 25172 106876 25182 106932
rect 3378 106764 3388 106820
rect 3444 106764 8540 106820
rect 8596 106764 8606 106820
rect 12898 106764 12908 106820
rect 12964 106764 14476 106820
rect 14532 106764 18396 106820
rect 18452 106764 18462 106820
rect 5506 106652 5516 106708
rect 5572 106652 6748 106708
rect 6804 106652 17948 106708
rect 18004 106652 18014 106708
rect 18722 106652 18732 106708
rect 18788 106652 20188 106708
rect 20244 106652 20254 106708
rect 0 106596 112 106624
rect 3794 106596 3804 106652
rect 3860 106596 3908 106652
rect 3964 106596 4012 106652
rect 4068 106596 4078 106652
rect 23794 106596 23804 106652
rect 23860 106596 23908 106652
rect 23964 106596 24012 106652
rect 24068 106596 24078 106652
rect 0 106540 1372 106596
rect 1428 106540 1596 106596
rect 1652 106540 1662 106596
rect 5394 106540 5404 106596
rect 5460 106540 6300 106596
rect 6356 106540 6366 106596
rect 11778 106540 11788 106596
rect 11844 106540 13356 106596
rect 13412 106540 13422 106596
rect 0 106512 112 106540
rect 2118 106428 2156 106484
rect 2212 106428 2222 106484
rect 2370 106428 2380 106484
rect 2436 106428 2716 106484
rect 2772 106428 2782 106484
rect 2930 106428 2940 106484
rect 2996 106428 11564 106484
rect 11620 106428 11630 106484
rect 13010 106428 13020 106484
rect 13076 106428 14028 106484
rect 14084 106428 17612 106484
rect 17668 106428 17678 106484
rect 18610 106428 18620 106484
rect 18676 106428 19852 106484
rect 19908 106428 19918 106484
rect 1922 106316 1932 106372
rect 1988 106316 3892 106372
rect 4498 106316 4508 106372
rect 4564 106316 15148 106372
rect 15204 106316 15214 106372
rect 19180 106316 23100 106372
rect 23156 106316 23166 106372
rect 3836 106260 3892 106316
rect 354 106204 364 106260
rect 420 106204 1260 106260
rect 1316 106204 1820 106260
rect 1876 106204 1886 106260
rect 2034 106204 2044 106260
rect 2100 106204 2156 106260
rect 2212 106204 2828 106260
rect 2884 106204 2894 106260
rect 3042 106204 3052 106260
rect 3108 106204 3612 106260
rect 3668 106204 3678 106260
rect 3836 106204 6468 106260
rect 7634 106204 7644 106260
rect 7700 106204 8428 106260
rect 8484 106204 13020 106260
rect 13076 106204 13086 106260
rect 13234 106204 13244 106260
rect 13300 106204 16716 106260
rect 16772 106204 18508 106260
rect 18564 106204 18574 106260
rect 0 106148 112 106176
rect 0 106092 1484 106148
rect 1540 106092 1550 106148
rect 2706 106092 2716 106148
rect 2772 106092 5516 106148
rect 5572 106092 5582 106148
rect 0 106064 112 106092
rect 1922 105980 1932 106036
rect 1988 105980 3276 106036
rect 3332 105980 3342 106036
rect 4162 105980 4172 106036
rect 4228 105980 4396 106036
rect 4452 105980 4462 106036
rect 2146 105868 2156 105924
rect 2212 105868 2604 105924
rect 2660 105868 2670 105924
rect 3490 105868 3500 105924
rect 3556 105868 4284 105924
rect 4340 105868 4350 105924
rect 5730 105868 5740 105924
rect 5796 105868 5964 105924
rect 6020 105868 6030 105924
rect 4454 105812 4464 105868
rect 4520 105812 4568 105868
rect 4624 105812 4672 105868
rect 4728 105812 4738 105868
rect 6412 105812 6468 106204
rect 19180 106148 19236 106316
rect 31584 106260 31696 106288
rect 21746 106204 21756 106260
rect 21812 106204 26124 106260
rect 26180 106204 26190 106260
rect 30594 106204 30604 106260
rect 30660 106204 31696 106260
rect 31584 106176 31696 106204
rect 7158 106092 7196 106148
rect 7252 106092 7262 106148
rect 9986 106092 9996 106148
rect 10052 106092 19236 106148
rect 22642 106092 22652 106148
rect 22708 106092 26236 106148
rect 26292 106092 26302 106148
rect 6962 105980 6972 106036
rect 7028 105980 7532 106036
rect 7588 105980 7598 106036
rect 10770 105980 10780 106036
rect 10836 105980 13132 106036
rect 13188 105980 13198 106036
rect 13458 105980 13468 106036
rect 13524 105980 29596 106036
rect 29652 105980 29662 106036
rect 6626 105868 6636 105924
rect 6692 105868 8316 105924
rect 8372 105868 8382 105924
rect 11218 105868 11228 105924
rect 11284 105868 13244 105924
rect 13300 105868 13310 105924
rect 24454 105812 24464 105868
rect 24520 105812 24568 105868
rect 24624 105812 24672 105868
rect 24728 105812 24738 105868
rect 1708 105756 4060 105812
rect 4116 105756 4126 105812
rect 6412 105756 6972 105812
rect 7028 105756 7038 105812
rect 9090 105756 9100 105812
rect 9156 105756 13132 105812
rect 13188 105756 13198 105812
rect 13356 105756 24220 105812
rect 24276 105756 24286 105812
rect 0 105700 112 105728
rect 1708 105700 1764 105756
rect 13356 105700 13412 105756
rect 0 105644 1764 105700
rect 2258 105644 2268 105700
rect 2324 105644 9044 105700
rect 9202 105644 9212 105700
rect 9268 105644 13412 105700
rect 13794 105644 13804 105700
rect 13860 105644 17948 105700
rect 18004 105644 18014 105700
rect 0 105616 112 105644
rect 2706 105532 2716 105588
rect 2772 105532 4732 105588
rect 4788 105532 4798 105588
rect 6962 105532 6972 105588
rect 7028 105532 8092 105588
rect 8148 105532 8158 105588
rect 8988 105476 9044 105644
rect 13458 105532 13468 105588
rect 13524 105532 14924 105588
rect 14980 105532 17948 105588
rect 18004 105532 18014 105588
rect 19030 105532 19068 105588
rect 19124 105532 19134 105588
rect 19394 105532 19404 105588
rect 19460 105532 30268 105588
rect 30324 105532 30334 105588
rect 2034 105420 2044 105476
rect 2100 105420 3388 105476
rect 3602 105420 3612 105476
rect 3668 105420 3836 105476
rect 3892 105420 3902 105476
rect 4050 105420 4060 105476
rect 4116 105420 6972 105476
rect 7028 105420 7038 105476
rect 8988 105420 21420 105476
rect 21476 105420 21486 105476
rect 3332 105364 3388 105420
rect 3332 105308 13804 105364
rect 13860 105308 13870 105364
rect 0 105252 112 105280
rect 0 105196 2716 105252
rect 2772 105196 3164 105252
rect 3220 105196 3230 105252
rect 3332 105196 4228 105252
rect 4498 105196 4508 105252
rect 4564 105196 5068 105252
rect 5124 105196 5134 105252
rect 5282 105196 5292 105252
rect 5348 105196 5516 105252
rect 5572 105196 5582 105252
rect 13570 105196 13580 105252
rect 13636 105196 13692 105252
rect 13748 105196 14364 105252
rect 14420 105196 16604 105252
rect 16660 105196 16670 105252
rect 17154 105196 17164 105252
rect 17220 105196 19068 105252
rect 19124 105196 19134 105252
rect 0 105168 112 105196
rect 3332 105028 3388 105196
rect 4172 105140 4228 105196
rect 31584 105140 31696 105168
rect 4172 105084 7980 105140
rect 8036 105084 20076 105140
rect 20132 105084 20142 105140
rect 30594 105084 30604 105140
rect 30660 105084 31696 105140
rect 3794 105028 3804 105084
rect 3860 105028 3908 105084
rect 3964 105028 4012 105084
rect 4068 105028 4078 105084
rect 23794 105028 23804 105084
rect 23860 105028 23908 105084
rect 23964 105028 24012 105084
rect 24068 105028 24078 105084
rect 31584 105056 31696 105084
rect 1708 104972 3388 105028
rect 5282 104972 5292 105028
rect 5348 104972 6860 105028
rect 6916 104972 6926 105028
rect 8082 104972 8092 105028
rect 8148 104972 14252 105028
rect 14308 104972 15820 105028
rect 15876 104972 15886 105028
rect 914 104860 924 104916
rect 980 104860 1260 104916
rect 1316 104860 1326 104916
rect 0 104804 112 104832
rect 1708 104804 1764 104972
rect 0 104748 1764 104804
rect 2492 104860 22876 104916
rect 22932 104860 22942 104916
rect 0 104720 112 104748
rect 2492 104692 2548 104860
rect 4050 104748 4060 104804
rect 4116 104748 4620 104804
rect 4676 104748 4686 104804
rect 10994 104748 11004 104804
rect 11060 104748 11452 104804
rect 11508 104748 11518 104804
rect 1586 104636 1596 104692
rect 1652 104636 2548 104692
rect 2604 104636 13468 104692
rect 13524 104636 13534 104692
rect 2604 104580 2660 104636
rect 1362 104524 1372 104580
rect 1428 104524 1708 104580
rect 1764 104524 2660 104580
rect 3714 104524 3724 104580
rect 3780 104524 5572 104580
rect 6962 104524 6972 104580
rect 7028 104524 8540 104580
rect 8596 104524 8606 104580
rect 12338 104524 12348 104580
rect 12404 104524 16156 104580
rect 16212 104524 16222 104580
rect 5516 104468 5572 104524
rect 4162 104412 4172 104468
rect 4228 104412 4844 104468
rect 4900 104412 4910 104468
rect 5516 104412 7420 104468
rect 7476 104412 7486 104468
rect 8054 104412 8092 104468
rect 8148 104412 9324 104468
rect 9380 104412 9390 104468
rect 9622 104412 9660 104468
rect 9716 104412 9726 104468
rect 11106 104412 11116 104468
rect 11172 104412 11340 104468
rect 11396 104412 11452 104468
rect 11508 104412 11518 104468
rect 11666 104412 11676 104468
rect 11732 104412 11770 104468
rect 16258 104412 16268 104468
rect 16324 104412 16716 104468
rect 16772 104412 16782 104468
rect 18162 104412 18172 104468
rect 18228 104412 19516 104468
rect 19572 104412 19582 104468
rect 0 104356 112 104384
rect 0 104300 2268 104356
rect 2324 104300 2334 104356
rect 7298 104300 7308 104356
rect 7364 104300 21868 104356
rect 21924 104300 21934 104356
rect 0 104272 112 104300
rect 4454 104244 4464 104300
rect 4520 104244 4568 104300
rect 4624 104244 4672 104300
rect 4728 104244 4738 104300
rect 24454 104244 24464 104300
rect 24520 104244 24568 104300
rect 24624 104244 24672 104300
rect 24728 104244 24738 104300
rect 2566 104188 2604 104244
rect 2660 104188 2670 104244
rect 4834 104188 4844 104244
rect 4900 104188 4910 104244
rect 6038 104188 6076 104244
rect 6132 104188 6142 104244
rect 6738 104188 6748 104244
rect 6804 104188 7420 104244
rect 7476 104188 17724 104244
rect 17780 104188 19068 104244
rect 19124 104188 19134 104244
rect 4844 104132 4900 104188
rect 2146 104076 2156 104132
rect 2212 104076 4004 104132
rect 4162 104076 4172 104132
rect 4228 104076 4900 104132
rect 6178 104076 6188 104132
rect 6244 104076 7140 104132
rect 11862 104076 11900 104132
rect 11956 104076 11966 104132
rect 13458 104076 13468 104132
rect 13524 104076 14700 104132
rect 14756 104076 16828 104132
rect 16884 104076 16894 104132
rect 20850 104076 20860 104132
rect 20916 104076 30268 104132
rect 30324 104076 30334 104132
rect 3948 104020 4004 104076
rect 7084 104020 7140 104076
rect 31584 104020 31696 104048
rect 1558 103964 1596 104020
rect 1652 103964 1662 104020
rect 2594 103964 2604 104020
rect 2660 103964 2716 104020
rect 2772 103964 2782 104020
rect 3948 103964 5404 104020
rect 5460 103964 5470 104020
rect 5954 103964 5964 104020
rect 6020 103964 6412 104020
rect 6468 103964 6478 104020
rect 7074 103964 7084 104020
rect 7140 103964 8092 104020
rect 8148 103964 8158 104020
rect 11666 103964 11676 104020
rect 11732 103964 15260 104020
rect 15316 103964 15326 104020
rect 18946 103964 18956 104020
rect 19012 103964 19628 104020
rect 19684 103964 19694 104020
rect 30594 103964 30604 104020
rect 30660 103964 31696 104020
rect 31584 103936 31696 103964
rect 0 103908 112 103936
rect 0 103852 1204 103908
rect 1362 103852 1372 103908
rect 1428 103852 7308 103908
rect 7364 103852 7374 103908
rect 11442 103852 11452 103908
rect 11508 103852 11676 103908
rect 11732 103852 11742 103908
rect 12002 103852 12012 103908
rect 12068 103852 15596 103908
rect 15652 103852 15662 103908
rect 0 103824 112 103852
rect 1148 103796 1204 103852
rect 1148 103740 2604 103796
rect 2660 103740 2670 103796
rect 4386 103740 4396 103796
rect 4452 103740 5068 103796
rect 5124 103740 6748 103796
rect 6804 103740 9772 103796
rect 9828 103740 11900 103796
rect 11956 103740 12908 103796
rect 12964 103740 12974 103796
rect 13682 103740 13692 103796
rect 13748 103740 14700 103796
rect 14756 103740 14766 103796
rect 15922 103740 15932 103796
rect 15988 103740 19964 103796
rect 20020 103740 20300 103796
rect 20356 103740 20366 103796
rect 3612 103628 4228 103684
rect 5394 103628 5404 103684
rect 5460 103628 6636 103684
rect 6692 103628 10108 103684
rect 10164 103628 10780 103684
rect 10836 103628 10846 103684
rect 11218 103628 11228 103684
rect 11284 103628 11676 103684
rect 11732 103628 11742 103684
rect 12114 103628 12124 103684
rect 12180 103628 13132 103684
rect 13188 103628 15372 103684
rect 15428 103628 15438 103684
rect 0 103460 112 103488
rect 3612 103460 3668 103628
rect 3794 103460 3804 103516
rect 3860 103460 3908 103516
rect 3964 103460 4012 103516
rect 4068 103460 4078 103516
rect 4172 103460 4228 103628
rect 5730 103516 5740 103572
rect 5796 103516 10444 103572
rect 10500 103516 10510 103572
rect 11732 103516 13580 103572
rect 13636 103516 17836 103572
rect 17892 103516 17902 103572
rect 11732 103460 11788 103516
rect 23794 103460 23804 103516
rect 23860 103460 23908 103516
rect 23964 103460 24012 103516
rect 24068 103460 24078 103516
rect 0 103404 1932 103460
rect 1988 103404 3668 103460
rect 4172 103404 11788 103460
rect 0 103376 112 103404
rect 3714 103292 3724 103348
rect 3780 103292 5068 103348
rect 5124 103292 5134 103348
rect 5730 103292 5740 103348
rect 5796 103292 5806 103348
rect 6290 103292 6300 103348
rect 6356 103292 8876 103348
rect 8932 103292 13804 103348
rect 13860 103292 13870 103348
rect 1026 103180 1036 103236
rect 1092 103180 3500 103236
rect 3556 103180 3948 103236
rect 4004 103180 4014 103236
rect 5740 103124 5796 103292
rect 11554 103180 11564 103236
rect 11620 103180 12908 103236
rect 12964 103180 12974 103236
rect 14130 103180 14140 103236
rect 14196 103180 17276 103236
rect 17332 103180 17342 103236
rect 2146 103068 2156 103124
rect 2212 103068 3836 103124
rect 3892 103068 3902 103124
rect 4172 103068 5796 103124
rect 6178 103068 6188 103124
rect 6244 103068 6748 103124
rect 6804 103068 6814 103124
rect 9286 103068 9324 103124
rect 9380 103068 9390 103124
rect 11442 103068 11452 103124
rect 11508 103068 11676 103124
rect 11732 103068 11742 103124
rect 16594 103068 16604 103124
rect 16660 103068 17052 103124
rect 17108 103068 17118 103124
rect 0 103012 112 103040
rect 4172 103012 4228 103068
rect 0 102956 4228 103012
rect 4386 102956 4396 103012
rect 4452 102956 5740 103012
rect 5796 102956 5806 103012
rect 0 102928 112 102956
rect 31584 102900 31696 102928
rect 1026 102844 1036 102900
rect 1092 102844 2380 102900
rect 2436 102844 4732 102900
rect 4788 102844 4798 102900
rect 5282 102844 5292 102900
rect 5348 102844 5628 102900
rect 5684 102844 5694 102900
rect 10434 102844 10444 102900
rect 10500 102844 10556 102900
rect 10612 102844 10622 102900
rect 16566 102844 16604 102900
rect 16660 102844 17724 102900
rect 17780 102844 17790 102900
rect 19506 102844 19516 102900
rect 19572 102844 30268 102900
rect 30324 102844 30334 102900
rect 30594 102844 30604 102900
rect 30660 102844 31696 102900
rect 31584 102816 31696 102844
rect 1474 102732 1484 102788
rect 1540 102732 1596 102788
rect 1652 102732 1662 102788
rect 3826 102732 3836 102788
rect 3892 102732 4060 102788
rect 4116 102732 4126 102788
rect 4844 102732 8092 102788
rect 8148 102732 8158 102788
rect 4454 102676 4464 102732
rect 4520 102676 4568 102732
rect 4624 102676 4672 102732
rect 4728 102676 4738 102732
rect 1708 102620 4340 102676
rect 0 102564 112 102592
rect 1708 102564 1764 102620
rect 0 102508 1764 102564
rect 4284 102564 4340 102620
rect 4844 102564 4900 102732
rect 24454 102676 24464 102732
rect 24520 102676 24568 102732
rect 24624 102676 24672 102732
rect 24728 102676 24738 102732
rect 6402 102620 6412 102676
rect 6468 102620 6478 102676
rect 4284 102508 4900 102564
rect 5394 102508 5404 102564
rect 5460 102508 5470 102564
rect 0 102480 112 102508
rect 5404 102452 5460 102508
rect 6412 102452 6468 102620
rect 9650 102508 9660 102564
rect 9716 102508 10668 102564
rect 10724 102508 10734 102564
rect 13244 102508 13692 102564
rect 13748 102508 13758 102564
rect 13244 102452 13300 102508
rect 1362 102396 1372 102452
rect 1428 102396 1708 102452
rect 1764 102396 1774 102452
rect 3266 102396 3276 102452
rect 3332 102396 5068 102452
rect 5124 102396 5134 102452
rect 5404 102396 5852 102452
rect 5908 102396 5918 102452
rect 6412 102396 8988 102452
rect 9044 102396 9054 102452
rect 10892 102396 12684 102452
rect 12740 102396 13300 102452
rect 13458 102396 13468 102452
rect 13524 102396 13916 102452
rect 13972 102396 13982 102452
rect 17602 102396 17612 102452
rect 17668 102396 30268 102452
rect 30324 102396 30334 102452
rect 1138 102284 1148 102340
rect 1204 102284 6076 102340
rect 6132 102284 6142 102340
rect 7186 102284 7196 102340
rect 7252 102284 8652 102340
rect 8708 102284 8718 102340
rect 10892 102228 10948 102396
rect 14578 102284 14588 102340
rect 14644 102284 15260 102340
rect 15316 102284 15326 102340
rect 802 102172 812 102228
rect 868 102172 5404 102228
rect 5460 102172 5470 102228
rect 5842 102172 5852 102228
rect 5908 102172 10892 102228
rect 10948 102172 10958 102228
rect 0 102116 112 102144
rect 0 102060 1876 102116
rect 2930 102060 2940 102116
rect 2996 102060 7644 102116
rect 7700 102060 7710 102116
rect 10994 102060 11004 102116
rect 11060 102060 17276 102116
rect 17332 102060 17342 102116
rect 0 102032 112 102060
rect 0 101668 112 101696
rect 0 101612 1764 101668
rect 0 101584 112 101612
rect 0 101220 112 101248
rect 1708 101220 1764 101612
rect 1820 101332 1876 102060
rect 5282 101948 5292 102004
rect 5348 101948 17388 102004
rect 17444 101948 17454 102004
rect 3794 101892 3804 101948
rect 3860 101892 3908 101948
rect 3964 101892 4012 101948
rect 4068 101892 4078 101948
rect 23794 101892 23804 101948
rect 23860 101892 23908 101948
rect 23964 101892 24012 101948
rect 24068 101892 24078 101948
rect 5170 101836 5180 101892
rect 5236 101836 10444 101892
rect 10500 101836 10510 101892
rect 12450 101836 12460 101892
rect 12516 101836 13244 101892
rect 13300 101836 13310 101892
rect 31584 101780 31696 101808
rect 2930 101724 2940 101780
rect 2996 101724 18844 101780
rect 18900 101724 18910 101780
rect 30594 101724 30604 101780
rect 30660 101724 31696 101780
rect 31584 101696 31696 101724
rect 3332 101612 14140 101668
rect 14196 101612 14206 101668
rect 3332 101332 3388 101612
rect 5394 101500 5404 101556
rect 5460 101500 6412 101556
rect 6468 101500 6478 101556
rect 3602 101388 3612 101444
rect 3668 101388 3678 101444
rect 4386 101388 4396 101444
rect 4452 101388 4844 101444
rect 4900 101388 4910 101444
rect 5394 101388 5404 101444
rect 5460 101388 5740 101444
rect 5796 101388 5806 101444
rect 6066 101388 6076 101444
rect 6132 101388 10108 101444
rect 10164 101388 10174 101444
rect 1820 101276 3388 101332
rect 3612 101332 3668 101388
rect 12684 101332 12740 101612
rect 12898 101500 12908 101556
rect 12964 101500 13580 101556
rect 13636 101500 13646 101556
rect 14914 101500 14924 101556
rect 14980 101500 15484 101556
rect 15540 101500 15550 101556
rect 13458 101388 13468 101444
rect 13524 101388 15260 101444
rect 15316 101388 15326 101444
rect 3612 101276 5292 101332
rect 5348 101276 5358 101332
rect 12684 101276 13580 101332
rect 13636 101276 13646 101332
rect 0 101164 1036 101220
rect 1092 101164 1102 101220
rect 1708 101164 3612 101220
rect 3668 101164 3678 101220
rect 5506 101164 5516 101220
rect 5572 101164 6076 101220
rect 6132 101164 6142 101220
rect 6626 101164 6636 101220
rect 6692 101164 17388 101220
rect 17444 101164 17454 101220
rect 0 101136 112 101164
rect 4454 101108 4464 101164
rect 4520 101108 4568 101164
rect 4624 101108 4672 101164
rect 4728 101108 4738 101164
rect 24454 101108 24464 101164
rect 24520 101108 24568 101164
rect 24624 101108 24672 101164
rect 24728 101108 24738 101164
rect 10098 101052 10108 101108
rect 10164 101052 11004 101108
rect 11060 101052 11070 101108
rect 11330 101052 11340 101108
rect 11396 101052 14924 101108
rect 14980 101052 18508 101108
rect 18564 101052 18574 101108
rect 2342 100940 2380 100996
rect 2436 100940 2446 100996
rect 4050 100940 4060 100996
rect 4116 100940 21084 100996
rect 21140 100940 21150 100996
rect 9538 100828 9548 100884
rect 9604 100828 10332 100884
rect 10388 100828 11116 100884
rect 11172 100828 11182 100884
rect 12338 100828 12348 100884
rect 12404 100828 13692 100884
rect 13748 100828 14028 100884
rect 14084 100828 14094 100884
rect 0 100772 112 100800
rect 0 100716 1092 100772
rect 1250 100716 1260 100772
rect 1316 100716 2380 100772
rect 2436 100716 2828 100772
rect 2884 100716 2894 100772
rect 3490 100716 3500 100772
rect 3556 100716 3836 100772
rect 3892 100716 3902 100772
rect 7270 100716 7308 100772
rect 7364 100716 7374 100772
rect 8194 100716 8204 100772
rect 8260 100716 9884 100772
rect 9940 100716 9950 100772
rect 14242 100716 14252 100772
rect 14308 100716 17276 100772
rect 17332 100716 17342 100772
rect 17826 100716 17836 100772
rect 17892 100716 29484 100772
rect 29540 100716 29550 100772
rect 0 100688 112 100716
rect 1036 100660 1092 100716
rect 31584 100660 31696 100688
rect 1036 100604 2716 100660
rect 2772 100604 2782 100660
rect 6626 100604 6636 100660
rect 6692 100604 16940 100660
rect 16996 100604 17006 100660
rect 30594 100604 30604 100660
rect 30660 100604 31696 100660
rect 31584 100576 31696 100604
rect 578 100492 588 100548
rect 644 100492 1260 100548
rect 1316 100492 1326 100548
rect 3602 100492 3612 100548
rect 3668 100492 5516 100548
rect 5572 100492 5582 100548
rect 6178 100492 6188 100548
rect 6244 100492 7420 100548
rect 7476 100492 7486 100548
rect 8642 100492 8652 100548
rect 8708 100492 9548 100548
rect 9604 100492 9614 100548
rect 17266 100492 17276 100548
rect 17332 100492 18060 100548
rect 18116 100492 18126 100548
rect 5618 100380 5628 100436
rect 5684 100380 7196 100436
rect 7252 100380 7262 100436
rect 7420 100380 16828 100436
rect 16884 100380 16894 100436
rect 0 100324 112 100352
rect 3794 100324 3804 100380
rect 3860 100324 3908 100380
rect 3964 100324 4012 100380
rect 4068 100324 4078 100380
rect 0 100268 1764 100324
rect 5058 100268 5068 100324
rect 5124 100268 5180 100324
rect 5236 100268 5404 100324
rect 5460 100268 5470 100324
rect 0 100240 112 100268
rect 1708 100100 1764 100268
rect 7420 100212 7476 100380
rect 23794 100324 23804 100380
rect 23860 100324 23908 100380
rect 23964 100324 24012 100380
rect 24068 100324 24078 100380
rect 7634 100268 7644 100324
rect 7700 100268 20972 100324
rect 21028 100268 21038 100324
rect 2930 100156 2940 100212
rect 2996 100156 7476 100212
rect 9426 100156 9436 100212
rect 9492 100156 9996 100212
rect 10052 100156 10062 100212
rect 10322 100156 10332 100212
rect 10388 100156 10668 100212
rect 10724 100156 10734 100212
rect 13122 100156 13132 100212
rect 13188 100156 13356 100212
rect 13412 100156 13422 100212
rect 13906 100156 13916 100212
rect 13972 100156 14476 100212
rect 14532 100156 14542 100212
rect 15092 100156 17836 100212
rect 17892 100156 17902 100212
rect 15092 100100 15148 100156
rect 1708 100044 3388 100100
rect 4050 100044 4060 100100
rect 4116 100044 15148 100100
rect 3332 99988 3388 100044
rect 242 99932 252 99988
rect 308 99932 1260 99988
rect 1316 99932 1326 99988
rect 3332 99932 5180 99988
rect 5236 99932 5246 99988
rect 8082 99932 8092 99988
rect 8148 99932 9324 99988
rect 9380 99932 10220 99988
rect 10276 99932 10286 99988
rect 10658 99932 10668 99988
rect 10724 99932 11452 99988
rect 11508 99932 11518 99988
rect 12114 99932 12124 99988
rect 12180 99932 14140 99988
rect 14196 99932 14206 99988
rect 0 99876 112 99904
rect 0 99820 4732 99876
rect 4788 99820 4798 99876
rect 9538 99820 9548 99876
rect 9604 99820 11228 99876
rect 11284 99820 13468 99876
rect 13524 99820 13534 99876
rect 17686 99820 17724 99876
rect 17780 99820 17790 99876
rect 0 99792 112 99820
rect 4172 99708 9884 99764
rect 9940 99708 9950 99764
rect 10098 99708 10108 99764
rect 10164 99708 10556 99764
rect 10612 99708 10622 99764
rect 11330 99708 11340 99764
rect 11396 99708 11406 99764
rect 17602 99708 17612 99764
rect 17668 99708 30268 99764
rect 30324 99708 30334 99764
rect 4172 99652 4228 99708
rect 11340 99652 11396 99708
rect 130 99596 140 99652
rect 196 99596 2156 99652
rect 2212 99596 2222 99652
rect 3602 99596 3612 99652
rect 3668 99596 4228 99652
rect 5842 99596 5852 99652
rect 5908 99596 6188 99652
rect 6244 99596 6254 99652
rect 9650 99596 9660 99652
rect 9716 99596 11396 99652
rect 4454 99540 4464 99596
rect 4520 99540 4568 99596
rect 4624 99540 4672 99596
rect 4728 99540 4738 99596
rect 24454 99540 24464 99596
rect 24520 99540 24568 99596
rect 24624 99540 24672 99596
rect 24728 99540 24738 99596
rect 31584 99540 31696 99568
rect 2818 99484 2828 99540
rect 2884 99484 3164 99540
rect 3220 99484 3230 99540
rect 7186 99484 7196 99540
rect 7252 99484 13916 99540
rect 13972 99484 14084 99540
rect 30594 99484 30604 99540
rect 30660 99484 31696 99540
rect 0 99428 112 99456
rect 14028 99428 14084 99484
rect 31584 99456 31696 99484
rect 0 99372 4284 99428
rect 4340 99372 11564 99428
rect 11620 99372 11900 99428
rect 11956 99372 11966 99428
rect 14018 99372 14028 99428
rect 14084 99372 18956 99428
rect 19012 99372 19022 99428
rect 0 99344 112 99372
rect 2258 99260 2268 99316
rect 2324 99260 3276 99316
rect 3332 99260 3342 99316
rect 3602 99260 3612 99316
rect 3668 99260 4396 99316
rect 4452 99260 9660 99316
rect 9716 99260 9726 99316
rect 19282 99260 19292 99316
rect 19348 99260 30268 99316
rect 30324 99260 30334 99316
rect 3154 99148 3164 99204
rect 3220 99148 3388 99204
rect 3444 99148 3454 99204
rect 5282 99148 5292 99204
rect 5348 99148 5964 99204
rect 6020 99148 6030 99204
rect 11666 99148 11676 99204
rect 11732 99148 12572 99204
rect 12628 99148 12908 99204
rect 12964 99148 12974 99204
rect 18834 99148 18844 99204
rect 18900 99148 19516 99204
rect 19572 99148 19964 99204
rect 20020 99148 20030 99204
rect 2370 99036 2380 99092
rect 2436 99036 6188 99092
rect 6244 99036 6254 99092
rect 19292 99036 29372 99092
rect 29428 99036 29438 99092
rect 0 98980 112 99008
rect 19292 98980 19348 99036
rect 0 98924 3276 98980
rect 3332 98924 3342 98980
rect 3612 98924 3836 98980
rect 3892 98924 3902 98980
rect 4274 98924 4284 98980
rect 4340 98924 5180 98980
rect 5236 98924 8204 98980
rect 8260 98924 8270 98980
rect 10108 98924 17388 98980
rect 17444 98924 19348 98980
rect 20066 98924 20076 98980
rect 20132 98924 29260 98980
rect 29316 98924 29326 98980
rect 0 98896 112 98924
rect 3612 98868 3668 98924
rect 1362 98812 1372 98868
rect 1428 98812 2268 98868
rect 2324 98812 3668 98868
rect 5058 98812 5068 98868
rect 5124 98812 6412 98868
rect 6468 98812 6478 98868
rect 7522 98812 7532 98868
rect 7588 98812 8092 98868
rect 8148 98812 8158 98868
rect 3794 98756 3804 98812
rect 3860 98756 3908 98812
rect 3964 98756 4012 98812
rect 4068 98756 4078 98812
rect 4386 98700 4396 98756
rect 4452 98700 6076 98756
rect 6132 98700 6142 98756
rect 6962 98700 6972 98756
rect 7028 98700 7308 98756
rect 7364 98700 7374 98756
rect 2370 98588 2380 98644
rect 2436 98588 5292 98644
rect 5348 98588 5358 98644
rect 0 98532 112 98560
rect 10108 98532 10164 98924
rect 10322 98812 10332 98868
rect 10388 98812 13020 98868
rect 13076 98812 13086 98868
rect 15708 98756 15764 98924
rect 18386 98812 18396 98868
rect 18452 98812 19852 98868
rect 19908 98812 19918 98868
rect 20290 98812 20300 98868
rect 20356 98812 21196 98868
rect 21252 98812 21262 98868
rect 23794 98756 23804 98812
rect 23860 98756 23908 98812
rect 23964 98756 24012 98812
rect 24068 98756 24078 98812
rect 15698 98700 15708 98756
rect 15764 98700 15774 98756
rect 10994 98588 11004 98644
rect 11060 98588 11228 98644
rect 11284 98588 13020 98644
rect 13076 98588 13086 98644
rect 0 98476 252 98532
rect 308 98476 318 98532
rect 690 98476 700 98532
rect 756 98476 10108 98532
rect 10164 98476 10174 98532
rect 12562 98476 12572 98532
rect 12628 98476 14364 98532
rect 14420 98476 14430 98532
rect 15474 98476 15484 98532
rect 15540 98476 16044 98532
rect 16100 98476 18844 98532
rect 18900 98476 18910 98532
rect 0 98448 112 98476
rect 31584 98420 31696 98448
rect 4722 98364 4732 98420
rect 4788 98364 4798 98420
rect 5282 98364 5292 98420
rect 5348 98364 7420 98420
rect 7476 98364 7486 98420
rect 18134 98364 18172 98420
rect 18228 98364 18238 98420
rect 18610 98364 18620 98420
rect 18676 98364 19292 98420
rect 19348 98364 19358 98420
rect 30594 98364 30604 98420
rect 30660 98364 31696 98420
rect 2370 98252 2380 98308
rect 2436 98252 2604 98308
rect 2660 98252 2670 98308
rect 4162 98252 4172 98308
rect 4228 98252 4396 98308
rect 4452 98252 4462 98308
rect 4732 98196 4788 98364
rect 31584 98336 31696 98364
rect 4946 98252 4956 98308
rect 5012 98252 5068 98308
rect 5124 98252 5134 98308
rect 5702 98252 5740 98308
rect 5796 98252 5806 98308
rect 6850 98252 6860 98308
rect 6916 98252 7980 98308
rect 8036 98252 8046 98308
rect 16118 98252 16156 98308
rect 16212 98252 16222 98308
rect 2258 98140 2268 98196
rect 2324 98140 2828 98196
rect 2884 98140 2894 98196
rect 3332 98140 5292 98196
rect 5348 98140 5358 98196
rect 6850 98140 6860 98196
rect 6916 98140 9548 98196
rect 9604 98140 9614 98196
rect 18274 98140 18284 98196
rect 18340 98140 19852 98196
rect 19908 98140 19918 98196
rect 0 98084 112 98112
rect 3332 98084 3388 98140
rect 0 98028 3388 98084
rect 6514 98028 6524 98084
rect 6580 98028 10276 98084
rect 14326 98028 14364 98084
rect 14420 98028 14430 98084
rect 14774 98028 14812 98084
rect 14868 98028 14878 98084
rect 0 98000 112 98028
rect 4454 97972 4464 98028
rect 4520 97972 4568 98028
rect 4624 97972 4672 98028
rect 4728 97972 4738 98028
rect 10220 97972 10276 98028
rect 24454 97972 24464 98028
rect 24520 97972 24568 98028
rect 24624 97972 24672 98028
rect 24728 97972 24738 98028
rect 10220 97916 11788 97972
rect 11844 97916 13692 97972
rect 13748 97916 15148 97972
rect 16370 97916 16380 97972
rect 16436 97916 17836 97972
rect 17892 97916 18060 97972
rect 18116 97916 18126 97972
rect 15092 97860 15148 97916
rect 466 97804 476 97860
rect 532 97804 1708 97860
rect 1764 97804 1774 97860
rect 4498 97804 4508 97860
rect 4564 97804 6524 97860
rect 6580 97804 14476 97860
rect 14532 97804 14542 97860
rect 15092 97804 20076 97860
rect 20132 97804 20142 97860
rect 4050 97692 4060 97748
rect 4116 97692 4956 97748
rect 5012 97692 5022 97748
rect 6178 97692 6188 97748
rect 6244 97692 7308 97748
rect 7364 97692 7374 97748
rect 7756 97692 10556 97748
rect 10612 97692 10622 97748
rect 14354 97692 14364 97748
rect 14420 97692 18396 97748
rect 18452 97692 22988 97748
rect 23044 97692 23054 97748
rect 0 97636 112 97664
rect 7756 97636 7812 97692
rect 0 97580 6412 97636
rect 6468 97580 6478 97636
rect 7410 97580 7420 97636
rect 7476 97580 7756 97636
rect 7812 97580 7822 97636
rect 8194 97580 8204 97636
rect 8260 97580 8652 97636
rect 8708 97580 9212 97636
rect 9268 97580 9278 97636
rect 11106 97580 11116 97636
rect 11172 97580 16940 97636
rect 16996 97580 17006 97636
rect 17154 97580 17164 97636
rect 17220 97580 18284 97636
rect 18340 97580 18350 97636
rect 0 97552 112 97580
rect 4498 97468 4508 97524
rect 4564 97468 4844 97524
rect 4900 97468 4910 97524
rect 6066 97468 6076 97524
rect 6132 97468 7084 97524
rect 7140 97468 7150 97524
rect 7634 97468 7644 97524
rect 7700 97468 8092 97524
rect 8148 97468 8158 97524
rect 13010 97468 13020 97524
rect 13076 97468 14476 97524
rect 14532 97468 14542 97524
rect 15922 97468 15932 97524
rect 15988 97468 16380 97524
rect 16436 97468 16446 97524
rect 16818 97468 16828 97524
rect 16884 97468 18732 97524
rect 18788 97468 18798 97524
rect 3332 97356 6244 97412
rect 7718 97356 7756 97412
rect 7812 97356 7822 97412
rect 9986 97356 9996 97412
rect 10052 97356 11340 97412
rect 11396 97356 11406 97412
rect 0 97188 112 97216
rect 3332 97188 3388 97356
rect 3794 97188 3804 97244
rect 3860 97188 3908 97244
rect 3964 97188 4012 97244
rect 4068 97188 4078 97244
rect 6188 97188 6244 97356
rect 31584 97300 31696 97328
rect 6402 97244 6412 97300
rect 6468 97244 8428 97300
rect 8484 97244 10332 97300
rect 10388 97244 10398 97300
rect 12114 97244 12124 97300
rect 12180 97244 12684 97300
rect 12740 97244 12908 97300
rect 12964 97244 12974 97300
rect 30594 97244 30604 97300
rect 30660 97244 31696 97300
rect 23794 97188 23804 97244
rect 23860 97188 23908 97244
rect 23964 97188 24012 97244
rect 24068 97188 24078 97244
rect 31584 97216 31696 97244
rect 0 97132 3388 97188
rect 6188 97132 7420 97188
rect 7476 97132 14364 97188
rect 14420 97132 14430 97188
rect 14578 97132 14588 97188
rect 14644 97132 14924 97188
rect 14980 97132 14990 97188
rect 0 97104 112 97132
rect 3266 97020 3276 97076
rect 3332 97020 12796 97076
rect 12852 97020 14700 97076
rect 14756 97020 14766 97076
rect 14924 97020 16716 97076
rect 16772 97020 19516 97076
rect 19572 97020 19582 97076
rect 14924 96964 14980 97020
rect 2146 96908 2156 96964
rect 2212 96908 3388 96964
rect 3490 96908 3500 96964
rect 3556 96908 5404 96964
rect 5460 96908 5516 96964
rect 5572 96908 5582 96964
rect 6626 96908 6636 96964
rect 6692 96908 13916 96964
rect 13972 96908 13982 96964
rect 14130 96908 14140 96964
rect 14196 96908 14980 96964
rect 3332 96852 3388 96908
rect 1586 96796 1596 96852
rect 1652 96796 2716 96852
rect 2772 96796 2782 96852
rect 3332 96796 8204 96852
rect 8260 96796 9884 96852
rect 9940 96796 9950 96852
rect 10882 96796 10892 96852
rect 10948 96796 11564 96852
rect 11620 96796 11630 96852
rect 12002 96796 12012 96852
rect 12068 96796 13692 96852
rect 13748 96796 13758 96852
rect 22194 96796 22204 96852
rect 22260 96796 29484 96852
rect 29540 96796 29550 96852
rect 0 96740 112 96768
rect 0 96684 3612 96740
rect 3668 96684 3678 96740
rect 6178 96684 6188 96740
rect 6244 96684 14140 96740
rect 14196 96684 14206 96740
rect 15484 96684 17836 96740
rect 17892 96684 17902 96740
rect 21746 96684 21756 96740
rect 21812 96684 22316 96740
rect 22372 96684 22382 96740
rect 0 96656 112 96684
rect 15484 96628 15540 96684
rect 3332 96572 10444 96628
rect 10500 96572 15540 96628
rect 15670 96572 15708 96628
rect 15764 96572 15774 96628
rect 21858 96572 21868 96628
rect 21924 96572 29484 96628
rect 29540 96572 29550 96628
rect 3332 96516 3388 96572
rect 21868 96516 21924 96572
rect 130 96460 140 96516
rect 196 96460 3388 96516
rect 5282 96460 5292 96516
rect 5348 96460 5740 96516
rect 5796 96460 5806 96516
rect 6402 96460 6412 96516
rect 6468 96460 18284 96516
rect 18340 96460 21924 96516
rect 4454 96404 4464 96460
rect 4520 96404 4568 96460
rect 4624 96404 4672 96460
rect 4728 96404 4738 96460
rect 24454 96404 24464 96460
rect 24520 96404 24568 96460
rect 24624 96404 24672 96460
rect 24728 96404 24738 96460
rect 2146 96348 2156 96404
rect 2212 96348 2940 96404
rect 2996 96348 3006 96404
rect 4946 96348 4956 96404
rect 5012 96348 7308 96404
rect 7364 96348 7374 96404
rect 11228 96348 15036 96404
rect 15092 96348 15102 96404
rect 15474 96348 15484 96404
rect 15540 96348 16492 96404
rect 16548 96348 16558 96404
rect 0 96292 112 96320
rect 11228 96292 11284 96348
rect 0 96236 1260 96292
rect 1316 96236 1326 96292
rect 2594 96236 2604 96292
rect 2660 96236 3164 96292
rect 3220 96236 11284 96292
rect 11442 96236 11452 96292
rect 11508 96236 12908 96292
rect 12964 96236 12974 96292
rect 13906 96236 13916 96292
rect 13972 96236 15932 96292
rect 15988 96236 19964 96292
rect 20020 96236 20030 96292
rect 0 96208 112 96236
rect 31584 96180 31696 96208
rect 1670 96124 1708 96180
rect 1764 96124 6412 96180
rect 6468 96124 6478 96180
rect 11666 96124 11676 96180
rect 11732 96124 13468 96180
rect 13524 96124 13534 96180
rect 15362 96124 15372 96180
rect 15428 96124 16492 96180
rect 16548 96124 17052 96180
rect 17108 96124 17118 96180
rect 17798 96124 17836 96180
rect 17892 96124 17902 96180
rect 18946 96124 18956 96180
rect 19012 96124 25676 96180
rect 25732 96124 25742 96180
rect 30594 96124 30604 96180
rect 30660 96124 31696 96180
rect 31584 96096 31696 96124
rect 3490 96012 3500 96068
rect 3556 96012 6748 96068
rect 6804 96012 7532 96068
rect 7588 96012 7598 96068
rect 10322 96012 10332 96068
rect 10388 96012 12460 96068
rect 12516 96012 12526 96068
rect 17714 96012 17724 96068
rect 17780 96012 18060 96068
rect 18116 96012 18172 96068
rect 18228 96012 18238 96068
rect 1362 95900 1372 95956
rect 1428 95900 1708 95956
rect 1764 95900 1774 95956
rect 2706 95900 2716 95956
rect 2772 95900 3500 95956
rect 3556 95900 3566 95956
rect 4610 95900 4620 95956
rect 4676 95900 5068 95956
rect 5124 95900 5134 95956
rect 14354 95900 14364 95956
rect 14420 95900 15260 95956
rect 15316 95900 15708 95956
rect 15764 95900 15774 95956
rect 18386 95900 18396 95956
rect 18452 95900 19516 95956
rect 19572 95900 20972 95956
rect 21028 95900 21756 95956
rect 21812 95900 21822 95956
rect 0 95844 112 95872
rect 0 95788 476 95844
rect 532 95788 542 95844
rect 1474 95788 1484 95844
rect 1540 95788 2380 95844
rect 2436 95788 2446 95844
rect 3602 95788 3612 95844
rect 3668 95788 5012 95844
rect 11778 95788 11788 95844
rect 11844 95788 13244 95844
rect 13300 95788 13310 95844
rect 14018 95788 14028 95844
rect 14084 95788 16828 95844
rect 16884 95788 16894 95844
rect 0 95760 112 95788
rect 4956 95732 5012 95788
rect 1922 95676 1932 95732
rect 1988 95676 3612 95732
rect 3668 95676 3678 95732
rect 4956 95676 8652 95732
rect 8708 95676 8718 95732
rect 8866 95676 8876 95732
rect 8932 95676 10444 95732
rect 10500 95676 10510 95732
rect 14018 95676 14028 95732
rect 14084 95676 17948 95732
rect 18004 95676 18014 95732
rect 3794 95620 3804 95676
rect 3860 95620 3908 95676
rect 3964 95620 4012 95676
rect 4068 95620 4078 95676
rect 23794 95620 23804 95676
rect 23860 95620 23908 95676
rect 23964 95620 24012 95676
rect 24068 95620 24078 95676
rect 7074 95564 7084 95620
rect 7140 95564 7308 95620
rect 7364 95564 7374 95620
rect 8530 95564 8540 95620
rect 8596 95564 9996 95620
rect 10052 95564 10062 95620
rect 5170 95452 5180 95508
rect 5236 95452 18956 95508
rect 19012 95452 19022 95508
rect 0 95396 112 95424
rect 0 95340 3612 95396
rect 3668 95340 3678 95396
rect 3948 95340 6076 95396
rect 6132 95340 6142 95396
rect 7074 95340 7084 95396
rect 7140 95340 10108 95396
rect 10164 95340 10174 95396
rect 10434 95340 10444 95396
rect 10500 95340 10780 95396
rect 10836 95340 10846 95396
rect 0 95312 112 95340
rect 3948 95284 4004 95340
rect 1474 95228 1484 95284
rect 1540 95228 2828 95284
rect 2884 95228 2894 95284
rect 3500 95228 4004 95284
rect 4162 95228 4172 95284
rect 4228 95228 4284 95284
rect 4340 95228 4350 95284
rect 8978 95228 8988 95284
rect 9044 95228 9548 95284
rect 9604 95228 9614 95284
rect 9874 95228 9884 95284
rect 9940 95228 11116 95284
rect 11172 95228 11182 95284
rect 19842 95228 19852 95284
rect 19908 95228 30380 95284
rect 30436 95228 30446 95284
rect 3500 95172 3556 95228
rect 2706 95116 2716 95172
rect 2772 95116 3500 95172
rect 3556 95116 3566 95172
rect 4050 95116 4060 95172
rect 4116 95116 4620 95172
rect 4676 95116 4686 95172
rect 6626 95116 6636 95172
rect 6692 95116 6972 95172
rect 7028 95116 7038 95172
rect 14130 95116 14140 95172
rect 14196 95116 14812 95172
rect 14868 95116 14878 95172
rect 31584 95060 31696 95088
rect 3332 95004 15148 95060
rect 23314 95004 23324 95060
rect 23380 95004 24892 95060
rect 24948 95004 24958 95060
rect 30594 95004 30604 95060
rect 30660 95004 31696 95060
rect 0 94948 112 94976
rect 3332 94948 3388 95004
rect 15092 94948 15148 95004
rect 31584 94976 31696 95004
rect 0 94892 3388 94948
rect 9090 94892 9100 94948
rect 9156 94892 14812 94948
rect 14868 94892 14878 94948
rect 15092 94892 20524 94948
rect 20580 94892 20590 94948
rect 0 94864 112 94892
rect 4454 94836 4464 94892
rect 4520 94836 4568 94892
rect 4624 94836 4672 94892
rect 4728 94836 4738 94892
rect 24454 94836 24464 94892
rect 24520 94836 24568 94892
rect 24624 94836 24672 94892
rect 24728 94836 24738 94892
rect 3490 94780 3500 94836
rect 3556 94780 4284 94836
rect 4340 94780 4350 94836
rect 8530 94780 8540 94836
rect 8596 94780 8764 94836
rect 8820 94780 10332 94836
rect 10388 94780 10398 94836
rect 10556 94780 23772 94836
rect 23828 94780 23838 94836
rect 10556 94724 10612 94780
rect 1810 94668 1820 94724
rect 1876 94668 4396 94724
rect 4452 94668 5740 94724
rect 5796 94668 5806 94724
rect 8642 94668 8652 94724
rect 8708 94668 8988 94724
rect 9044 94668 10612 94724
rect 12226 94668 12236 94724
rect 12292 94668 18172 94724
rect 18228 94668 18238 94724
rect 19618 94668 19628 94724
rect 19684 94668 20076 94724
rect 20132 94668 20142 94724
rect 23650 94668 23660 94724
rect 23716 94668 30268 94724
rect 30324 94668 30334 94724
rect 1250 94556 1260 94612
rect 1316 94556 4844 94612
rect 4900 94556 4910 94612
rect 6962 94556 6972 94612
rect 7028 94556 10892 94612
rect 10948 94556 10958 94612
rect 11862 94556 11900 94612
rect 11956 94556 11966 94612
rect 18844 94556 23324 94612
rect 23380 94556 23390 94612
rect 0 94500 112 94528
rect 18844 94500 18900 94556
rect 0 94444 1932 94500
rect 1988 94444 1998 94500
rect 2482 94444 2492 94500
rect 2548 94444 4060 94500
rect 4116 94444 4126 94500
rect 5394 94444 5404 94500
rect 5460 94444 6188 94500
rect 6244 94444 7084 94500
rect 7140 94444 7150 94500
rect 8194 94444 8204 94500
rect 8260 94444 14700 94500
rect 14756 94444 14766 94500
rect 17490 94444 17500 94500
rect 17556 94444 18172 94500
rect 18228 94444 18844 94500
rect 18900 94444 18910 94500
rect 19954 94444 19964 94500
rect 20020 94444 20188 94500
rect 20244 94444 22092 94500
rect 22148 94444 22158 94500
rect 0 94416 112 94444
rect 1474 94332 1484 94388
rect 1540 94332 2156 94388
rect 2212 94332 3388 94388
rect 3444 94332 3454 94388
rect 5506 94332 5516 94388
rect 5572 94332 8428 94388
rect 8484 94332 8494 94388
rect 13878 94332 13916 94388
rect 13972 94332 13982 94388
rect 15810 94332 15820 94388
rect 15876 94332 27804 94388
rect 27860 94332 27870 94388
rect 2034 94220 2044 94276
rect 2100 94220 6972 94276
rect 7028 94220 7038 94276
rect 10210 94220 10220 94276
rect 10276 94220 17164 94276
rect 17220 94220 17230 94276
rect 19282 94220 19292 94276
rect 19348 94220 20188 94276
rect 20244 94220 22204 94276
rect 22260 94220 22270 94276
rect 22418 94220 22428 94276
rect 22484 94220 22764 94276
rect 22820 94220 22830 94276
rect 23212 94220 26348 94276
rect 26404 94220 26414 94276
rect 23212 94164 23268 94220
rect 2146 94108 2156 94164
rect 2212 94108 2492 94164
rect 2548 94108 2558 94164
rect 4834 94108 4844 94164
rect 4900 94108 5572 94164
rect 6290 94108 6300 94164
rect 6356 94108 9996 94164
rect 10052 94108 11004 94164
rect 11060 94108 11070 94164
rect 13570 94108 13580 94164
rect 13636 94108 13916 94164
rect 13972 94108 13982 94164
rect 17154 94108 17164 94164
rect 17220 94108 23268 94164
rect 0 94052 112 94080
rect 3794 94052 3804 94108
rect 3860 94052 3908 94108
rect 3964 94052 4012 94108
rect 4068 94052 4078 94108
rect 5516 94052 5572 94108
rect 23794 94052 23804 94108
rect 23860 94052 23908 94108
rect 23964 94052 24012 94108
rect 24068 94052 24078 94108
rect 0 93996 3388 94052
rect 3490 93996 3500 94052
rect 3556 93996 3612 94052
rect 3668 93996 3678 94052
rect 5506 93996 5516 94052
rect 5572 93996 5582 94052
rect 7868 93996 8876 94052
rect 8932 93996 8942 94052
rect 10770 93996 10780 94052
rect 10836 93996 10892 94052
rect 10948 93996 10958 94052
rect 13458 93996 13468 94052
rect 13524 93996 14140 94052
rect 14196 93996 14206 94052
rect 17714 93996 17724 94052
rect 17780 93996 18396 94052
rect 18452 93996 18462 94052
rect 0 93968 112 93996
rect 3332 93940 3388 93996
rect 7868 93940 7924 93996
rect 31584 93940 31696 93968
rect 3332 93884 7924 93940
rect 8418 93884 8428 93940
rect 8484 93884 9324 93940
rect 9380 93884 10444 93940
rect 10500 93884 10510 93940
rect 17826 93884 17836 93940
rect 17892 93884 21084 93940
rect 21140 93884 21150 93940
rect 30594 93884 30604 93940
rect 30660 93884 31696 93940
rect 31584 93856 31696 93884
rect 3154 93772 3164 93828
rect 3220 93772 3276 93828
rect 3332 93772 3342 93828
rect 3490 93772 3500 93828
rect 3556 93772 4284 93828
rect 4340 93772 4350 93828
rect 9212 93772 16380 93828
rect 16436 93772 16446 93828
rect 2370 93660 2380 93716
rect 2436 93660 3948 93716
rect 4004 93660 4014 93716
rect 5730 93660 5740 93716
rect 5796 93660 6188 93716
rect 6244 93660 6254 93716
rect 0 93604 112 93632
rect 9212 93604 9268 93772
rect 10770 93660 10780 93716
rect 10836 93660 11228 93716
rect 11284 93660 11294 93716
rect 11554 93660 11564 93716
rect 11620 93660 11900 93716
rect 11956 93660 13132 93716
rect 13188 93660 13198 93716
rect 15138 93660 15148 93716
rect 15204 93660 17052 93716
rect 17108 93660 17118 93716
rect 17798 93660 17836 93716
rect 17892 93660 17902 93716
rect 0 93548 9268 93604
rect 9538 93548 9548 93604
rect 9604 93548 15484 93604
rect 15540 93548 15550 93604
rect 0 93520 112 93548
rect 466 93436 476 93492
rect 532 93436 5740 93492
rect 5796 93436 5806 93492
rect 8754 93436 8764 93492
rect 8820 93436 9324 93492
rect 9380 93436 13468 93492
rect 13524 93436 13534 93492
rect 17938 93436 17948 93492
rect 18004 93436 19180 93492
rect 19236 93436 19246 93492
rect 19506 93436 19516 93492
rect 19572 93436 30268 93492
rect 30324 93436 30334 93492
rect 5058 93324 5068 93380
rect 5124 93324 5964 93380
rect 6020 93324 10780 93380
rect 10836 93324 14028 93380
rect 14084 93324 14476 93380
rect 14532 93324 14542 93380
rect 15474 93324 15484 93380
rect 15540 93324 15932 93380
rect 15988 93324 15998 93380
rect 4454 93268 4464 93324
rect 4520 93268 4568 93324
rect 4624 93268 4672 93324
rect 4728 93268 4738 93324
rect 24454 93268 24464 93324
rect 24520 93268 24568 93324
rect 24624 93268 24672 93324
rect 24728 93268 24738 93324
rect 7046 93212 7084 93268
rect 7140 93212 7150 93268
rect 8306 93212 8316 93268
rect 8372 93212 10668 93268
rect 10724 93212 13580 93268
rect 13636 93212 13646 93268
rect 0 93156 112 93184
rect 0 93100 19740 93156
rect 19796 93100 19806 93156
rect 0 93072 112 93100
rect 1586 92988 1596 93044
rect 1652 92988 2044 93044
rect 2100 92988 2110 93044
rect 8530 92988 8540 93044
rect 8596 92988 8876 93044
rect 8932 92988 8942 93044
rect 10322 92988 10332 93044
rect 10388 92988 11676 93044
rect 11732 92988 11742 93044
rect 14802 92988 14812 93044
rect 14868 92988 15036 93044
rect 15092 92988 15102 93044
rect 15586 92988 15596 93044
rect 15652 92988 20580 93044
rect 20850 92988 20860 93044
rect 20916 92988 24668 93044
rect 24724 92988 24734 93044
rect 5058 92876 5068 92932
rect 5124 92876 5628 92932
rect 5684 92876 5694 92932
rect 6626 92876 6636 92932
rect 6692 92876 8316 92932
rect 8372 92876 8382 92932
rect 8754 92876 8764 92932
rect 8820 92876 9660 92932
rect 9716 92876 9726 92932
rect 10882 92876 10892 92932
rect 10948 92876 11004 92932
rect 11060 92876 11070 92932
rect 13570 92876 13580 92932
rect 13636 92876 14476 92932
rect 14532 92876 17052 92932
rect 17108 92876 17724 92932
rect 17780 92876 17790 92932
rect 20524 92820 20580 92988
rect 21634 92876 21644 92932
rect 21700 92876 22316 92932
rect 22372 92876 22382 92932
rect 31584 92820 31696 92848
rect 466 92764 476 92820
rect 532 92764 2100 92820
rect 5954 92764 5964 92820
rect 6020 92764 18508 92820
rect 18564 92764 18574 92820
rect 20524 92764 20860 92820
rect 20916 92764 20926 92820
rect 30594 92764 30604 92820
rect 30660 92764 31696 92820
rect 0 92708 112 92736
rect 2044 92708 2100 92764
rect 31584 92736 31696 92764
rect 0 92652 1036 92708
rect 1092 92652 1102 92708
rect 2044 92652 4956 92708
rect 5012 92652 5124 92708
rect 5282 92652 5292 92708
rect 5348 92652 11788 92708
rect 11844 92652 11854 92708
rect 14690 92652 14700 92708
rect 14756 92652 16268 92708
rect 16324 92652 16334 92708
rect 18722 92652 18732 92708
rect 18788 92652 19404 92708
rect 19460 92652 19470 92708
rect 21634 92652 21644 92708
rect 21700 92652 25452 92708
rect 25508 92652 25518 92708
rect 25778 92652 25788 92708
rect 25844 92652 28028 92708
rect 28084 92652 28094 92708
rect 0 92624 112 92652
rect 5068 92596 5124 92652
rect 5068 92540 6076 92596
rect 6132 92540 6300 92596
rect 6356 92540 6366 92596
rect 6738 92540 6748 92596
rect 6804 92540 7084 92596
rect 7140 92540 7150 92596
rect 15026 92540 15036 92596
rect 15092 92540 15596 92596
rect 15652 92540 15662 92596
rect 16044 92540 17500 92596
rect 17556 92540 17566 92596
rect 18498 92540 18508 92596
rect 18564 92540 19852 92596
rect 19908 92540 19918 92596
rect 3794 92484 3804 92540
rect 3860 92484 3908 92540
rect 3964 92484 4012 92540
rect 4068 92484 4078 92540
rect 4834 92428 4844 92484
rect 4900 92428 5404 92484
rect 5460 92428 5470 92484
rect 5730 92428 5740 92484
rect 5796 92428 5964 92484
rect 6020 92428 11900 92484
rect 11956 92428 11966 92484
rect 12898 92428 12908 92484
rect 12964 92428 13916 92484
rect 13972 92428 13982 92484
rect 16044 92372 16100 92540
rect 23794 92484 23804 92540
rect 23860 92484 23908 92540
rect 23964 92484 24012 92540
rect 24068 92484 24078 92540
rect 16594 92428 16604 92484
rect 16660 92428 19292 92484
rect 19348 92428 19358 92484
rect 3332 92316 8204 92372
rect 8260 92316 8270 92372
rect 9314 92316 9324 92372
rect 9380 92316 16100 92372
rect 16258 92316 16268 92372
rect 16324 92316 16492 92372
rect 16548 92316 16558 92372
rect 17798 92316 17836 92372
rect 17892 92316 17902 92372
rect 20066 92316 20076 92372
rect 20132 92316 21532 92372
rect 21588 92316 21598 92372
rect 0 92260 112 92288
rect 3332 92260 3388 92316
rect 0 92204 3388 92260
rect 5394 92204 5404 92260
rect 5460 92204 7980 92260
rect 8036 92204 8046 92260
rect 9426 92204 9436 92260
rect 9492 92204 9660 92260
rect 9716 92204 9726 92260
rect 15586 92204 15596 92260
rect 15652 92204 15662 92260
rect 15820 92204 21868 92260
rect 21924 92204 21934 92260
rect 0 92176 112 92204
rect 15596 92148 15652 92204
rect 15820 92148 15876 92204
rect 2258 92092 2268 92148
rect 2324 92092 5068 92148
rect 5124 92092 5134 92148
rect 9212 92092 15652 92148
rect 15708 92092 15876 92148
rect 16034 92092 16044 92148
rect 16100 92092 17052 92148
rect 17108 92092 17118 92148
rect 17266 92092 17276 92148
rect 17332 92092 17948 92148
rect 18004 92092 18014 92148
rect 21074 92092 21084 92148
rect 21140 92092 21308 92148
rect 21364 92092 21374 92148
rect 21746 92092 21756 92148
rect 21812 92092 22652 92148
rect 22708 92092 22718 92148
rect 1474 91980 1484 92036
rect 1540 91980 5740 92036
rect 5796 91980 6636 92036
rect 6692 91980 6702 92036
rect 3332 91868 4900 91924
rect 6486 91868 6524 91924
rect 6580 91868 6590 91924
rect 7746 91868 7756 91924
rect 7812 91868 8316 91924
rect 8372 91868 8382 91924
rect 8530 91868 8540 91924
rect 8596 91868 8764 91924
rect 8820 91868 8830 91924
rect 0 91812 112 91840
rect 3332 91812 3388 91868
rect 0 91756 3388 91812
rect 4844 91812 4900 91868
rect 9212 91812 9268 92092
rect 15708 92036 15764 92092
rect 4844 91756 9268 91812
rect 12908 91980 15764 92036
rect 15922 91980 15932 92036
rect 15988 91980 17164 92036
rect 17220 91980 17230 92036
rect 0 91728 112 91756
rect 4454 91700 4464 91756
rect 4520 91700 4568 91756
rect 4624 91700 4672 91756
rect 4728 91700 4738 91756
rect 7074 91532 7084 91588
rect 7140 91532 7420 91588
rect 7476 91532 7486 91588
rect 8194 91532 8204 91588
rect 8260 91532 12684 91588
rect 12740 91532 12750 91588
rect 12908 91476 12964 91980
rect 15932 91924 15988 91980
rect 15138 91868 15148 91924
rect 15204 91868 15988 91924
rect 19506 91868 19516 91924
rect 19572 91868 30268 91924
rect 30324 91868 30334 91924
rect 24454 91700 24464 91756
rect 24520 91700 24568 91756
rect 24624 91700 24672 91756
rect 24728 91700 24738 91756
rect 31584 91700 31696 91728
rect 19282 91644 19292 91700
rect 19348 91644 19516 91700
rect 19572 91644 19582 91700
rect 21942 91644 21980 91700
rect 22036 91644 22046 91700
rect 30594 91644 30604 91700
rect 30660 91644 31696 91700
rect 31584 91616 31696 91644
rect 14802 91532 14812 91588
rect 14868 91532 18620 91588
rect 18676 91532 18686 91588
rect 2370 91420 2380 91476
rect 2436 91420 2828 91476
rect 2884 91420 2894 91476
rect 4610 91420 4620 91476
rect 4676 91420 4956 91476
rect 5012 91420 5022 91476
rect 6178 91420 6188 91476
rect 6244 91420 6524 91476
rect 6580 91420 6590 91476
rect 7074 91420 7084 91476
rect 7140 91420 7980 91476
rect 8036 91420 10892 91476
rect 10948 91420 10958 91476
rect 11116 91420 12964 91476
rect 17714 91420 17724 91476
rect 17780 91420 20188 91476
rect 20244 91420 20254 91476
rect 0 91364 112 91392
rect 11116 91364 11172 91420
rect 0 91308 11172 91364
rect 12114 91308 12124 91364
rect 12180 91308 13244 91364
rect 13300 91308 14364 91364
rect 14420 91308 14430 91364
rect 15250 91308 15260 91364
rect 15316 91308 16156 91364
rect 16212 91308 18172 91364
rect 18228 91308 18238 91364
rect 18834 91308 18844 91364
rect 18900 91308 19740 91364
rect 19796 91308 19806 91364
rect 0 91280 112 91308
rect 802 91196 812 91252
rect 868 91196 1260 91252
rect 1316 91196 1484 91252
rect 1540 91196 4956 91252
rect 5012 91196 5022 91252
rect 14018 91196 14028 91252
rect 14084 91196 14476 91252
rect 14532 91196 14542 91252
rect 15922 91196 15932 91252
rect 15988 91196 17948 91252
rect 18004 91196 18014 91252
rect 2716 91140 2772 91196
rect 2706 91084 2716 91140
rect 2772 91084 2782 91140
rect 3042 91084 3052 91140
rect 3108 91084 3118 91140
rect 6486 91084 6524 91140
rect 6580 91084 6590 91140
rect 13794 91084 13804 91140
rect 13860 91084 16828 91140
rect 16884 91084 17724 91140
rect 17780 91084 18732 91140
rect 18788 91084 18798 91140
rect 22082 91084 22092 91140
rect 22148 91084 22764 91140
rect 22820 91084 22830 91140
rect 0 90916 112 90944
rect 3052 90916 3108 91084
rect 3266 90972 3276 91028
rect 3332 90972 3342 91028
rect 15698 90972 15708 91028
rect 15764 90972 16716 91028
rect 16772 90972 16782 91028
rect 0 90860 3108 90916
rect 0 90832 112 90860
rect 578 90636 588 90692
rect 644 90636 1484 90692
rect 1540 90636 1550 90692
rect 3276 90580 3332 90972
rect 3794 90916 3804 90972
rect 3860 90916 3908 90972
rect 3964 90916 4012 90972
rect 4068 90916 4078 90972
rect 23794 90916 23804 90972
rect 23860 90916 23908 90972
rect 23964 90916 24012 90972
rect 24068 90916 24078 90972
rect 5730 90860 5740 90916
rect 5796 90860 11900 90916
rect 11956 90860 19180 90916
rect 19236 90860 19246 90916
rect 19852 90860 21532 90916
rect 21588 90860 21598 90916
rect 21858 90860 21868 90916
rect 21924 90860 22204 90916
rect 22260 90860 22270 90916
rect 19852 90804 19908 90860
rect 5954 90748 5964 90804
rect 6020 90748 7084 90804
rect 7140 90748 7150 90804
rect 12450 90748 12460 90804
rect 12516 90748 19908 90804
rect 20066 90748 20076 90804
rect 20132 90748 20412 90804
rect 20468 90748 20478 90804
rect 20850 90748 20860 90804
rect 20916 90748 21756 90804
rect 21812 90748 21822 90804
rect 7410 90636 7420 90692
rect 7476 90636 13020 90692
rect 13076 90636 13086 90692
rect 15474 90636 15484 90692
rect 15540 90636 15820 90692
rect 15876 90636 15886 90692
rect 18722 90636 18732 90692
rect 18788 90636 20972 90692
rect 21028 90636 21038 90692
rect 21186 90636 21196 90692
rect 21252 90636 21532 90692
rect 21588 90636 21598 90692
rect 31584 90580 31696 90608
rect 3154 90524 3164 90580
rect 3220 90524 3332 90580
rect 3602 90524 3612 90580
rect 3668 90524 12124 90580
rect 12180 90524 18844 90580
rect 18900 90524 18910 90580
rect 20626 90524 20636 90580
rect 20692 90524 22204 90580
rect 22260 90524 22270 90580
rect 30594 90524 30604 90580
rect 30660 90524 31696 90580
rect 31584 90496 31696 90524
rect 0 90468 112 90496
rect 0 90412 10220 90468
rect 10276 90412 10286 90468
rect 11732 90412 12796 90468
rect 12852 90412 12862 90468
rect 13122 90412 13132 90468
rect 13188 90412 30268 90468
rect 30324 90412 30334 90468
rect 0 90384 112 90412
rect 11732 90356 11788 90412
rect 578 90300 588 90356
rect 644 90300 1148 90356
rect 1204 90300 1214 90356
rect 2370 90300 2380 90356
rect 2436 90300 4060 90356
rect 4116 90300 4126 90356
rect 4284 90300 6860 90356
rect 6916 90300 6926 90356
rect 11106 90300 11116 90356
rect 11172 90300 11228 90356
rect 11284 90300 11788 90356
rect 13458 90300 13468 90356
rect 13524 90300 13916 90356
rect 13972 90300 13982 90356
rect 14578 90300 14588 90356
rect 14644 90300 15148 90356
rect 15204 90300 15214 90356
rect 16706 90300 16716 90356
rect 16772 90300 18172 90356
rect 18228 90300 18238 90356
rect 22642 90300 22652 90356
rect 22708 90300 27916 90356
rect 27972 90300 27982 90356
rect 4284 90132 4340 90300
rect 5394 90188 5404 90244
rect 5460 90188 6188 90244
rect 6244 90188 9660 90244
rect 9716 90188 9726 90244
rect 11638 90188 11676 90244
rect 11732 90188 13580 90244
rect 13636 90188 13646 90244
rect 16034 90188 16044 90244
rect 16100 90188 16492 90244
rect 16548 90188 17500 90244
rect 17556 90188 17724 90244
rect 17780 90188 17790 90244
rect 4454 90132 4464 90188
rect 4520 90132 4568 90188
rect 4624 90132 4672 90188
rect 4728 90132 4738 90188
rect 24454 90132 24464 90188
rect 24520 90132 24568 90188
rect 24624 90132 24672 90188
rect 24728 90132 24738 90188
rect 1138 90076 1148 90132
rect 1204 90076 1708 90132
rect 1764 90076 1774 90132
rect 2706 90076 2716 90132
rect 2772 90076 4340 90132
rect 9874 90076 9884 90132
rect 9940 90076 12236 90132
rect 12292 90076 12302 90132
rect 13346 90076 13356 90132
rect 13412 90076 14364 90132
rect 14420 90076 14430 90132
rect 0 90020 112 90048
rect 0 89964 17836 90020
rect 17892 89964 17902 90020
rect 0 89936 112 89964
rect 242 89852 252 89908
rect 308 89852 7028 89908
rect 7186 89852 7196 89908
rect 7252 89852 7644 89908
rect 7700 89852 7710 89908
rect 7858 89852 7868 89908
rect 7924 89852 9324 89908
rect 9380 89852 10108 89908
rect 10164 89852 10174 89908
rect 12562 89852 12572 89908
rect 12628 89852 30268 89908
rect 30324 89852 30334 89908
rect 0 89572 112 89600
rect 2940 89572 2996 89852
rect 6972 89796 7028 89852
rect 3378 89740 3388 89796
rect 3444 89740 3724 89796
rect 3780 89740 3790 89796
rect 6972 89740 8372 89796
rect 13682 89740 13692 89796
rect 13748 89740 14140 89796
rect 14196 89740 14206 89796
rect 15026 89740 15036 89796
rect 15092 89740 16940 89796
rect 16996 89740 17006 89796
rect 8316 89684 8372 89740
rect 3154 89628 3164 89684
rect 3220 89628 7532 89684
rect 7588 89628 7598 89684
rect 8316 89628 15148 89684
rect 0 89516 1764 89572
rect 2566 89516 2604 89572
rect 2660 89516 2670 89572
rect 2940 89516 3052 89572
rect 3108 89516 3118 89572
rect 7830 89516 7868 89572
rect 7924 89516 7934 89572
rect 11218 89516 11228 89572
rect 11284 89516 11788 89572
rect 11844 89516 11854 89572
rect 0 89488 112 89516
rect 1708 89460 1764 89516
rect 15092 89460 15148 89628
rect 31584 89460 31696 89488
rect 1708 89404 3388 89460
rect 15092 89404 20636 89460
rect 20692 89404 20702 89460
rect 30594 89404 30604 89460
rect 30660 89404 31696 89460
rect 3332 89236 3388 89404
rect 3794 89348 3804 89404
rect 3860 89348 3908 89404
rect 3964 89348 4012 89404
rect 4068 89348 4078 89404
rect 23794 89348 23804 89404
rect 23860 89348 23908 89404
rect 23964 89348 24012 89404
rect 24068 89348 24078 89404
rect 31584 89376 31696 89404
rect 5842 89292 5852 89348
rect 5908 89292 6188 89348
rect 6244 89292 6254 89348
rect 8082 89292 8092 89348
rect 8148 89292 8204 89348
rect 8260 89292 8270 89348
rect 17266 89292 17276 89348
rect 17332 89292 18060 89348
rect 18116 89292 18126 89348
rect 2258 89180 2268 89236
rect 2324 89180 2716 89236
rect 2772 89180 2782 89236
rect 3332 89180 20636 89236
rect 20692 89180 22876 89236
rect 22932 89180 22942 89236
rect 0 89124 112 89152
rect 0 89068 4172 89124
rect 4228 89068 4238 89124
rect 4396 89068 5068 89124
rect 5124 89068 5134 89124
rect 9650 89068 9660 89124
rect 9716 89068 10556 89124
rect 10612 89068 13020 89124
rect 13076 89068 13086 89124
rect 26226 89068 26236 89124
rect 26292 89068 27132 89124
rect 27188 89068 27198 89124
rect 0 89040 112 89068
rect 4396 89012 4452 89068
rect 1026 88956 1036 89012
rect 1092 88956 1708 89012
rect 1764 88956 2604 89012
rect 2660 88956 2670 89012
rect 3154 88956 3164 89012
rect 3220 88956 4452 89012
rect 5058 88956 5068 89012
rect 5124 88956 6636 89012
rect 6692 88956 6702 89012
rect 6962 88956 6972 89012
rect 7028 88956 8764 89012
rect 8820 88956 8830 89012
rect 8978 88956 8988 89012
rect 9044 88956 9324 89012
rect 9380 88956 9390 89012
rect 11004 88956 11116 89012
rect 11172 88956 11182 89012
rect 14466 88956 14476 89012
rect 14532 88956 18732 89012
rect 18788 88956 21980 89012
rect 22036 88956 24332 89012
rect 24388 88956 24398 89012
rect 4834 88844 4844 88900
rect 4900 88844 6860 88900
rect 6916 88844 6926 88900
rect 3332 88732 5684 88788
rect 5842 88732 5852 88788
rect 5908 88732 8988 88788
rect 9044 88732 9054 88788
rect 0 88676 112 88704
rect 3332 88676 3388 88732
rect 0 88620 3388 88676
rect 5628 88676 5684 88732
rect 11004 88676 11060 88956
rect 16594 88844 16604 88900
rect 16660 88844 17388 88900
rect 17444 88844 17454 88900
rect 17490 88732 17500 88788
rect 17556 88732 18284 88788
rect 18340 88732 18350 88788
rect 18498 88732 18508 88788
rect 18564 88732 24892 88788
rect 24948 88732 24958 88788
rect 5628 88620 11060 88676
rect 13346 88620 13356 88676
rect 13412 88620 13422 88676
rect 0 88592 112 88620
rect 4454 88564 4464 88620
rect 4520 88564 4568 88620
rect 4624 88564 4672 88620
rect 4728 88564 4738 88620
rect 13356 88564 13412 88620
rect 24454 88564 24464 88620
rect 24520 88564 24568 88620
rect 24624 88564 24672 88620
rect 24728 88564 24738 88620
rect 5730 88508 5740 88564
rect 5796 88508 6636 88564
rect 6692 88508 13412 88564
rect 3332 88396 14812 88452
rect 14868 88396 14878 88452
rect 0 88228 112 88256
rect 3332 88228 3388 88396
rect 31584 88340 31696 88368
rect 9846 88284 9884 88340
rect 9940 88284 9950 88340
rect 11218 88284 11228 88340
rect 11284 88284 11452 88340
rect 11508 88284 11518 88340
rect 13682 88284 13692 88340
rect 13748 88284 14028 88340
rect 14084 88284 18396 88340
rect 18452 88284 18462 88340
rect 30594 88284 30604 88340
rect 30660 88284 31696 88340
rect 31584 88256 31696 88284
rect 0 88172 3388 88228
rect 3490 88172 3500 88228
rect 3556 88172 3612 88228
rect 3668 88172 3678 88228
rect 12674 88172 12684 88228
rect 12740 88172 13244 88228
rect 13300 88172 13310 88228
rect 14914 88172 14924 88228
rect 14980 88172 21196 88228
rect 21252 88172 21420 88228
rect 21476 88172 21486 88228
rect 0 88144 112 88172
rect 3238 88060 3276 88116
rect 3332 88060 3342 88116
rect 3714 88060 3724 88116
rect 3780 88060 4060 88116
rect 4116 88060 13804 88116
rect 13860 88060 13870 88116
rect 3332 87948 5292 88004
rect 5348 87948 5358 88004
rect 19282 87948 19292 88004
rect 19348 87948 19628 88004
rect 19684 87948 19694 88004
rect 0 87780 112 87808
rect 3332 87780 3388 87948
rect 3794 87780 3804 87836
rect 3860 87780 3908 87836
rect 3964 87780 4012 87836
rect 4068 87780 4078 87836
rect 23794 87780 23804 87836
rect 23860 87780 23908 87836
rect 23964 87780 24012 87836
rect 24068 87780 24078 87836
rect 0 87724 3388 87780
rect 10546 87724 10556 87780
rect 10612 87724 12796 87780
rect 12852 87724 12862 87780
rect 0 87696 112 87724
rect 3378 87612 3388 87668
rect 3444 87612 3482 87668
rect 13122 87612 13132 87668
rect 13188 87612 15036 87668
rect 15092 87612 18060 87668
rect 18116 87612 22316 87668
rect 22372 87612 22382 87668
rect 1698 87500 1708 87556
rect 1764 87500 1820 87556
rect 1876 87500 2716 87556
rect 2772 87500 2782 87556
rect 6290 87500 6300 87556
rect 6356 87500 7084 87556
rect 7140 87500 7150 87556
rect 11442 87500 11452 87556
rect 11508 87500 15372 87556
rect 15428 87500 16716 87556
rect 16772 87500 16782 87556
rect 20514 87500 20524 87556
rect 20580 87500 22652 87556
rect 22708 87500 22718 87556
rect 23874 87500 23884 87556
rect 23940 87500 25900 87556
rect 25956 87500 25966 87556
rect 1362 87388 1372 87444
rect 1428 87388 4284 87444
rect 4340 87388 4350 87444
rect 8418 87388 8428 87444
rect 8484 87388 11228 87444
rect 11284 87388 11294 87444
rect 11554 87388 11564 87444
rect 11620 87388 11788 87444
rect 11844 87388 11854 87444
rect 14690 87388 14700 87444
rect 14756 87388 15484 87444
rect 15540 87388 16492 87444
rect 16548 87388 16558 87444
rect 17490 87388 17500 87444
rect 17556 87388 22876 87444
rect 22932 87388 22942 87444
rect 23202 87388 23212 87444
rect 23268 87388 30268 87444
rect 30324 87388 30334 87444
rect 0 87332 112 87360
rect 0 87276 140 87332
rect 196 87276 206 87332
rect 2146 87276 2156 87332
rect 2212 87276 6188 87332
rect 6244 87276 6254 87332
rect 9426 87276 9436 87332
rect 9492 87276 11004 87332
rect 11060 87276 14364 87332
rect 14420 87276 14924 87332
rect 14980 87276 14990 87332
rect 21298 87276 21308 87332
rect 21364 87276 21756 87332
rect 21812 87276 21822 87332
rect 0 87248 112 87276
rect 31584 87220 31696 87248
rect 1138 87164 1148 87220
rect 1204 87164 2604 87220
rect 2660 87164 2670 87220
rect 18806 87164 18844 87220
rect 18900 87164 18910 87220
rect 20514 87164 20524 87220
rect 20580 87164 20748 87220
rect 20804 87164 20814 87220
rect 30594 87164 30604 87220
rect 30660 87164 31696 87220
rect 31584 87136 31696 87164
rect 1698 87052 1708 87108
rect 1764 87052 4340 87108
rect 14354 87052 14364 87108
rect 14420 87052 19628 87108
rect 19684 87052 19852 87108
rect 19908 87052 20188 87108
rect 20244 87052 20254 87108
rect 0 86884 112 86912
rect 4284 86884 4340 87052
rect 4454 86996 4464 87052
rect 4520 86996 4568 87052
rect 4624 86996 4672 87052
rect 4728 86996 4738 87052
rect 24454 86996 24464 87052
rect 24520 86996 24568 87052
rect 24624 86996 24672 87052
rect 24728 86996 24738 87052
rect 6290 86940 6300 86996
rect 6356 86940 6412 86996
rect 6468 86940 6478 86996
rect 7084 86940 23548 86996
rect 23604 86940 23614 86996
rect 0 86828 2044 86884
rect 2100 86828 2110 86884
rect 2594 86828 2604 86884
rect 2660 86828 3948 86884
rect 4004 86828 4014 86884
rect 4284 86828 6748 86884
rect 6804 86828 6814 86884
rect 0 86800 112 86828
rect 7084 86772 7140 86940
rect 7298 86828 7308 86884
rect 7364 86828 11340 86884
rect 11396 86828 11406 86884
rect 17378 86828 17388 86884
rect 17444 86828 21868 86884
rect 21924 86828 21934 86884
rect 690 86716 700 86772
rect 756 86716 1484 86772
rect 1540 86716 1596 86772
rect 1652 86716 1662 86772
rect 2706 86716 2716 86772
rect 2772 86716 7084 86772
rect 7140 86716 7150 86772
rect 9986 86716 9996 86772
rect 10052 86716 11004 86772
rect 11060 86716 12460 86772
rect 12516 86716 12526 86772
rect 18722 86716 18732 86772
rect 18788 86716 19852 86772
rect 19908 86716 19918 86772
rect 23090 86716 23100 86772
rect 23156 86716 23436 86772
rect 23492 86716 23502 86772
rect 3714 86604 3724 86660
rect 3780 86604 5404 86660
rect 5460 86604 5470 86660
rect 10994 86604 11004 86660
rect 11060 86604 11788 86660
rect 11844 86604 11854 86660
rect 13430 86604 13468 86660
rect 13524 86604 13534 86660
rect 18946 86604 18956 86660
rect 19012 86604 22652 86660
rect 22708 86604 22718 86660
rect 1362 86492 1372 86548
rect 1428 86492 1596 86548
rect 1652 86492 1662 86548
rect 3938 86492 3948 86548
rect 4004 86492 13916 86548
rect 13972 86492 14700 86548
rect 14756 86492 14766 86548
rect 0 86436 112 86464
rect 0 86380 10220 86436
rect 10276 86380 20860 86436
rect 20916 86380 23996 86436
rect 24052 86380 24062 86436
rect 0 86352 112 86380
rect 1250 86268 1260 86324
rect 1316 86268 1932 86324
rect 1988 86268 1998 86324
rect 11330 86268 11340 86324
rect 11396 86268 13468 86324
rect 13524 86268 13534 86324
rect 3794 86212 3804 86268
rect 3860 86212 3908 86268
rect 3964 86212 4012 86268
rect 4068 86212 4078 86268
rect 23794 86212 23804 86268
rect 23860 86212 23908 86268
rect 23964 86212 24012 86268
rect 24068 86212 24078 86268
rect 2370 86156 2380 86212
rect 2436 86156 2716 86212
rect 2772 86156 2782 86212
rect 6738 86156 6748 86212
rect 6804 86156 13580 86212
rect 13636 86156 13646 86212
rect 14242 86156 14252 86212
rect 14308 86156 20860 86212
rect 20916 86156 20926 86212
rect 21858 86156 21868 86212
rect 21924 86156 22540 86212
rect 22596 86156 22606 86212
rect 21868 86100 21924 86156
rect 31584 86100 31696 86128
rect 1586 86044 1596 86100
rect 1652 86044 3948 86100
rect 4004 86044 4014 86100
rect 5068 86044 9716 86100
rect 10994 86044 11004 86100
rect 11060 86044 21924 86100
rect 22866 86044 22876 86100
rect 22932 86044 23324 86100
rect 23380 86044 23390 86100
rect 23510 86044 23548 86100
rect 23604 86044 23614 86100
rect 30594 86044 30604 86100
rect 30660 86044 31696 86100
rect 0 85988 112 86016
rect 5068 85988 5124 86044
rect 9660 85988 9716 86044
rect 31584 86016 31696 86044
rect 0 85932 5124 85988
rect 5282 85932 5292 85988
rect 5348 85932 9436 85988
rect 9492 85932 9502 85988
rect 9660 85932 11116 85988
rect 11172 85932 11182 85988
rect 13570 85932 13580 85988
rect 13636 85932 13804 85988
rect 13860 85932 13870 85988
rect 14242 85932 14252 85988
rect 14308 85932 14700 85988
rect 14756 85932 14766 85988
rect 15138 85932 15148 85988
rect 15204 85932 15708 85988
rect 15764 85932 15774 85988
rect 16034 85932 16044 85988
rect 16100 85932 16828 85988
rect 16884 85932 17836 85988
rect 17892 85932 17902 85988
rect 19170 85932 19180 85988
rect 19236 85932 19404 85988
rect 19460 85932 19470 85988
rect 22978 85932 22988 85988
rect 23044 85932 23436 85988
rect 23492 85932 23502 85988
rect 0 85904 112 85932
rect 1810 85820 1820 85876
rect 1876 85820 5628 85876
rect 5684 85820 5694 85876
rect 6178 85820 6188 85876
rect 6244 85820 12012 85876
rect 12068 85820 13468 85876
rect 13524 85820 13534 85876
rect 14130 85820 14140 85876
rect 14196 85820 14812 85876
rect 14868 85820 14878 85876
rect 16370 85820 16380 85876
rect 16436 85820 17164 85876
rect 17220 85820 17230 85876
rect 21522 85820 21532 85876
rect 21588 85820 22540 85876
rect 22596 85820 22606 85876
rect 22754 85820 22764 85876
rect 22820 85820 23548 85876
rect 23604 85820 23614 85876
rect 130 85708 140 85764
rect 196 85708 1036 85764
rect 1092 85708 1102 85764
rect 1474 85708 1484 85764
rect 1540 85708 3388 85764
rect 3444 85708 3454 85764
rect 8866 85708 8876 85764
rect 8932 85708 14140 85764
rect 14196 85708 14364 85764
rect 14420 85708 14430 85764
rect 14578 85708 14588 85764
rect 14644 85708 15372 85764
rect 15428 85708 16604 85764
rect 16660 85708 16670 85764
rect 19394 85708 19404 85764
rect 19460 85708 20748 85764
rect 20804 85708 20814 85764
rect 21298 85708 21308 85764
rect 21364 85708 24108 85764
rect 24164 85708 24174 85764
rect 24434 85708 24444 85764
rect 24500 85708 30268 85764
rect 30324 85708 30334 85764
rect 690 85596 700 85652
rect 756 85596 1484 85652
rect 1540 85596 1550 85652
rect 2594 85596 2604 85652
rect 2660 85596 3164 85652
rect 3220 85596 3230 85652
rect 4274 85596 4284 85652
rect 4340 85596 6524 85652
rect 6580 85596 6590 85652
rect 13794 85596 13804 85652
rect 13860 85596 17052 85652
rect 17108 85596 17118 85652
rect 21942 85596 21980 85652
rect 22036 85596 22046 85652
rect 23874 85596 23884 85652
rect 23940 85596 28140 85652
rect 28196 85596 28206 85652
rect 0 85540 112 85568
rect 0 85484 3388 85540
rect 14018 85484 14028 85540
rect 14084 85484 14140 85540
rect 14196 85484 14206 85540
rect 14364 85484 16044 85540
rect 16100 85484 16110 85540
rect 16594 85484 16604 85540
rect 16660 85484 23548 85540
rect 23604 85484 23614 85540
rect 0 85456 112 85484
rect 1446 85372 1484 85428
rect 1540 85372 1550 85428
rect 2034 85372 2044 85428
rect 2100 85372 2380 85428
rect 2436 85372 2446 85428
rect 3332 85316 3388 85484
rect 4454 85428 4464 85484
rect 4520 85428 4568 85484
rect 4624 85428 4672 85484
rect 4728 85428 4738 85484
rect 14364 85428 14420 85484
rect 24454 85428 24464 85484
rect 24520 85428 24568 85484
rect 24624 85428 24672 85484
rect 24728 85428 24738 85484
rect 12786 85372 12796 85428
rect 12852 85372 14420 85428
rect 17154 85372 17164 85428
rect 17220 85372 17276 85428
rect 17332 85372 17342 85428
rect 2258 85260 2268 85316
rect 2324 85260 2334 85316
rect 3332 85260 8092 85316
rect 8148 85260 8158 85316
rect 10882 85260 10892 85316
rect 10948 85260 13244 85316
rect 13300 85260 13356 85316
rect 13412 85260 13422 85316
rect 16604 85260 17388 85316
rect 17444 85260 17454 85316
rect 19618 85260 19628 85316
rect 19684 85260 20412 85316
rect 20468 85260 20478 85316
rect 23062 85260 23100 85316
rect 23156 85260 23166 85316
rect 23538 85260 23548 85316
rect 23604 85260 24332 85316
rect 24388 85260 24398 85316
rect 0 85092 112 85120
rect 2268 85092 2324 85260
rect 16604 85204 16660 85260
rect 2818 85148 2828 85204
rect 2884 85148 2940 85204
rect 2996 85148 3006 85204
rect 6402 85148 6412 85204
rect 6468 85148 11228 85204
rect 11284 85148 16660 85204
rect 23874 85148 23884 85204
rect 23940 85148 30268 85204
rect 30324 85148 30334 85204
rect 0 85036 980 85092
rect 2034 85036 2044 85092
rect 2100 85036 2604 85092
rect 2660 85036 2670 85092
rect 3490 85036 3500 85092
rect 3556 85036 8988 85092
rect 9044 85036 9054 85092
rect 12450 85036 12460 85092
rect 12516 85036 13244 85092
rect 13300 85036 13310 85092
rect 14914 85036 14924 85092
rect 14980 85036 15148 85092
rect 15204 85036 15214 85092
rect 16034 85036 16044 85092
rect 16100 85036 16828 85092
rect 16884 85036 16894 85092
rect 19730 85036 19740 85092
rect 19796 85036 19964 85092
rect 20020 85036 20972 85092
rect 21028 85036 21038 85092
rect 22530 85036 22540 85092
rect 22596 85036 23436 85092
rect 23492 85036 23502 85092
rect 0 85008 112 85036
rect 924 84868 980 85036
rect 31584 84980 31696 85008
rect 1138 84924 1148 84980
rect 1204 84924 1820 84980
rect 1876 84924 1886 84980
rect 2258 84924 2268 84980
rect 2324 84924 2492 84980
rect 2548 84924 2558 84980
rect 2716 84924 8204 84980
rect 8260 84924 8270 84980
rect 11218 84924 11228 84980
rect 11284 84924 11452 84980
rect 11508 84924 11518 84980
rect 13346 84924 13356 84980
rect 13412 84924 15148 84980
rect 15204 84924 15214 84980
rect 16146 84924 16156 84980
rect 16212 84924 18004 84980
rect 21186 84924 21196 84980
rect 21252 84924 21420 84980
rect 21476 84924 21486 84980
rect 30594 84924 30604 84980
rect 30660 84924 31696 84980
rect 2716 84868 2772 84924
rect 924 84812 2772 84868
rect 3826 84812 3836 84868
rect 3892 84812 8204 84868
rect 8260 84812 8270 84868
rect 9884 84812 12460 84868
rect 12516 84812 12526 84868
rect 14354 84812 14364 84868
rect 14420 84812 16828 84868
rect 16884 84812 16894 84868
rect 9884 84756 9940 84812
rect 1362 84700 1372 84756
rect 1428 84700 3444 84756
rect 6178 84700 6188 84756
rect 6244 84700 9940 84756
rect 10098 84700 10108 84756
rect 10164 84700 15596 84756
rect 15652 84700 15662 84756
rect 0 84644 112 84672
rect 0 84588 1540 84644
rect 0 84560 112 84588
rect 1484 84420 1540 84588
rect 3388 84532 3444 84700
rect 3794 84644 3804 84700
rect 3860 84644 3908 84700
rect 3964 84644 4012 84700
rect 4068 84644 4078 84700
rect 17948 84644 18004 84924
rect 31584 84896 31696 84924
rect 18610 84812 18620 84868
rect 18676 84812 19852 84868
rect 19908 84812 19918 84868
rect 19394 84700 19404 84756
rect 19460 84700 20076 84756
rect 20132 84700 20142 84756
rect 21410 84700 21420 84756
rect 21476 84700 21644 84756
rect 21700 84700 21710 84756
rect 23794 84644 23804 84700
rect 23860 84644 23908 84700
rect 23964 84644 24012 84700
rect 24068 84644 24078 84700
rect 4946 84588 4956 84644
rect 5012 84588 7420 84644
rect 7476 84588 7486 84644
rect 9090 84588 9100 84644
rect 9156 84588 9884 84644
rect 9940 84588 9950 84644
rect 10882 84588 10892 84644
rect 10948 84588 11228 84644
rect 11284 84588 11294 84644
rect 17948 84588 19628 84644
rect 19684 84588 19694 84644
rect 3126 84476 3164 84532
rect 3220 84476 3230 84532
rect 3388 84476 11900 84532
rect 11956 84476 11966 84532
rect 16930 84476 16940 84532
rect 16996 84476 17276 84532
rect 17332 84476 17342 84532
rect 19058 84476 19068 84532
rect 19124 84476 21644 84532
rect 21700 84476 21710 84532
rect 1484 84364 10108 84420
rect 10164 84364 10174 84420
rect 10546 84364 10556 84420
rect 10612 84364 11004 84420
rect 11060 84364 11340 84420
rect 11396 84364 11406 84420
rect 13122 84364 13132 84420
rect 13188 84364 13468 84420
rect 13524 84364 15036 84420
rect 15092 84364 15102 84420
rect 19282 84364 19292 84420
rect 19348 84364 19740 84420
rect 19796 84364 19806 84420
rect 2818 84252 2828 84308
rect 2884 84252 3276 84308
rect 3332 84252 3342 84308
rect 4162 84252 4172 84308
rect 4228 84252 4844 84308
rect 4900 84252 4910 84308
rect 5842 84252 5852 84308
rect 5908 84252 6188 84308
rect 6244 84252 6254 84308
rect 7522 84252 7532 84308
rect 7588 84252 8876 84308
rect 8932 84252 8942 84308
rect 9650 84252 9660 84308
rect 9716 84252 12348 84308
rect 12404 84252 12414 84308
rect 13906 84252 13916 84308
rect 13972 84252 15932 84308
rect 15988 84252 16604 84308
rect 16660 84252 16670 84308
rect 17714 84252 17724 84308
rect 17780 84252 18060 84308
rect 18116 84252 18126 84308
rect 21074 84252 21084 84308
rect 21140 84252 22092 84308
rect 22148 84252 22158 84308
rect 0 84196 112 84224
rect 0 84140 6300 84196
rect 6356 84140 6366 84196
rect 6850 84140 6860 84196
rect 6916 84140 9884 84196
rect 9940 84140 9950 84196
rect 13010 84140 13020 84196
rect 13076 84140 13692 84196
rect 13748 84140 14924 84196
rect 14980 84140 14990 84196
rect 16034 84140 16044 84196
rect 16100 84140 19068 84196
rect 19124 84140 19134 84196
rect 0 84112 112 84140
rect 1138 84028 1148 84084
rect 1204 84028 1484 84084
rect 1540 84028 1550 84084
rect 2034 84028 2044 84084
rect 2100 84028 2156 84084
rect 2212 84028 2222 84084
rect 3042 84028 3052 84084
rect 3108 84028 3164 84084
rect 3220 84028 3230 84084
rect 4386 84028 4396 84084
rect 4452 84028 4900 84084
rect 5618 84028 5628 84084
rect 5684 84028 5964 84084
rect 6020 84028 6030 84084
rect 8082 84028 8092 84084
rect 8148 84028 8484 84084
rect 9650 84028 9660 84084
rect 9716 84028 13916 84084
rect 13972 84028 13982 84084
rect 16146 84028 16156 84084
rect 16212 84028 16716 84084
rect 16772 84028 16782 84084
rect 17826 84028 17836 84084
rect 17892 84028 19292 84084
rect 19348 84028 19358 84084
rect 23650 84028 23660 84084
rect 23716 84028 30268 84084
rect 30324 84028 30334 84084
rect 4844 83972 4900 84028
rect 4844 83916 5404 83972
rect 5460 83916 5470 83972
rect 7858 83916 7868 83972
rect 7924 83916 8204 83972
rect 8260 83916 8270 83972
rect 4454 83860 4464 83916
rect 4520 83860 4568 83916
rect 4624 83860 4672 83916
rect 4728 83860 4738 83916
rect 8428 83860 8484 84028
rect 12796 83860 12852 84028
rect 15026 83916 15036 83972
rect 15092 83916 17500 83972
rect 17556 83916 17566 83972
rect 24454 83860 24464 83916
rect 24520 83860 24568 83916
rect 24624 83860 24672 83916
rect 24728 83860 24738 83916
rect 31584 83860 31696 83888
rect 8418 83804 8428 83860
rect 8484 83804 8494 83860
rect 12786 83804 12796 83860
rect 12852 83804 12862 83860
rect 30594 83804 30604 83860
rect 30660 83804 31696 83860
rect 31584 83776 31696 83804
rect 0 83748 112 83776
rect 0 83692 252 83748
rect 308 83692 318 83748
rect 1810 83692 1820 83748
rect 1876 83692 5404 83748
rect 5460 83692 5470 83748
rect 5618 83692 5628 83748
rect 5684 83692 9884 83748
rect 9940 83692 9950 83748
rect 13010 83692 13020 83748
rect 13076 83692 13244 83748
rect 13300 83692 13310 83748
rect 0 83664 112 83692
rect 2370 83580 2380 83636
rect 2436 83580 2716 83636
rect 2772 83580 2782 83636
rect 5058 83580 5068 83636
rect 5124 83580 5134 83636
rect 8866 83580 8876 83636
rect 8932 83580 8988 83636
rect 9044 83580 9054 83636
rect 690 83468 700 83524
rect 756 83468 3948 83524
rect 4004 83468 4014 83524
rect 1922 83356 1932 83412
rect 1988 83356 3388 83412
rect 0 83300 112 83328
rect 3332 83300 3388 83356
rect 5068 83300 5124 83580
rect 6962 83468 6972 83524
rect 7028 83468 9212 83524
rect 9268 83468 9278 83524
rect 9874 83468 9884 83524
rect 9940 83468 10332 83524
rect 10388 83468 10398 83524
rect 16034 83468 16044 83524
rect 16100 83468 17052 83524
rect 17108 83468 17118 83524
rect 8866 83356 8876 83412
rect 8932 83356 9772 83412
rect 9828 83356 9838 83412
rect 14354 83356 14364 83412
rect 14420 83356 14476 83412
rect 14532 83356 14812 83412
rect 14868 83356 14878 83412
rect 0 83244 364 83300
rect 420 83244 430 83300
rect 3332 83244 5852 83300
rect 5908 83244 9212 83300
rect 9268 83244 9278 83300
rect 12002 83244 12012 83300
rect 12068 83244 13468 83300
rect 13524 83244 13534 83300
rect 18834 83244 18844 83300
rect 18900 83244 19516 83300
rect 19572 83244 19582 83300
rect 0 83216 112 83244
rect 5394 83132 5404 83188
rect 5460 83132 11340 83188
rect 11396 83132 11676 83188
rect 11732 83132 11742 83188
rect 12450 83132 12460 83188
rect 12516 83132 14588 83188
rect 14644 83132 14654 83188
rect 3794 83076 3804 83132
rect 3860 83076 3908 83132
rect 3964 83076 4012 83132
rect 4068 83076 4078 83132
rect 23794 83076 23804 83132
rect 23860 83076 23908 83132
rect 23964 83076 24012 83132
rect 24068 83076 24078 83132
rect 3332 82908 11004 82964
rect 11060 82908 11070 82964
rect 14466 82908 14476 82964
rect 14532 82908 16044 82964
rect 16100 82908 16110 82964
rect 0 82852 112 82880
rect 3332 82852 3388 82908
rect 0 82796 3388 82852
rect 5618 82796 5628 82852
rect 5684 82796 5852 82852
rect 5908 82796 5918 82852
rect 8754 82796 8764 82852
rect 8820 82796 16940 82852
rect 16996 82796 18060 82852
rect 18116 82796 18126 82852
rect 0 82768 112 82796
rect 31584 82740 31696 82768
rect 1698 82684 1708 82740
rect 1764 82684 1820 82740
rect 1876 82684 1886 82740
rect 2818 82684 2828 82740
rect 2884 82684 3052 82740
rect 3108 82684 3118 82740
rect 5282 82684 5292 82740
rect 5348 82684 8316 82740
rect 8372 82684 8382 82740
rect 10210 82684 10220 82740
rect 10276 82684 14028 82740
rect 14084 82684 14924 82740
rect 14980 82684 14990 82740
rect 30594 82684 30604 82740
rect 30660 82684 31696 82740
rect 31584 82656 31696 82684
rect 1708 82572 12012 82628
rect 12068 82572 12078 82628
rect 16706 82572 16716 82628
rect 16772 82572 22428 82628
rect 22484 82572 22494 82628
rect 22866 82572 22876 82628
rect 22932 82572 30268 82628
rect 30324 82572 30334 82628
rect 0 82404 112 82432
rect 1708 82404 1764 82572
rect 2258 82460 2268 82516
rect 2324 82460 8092 82516
rect 8148 82460 8158 82516
rect 8306 82460 8316 82516
rect 8372 82460 10108 82516
rect 10164 82460 10174 82516
rect 10322 82460 10332 82516
rect 10388 82460 10556 82516
rect 10612 82460 13020 82516
rect 13076 82460 14476 82516
rect 14532 82460 14542 82516
rect 15922 82460 15932 82516
rect 15988 82460 16604 82516
rect 16660 82460 16670 82516
rect 18498 82460 18508 82516
rect 18564 82460 26460 82516
rect 26516 82460 26526 82516
rect 0 82348 1764 82404
rect 5282 82348 5292 82404
rect 5348 82348 5460 82404
rect 7074 82348 7084 82404
rect 7140 82348 11004 82404
rect 11060 82348 11070 82404
rect 11890 82348 11900 82404
rect 11956 82348 17388 82404
rect 17444 82348 17454 82404
rect 0 82320 112 82348
rect 4454 82292 4464 82348
rect 4520 82292 4568 82348
rect 4624 82292 4672 82348
rect 4728 82292 4738 82348
rect 5404 82292 5460 82348
rect 24454 82292 24464 82348
rect 24520 82292 24568 82348
rect 24624 82292 24672 82348
rect 24728 82292 24738 82348
rect 1586 82236 1596 82292
rect 1652 82236 2156 82292
rect 2212 82236 2222 82292
rect 2370 82236 2380 82292
rect 2436 82236 2716 82292
rect 2772 82236 2782 82292
rect 5404 82236 8316 82292
rect 8372 82236 8382 82292
rect 14018 82236 14028 82292
rect 14084 82236 15036 82292
rect 15092 82236 18172 82292
rect 18228 82236 18238 82292
rect 2034 82124 2044 82180
rect 2100 82124 6748 82180
rect 6804 82124 6814 82180
rect 7074 82124 7084 82180
rect 7140 82124 8540 82180
rect 8596 82124 8606 82180
rect 10098 82124 10108 82180
rect 10164 82124 14308 82180
rect 14466 82124 14476 82180
rect 14532 82124 15764 82180
rect 20514 82124 20524 82180
rect 20580 82124 21196 82180
rect 21252 82124 21262 82180
rect 14252 82068 14308 82124
rect 15708 82068 15764 82124
rect 1138 82012 1148 82068
rect 1204 82012 1484 82068
rect 1540 82012 3724 82068
rect 3780 82012 5068 82068
rect 5124 82012 5134 82068
rect 7858 82012 7868 82068
rect 7924 82012 8428 82068
rect 8484 82012 8494 82068
rect 12898 82012 12908 82068
rect 12964 82012 13468 82068
rect 13524 82012 13534 82068
rect 14252 82012 15540 82068
rect 15698 82012 15708 82068
rect 15764 82012 15774 82068
rect 19954 82012 19964 82068
rect 20020 82012 22540 82068
rect 22596 82012 22606 82068
rect 0 81956 112 81984
rect 15484 81956 15540 82012
rect 0 81900 9324 81956
rect 9380 81900 9390 81956
rect 11106 81900 11116 81956
rect 11172 81900 14252 81956
rect 14308 81900 14318 81956
rect 15484 81900 19404 81956
rect 19460 81900 20412 81956
rect 20468 81900 20478 81956
rect 21186 81900 21196 81956
rect 21252 81900 29484 81956
rect 29540 81900 29550 81956
rect 0 81872 112 81900
rect 20412 81844 20468 81900
rect 2118 81788 2156 81844
rect 2212 81788 2492 81844
rect 2548 81788 14924 81844
rect 14980 81788 14990 81844
rect 20412 81788 23212 81844
rect 23268 81788 23278 81844
rect 14476 81732 14532 81788
rect 3042 81676 3052 81732
rect 3108 81676 3276 81732
rect 3332 81676 3342 81732
rect 3602 81676 3612 81732
rect 3668 81676 4508 81732
rect 4564 81676 4574 81732
rect 5394 81676 5404 81732
rect 5460 81676 14028 81732
rect 14084 81676 14094 81732
rect 14466 81676 14476 81732
rect 14532 81676 14542 81732
rect 14802 81676 14812 81732
rect 14868 81676 15484 81732
rect 15540 81676 15550 81732
rect 3612 81620 3668 81676
rect 31584 81620 31696 81648
rect 3378 81564 3388 81620
rect 3444 81564 3668 81620
rect 6402 81564 6412 81620
rect 6468 81564 15148 81620
rect 30594 81564 30604 81620
rect 30660 81564 31696 81620
rect 0 81508 112 81536
rect 3794 81508 3804 81564
rect 3860 81508 3908 81564
rect 3964 81508 4012 81564
rect 4068 81508 4078 81564
rect 0 81452 3388 81508
rect 4834 81452 4844 81508
rect 4900 81452 9100 81508
rect 9156 81452 9166 81508
rect 9314 81452 9324 81508
rect 9380 81452 10668 81508
rect 10724 81452 10734 81508
rect 14354 81452 14364 81508
rect 14420 81452 14588 81508
rect 14644 81452 14654 81508
rect 0 81424 112 81452
rect 3332 81396 3388 81452
rect 15092 81396 15148 81564
rect 23794 81508 23804 81564
rect 23860 81508 23908 81564
rect 23964 81508 24012 81564
rect 24068 81508 24078 81564
rect 31584 81536 31696 81564
rect 15922 81452 15932 81508
rect 15988 81452 16156 81508
rect 16212 81452 16222 81508
rect 3332 81340 7420 81396
rect 7476 81340 9100 81396
rect 9156 81340 9166 81396
rect 13010 81340 13020 81396
rect 13076 81340 13132 81396
rect 13188 81340 13198 81396
rect 13906 81340 13916 81396
rect 13972 81340 14700 81396
rect 14756 81340 14766 81396
rect 15092 81340 18396 81396
rect 18452 81340 20916 81396
rect 20860 81284 20916 81340
rect 4162 81228 4172 81284
rect 4228 81228 6748 81284
rect 6804 81228 8092 81284
rect 8148 81228 8158 81284
rect 10108 81228 14868 81284
rect 15110 81228 15148 81284
rect 15204 81228 15214 81284
rect 15474 81228 15484 81284
rect 15540 81228 15708 81284
rect 15764 81228 19292 81284
rect 19348 81228 19358 81284
rect 20850 81228 20860 81284
rect 20916 81228 21980 81284
rect 22036 81228 22046 81284
rect 3332 81116 9884 81172
rect 9940 81116 9950 81172
rect 0 81060 112 81088
rect 3332 81060 3388 81116
rect 10108 81060 10164 81228
rect 14812 81172 14868 81228
rect 12338 81116 12348 81172
rect 12404 81116 12908 81172
rect 12964 81116 12974 81172
rect 13682 81116 13692 81172
rect 13748 81116 14588 81172
rect 14644 81116 14654 81172
rect 14802 81116 14812 81172
rect 14868 81116 21196 81172
rect 21252 81116 21262 81172
rect 0 81004 3388 81060
rect 4284 81004 6412 81060
rect 6468 81004 6478 81060
rect 6626 81004 6636 81060
rect 6692 81004 7756 81060
rect 7812 81004 7822 81060
rect 7980 81004 8540 81060
rect 8596 81004 9492 81060
rect 9650 81004 9660 81060
rect 9716 81004 10164 81060
rect 0 80976 112 81004
rect 802 80892 812 80948
rect 868 80892 3948 80948
rect 4004 80892 4014 80948
rect 4284 80836 4340 81004
rect 4498 80892 4508 80948
rect 4564 80892 4844 80948
rect 4900 80892 4910 80948
rect 7980 80836 8036 81004
rect 9436 80948 9492 81004
rect 12908 80948 12964 81116
rect 14588 81060 14644 81116
rect 14588 81004 15036 81060
rect 15092 81004 15102 81060
rect 21298 81004 21308 81060
rect 21364 81004 21532 81060
rect 21588 81004 21598 81060
rect 9436 80892 10332 80948
rect 10388 80892 10398 80948
rect 10770 80892 10780 80948
rect 10836 80892 12236 80948
rect 12292 80892 12302 80948
rect 12908 80892 15484 80948
rect 15540 80892 15550 80948
rect 22390 80892 22428 80948
rect 22484 80892 22494 80948
rect 914 80780 924 80836
rect 980 80780 4340 80836
rect 6178 80780 6188 80836
rect 6244 80780 6636 80836
rect 6692 80780 8036 80836
rect 8194 80780 8204 80836
rect 8260 80780 13468 80836
rect 13524 80780 18844 80836
rect 18900 80780 19964 80836
rect 20020 80780 20030 80836
rect 22194 80780 22204 80836
rect 22260 80780 22652 80836
rect 22708 80780 22718 80836
rect 4454 80724 4464 80780
rect 4520 80724 4568 80780
rect 4624 80724 4672 80780
rect 4728 80724 4738 80780
rect 24454 80724 24464 80780
rect 24520 80724 24568 80780
rect 24624 80724 24672 80780
rect 24728 80724 24738 80780
rect 5058 80668 5068 80724
rect 5124 80668 5740 80724
rect 5796 80668 5806 80724
rect 13346 80668 13356 80724
rect 13412 80668 14812 80724
rect 14868 80668 14878 80724
rect 15026 80668 15036 80724
rect 15092 80668 15130 80724
rect 21858 80668 21868 80724
rect 21924 80668 22876 80724
rect 22932 80668 22942 80724
rect 0 80612 112 80640
rect 0 80556 8260 80612
rect 0 80528 112 80556
rect 2482 80444 2492 80500
rect 2548 80444 3612 80500
rect 3668 80444 3678 80500
rect 6514 80444 6524 80500
rect 6580 80444 7196 80500
rect 7252 80444 7262 80500
rect 8204 80388 8260 80556
rect 10220 80556 11228 80612
rect 11284 80556 12908 80612
rect 12964 80556 12974 80612
rect 15138 80556 15148 80612
rect 15204 80556 15820 80612
rect 15876 80556 15886 80612
rect 20290 80556 20300 80612
rect 20356 80556 21420 80612
rect 21476 80556 21486 80612
rect 10220 80500 10276 80556
rect 12908 80500 12964 80556
rect 31584 80500 31696 80528
rect 10210 80444 10220 80500
rect 10276 80444 10286 80500
rect 12908 80444 21980 80500
rect 22036 80444 22764 80500
rect 22820 80444 22830 80500
rect 30594 80444 30604 80500
rect 30660 80444 31696 80500
rect 31584 80416 31696 80444
rect 2034 80332 2044 80388
rect 2100 80332 2380 80388
rect 2436 80332 2828 80388
rect 2884 80332 2894 80388
rect 3266 80332 3276 80388
rect 3332 80332 3612 80388
rect 3668 80332 3678 80388
rect 8204 80332 23548 80388
rect 23604 80332 23614 80388
rect 1026 80220 1036 80276
rect 1092 80220 6076 80276
rect 6132 80220 6142 80276
rect 6738 80220 6748 80276
rect 6804 80220 14700 80276
rect 14756 80220 14766 80276
rect 0 80164 112 80192
rect 0 80108 1708 80164
rect 1764 80108 1774 80164
rect 2258 80108 2268 80164
rect 2324 80108 3164 80164
rect 3220 80108 5852 80164
rect 5908 80108 6188 80164
rect 6244 80108 10556 80164
rect 10612 80108 10622 80164
rect 14914 80108 14924 80164
rect 14980 80108 22204 80164
rect 22260 80108 22270 80164
rect 0 80080 112 80108
rect 578 79996 588 80052
rect 644 79996 1932 80052
rect 1988 79996 1998 80052
rect 9874 79996 9884 80052
rect 9940 79996 10332 80052
rect 10388 79996 10398 80052
rect 26534 79996 26572 80052
rect 26628 79996 26638 80052
rect 3794 79940 3804 79996
rect 3860 79940 3908 79996
rect 3964 79940 4012 79996
rect 4068 79940 4078 79996
rect 23794 79940 23804 79996
rect 23860 79940 23908 79996
rect 23964 79940 24012 79996
rect 24068 79940 24078 79996
rect 9090 79884 9100 79940
rect 9156 79884 10556 79940
rect 10612 79884 10622 79940
rect 10882 79884 10892 79940
rect 10948 79884 11452 79940
rect 11508 79884 11518 79940
rect 578 79772 588 79828
rect 644 79772 4956 79828
rect 5012 79772 5022 79828
rect 8642 79772 8652 79828
rect 8708 79772 9100 79828
rect 9156 79772 9166 79828
rect 10434 79772 10444 79828
rect 10500 79772 10510 79828
rect 22082 79772 22092 79828
rect 22148 79772 22428 79828
rect 22484 79772 22494 79828
rect 0 79716 112 79744
rect 10444 79716 10500 79772
rect 0 79660 11452 79716
rect 11508 79660 11518 79716
rect 11732 79660 29484 79716
rect 29540 79660 29550 79716
rect 0 79632 112 79660
rect 11732 79604 11788 79660
rect 1698 79548 1708 79604
rect 1764 79548 7532 79604
rect 7588 79548 7598 79604
rect 7858 79548 7868 79604
rect 7924 79548 8764 79604
rect 8820 79548 8830 79604
rect 10322 79548 10332 79604
rect 10388 79548 11788 79604
rect 14354 79548 14364 79604
rect 14420 79548 15148 79604
rect 15204 79548 15214 79604
rect 15586 79548 15596 79604
rect 15652 79548 16716 79604
rect 16772 79548 16782 79604
rect 17826 79548 17836 79604
rect 17892 79548 18732 79604
rect 18788 79548 18798 79604
rect 19954 79548 19964 79604
rect 20020 79548 20748 79604
rect 20804 79548 20972 79604
rect 21028 79548 21038 79604
rect 22306 79548 22316 79604
rect 22372 79548 22428 79604
rect 22484 79548 22494 79604
rect 23762 79548 23772 79604
rect 23828 79548 25004 79604
rect 25060 79548 25070 79604
rect 1250 79436 1260 79492
rect 1316 79436 1932 79492
rect 1988 79436 1998 79492
rect 6738 79436 6748 79492
rect 6804 79436 6860 79492
rect 6916 79436 6926 79492
rect 8418 79436 8428 79492
rect 8484 79436 12124 79492
rect 12180 79436 12190 79492
rect 12898 79436 12908 79492
rect 12964 79436 13132 79492
rect 13188 79436 16604 79492
rect 16660 79436 16670 79492
rect 31584 79380 31696 79408
rect 2482 79324 2492 79380
rect 2548 79324 2828 79380
rect 2884 79324 2894 79380
rect 3378 79324 3388 79380
rect 3444 79324 3482 79380
rect 4284 79324 5404 79380
rect 5460 79324 5470 79380
rect 5842 79324 5852 79380
rect 5908 79324 6412 79380
rect 6468 79324 7196 79380
rect 7252 79324 7262 79380
rect 9090 79324 9100 79380
rect 9156 79324 9436 79380
rect 9492 79324 9502 79380
rect 10098 79324 10108 79380
rect 10164 79324 10332 79380
rect 10388 79324 10398 79380
rect 10546 79324 10556 79380
rect 10612 79324 11228 79380
rect 11284 79324 17948 79380
rect 18004 79324 18014 79380
rect 30594 79324 30604 79380
rect 30660 79324 31696 79380
rect 0 79268 112 79296
rect 4284 79268 4340 79324
rect 31584 79296 31696 79324
rect 0 79212 4340 79268
rect 8082 79212 8092 79268
rect 8148 79212 20076 79268
rect 20132 79212 20142 79268
rect 0 79184 112 79212
rect 4454 79156 4464 79212
rect 4520 79156 4568 79212
rect 4624 79156 4672 79212
rect 4728 79156 4738 79212
rect 24454 79156 24464 79212
rect 24520 79156 24568 79212
rect 24624 79156 24672 79212
rect 24728 79156 24738 79212
rect 914 79100 924 79156
rect 980 79100 4060 79156
rect 4116 79100 4126 79156
rect 6850 79100 6860 79156
rect 6916 79100 8428 79156
rect 8484 79100 8494 79156
rect 14914 79100 14924 79156
rect 14980 79100 17612 79156
rect 17668 79100 17678 79156
rect 1474 78988 1484 79044
rect 1540 78988 1708 79044
rect 1764 78988 1774 79044
rect 2706 78988 2716 79044
rect 2772 78988 8540 79044
rect 8596 78988 8606 79044
rect 11442 78988 11452 79044
rect 11508 78988 11676 79044
rect 11732 78988 11742 79044
rect 12562 78988 12572 79044
rect 12628 78988 13132 79044
rect 13188 78988 13198 79044
rect 16370 78988 16380 79044
rect 16436 78988 17276 79044
rect 17332 78988 17500 79044
rect 17556 78988 17566 79044
rect 690 78876 700 78932
rect 756 78876 1708 78932
rect 1764 78876 1774 78932
rect 3332 78876 7308 78932
rect 7364 78876 7374 78932
rect 8306 78876 8316 78932
rect 8372 78876 9548 78932
rect 9604 78876 9614 78932
rect 11218 78876 11228 78932
rect 11284 78876 11676 78932
rect 11732 78876 11742 78932
rect 12002 78876 12012 78932
rect 12068 78876 12348 78932
rect 12404 78876 14252 78932
rect 14308 78876 14318 78932
rect 17602 78876 17612 78932
rect 17668 78876 20188 78932
rect 20244 78876 20254 78932
rect 22082 78876 22092 78932
rect 22148 78876 22876 78932
rect 22932 78876 29484 78932
rect 29540 78876 29550 78932
rect 0 78820 112 78848
rect 3332 78820 3388 78876
rect 0 78764 3388 78820
rect 3938 78764 3948 78820
rect 4004 78764 15148 78820
rect 16034 78764 16044 78820
rect 16100 78764 17052 78820
rect 17108 78764 17118 78820
rect 17602 78764 17612 78820
rect 17668 78764 18172 78820
rect 18228 78764 18238 78820
rect 20514 78764 20524 78820
rect 20580 78764 22316 78820
rect 22372 78764 22382 78820
rect 0 78736 112 78764
rect 2370 78652 2380 78708
rect 2436 78652 2940 78708
rect 2996 78652 6076 78708
rect 6132 78652 6142 78708
rect 10770 78652 10780 78708
rect 10836 78652 11228 78708
rect 11284 78652 11294 78708
rect 11666 78652 11676 78708
rect 11732 78652 12628 78708
rect 15092 78652 15148 78764
rect 15204 78652 16156 78708
rect 16212 78652 16222 78708
rect 12572 78596 12628 78652
rect 1698 78540 1708 78596
rect 1764 78540 9324 78596
rect 9380 78540 9390 78596
rect 11442 78540 11452 78596
rect 11508 78540 12236 78596
rect 12292 78540 12302 78596
rect 12562 78540 12572 78596
rect 12628 78540 12638 78596
rect 15810 78540 15820 78596
rect 15876 78540 20300 78596
rect 20356 78540 21084 78596
rect 21140 78540 21150 78596
rect 7074 78428 7084 78484
rect 7140 78428 7980 78484
rect 8036 78428 8046 78484
rect 9650 78428 9660 78484
rect 9716 78428 12012 78484
rect 12068 78428 12078 78484
rect 0 78372 112 78400
rect 3794 78372 3804 78428
rect 3860 78372 3908 78428
rect 3964 78372 4012 78428
rect 4068 78372 4078 78428
rect 23794 78372 23804 78428
rect 23860 78372 23908 78428
rect 23964 78372 24012 78428
rect 24068 78372 24078 78428
rect 0 78316 1820 78372
rect 1876 78316 1886 78372
rect 3490 78316 3500 78372
rect 3556 78316 3566 78372
rect 4162 78316 4172 78372
rect 4228 78316 5404 78372
rect 5460 78316 5470 78372
rect 6066 78316 6076 78372
rect 6132 78316 10892 78372
rect 10948 78316 10958 78372
rect 11218 78316 11228 78372
rect 11284 78316 12348 78372
rect 12404 78316 12414 78372
rect 14578 78316 14588 78372
rect 14644 78316 14812 78372
rect 14868 78316 14878 78372
rect 0 78288 112 78316
rect 3500 78260 3556 78316
rect 31584 78260 31696 78288
rect 1922 78204 1932 78260
rect 1988 78204 5628 78260
rect 5684 78204 5694 78260
rect 5852 78204 8932 78260
rect 9090 78204 9100 78260
rect 9156 78204 10108 78260
rect 10164 78204 10444 78260
rect 10500 78204 11340 78260
rect 11396 78204 13020 78260
rect 13076 78204 13086 78260
rect 13244 78204 18732 78260
rect 18788 78204 18798 78260
rect 30594 78204 30604 78260
rect 30660 78204 31696 78260
rect 5852 78148 5908 78204
rect 1250 78092 1260 78148
rect 1316 78092 1820 78148
rect 1876 78092 2716 78148
rect 2772 78092 2782 78148
rect 5394 78092 5404 78148
rect 5460 78092 5908 78148
rect 6850 78092 6860 78148
rect 6916 78092 8316 78148
rect 8372 78092 8382 78148
rect 1708 77980 7084 78036
rect 7140 77980 7150 78036
rect 7858 77980 7868 78036
rect 7924 77980 8148 78036
rect 0 77924 112 77952
rect 1708 77924 1764 77980
rect 0 77868 1764 77924
rect 3042 77868 3052 77924
rect 3108 77868 3388 77924
rect 3444 77868 3454 77924
rect 5590 77868 5628 77924
rect 5684 77868 6412 77924
rect 6468 77868 6478 77924
rect 0 77840 112 77868
rect 3154 77756 3164 77812
rect 3220 77756 3276 77812
rect 3332 77756 3342 77812
rect 3602 77756 3612 77812
rect 3668 77756 4172 77812
rect 4228 77756 4238 77812
rect 7410 77756 7420 77812
rect 7476 77756 7868 77812
rect 7924 77756 7934 77812
rect 8092 77700 8148 77980
rect 8876 77924 8932 78204
rect 9426 78092 9436 78148
rect 9492 78092 12236 78148
rect 12292 78092 12302 78148
rect 13244 78036 13300 78204
rect 31584 78176 31696 78204
rect 13682 78092 13692 78148
rect 13748 78092 15820 78148
rect 15876 78092 15886 78148
rect 9538 77980 9548 78036
rect 9604 77980 13300 78036
rect 15138 77980 15148 78036
rect 15204 77980 15484 78036
rect 15540 77980 16828 78036
rect 16884 77980 16894 78036
rect 8876 77868 9772 77924
rect 9828 77868 9838 77924
rect 10322 77868 10332 77924
rect 10388 77868 10556 77924
rect 10612 77868 10622 77924
rect 15922 77868 15932 77924
rect 15988 77868 19628 77924
rect 19684 77868 29484 77924
rect 29540 77868 29550 77924
rect 15932 77812 15988 77868
rect 8530 77756 8540 77812
rect 8596 77756 10892 77812
rect 10948 77756 15988 77812
rect 18722 77756 18732 77812
rect 18788 77756 29372 77812
rect 29428 77756 29438 77812
rect 8092 77644 8988 77700
rect 9044 77644 9660 77700
rect 9716 77644 9726 77700
rect 20178 77644 20188 77700
rect 20244 77644 22988 77700
rect 23044 77644 23054 77700
rect 4454 77588 4464 77644
rect 4520 77588 4568 77644
rect 4624 77588 4672 77644
rect 4728 77588 4738 77644
rect 24454 77588 24464 77644
rect 24520 77588 24568 77644
rect 24624 77588 24672 77644
rect 24728 77588 24738 77644
rect 2034 77532 2044 77588
rect 2100 77532 3052 77588
rect 3108 77532 3118 77588
rect 5516 77532 7756 77588
rect 7812 77532 7822 77588
rect 8418 77532 8428 77588
rect 8484 77532 9548 77588
rect 9604 77532 9614 77588
rect 20738 77532 20748 77588
rect 20804 77532 21196 77588
rect 21252 77532 21262 77588
rect 0 77476 112 77504
rect 5516 77476 5572 77532
rect 0 77420 5572 77476
rect 6598 77420 6636 77476
rect 6692 77420 6702 77476
rect 9426 77420 9436 77476
rect 9492 77420 15148 77476
rect 0 77392 112 77420
rect 15092 77364 15148 77420
rect 17388 77420 22092 77476
rect 22148 77420 22158 77476
rect 17388 77364 17444 77420
rect 1586 77308 1596 77364
rect 1652 77308 3948 77364
rect 4004 77308 4014 77364
rect 4834 77308 4844 77364
rect 4900 77308 5068 77364
rect 5124 77308 5134 77364
rect 5282 77308 5292 77364
rect 5348 77308 11676 77364
rect 11732 77308 11742 77364
rect 15092 77308 17388 77364
rect 17444 77308 17454 77364
rect 17602 77308 17612 77364
rect 17668 77308 20412 77364
rect 20468 77308 20478 77364
rect 20738 77308 20748 77364
rect 20804 77308 21420 77364
rect 21476 77308 21486 77364
rect 2146 77196 2156 77252
rect 2212 77196 2380 77252
rect 2436 77196 2446 77252
rect 3378 77196 3388 77252
rect 3444 77196 5180 77252
rect 5236 77196 5246 77252
rect 8082 77196 8092 77252
rect 8148 77196 9324 77252
rect 9380 77196 9390 77252
rect 9538 77196 9548 77252
rect 9604 77196 10892 77252
rect 10948 77196 10958 77252
rect 11442 77196 11452 77252
rect 11508 77196 12124 77252
rect 12180 77196 12190 77252
rect 19954 77196 19964 77252
rect 20020 77196 20636 77252
rect 20692 77196 20702 77252
rect 0 77028 112 77056
rect 2380 77028 2436 77196
rect 4274 77084 4284 77140
rect 4340 77084 4396 77140
rect 4452 77084 4462 77140
rect 7522 77084 7532 77140
rect 7588 77084 13468 77140
rect 13524 77084 13534 77140
rect 0 76972 588 77028
rect 644 76972 654 77028
rect 2380 76972 4172 77028
rect 4228 76972 4238 77028
rect 9202 76972 9212 77028
rect 9268 76972 10668 77028
rect 10724 76972 10734 77028
rect 18162 76972 18172 77028
rect 18228 76972 18508 77028
rect 18564 76972 18574 77028
rect 0 76944 112 76972
rect 2706 76860 2716 76916
rect 2772 76860 3164 76916
rect 3220 76860 3230 76916
rect 5842 76860 5852 76916
rect 5908 76860 15148 76916
rect 15474 76860 15484 76916
rect 15540 76860 16492 76916
rect 16548 76860 21588 76916
rect 3794 76804 3804 76860
rect 3860 76804 3908 76860
rect 3964 76804 4012 76860
rect 4068 76804 4078 76860
rect 15092 76804 15148 76860
rect 21532 76804 21588 76860
rect 23794 76804 23804 76860
rect 23860 76804 23908 76860
rect 23964 76804 24012 76860
rect 24068 76804 24078 76860
rect 242 76748 252 76804
rect 308 76748 1036 76804
rect 1092 76748 1102 76804
rect 3332 76748 3612 76804
rect 3668 76748 3678 76804
rect 6626 76748 6636 76804
rect 6692 76748 12908 76804
rect 12964 76748 12974 76804
rect 15092 76748 19404 76804
rect 19460 76748 19470 76804
rect 21522 76748 21532 76804
rect 21588 76748 21598 76804
rect 3332 76692 3388 76748
rect 914 76636 924 76692
rect 980 76636 990 76692
rect 2594 76636 2604 76692
rect 2660 76636 3388 76692
rect 0 76580 112 76608
rect 0 76524 140 76580
rect 196 76524 206 76580
rect 0 76496 112 76524
rect 0 76132 112 76160
rect 924 76132 980 76636
rect 1698 76524 1708 76580
rect 1764 76524 2156 76580
rect 2212 76524 6636 76580
rect 6692 76524 6702 76580
rect 6962 76524 6972 76580
rect 7028 76524 11900 76580
rect 11956 76524 11966 76580
rect 12674 76524 12684 76580
rect 12740 76524 12908 76580
rect 12964 76524 17724 76580
rect 17780 76524 17790 76580
rect 26226 76524 26236 76580
rect 26292 76524 26684 76580
rect 26740 76524 26750 76580
rect 3154 76412 3164 76468
rect 3220 76412 3388 76468
rect 3444 76412 3454 76468
rect 3602 76412 3612 76468
rect 3668 76412 5740 76468
rect 5796 76412 5806 76468
rect 8866 76412 8876 76468
rect 8932 76412 9884 76468
rect 9940 76412 9950 76468
rect 12114 76412 12124 76468
rect 12180 76412 13244 76468
rect 13300 76412 13310 76468
rect 17938 76412 17948 76468
rect 18004 76412 18396 76468
rect 18452 76412 19516 76468
rect 19572 76412 19582 76468
rect 21410 76412 21420 76468
rect 21476 76412 22316 76468
rect 22372 76412 22382 76468
rect 26534 76412 26572 76468
rect 26628 76412 26638 76468
rect 2370 76300 2380 76356
rect 2436 76300 2716 76356
rect 2772 76300 2782 76356
rect 5058 76300 5068 76356
rect 5124 76300 7644 76356
rect 7700 76300 7710 76356
rect 10210 76300 10220 76356
rect 10276 76300 10892 76356
rect 10948 76300 11228 76356
rect 11284 76300 11294 76356
rect 17266 76300 17276 76356
rect 17332 76300 18844 76356
rect 18900 76300 18910 76356
rect 20514 76300 20524 76356
rect 20580 76300 21308 76356
rect 21364 76300 21868 76356
rect 21924 76300 21934 76356
rect 1250 76188 1260 76244
rect 1316 76188 1372 76244
rect 1428 76188 1438 76244
rect 5954 76188 5964 76244
rect 6020 76188 8092 76244
rect 8148 76188 8158 76244
rect 20738 76188 20748 76244
rect 20804 76188 21084 76244
rect 21140 76188 21150 76244
rect 0 76076 980 76132
rect 6290 76076 6300 76132
rect 6356 76076 10556 76132
rect 10612 76076 10622 76132
rect 0 76048 112 76076
rect 4454 76020 4464 76076
rect 4520 76020 4568 76076
rect 4624 76020 4672 76076
rect 4728 76020 4738 76076
rect 24454 76020 24464 76076
rect 24520 76020 24568 76076
rect 24624 76020 24672 76076
rect 24728 76020 24738 76076
rect 13570 75964 13580 76020
rect 13636 75964 14028 76020
rect 14084 75964 14094 76020
rect 1474 75852 1484 75908
rect 1540 75852 1550 75908
rect 6178 75852 6188 75908
rect 6244 75852 6524 75908
rect 6580 75852 6692 75908
rect 7046 75852 7084 75908
rect 7140 75852 7980 75908
rect 8036 75852 8046 75908
rect 17490 75852 17500 75908
rect 17556 75852 18060 75908
rect 18116 75852 18126 75908
rect 0 75684 112 75712
rect 0 75628 1260 75684
rect 1316 75628 1326 75684
rect 0 75600 112 75628
rect 1484 75572 1540 75852
rect 6636 75796 6692 75852
rect 1922 75740 1932 75796
rect 1988 75740 5852 75796
rect 5908 75740 5918 75796
rect 6626 75740 6636 75796
rect 6692 75740 12348 75796
rect 12404 75740 12414 75796
rect 20402 75740 20412 75796
rect 20468 75740 21756 75796
rect 21812 75740 21822 75796
rect 2258 75628 2268 75684
rect 2324 75628 2940 75684
rect 2996 75628 3006 75684
rect 3938 75628 3948 75684
rect 4004 75628 6188 75684
rect 6244 75628 6254 75684
rect 8194 75628 8204 75684
rect 8260 75628 8540 75684
rect 8596 75628 8606 75684
rect 1260 75516 1540 75572
rect 2146 75516 2156 75572
rect 2212 75516 2492 75572
rect 2548 75516 2558 75572
rect 12226 75516 12236 75572
rect 12292 75516 12572 75572
rect 12628 75516 12638 75572
rect 16146 75516 16156 75572
rect 16212 75516 17388 75572
rect 17444 75516 17454 75572
rect 1260 75460 1316 75516
rect 18 75404 28 75460
rect 84 75404 924 75460
rect 980 75404 990 75460
rect 1250 75404 1260 75460
rect 1316 75404 1326 75460
rect 4162 75404 4172 75460
rect 4228 75404 4956 75460
rect 5012 75404 5022 75460
rect 20178 75404 20188 75460
rect 20244 75404 22988 75460
rect 23044 75404 23054 75460
rect 0 75236 112 75264
rect 3794 75236 3804 75292
rect 3860 75236 3908 75292
rect 3964 75236 4012 75292
rect 4068 75236 4078 75292
rect 23794 75236 23804 75292
rect 23860 75236 23908 75292
rect 23964 75236 24012 75292
rect 24068 75236 24078 75292
rect 0 75180 812 75236
rect 868 75180 878 75236
rect 8194 75180 8204 75236
rect 8260 75180 8428 75236
rect 8484 75180 8494 75236
rect 0 75152 112 75180
rect 4274 75068 4284 75124
rect 4340 75068 5852 75124
rect 5908 75068 5918 75124
rect 10994 75068 11004 75124
rect 11060 75068 11676 75124
rect 11732 75068 16268 75124
rect 16324 75068 16334 75124
rect 16818 75068 16828 75124
rect 16884 75068 17052 75124
rect 17108 75068 17118 75124
rect 17826 75068 17836 75124
rect 17892 75068 18732 75124
rect 18788 75068 19740 75124
rect 19796 75068 19806 75124
rect 4386 74956 4396 75012
rect 4452 74956 20524 75012
rect 20580 74956 20590 75012
rect 2258 74844 2268 74900
rect 2324 74844 3836 74900
rect 3892 74844 3902 74900
rect 4246 74844 4284 74900
rect 4340 74844 4350 74900
rect 12114 74844 12124 74900
rect 12180 74844 13132 74900
rect 13188 74844 13198 74900
rect 16034 74844 16044 74900
rect 16100 74844 17052 74900
rect 17108 74844 17118 74900
rect 0 74788 112 74816
rect 0 74732 700 74788
rect 756 74732 766 74788
rect 2930 74732 2940 74788
rect 2996 74732 4956 74788
rect 5012 74732 5022 74788
rect 12002 74732 12012 74788
rect 12068 74732 13804 74788
rect 13860 74732 13870 74788
rect 14354 74732 14364 74788
rect 14420 74732 14812 74788
rect 14868 74732 14878 74788
rect 16706 74732 16716 74788
rect 16772 74732 17612 74788
rect 17668 74732 17678 74788
rect 0 74704 112 74732
rect 31584 74676 31696 74704
rect 3826 74620 3836 74676
rect 3892 74620 6524 74676
rect 6580 74620 6590 74676
rect 12338 74620 12348 74676
rect 12404 74620 13020 74676
rect 13076 74620 13086 74676
rect 17042 74620 17052 74676
rect 17108 74620 17724 74676
rect 17780 74620 17790 74676
rect 23314 74620 23324 74676
rect 23380 74620 30268 74676
rect 30324 74620 30334 74676
rect 30594 74620 30604 74676
rect 30660 74620 31696 74676
rect 31584 74592 31696 74620
rect 914 74508 924 74564
rect 980 74508 4060 74564
rect 4116 74508 4126 74564
rect 4454 74452 4464 74508
rect 4520 74452 4568 74508
rect 4624 74452 4672 74508
rect 4728 74452 4738 74508
rect 24454 74452 24464 74508
rect 24520 74452 24568 74508
rect 24624 74452 24672 74508
rect 24728 74452 24738 74508
rect 3154 74396 3164 74452
rect 3220 74396 3948 74452
rect 4004 74396 4014 74452
rect 12898 74396 12908 74452
rect 12964 74396 16380 74452
rect 16436 74396 16446 74452
rect 0 74340 112 74368
rect 0 74284 5628 74340
rect 5684 74284 5694 74340
rect 7522 74284 7532 74340
rect 7588 74284 16716 74340
rect 16772 74284 16782 74340
rect 22418 74284 22428 74340
rect 22484 74284 22988 74340
rect 23044 74284 23054 74340
rect 0 74256 112 74284
rect 242 74172 252 74228
rect 308 74172 1036 74228
rect 1092 74172 1102 74228
rect 3490 74172 3500 74228
rect 3556 74172 3836 74228
rect 3892 74172 7420 74228
rect 7476 74172 7486 74228
rect 13682 74172 13692 74228
rect 13748 74172 18396 74228
rect 18452 74172 18462 74228
rect 1334 74060 1372 74116
rect 1428 74060 1438 74116
rect 4274 74060 4284 74116
rect 4340 74060 5068 74116
rect 5124 74060 5134 74116
rect 7970 74060 7980 74116
rect 8036 74060 9884 74116
rect 9940 74060 9950 74116
rect 10658 74060 10668 74116
rect 10724 74060 11452 74116
rect 11508 74060 12236 74116
rect 12292 74060 13468 74116
rect 13524 74060 14476 74116
rect 14532 74060 16604 74116
rect 16660 74060 16670 74116
rect 17042 74060 17052 74116
rect 17108 74060 17388 74116
rect 17444 74060 17454 74116
rect 17714 74060 17724 74116
rect 17780 74060 18620 74116
rect 18676 74060 18686 74116
rect 19730 74060 19740 74116
rect 19796 74060 20188 74116
rect 20244 74060 20254 74116
rect 21074 74060 21084 74116
rect 21140 74060 21420 74116
rect 21476 74060 21486 74116
rect 23426 74060 23436 74116
rect 23492 74060 30268 74116
rect 30324 74060 30334 74116
rect 1250 73948 1260 74004
rect 1316 73948 3612 74004
rect 3668 73948 3678 74004
rect 6850 73948 6860 74004
rect 6916 73948 11788 74004
rect 11844 73948 11854 74004
rect 17574 73948 17612 74004
rect 17668 73948 18172 74004
rect 18228 73948 18238 74004
rect 0 73892 112 73920
rect 0 73836 7084 73892
rect 7140 73836 7150 73892
rect 9538 73836 9548 73892
rect 9604 73836 10668 73892
rect 10724 73836 11340 73892
rect 11396 73836 11406 73892
rect 0 73808 112 73836
rect 7186 73724 7196 73780
rect 7252 73724 7532 73780
rect 7588 73724 7598 73780
rect 3794 73668 3804 73724
rect 3860 73668 3908 73724
rect 3964 73668 4012 73724
rect 4068 73668 4078 73724
rect 23794 73668 23804 73724
rect 23860 73668 23908 73724
rect 23964 73668 24012 73724
rect 24068 73668 24078 73724
rect 7410 73612 7420 73668
rect 7476 73612 10556 73668
rect 10612 73612 10622 73668
rect 31584 73556 31696 73584
rect 2258 73500 2268 73556
rect 2324 73500 2716 73556
rect 2772 73500 2782 73556
rect 9314 73500 9324 73556
rect 9380 73500 10780 73556
rect 10836 73500 10846 73556
rect 18050 73500 18060 73556
rect 18116 73500 18396 73556
rect 18452 73500 18462 73556
rect 30594 73500 30604 73556
rect 30660 73500 31696 73556
rect 31584 73472 31696 73500
rect 0 73444 112 73472
rect 0 73388 6524 73444
rect 6580 73388 6590 73444
rect 8194 73388 8204 73444
rect 8260 73388 10220 73444
rect 10276 73388 10286 73444
rect 12674 73388 12684 73444
rect 12740 73388 12796 73444
rect 12852 73388 12862 73444
rect 20626 73388 20636 73444
rect 20692 73388 20702 73444
rect 0 73360 112 73388
rect 20636 73332 20692 73388
rect 2818 73276 2828 73332
rect 2884 73276 2940 73332
rect 2996 73276 7588 73332
rect 7746 73276 7756 73332
rect 7812 73276 9772 73332
rect 9828 73276 9838 73332
rect 13234 73276 13244 73332
rect 13300 73276 13692 73332
rect 13748 73276 13758 73332
rect 15026 73276 15036 73332
rect 15092 73276 15932 73332
rect 15988 73276 16716 73332
rect 16772 73276 22652 73332
rect 22708 73276 22718 73332
rect 2034 73164 2044 73220
rect 2100 73164 4956 73220
rect 5012 73164 5022 73220
rect 7532 73108 7588 73276
rect 8306 73164 8316 73220
rect 8372 73164 10780 73220
rect 10836 73164 11228 73220
rect 11284 73164 11294 73220
rect 11666 73164 11676 73220
rect 11732 73164 20076 73220
rect 20132 73164 20142 73220
rect 2604 73052 5180 73108
rect 5236 73052 5246 73108
rect 7532 73052 9324 73108
rect 9380 73052 9390 73108
rect 12226 73052 12236 73108
rect 12292 73052 13804 73108
rect 13860 73052 13870 73108
rect 20962 73052 20972 73108
rect 21028 73052 21532 73108
rect 21588 73052 21598 73108
rect 0 72996 112 73024
rect 2604 72996 2660 73052
rect 0 72940 2660 72996
rect 5618 72940 5628 72996
rect 5684 72940 5852 72996
rect 5908 72940 11340 72996
rect 11396 72940 11406 72996
rect 14578 72940 14588 72996
rect 14644 72940 14924 72996
rect 14980 72940 14990 72996
rect 0 72912 112 72940
rect 4454 72884 4464 72940
rect 4520 72884 4568 72940
rect 4624 72884 4672 72940
rect 4728 72884 4738 72940
rect 7196 72884 7252 72940
rect 24454 72884 24464 72940
rect 24520 72884 24568 72940
rect 24624 72884 24672 72940
rect 24728 72884 24738 72940
rect 1782 72828 1820 72884
rect 1876 72828 1886 72884
rect 7186 72828 7196 72884
rect 7252 72828 7262 72884
rect 8866 72828 8876 72884
rect 8932 72828 9212 72884
rect 9268 72828 9278 72884
rect 11106 72828 11116 72884
rect 11172 72828 11676 72884
rect 11732 72828 11742 72884
rect 13570 72828 13580 72884
rect 13636 72828 14980 72884
rect 2034 72716 2044 72772
rect 2100 72716 2492 72772
rect 2548 72716 2558 72772
rect 3042 72716 3052 72772
rect 3108 72716 5292 72772
rect 5348 72716 5358 72772
rect 10322 72716 10332 72772
rect 10388 72716 11452 72772
rect 11508 72716 11518 72772
rect 12786 72716 12796 72772
rect 12852 72716 14252 72772
rect 14308 72716 14318 72772
rect 14924 72660 14980 72828
rect 17350 72716 17388 72772
rect 17444 72716 17454 72772
rect 2258 72604 2268 72660
rect 2324 72604 6300 72660
rect 6356 72604 6366 72660
rect 6626 72604 6636 72660
rect 6692 72604 13804 72660
rect 13860 72604 13870 72660
rect 14914 72604 14924 72660
rect 14980 72604 21308 72660
rect 21364 72604 21374 72660
rect 0 72548 112 72576
rect 0 72492 1596 72548
rect 1652 72492 1662 72548
rect 2594 72492 2604 72548
rect 2660 72492 2828 72548
rect 2884 72492 2894 72548
rect 4386 72492 4396 72548
rect 4452 72492 5068 72548
rect 5124 72492 7756 72548
rect 7812 72492 7822 72548
rect 9426 72492 9436 72548
rect 9492 72492 10332 72548
rect 10388 72492 10398 72548
rect 10770 72492 10780 72548
rect 10836 72492 11228 72548
rect 11284 72492 11788 72548
rect 11844 72492 11854 72548
rect 20066 72492 20076 72548
rect 20132 72492 20860 72548
rect 20916 72492 20926 72548
rect 0 72464 112 72492
rect 31584 72436 31696 72464
rect 1138 72380 1148 72436
rect 1204 72380 1820 72436
rect 1876 72380 1886 72436
rect 2146 72380 2156 72436
rect 2212 72380 8316 72436
rect 8372 72380 8382 72436
rect 9314 72380 9324 72436
rect 9380 72380 9772 72436
rect 9828 72380 10108 72436
rect 10164 72380 10174 72436
rect 11666 72380 11676 72436
rect 11732 72380 16044 72436
rect 16100 72380 16110 72436
rect 30594 72380 30604 72436
rect 30660 72380 31696 72436
rect 31584 72352 31696 72380
rect 6626 72268 6636 72324
rect 6692 72268 7420 72324
rect 7476 72268 7486 72324
rect 8082 72268 8092 72324
rect 8148 72268 9100 72324
rect 9156 72268 9166 72324
rect 10108 72268 13356 72324
rect 13412 72268 13916 72324
rect 13972 72268 13982 72324
rect 10108 72212 10164 72268
rect 10098 72156 10108 72212
rect 10164 72156 10174 72212
rect 15810 72156 15820 72212
rect 15876 72156 17612 72212
rect 17668 72156 17678 72212
rect 0 72100 112 72128
rect 3794 72100 3804 72156
rect 3860 72100 3908 72156
rect 3964 72100 4012 72156
rect 4068 72100 4078 72156
rect 23794 72100 23804 72156
rect 23860 72100 23908 72156
rect 23964 72100 24012 72156
rect 24068 72100 24078 72156
rect 0 72044 924 72100
rect 980 72044 990 72100
rect 0 72016 112 72044
rect 4834 71932 4844 71988
rect 4900 71932 14476 71988
rect 14532 71932 14542 71988
rect 19282 71932 19292 71988
rect 19348 71932 19964 71988
rect 20020 71932 20030 71988
rect 2034 71820 2044 71876
rect 2100 71820 5180 71876
rect 5236 71820 5852 71876
rect 5908 71820 5918 71876
rect 6038 71820 6076 71876
rect 6132 71820 6142 71876
rect 8978 71820 8988 71876
rect 9044 71820 11340 71876
rect 11396 71820 11406 71876
rect 19618 71820 19628 71876
rect 19684 71820 22988 71876
rect 23044 71820 23054 71876
rect 4274 71708 4284 71764
rect 4340 71708 6412 71764
rect 6468 71708 6478 71764
rect 16818 71708 16828 71764
rect 16884 71708 18284 71764
rect 18340 71708 21084 71764
rect 21140 71708 21150 71764
rect 0 71652 112 71680
rect 0 71596 6300 71652
rect 6356 71596 6366 71652
rect 10854 71596 10892 71652
rect 10948 71596 10958 71652
rect 15250 71596 15260 71652
rect 15316 71596 15708 71652
rect 15764 71596 15774 71652
rect 20850 71596 20860 71652
rect 20916 71596 21196 71652
rect 21252 71596 21420 71652
rect 21476 71596 21486 71652
rect 0 71568 112 71596
rect 1250 71484 1260 71540
rect 1316 71484 2156 71540
rect 2212 71484 2222 71540
rect 7746 71484 7756 71540
rect 7812 71484 8092 71540
rect 8148 71484 8158 71540
rect 14242 71484 14252 71540
rect 14308 71484 15596 71540
rect 15652 71484 15662 71540
rect 6290 71372 6300 71428
rect 6356 71372 8876 71428
rect 8932 71372 8942 71428
rect 16930 71372 16940 71428
rect 16996 71372 21196 71428
rect 21252 71372 21262 71428
rect 4454 71316 4464 71372
rect 4520 71316 4568 71372
rect 4624 71316 4672 71372
rect 4728 71316 4738 71372
rect 24454 71316 24464 71372
rect 24520 71316 24568 71372
rect 24624 71316 24672 71372
rect 24728 71316 24738 71372
rect 31584 71316 31696 71344
rect 5282 71260 5292 71316
rect 5348 71260 15708 71316
rect 15764 71260 15774 71316
rect 30594 71260 30604 71316
rect 30660 71260 31696 71316
rect 31584 71232 31696 71260
rect 0 71204 112 71232
rect 0 71148 5628 71204
rect 5684 71148 5694 71204
rect 0 71120 112 71148
rect 1474 71036 1484 71092
rect 1540 71036 7756 71092
rect 7812 71036 7822 71092
rect 10994 71036 11004 71092
rect 11060 71036 14812 71092
rect 14868 71036 14878 71092
rect 2258 70924 2268 70980
rect 2324 70924 2940 70980
rect 2996 70924 3006 70980
rect 3462 70924 3500 70980
rect 3556 70924 3566 70980
rect 4498 70924 4508 70980
rect 4564 70924 4956 70980
rect 5012 70924 5022 70980
rect 15092 70924 29484 70980
rect 29540 70924 29550 70980
rect 15092 70868 15148 70924
rect 812 70812 1932 70868
rect 1988 70812 1998 70868
rect 2594 70812 2604 70868
rect 2660 70812 2828 70868
rect 2884 70812 5852 70868
rect 5908 70812 5918 70868
rect 6850 70812 6860 70868
rect 6916 70812 15148 70868
rect 0 70756 112 70784
rect 812 70756 868 70812
rect 0 70700 868 70756
rect 1362 70700 1372 70756
rect 1428 70700 3276 70756
rect 3332 70700 3342 70756
rect 5058 70700 5068 70756
rect 5124 70700 6972 70756
rect 7028 70700 7038 70756
rect 9762 70700 9772 70756
rect 9828 70700 10444 70756
rect 10500 70700 10510 70756
rect 0 70672 112 70700
rect 1250 70588 1260 70644
rect 1316 70588 1484 70644
rect 1540 70588 1820 70644
rect 1876 70588 1886 70644
rect 2482 70588 2492 70644
rect 2548 70588 3500 70644
rect 3556 70588 3566 70644
rect 5282 70588 5292 70644
rect 5348 70588 8876 70644
rect 8932 70588 8942 70644
rect 12450 70588 12460 70644
rect 12516 70588 13020 70644
rect 13076 70588 13086 70644
rect 3794 70532 3804 70588
rect 3860 70532 3908 70588
rect 3964 70532 4012 70588
rect 4068 70532 4078 70588
rect 23794 70532 23804 70588
rect 23860 70532 23908 70588
rect 23964 70532 24012 70588
rect 24068 70532 24078 70588
rect 914 70476 924 70532
rect 980 70476 2044 70532
rect 2100 70476 2110 70532
rect 4274 70476 4284 70532
rect 4340 70476 9100 70532
rect 9156 70476 9166 70532
rect 14354 70476 14364 70532
rect 14420 70476 15372 70532
rect 15428 70476 16828 70532
rect 16884 70476 16894 70532
rect 18946 70476 18956 70532
rect 19012 70476 19852 70532
rect 19908 70476 19918 70532
rect 1250 70364 1260 70420
rect 1316 70364 1820 70420
rect 1876 70364 1886 70420
rect 0 70308 112 70336
rect 0 70252 5404 70308
rect 5460 70252 5470 70308
rect 0 70224 112 70252
rect 31584 70196 31696 70224
rect 1698 70140 1708 70196
rect 1764 70140 2044 70196
rect 2100 70140 2110 70196
rect 17714 70140 17724 70196
rect 17780 70140 19180 70196
rect 19236 70140 19246 70196
rect 20178 70140 20188 70196
rect 20244 70140 20692 70196
rect 30594 70140 30604 70196
rect 30660 70140 31696 70196
rect 20636 70084 20692 70140
rect 31584 70112 31696 70140
rect 2930 70028 2940 70084
rect 2996 70028 8092 70084
rect 8148 70028 8158 70084
rect 17266 70028 17276 70084
rect 17332 70028 18172 70084
rect 18228 70028 18238 70084
rect 20626 70028 20636 70084
rect 20692 70028 20702 70084
rect 2482 69916 2492 69972
rect 2548 69916 2828 69972
rect 2884 69916 2894 69972
rect 3332 69916 7868 69972
rect 7924 69916 7934 69972
rect 9762 69916 9772 69972
rect 9828 69916 9996 69972
rect 10052 69916 10062 69972
rect 20066 69916 20076 69972
rect 20132 69916 21644 69972
rect 21700 69916 21710 69972
rect 0 69860 112 69888
rect 3332 69860 3388 69916
rect 0 69804 3388 69860
rect 18722 69804 18732 69860
rect 18788 69804 21756 69860
rect 21812 69804 22428 69860
rect 22484 69804 22494 69860
rect 0 69776 112 69804
rect 4454 69748 4464 69804
rect 4520 69748 4568 69804
rect 4624 69748 4672 69804
rect 4728 69748 4738 69804
rect 24454 69748 24464 69804
rect 24520 69748 24568 69804
rect 24624 69748 24672 69804
rect 24728 69748 24738 69804
rect 1698 69580 1708 69636
rect 1764 69580 6748 69636
rect 6804 69580 6814 69636
rect 8194 69580 8204 69636
rect 8260 69580 11900 69636
rect 11956 69580 11966 69636
rect 9986 69468 9996 69524
rect 10052 69468 17276 69524
rect 17332 69468 18844 69524
rect 18900 69468 19516 69524
rect 19572 69468 19582 69524
rect 0 69412 112 69440
rect 0 69356 140 69412
rect 196 69356 206 69412
rect 1362 69356 1372 69412
rect 1428 69356 3276 69412
rect 3332 69356 3342 69412
rect 12226 69356 12236 69412
rect 12292 69356 13132 69412
rect 13188 69356 13198 69412
rect 14466 69356 14476 69412
rect 14532 69356 16940 69412
rect 16996 69356 21084 69412
rect 21140 69356 22876 69412
rect 22932 69356 22942 69412
rect 0 69328 112 69356
rect 1250 69244 1260 69300
rect 1316 69244 2940 69300
rect 2996 69244 3388 69300
rect 3444 69244 3454 69300
rect 3612 69244 8876 69300
rect 8932 69244 8942 69300
rect 0 68964 112 68992
rect 3612 68964 3668 69244
rect 3826 69132 3836 69188
rect 3892 69132 5740 69188
rect 5796 69132 5806 69188
rect 6626 69132 6636 69188
rect 6692 69132 7308 69188
rect 7364 69132 7374 69188
rect 19282 69132 19292 69188
rect 19348 69132 24276 69188
rect 5740 69076 5796 69132
rect 5740 69020 10556 69076
rect 10612 69020 11340 69076
rect 11396 69020 14476 69076
rect 14532 69020 14542 69076
rect 3794 68964 3804 69020
rect 3860 68964 3908 69020
rect 3964 68964 4012 69020
rect 4068 68964 4078 69020
rect 23794 68964 23804 69020
rect 23860 68964 23908 69020
rect 23964 68964 24012 69020
rect 24068 68964 24078 69020
rect 24220 68964 24276 69132
rect 31584 69076 31696 69104
rect 30594 69020 30604 69076
rect 30660 69020 31696 69076
rect 31584 68992 31696 69020
rect 0 68908 3668 68964
rect 5170 68908 5180 68964
rect 5236 68908 6580 68964
rect 7074 68908 7084 68964
rect 7140 68908 9996 68964
rect 10052 68908 10062 68964
rect 17266 68908 17276 68964
rect 17332 68908 18284 68964
rect 18340 68908 18956 68964
rect 19012 68908 19022 68964
rect 21074 68908 21084 68964
rect 21140 68908 21308 68964
rect 21364 68908 21374 68964
rect 24210 68908 24220 68964
rect 24276 68908 24286 68964
rect 0 68880 112 68908
rect 6524 68852 6580 68908
rect 4162 68796 4172 68852
rect 4228 68796 5964 68852
rect 6020 68796 6030 68852
rect 6514 68796 6524 68852
rect 6580 68796 7308 68852
rect 7364 68796 7374 68852
rect 7746 68796 7756 68852
rect 7812 68796 13356 68852
rect 13412 68796 14588 68852
rect 14644 68796 14654 68852
rect 17602 68796 17612 68852
rect 17668 68796 18172 68852
rect 18228 68796 18238 68852
rect 20962 68796 20972 68852
rect 21028 68796 21756 68852
rect 21812 68796 24332 68852
rect 24388 68796 24398 68852
rect 1362 68684 1372 68740
rect 1428 68684 3220 68740
rect 5618 68684 5628 68740
rect 5684 68684 12348 68740
rect 12404 68684 14140 68740
rect 14196 68684 14206 68740
rect 19954 68684 19964 68740
rect 20020 68684 23100 68740
rect 23156 68684 23166 68740
rect 3164 68628 3220 68684
rect 998 68572 1036 68628
rect 1092 68572 1102 68628
rect 1922 68572 1932 68628
rect 1988 68572 2940 68628
rect 2996 68572 3006 68628
rect 3164 68572 11788 68628
rect 11844 68572 11854 68628
rect 12786 68572 12796 68628
rect 12852 68572 15260 68628
rect 15316 68572 15326 68628
rect 20066 68572 20076 68628
rect 20132 68572 24668 68628
rect 24724 68572 24734 68628
rect 0 68516 112 68544
rect 0 68460 4844 68516
rect 4900 68460 4910 68516
rect 7718 68460 7756 68516
rect 7812 68460 7822 68516
rect 9314 68460 9324 68516
rect 9380 68460 11228 68516
rect 11284 68460 11294 68516
rect 14802 68460 14812 68516
rect 14868 68460 16268 68516
rect 16324 68460 16334 68516
rect 19058 68460 19068 68516
rect 19124 68460 23212 68516
rect 23268 68460 23436 68516
rect 23492 68460 23502 68516
rect 0 68432 112 68460
rect 354 68348 364 68404
rect 420 68348 1036 68404
rect 1092 68348 1102 68404
rect 3332 68348 7980 68404
rect 8036 68348 8046 68404
rect 8194 68348 8204 68404
rect 8260 68348 9436 68404
rect 9492 68348 9502 68404
rect 12898 68348 12908 68404
rect 12964 68348 13580 68404
rect 13636 68348 13646 68404
rect 20626 68348 20636 68404
rect 20692 68348 21420 68404
rect 21476 68348 21486 68404
rect 22642 68348 22652 68404
rect 22708 68348 24444 68404
rect 24500 68348 24510 68404
rect 28690 68348 28700 68404
rect 28756 68348 29484 68404
rect 29540 68348 29550 68404
rect 0 68068 112 68096
rect 0 68012 140 68068
rect 196 68012 206 68068
rect 1362 68012 1372 68068
rect 1428 68012 1820 68068
rect 1876 68012 1886 68068
rect 0 67984 112 68012
rect 466 67900 476 67956
rect 532 67900 1036 67956
rect 1092 67900 1102 67956
rect 130 67788 140 67844
rect 196 67788 1036 67844
rect 1092 67788 1102 67844
rect 3332 67732 3388 68348
rect 18386 68236 18396 68292
rect 18452 68236 20188 68292
rect 20244 68236 20972 68292
rect 21028 68236 22428 68292
rect 22484 68236 22494 68292
rect 4454 68180 4464 68236
rect 4520 68180 4568 68236
rect 4624 68180 4672 68236
rect 4728 68180 4738 68236
rect 24454 68180 24464 68236
rect 24520 68180 24568 68236
rect 24624 68180 24672 68236
rect 24728 68180 24738 68236
rect 6178 68124 6188 68180
rect 6244 68124 18844 68180
rect 18900 68124 18910 68180
rect 8082 68012 8092 68068
rect 8148 68012 12012 68068
rect 12068 68012 12348 68068
rect 12404 68012 15148 68068
rect 16818 68012 16828 68068
rect 16884 68012 18060 68068
rect 18116 68012 19180 68068
rect 19236 68012 19246 68068
rect 20738 68012 20748 68068
rect 20804 68012 21868 68068
rect 21924 68012 21934 68068
rect 15092 67956 15148 68012
rect 31584 67956 31696 67984
rect 4918 67900 4956 67956
rect 5012 67900 5022 67956
rect 12114 67900 12124 67956
rect 12180 67900 12796 67956
rect 12852 67900 12862 67956
rect 15092 67900 15260 67956
rect 15316 67900 15326 67956
rect 16146 67900 16156 67956
rect 16212 67900 17836 67956
rect 17892 67900 17902 67956
rect 20402 67900 20412 67956
rect 20468 67900 20636 67956
rect 20692 67900 21308 67956
rect 21364 67900 21374 67956
rect 30594 67900 30604 67956
rect 30660 67900 31696 67956
rect 31584 67872 31696 67900
rect 4498 67788 4508 67844
rect 4564 67788 5292 67844
rect 5348 67788 5358 67844
rect 11218 67788 11228 67844
rect 11284 67788 14140 67844
rect 14196 67788 14206 67844
rect 19394 67788 19404 67844
rect 19460 67788 20748 67844
rect 20804 67788 20814 67844
rect 14140 67732 14196 67788
rect 1708 67676 3388 67732
rect 3490 67676 3500 67732
rect 3556 67676 3948 67732
rect 4004 67676 4014 67732
rect 12898 67676 12908 67732
rect 12964 67676 13244 67732
rect 13300 67676 13310 67732
rect 14140 67676 16156 67732
rect 16212 67676 16716 67732
rect 16772 67676 18844 67732
rect 18900 67676 22876 67732
rect 22932 67676 22942 67732
rect 0 67620 112 67648
rect 1708 67620 1764 67676
rect 0 67564 1764 67620
rect 2146 67564 2156 67620
rect 2212 67564 6076 67620
rect 6132 67564 6142 67620
rect 9314 67564 9324 67620
rect 9380 67564 14924 67620
rect 14980 67564 15148 67620
rect 20738 67564 20748 67620
rect 20804 67564 21196 67620
rect 21252 67564 21262 67620
rect 0 67536 112 67564
rect 15092 67508 15148 67564
rect 9426 67452 9436 67508
rect 9492 67452 10220 67508
rect 10276 67452 10286 67508
rect 15092 67452 17612 67508
rect 17668 67452 17678 67508
rect 17836 67452 18172 67508
rect 18228 67452 19964 67508
rect 20020 67452 21868 67508
rect 21924 67452 23660 67508
rect 23716 67452 23726 67508
rect 3794 67396 3804 67452
rect 3860 67396 3908 67452
rect 3964 67396 4012 67452
rect 4068 67396 4078 67452
rect 17836 67396 17892 67452
rect 23794 67396 23804 67452
rect 23860 67396 23908 67452
rect 23964 67396 24012 67452
rect 24068 67396 24078 67452
rect 4162 67340 4172 67396
rect 4228 67340 7644 67396
rect 7700 67340 7710 67396
rect 14130 67340 14140 67396
rect 14196 67340 16044 67396
rect 16100 67340 16110 67396
rect 16940 67340 17892 67396
rect 19730 67340 19740 67396
rect 19796 67340 22652 67396
rect 22708 67340 22718 67396
rect 16940 67284 16996 67340
rect 1138 67228 1148 67284
rect 1204 67228 1820 67284
rect 1876 67228 1886 67284
rect 3378 67228 3388 67284
rect 3444 67228 3482 67284
rect 5404 67228 7084 67284
rect 7140 67228 7150 67284
rect 10658 67228 10668 67284
rect 10724 67228 11116 67284
rect 11172 67228 11182 67284
rect 15250 67228 15260 67284
rect 15316 67228 16996 67284
rect 19618 67228 19628 67284
rect 19684 67228 21196 67284
rect 21252 67228 23436 67284
rect 23492 67228 23502 67284
rect 0 67172 112 67200
rect 3388 67172 3444 67228
rect 5404 67172 5460 67228
rect 0 67116 588 67172
rect 644 67116 654 67172
rect 2380 67116 3444 67172
rect 3500 67116 5460 67172
rect 6514 67116 6524 67172
rect 6580 67116 6972 67172
rect 7028 67116 7038 67172
rect 8642 67116 8652 67172
rect 8708 67116 9996 67172
rect 10052 67116 14700 67172
rect 14756 67116 15932 67172
rect 15988 67116 15998 67172
rect 0 67088 112 67116
rect 2380 67060 2436 67116
rect 3500 67060 3556 67116
rect 2370 67004 2380 67060
rect 2436 67004 2446 67060
rect 2604 67004 3556 67060
rect 6626 67004 6636 67060
rect 6692 67004 7308 67060
rect 7364 67004 7374 67060
rect 8978 67004 8988 67060
rect 9044 67004 9548 67060
rect 9604 67004 9614 67060
rect 9874 67004 9884 67060
rect 9940 67004 14924 67060
rect 14980 67004 15484 67060
rect 15540 67004 15550 67060
rect 2604 66948 2660 67004
rect 16940 66948 16996 67228
rect 17154 67172 17164 67228
rect 17220 67172 17230 67228
rect 17164 67060 17220 67172
rect 18274 67116 18284 67172
rect 18340 67116 19292 67172
rect 19348 67116 19358 67172
rect 20738 67116 20748 67172
rect 20804 67116 21084 67172
rect 21140 67116 21150 67172
rect 17164 67004 18172 67060
rect 18228 67004 18844 67060
rect 18900 67004 20412 67060
rect 20468 67004 20478 67060
rect 914 66892 924 66948
rect 980 66892 1484 66948
rect 1540 66892 1550 66948
rect 2482 66892 2492 66948
rect 2548 66892 2660 66948
rect 3042 66892 3052 66948
rect 3108 66892 10892 66948
rect 10948 66892 10958 66948
rect 16940 66892 17164 66948
rect 17220 66892 17230 66948
rect 31584 66836 31696 66864
rect 578 66780 588 66836
rect 644 66780 1148 66836
rect 1204 66780 1214 66836
rect 4274 66780 4284 66836
rect 4340 66780 5404 66836
rect 5460 66780 5470 66836
rect 6962 66780 6972 66836
rect 7028 66780 9660 66836
rect 9716 66780 9726 66836
rect 13794 66780 13804 66836
rect 13860 66780 15148 66836
rect 15204 66780 15214 66836
rect 30594 66780 30604 66836
rect 30660 66780 31696 66836
rect 31584 66752 31696 66780
rect 0 66724 112 66752
rect 0 66668 252 66724
rect 308 66668 318 66724
rect 812 66668 2044 66724
rect 2100 66668 2110 66724
rect 7298 66668 7308 66724
rect 7364 66668 16268 66724
rect 16324 66668 17388 66724
rect 17444 66668 17454 66724
rect 0 66640 112 66668
rect 0 66276 112 66304
rect 812 66276 868 66668
rect 4454 66612 4464 66668
rect 4520 66612 4568 66668
rect 4624 66612 4672 66668
rect 4728 66612 4738 66668
rect 24454 66612 24464 66668
rect 24520 66612 24568 66668
rect 24624 66612 24672 66668
rect 24728 66612 24738 66668
rect 2146 66556 2156 66612
rect 2212 66556 3052 66612
rect 3108 66556 3118 66612
rect 5954 66556 5964 66612
rect 6020 66556 15036 66612
rect 15092 66556 15102 66612
rect 5964 66500 6020 66556
rect 1586 66444 1596 66500
rect 1652 66444 6020 66500
rect 18498 66444 18508 66500
rect 18564 66444 18956 66500
rect 19012 66444 19964 66500
rect 20020 66444 20748 66500
rect 20804 66444 20814 66500
rect 20962 66444 20972 66500
rect 21028 66444 30268 66500
rect 30324 66444 30334 66500
rect 1250 66332 1260 66388
rect 1316 66332 1820 66388
rect 1876 66332 2716 66388
rect 2772 66332 2782 66388
rect 3602 66332 3612 66388
rect 3668 66332 5964 66388
rect 6020 66332 6030 66388
rect 0 66220 868 66276
rect 2146 66220 2156 66276
rect 2212 66220 3948 66276
rect 4004 66220 4014 66276
rect 5142 66220 5180 66276
rect 5236 66220 5246 66276
rect 5842 66220 5852 66276
rect 5908 66220 6412 66276
rect 6468 66220 6478 66276
rect 17826 66220 17836 66276
rect 17892 66220 18508 66276
rect 18564 66220 18574 66276
rect 0 66192 112 66220
rect 3378 66108 3388 66164
rect 3444 66108 13916 66164
rect 13972 66108 13982 66164
rect 242 65996 252 66052
rect 308 65996 9100 66052
rect 9156 65996 9166 66052
rect 18498 65996 18508 66052
rect 18564 65996 18732 66052
rect 18788 65996 19068 66052
rect 19124 65996 19134 66052
rect 6066 65884 6076 65940
rect 6132 65884 6300 65940
rect 6356 65884 6366 65940
rect 0 65828 112 65856
rect 3794 65828 3804 65884
rect 3860 65828 3908 65884
rect 3964 65828 4012 65884
rect 4068 65828 4078 65884
rect 23794 65828 23804 65884
rect 23860 65828 23908 65884
rect 23964 65828 24012 65884
rect 24068 65828 24078 65884
rect 0 65772 700 65828
rect 756 65772 766 65828
rect 13570 65772 13580 65828
rect 13636 65772 13916 65828
rect 13972 65772 13982 65828
rect 0 65744 112 65772
rect 31584 65716 31696 65744
rect 1250 65660 1260 65716
rect 1316 65660 13468 65716
rect 13524 65660 13534 65716
rect 16146 65660 16156 65716
rect 16212 65660 16268 65716
rect 16324 65660 16334 65716
rect 30594 65660 30604 65716
rect 30660 65660 31696 65716
rect 31584 65632 31696 65660
rect 1922 65548 1932 65604
rect 1988 65548 5852 65604
rect 5908 65548 6524 65604
rect 6580 65548 8876 65604
rect 8932 65548 8942 65604
rect 13010 65548 13020 65604
rect 13076 65548 14252 65604
rect 14308 65548 15820 65604
rect 15876 65548 16940 65604
rect 16996 65548 18172 65604
rect 18228 65548 18238 65604
rect 4386 65436 4396 65492
rect 4452 65436 8204 65492
rect 8260 65436 8270 65492
rect 8530 65436 8540 65492
rect 8596 65436 9324 65492
rect 9380 65436 9390 65492
rect 0 65380 112 65408
rect 0 65324 3500 65380
rect 3556 65324 3566 65380
rect 0 65296 112 65324
rect 6290 65100 6300 65156
rect 6356 65100 13692 65156
rect 13748 65100 18732 65156
rect 18788 65100 21308 65156
rect 21364 65100 21374 65156
rect 4454 65044 4464 65100
rect 4520 65044 4568 65100
rect 4624 65044 4672 65100
rect 4728 65044 4738 65100
rect 24454 65044 24464 65100
rect 24520 65044 24568 65100
rect 24624 65044 24672 65100
rect 24728 65044 24738 65100
rect 2482 64988 2492 65044
rect 2548 64988 2828 65044
rect 2884 64988 2894 65044
rect 9202 64988 9212 65044
rect 9268 64988 9996 65044
rect 10052 64988 10062 65044
rect 0 64932 112 64960
rect 0 64876 4956 64932
rect 5012 64876 5022 64932
rect 0 64848 112 64876
rect 3602 64764 3612 64820
rect 3668 64764 5180 64820
rect 5236 64764 5246 64820
rect 8306 64764 8316 64820
rect 8372 64764 9996 64820
rect 10052 64764 10062 64820
rect 19058 64764 19068 64820
rect 19124 64764 30380 64820
rect 30436 64764 30446 64820
rect 4274 64652 4284 64708
rect 4340 64652 5740 64708
rect 5796 64652 5806 64708
rect 8194 64652 8204 64708
rect 8260 64652 9324 64708
rect 9380 64652 9390 64708
rect 31584 64596 31696 64624
rect 1586 64540 1596 64596
rect 1652 64540 4956 64596
rect 5012 64540 5022 64596
rect 7522 64540 7532 64596
rect 7588 64540 11004 64596
rect 11060 64540 11070 64596
rect 30594 64540 30604 64596
rect 30660 64540 31696 64596
rect 31584 64512 31696 64540
rect 0 64484 112 64512
rect 0 64428 3948 64484
rect 4004 64428 4014 64484
rect 0 64400 112 64428
rect 5058 64316 5068 64372
rect 5124 64316 13580 64372
rect 13636 64316 13646 64372
rect 3794 64260 3804 64316
rect 3860 64260 3908 64316
rect 3964 64260 4012 64316
rect 4068 64260 4078 64316
rect 23794 64260 23804 64316
rect 23860 64260 23908 64316
rect 23964 64260 24012 64316
rect 24068 64260 24078 64316
rect 1250 64092 1260 64148
rect 1316 64092 8036 64148
rect 8194 64092 8204 64148
rect 8260 64092 10444 64148
rect 10500 64092 10510 64148
rect 0 64036 112 64064
rect 7980 64036 8036 64092
rect 0 63980 812 64036
rect 868 63980 878 64036
rect 1698 63980 1708 64036
rect 1764 63980 4172 64036
rect 4228 63980 4238 64036
rect 7980 63980 8764 64036
rect 8820 63980 8830 64036
rect 10770 63980 10780 64036
rect 10836 63980 12572 64036
rect 12628 63980 12638 64036
rect 13122 63980 13132 64036
rect 13188 63980 14252 64036
rect 14308 63980 19628 64036
rect 19684 63980 20972 64036
rect 21028 63980 21038 64036
rect 0 63952 112 63980
rect 2818 63868 2828 63924
rect 2884 63868 3500 63924
rect 3556 63868 3566 63924
rect 9538 63868 9548 63924
rect 9604 63868 10332 63924
rect 10388 63868 10398 63924
rect 11778 63868 11788 63924
rect 11844 63868 17388 63924
rect 17444 63868 17454 63924
rect 25106 63868 25116 63924
rect 25172 63868 30492 63924
rect 30548 63868 30558 63924
rect 2370 63756 2380 63812
rect 2436 63756 2492 63812
rect 2548 63756 2558 63812
rect 7634 63756 7644 63812
rect 7700 63756 7980 63812
rect 8036 63756 8046 63812
rect 8418 63756 8428 63812
rect 8484 63756 9324 63812
rect 9380 63756 9884 63812
rect 9940 63756 9950 63812
rect 15092 63756 15484 63812
rect 15540 63756 15550 63812
rect 16818 63756 16828 63812
rect 16884 63756 18732 63812
rect 18788 63756 18798 63812
rect 20738 63756 20748 63812
rect 20804 63756 20972 63812
rect 21028 63756 21038 63812
rect 15092 63700 15148 63756
rect 3332 63644 5628 63700
rect 5684 63644 5694 63700
rect 6290 63644 6300 63700
rect 6356 63644 10892 63700
rect 10948 63644 15148 63700
rect 17714 63644 17724 63700
rect 17780 63644 19180 63700
rect 19236 63644 19246 63700
rect 0 63588 112 63616
rect 3332 63588 3388 63644
rect 0 63532 3388 63588
rect 17378 63532 17388 63588
rect 17444 63532 20076 63588
rect 20132 63532 20142 63588
rect 0 63504 112 63532
rect 4454 63476 4464 63532
rect 4520 63476 4568 63532
rect 4624 63476 4672 63532
rect 4728 63476 4738 63532
rect 24454 63476 24464 63532
rect 24520 63476 24568 63532
rect 24624 63476 24672 63532
rect 24728 63476 24738 63532
rect 31584 63476 31696 63504
rect 9874 63420 9884 63476
rect 9940 63420 21308 63476
rect 21364 63420 21374 63476
rect 30594 63420 30604 63476
rect 30660 63420 31696 63476
rect 31584 63392 31696 63420
rect 1362 63308 1372 63364
rect 1428 63308 2940 63364
rect 2996 63308 3006 63364
rect 5282 63308 5292 63364
rect 5348 63308 7980 63364
rect 8036 63308 8046 63364
rect 11732 63308 11900 63364
rect 11956 63308 12908 63364
rect 12964 63308 12974 63364
rect 13458 63308 13468 63364
rect 13524 63308 14476 63364
rect 14532 63308 17500 63364
rect 17556 63308 18396 63364
rect 18452 63308 18462 63364
rect 11732 63252 11788 63308
rect 5170 63196 5180 63252
rect 5236 63196 5628 63252
rect 5684 63196 11788 63252
rect 12908 63252 12964 63308
rect 12908 63196 15148 63252
rect 0 63140 112 63168
rect 0 63084 140 63140
rect 196 63084 206 63140
rect 1810 63084 1820 63140
rect 1876 63084 2940 63140
rect 2996 63084 3164 63140
rect 3220 63084 5740 63140
rect 5796 63084 6524 63140
rect 6580 63084 6590 63140
rect 7970 63084 7980 63140
rect 8036 63084 13916 63140
rect 13972 63084 13982 63140
rect 0 63056 112 63084
rect 15092 63028 15148 63196
rect 15250 63084 15260 63140
rect 15316 63084 15932 63140
rect 15988 63084 15998 63140
rect 16818 63084 16828 63140
rect 16884 63084 17500 63140
rect 17556 63084 17566 63140
rect 21410 63084 21420 63140
rect 21476 63084 22092 63140
rect 22148 63084 22158 63140
rect 28802 63084 28812 63140
rect 28868 63084 29484 63140
rect 29540 63084 29550 63140
rect 15092 62972 15708 63028
rect 15764 62972 15774 63028
rect 3378 62860 3388 62916
rect 3444 62860 4172 62916
rect 4228 62860 4238 62916
rect 6514 62860 6524 62916
rect 6580 62860 7420 62916
rect 7476 62860 7486 62916
rect 10434 62860 10444 62916
rect 10500 62860 11900 62916
rect 11956 62860 11966 62916
rect 12562 62860 12572 62916
rect 12628 62860 12908 62916
rect 12964 62860 12974 62916
rect 19618 62860 19628 62916
rect 19684 62860 19852 62916
rect 19908 62860 19918 62916
rect 9660 62748 13468 62804
rect 13524 62748 13534 62804
rect 0 62692 112 62720
rect 3794 62692 3804 62748
rect 3860 62692 3908 62748
rect 3964 62692 4012 62748
rect 4068 62692 4078 62748
rect 9660 62692 9716 62748
rect 23794 62692 23804 62748
rect 23860 62692 23908 62748
rect 23964 62692 24012 62748
rect 24068 62692 24078 62748
rect 0 62636 364 62692
rect 420 62636 430 62692
rect 4162 62636 4172 62692
rect 4228 62636 9716 62692
rect 9874 62636 9884 62692
rect 9940 62636 16268 62692
rect 16324 62636 16828 62692
rect 16884 62636 16894 62692
rect 19954 62636 19964 62692
rect 20020 62636 21420 62692
rect 21476 62636 21486 62692
rect 0 62608 112 62636
rect 2482 62524 2492 62580
rect 2548 62524 9996 62580
rect 10052 62524 10062 62580
rect 21074 62524 21084 62580
rect 21140 62524 21756 62580
rect 21812 62524 21822 62580
rect 3266 62412 3276 62468
rect 3332 62412 4956 62468
rect 5012 62412 5022 62468
rect 6066 62412 6076 62468
rect 6132 62412 6468 62468
rect 10882 62412 10892 62468
rect 10948 62412 11676 62468
rect 11732 62412 11742 62468
rect 14242 62412 14252 62468
rect 14308 62412 15148 62468
rect 15204 62412 15214 62468
rect 21186 62412 21196 62468
rect 21252 62412 21644 62468
rect 21700 62412 21710 62468
rect 6412 62356 6468 62412
rect 31584 62356 31696 62384
rect 2034 62300 2044 62356
rect 2100 62300 2716 62356
rect 2772 62300 2782 62356
rect 4172 62300 5964 62356
rect 6020 62300 6030 62356
rect 6402 62300 6412 62356
rect 6468 62300 15092 62356
rect 17266 62300 17276 62356
rect 17332 62300 23772 62356
rect 23828 62300 25004 62356
rect 25060 62300 25070 62356
rect 30594 62300 30604 62356
rect 30660 62300 31696 62356
rect 0 62244 112 62272
rect 0 62188 476 62244
rect 532 62188 542 62244
rect 1260 62188 1932 62244
rect 1988 62188 1998 62244
rect 0 62160 112 62188
rect 1260 62132 1316 62188
rect 1138 62076 1148 62132
rect 1204 62076 1316 62132
rect 4172 62132 4228 62300
rect 15036 62244 15092 62300
rect 31584 62272 31696 62300
rect 5282 62188 5292 62244
rect 5348 62188 6636 62244
rect 6692 62188 6702 62244
rect 15026 62188 15036 62244
rect 15092 62188 18956 62244
rect 19012 62188 20188 62244
rect 20244 62188 20254 62244
rect 21634 62188 21644 62244
rect 21700 62188 21756 62244
rect 21812 62188 21822 62244
rect 4172 62076 4284 62132
rect 4340 62076 4350 62132
rect 15250 62076 15260 62132
rect 15316 62076 16156 62132
rect 16212 62076 16222 62132
rect 16930 62076 16940 62132
rect 16996 62076 19068 62132
rect 19124 62076 19134 62132
rect 21158 62076 21196 62132
rect 21252 62076 21262 62132
rect 578 61964 588 62020
rect 644 61964 4340 62020
rect 5058 61964 5068 62020
rect 5124 61964 5628 62020
rect 5684 61964 5694 62020
rect 20626 61964 20636 62020
rect 20692 61964 21644 62020
rect 21700 61964 21710 62020
rect 1820 61852 3612 61908
rect 3668 61852 3678 61908
rect 0 61796 112 61824
rect 1820 61796 1876 61852
rect 4284 61796 4340 61964
rect 4454 61908 4464 61964
rect 4520 61908 4568 61964
rect 4624 61908 4672 61964
rect 4728 61908 4738 61964
rect 24454 61908 24464 61964
rect 24520 61908 24568 61964
rect 24624 61908 24672 61964
rect 24728 61908 24738 61964
rect 9986 61852 9996 61908
rect 10052 61852 11004 61908
rect 11060 61852 17276 61908
rect 17332 61852 17342 61908
rect 17714 61852 17724 61908
rect 17780 61852 17948 61908
rect 18004 61852 18014 61908
rect 0 61740 1876 61796
rect 2034 61740 2044 61796
rect 2100 61740 2156 61796
rect 2212 61740 2222 61796
rect 4284 61740 6076 61796
rect 6132 61740 6142 61796
rect 8978 61740 8988 61796
rect 9044 61740 9436 61796
rect 9492 61740 9502 61796
rect 15922 61740 15932 61796
rect 15988 61740 17612 61796
rect 17668 61740 17678 61796
rect 19058 61740 19068 61796
rect 19124 61740 20636 61796
rect 20692 61740 20702 61796
rect 0 61712 112 61740
rect 1362 61628 1372 61684
rect 1428 61628 1820 61684
rect 1876 61628 1886 61684
rect 3490 61628 3500 61684
rect 3556 61628 12348 61684
rect 12404 61628 12414 61684
rect 17154 61628 17164 61684
rect 17220 61628 18172 61684
rect 18228 61628 20524 61684
rect 20580 61628 20590 61684
rect 4610 61516 4620 61572
rect 4676 61516 5404 61572
rect 5460 61516 5470 61572
rect 6962 61516 6972 61572
rect 7028 61516 10948 61572
rect 11106 61516 11116 61572
rect 11172 61516 13020 61572
rect 13076 61516 13086 61572
rect 15586 61516 15596 61572
rect 15652 61516 15820 61572
rect 15876 61516 17052 61572
rect 17108 61516 17118 61572
rect 10892 61460 10948 61516
rect 1474 61404 1484 61460
rect 1540 61404 9212 61460
rect 9268 61404 9278 61460
rect 10892 61404 15036 61460
rect 15092 61404 18732 61460
rect 18788 61404 18798 61460
rect 0 61348 112 61376
rect 0 61292 700 61348
rect 756 61292 766 61348
rect 1586 61292 1596 61348
rect 1652 61292 10556 61348
rect 10612 61292 13132 61348
rect 13188 61292 13198 61348
rect 15922 61292 15932 61348
rect 15988 61292 16716 61348
rect 16772 61292 16782 61348
rect 0 61264 112 61292
rect 31584 61236 31696 61264
rect 12338 61180 12348 61236
rect 12404 61180 17388 61236
rect 17444 61180 17454 61236
rect 21522 61180 21532 61236
rect 21588 61180 22764 61236
rect 22820 61180 22830 61236
rect 30594 61180 30604 61236
rect 30660 61180 31696 61236
rect 3794 61124 3804 61180
rect 3860 61124 3908 61180
rect 3964 61124 4012 61180
rect 4068 61124 4078 61180
rect 23794 61124 23804 61180
rect 23860 61124 23908 61180
rect 23964 61124 24012 61180
rect 24068 61124 24078 61180
rect 31584 61152 31696 61180
rect 9538 61068 9548 61124
rect 9604 61068 10556 61124
rect 10612 61068 13804 61124
rect 13860 61068 17612 61124
rect 17668 61068 19068 61124
rect 19124 61068 20972 61124
rect 21028 61068 21038 61124
rect 14802 60956 14812 61012
rect 14868 60956 17164 61012
rect 17220 60956 17724 61012
rect 17780 60956 17790 61012
rect 0 60900 112 60928
rect 0 60844 700 60900
rect 756 60844 766 60900
rect 12450 60844 12460 60900
rect 12516 60844 16268 60900
rect 16324 60844 17836 60900
rect 17892 60844 20412 60900
rect 20468 60844 22428 60900
rect 22484 60844 22494 60900
rect 0 60816 112 60844
rect 11116 60732 14812 60788
rect 14868 60732 18508 60788
rect 18564 60732 18574 60788
rect 19282 60732 19292 60788
rect 19348 60732 20972 60788
rect 21028 60732 21038 60788
rect 21746 60732 21756 60788
rect 21812 60732 22204 60788
rect 22260 60732 23660 60788
rect 23716 60732 23726 60788
rect 2146 60620 2156 60676
rect 2212 60620 6636 60676
rect 6692 60620 6702 60676
rect 7746 60620 7756 60676
rect 7812 60620 10780 60676
rect 10836 60620 10846 60676
rect 11116 60564 11172 60732
rect 13122 60620 13132 60676
rect 13188 60620 14252 60676
rect 14308 60620 14318 60676
rect 15586 60620 15596 60676
rect 15652 60620 15932 60676
rect 15988 60620 15998 60676
rect 18162 60620 18172 60676
rect 18228 60620 18732 60676
rect 18788 60620 18798 60676
rect 20402 60620 20412 60676
rect 20468 60620 21868 60676
rect 21924 60620 22652 60676
rect 22708 60620 22718 60676
rect 1362 60508 1372 60564
rect 1428 60508 1820 60564
rect 1876 60508 1886 60564
rect 3154 60508 3164 60564
rect 3220 60508 11172 60564
rect 0 60452 112 60480
rect 0 60396 812 60452
rect 868 60396 878 60452
rect 0 60368 112 60396
rect 4454 60340 4464 60396
rect 4520 60340 4568 60396
rect 4624 60340 4672 60396
rect 4728 60340 4738 60396
rect 24454 60340 24464 60396
rect 24520 60340 24568 60396
rect 24624 60340 24672 60396
rect 24728 60340 24738 60396
rect 17714 60284 17724 60340
rect 17780 60284 17948 60340
rect 18004 60284 18014 60340
rect 5170 60172 5180 60228
rect 5236 60172 5964 60228
rect 6020 60172 6030 60228
rect 13570 60172 13580 60228
rect 13636 60172 16604 60228
rect 16660 60172 16670 60228
rect 19282 60172 19292 60228
rect 19348 60172 29596 60228
rect 29652 60172 29662 60228
rect 31584 60116 31696 60144
rect 6290 60060 6300 60116
rect 6356 60060 17500 60116
rect 17556 60060 20188 60116
rect 30594 60060 30604 60116
rect 30660 60060 31696 60116
rect 0 60004 112 60032
rect 20132 60004 20188 60060
rect 31584 60032 31696 60060
rect 0 59948 924 60004
rect 980 59948 990 60004
rect 2370 59948 2380 60004
rect 2436 59948 9884 60004
rect 9940 59948 9950 60004
rect 16594 59948 16604 60004
rect 16660 59948 18732 60004
rect 18788 59948 18956 60004
rect 19012 59948 19022 60004
rect 20132 59948 21868 60004
rect 21924 59948 21934 60004
rect 0 59920 112 59948
rect 2594 59836 2604 59892
rect 2660 59836 3612 59892
rect 3668 59836 5852 59892
rect 5908 59836 9436 59892
rect 9492 59836 9502 59892
rect 10098 59836 10108 59892
rect 10164 59836 18284 59892
rect 18340 59836 22204 59892
rect 22260 59836 22270 59892
rect 8754 59724 8764 59780
rect 8820 59724 14812 59780
rect 14868 59724 29708 59780
rect 29764 59724 29774 59780
rect 0 59556 112 59584
rect 3794 59556 3804 59612
rect 3860 59556 3908 59612
rect 3964 59556 4012 59612
rect 4068 59556 4078 59612
rect 23794 59556 23804 59612
rect 23860 59556 23908 59612
rect 23964 59556 24012 59612
rect 24068 59556 24078 59612
rect 0 59500 1036 59556
rect 1092 59500 1102 59556
rect 18722 59500 18732 59556
rect 18788 59500 19180 59556
rect 19236 59500 19246 59556
rect 20178 59500 20188 59556
rect 20244 59500 21644 59556
rect 21700 59500 21710 59556
rect 0 59472 112 59500
rect 10770 59388 10780 59444
rect 10836 59388 29484 59444
rect 29540 59388 29550 59444
rect 18946 59276 18956 59332
rect 19012 59276 19964 59332
rect 20020 59276 20030 59332
rect 20626 59276 20636 59332
rect 20692 59276 22092 59332
rect 22148 59276 22158 59332
rect 9426 59164 9436 59220
rect 9492 59164 13692 59220
rect 13748 59164 14700 59220
rect 14756 59164 14924 59220
rect 14980 59164 15372 59220
rect 15428 59164 16828 59220
rect 16884 59164 16894 59220
rect 0 59108 112 59136
rect 0 59052 2492 59108
rect 2548 59052 2558 59108
rect 2818 59052 2828 59108
rect 2884 59052 16716 59108
rect 16772 59052 16782 59108
rect 0 59024 112 59052
rect 31584 58996 31696 59024
rect 1362 58940 1372 58996
rect 1428 58940 1820 58996
rect 1876 58940 1886 58996
rect 30594 58940 30604 58996
rect 30660 58940 31696 58996
rect 31584 58912 31696 58940
rect 14578 58828 14588 58884
rect 14644 58828 16492 58884
rect 16548 58828 16558 58884
rect 4454 58772 4464 58828
rect 4520 58772 4568 58828
rect 4624 58772 4672 58828
rect 4728 58772 4738 58828
rect 24454 58772 24464 58828
rect 24520 58772 24568 58828
rect 24624 58772 24672 58828
rect 24728 58772 24738 58828
rect 1586 58716 1596 58772
rect 1652 58716 2268 58772
rect 2324 58716 2334 58772
rect 8306 58716 8316 58772
rect 8372 58716 9324 58772
rect 9380 58716 10108 58772
rect 10164 58716 10332 58772
rect 10388 58716 10398 58772
rect 0 58660 112 58688
rect 0 58604 924 58660
rect 980 58604 990 58660
rect 1362 58604 1372 58660
rect 1428 58604 11564 58660
rect 11620 58604 11630 58660
rect 17042 58604 17052 58660
rect 17108 58604 17948 58660
rect 18004 58604 18014 58660
rect 0 58576 112 58604
rect 7186 58492 7196 58548
rect 7252 58492 14028 58548
rect 14084 58492 19404 58548
rect 19460 58492 20860 58548
rect 20916 58492 20926 58548
rect 2034 58380 2044 58436
rect 2100 58380 13916 58436
rect 13972 58380 13982 58436
rect 0 58212 112 58240
rect 0 58156 1036 58212
rect 1092 58156 1102 58212
rect 1362 58156 1372 58212
rect 1428 58156 1932 58212
rect 1988 58156 1998 58212
rect 2156 58156 9996 58212
rect 10052 58156 14028 58212
rect 14084 58156 28700 58212
rect 28756 58156 28766 58212
rect 0 58128 112 58156
rect 2156 58100 2212 58156
rect 1922 58044 1932 58100
rect 1988 58044 2212 58100
rect 3794 57988 3804 58044
rect 3860 57988 3908 58044
rect 3964 57988 4012 58044
rect 4068 57988 4078 58044
rect 23794 57988 23804 58044
rect 23860 57988 23908 58044
rect 23964 57988 24012 58044
rect 24068 57988 24078 58044
rect 10658 57932 10668 57988
rect 10724 57932 11228 57988
rect 11284 57932 11294 57988
rect 31584 57876 31696 57904
rect 7746 57820 7756 57876
rect 7812 57820 15372 57876
rect 15428 57820 23436 57876
rect 23492 57820 23502 57876
rect 30594 57820 30604 57876
rect 30660 57820 31696 57876
rect 31584 57792 31696 57820
rect 0 57764 112 57792
rect 0 57708 1708 57764
rect 1764 57708 1774 57764
rect 3154 57708 3164 57764
rect 3220 57708 8540 57764
rect 8596 57708 29484 57764
rect 29540 57708 29550 57764
rect 0 57680 112 57708
rect 13570 57484 13580 57540
rect 13636 57484 25116 57540
rect 25172 57484 25182 57540
rect 3332 57372 4900 57428
rect 14242 57372 14252 57428
rect 14308 57372 15596 57428
rect 15652 57372 15662 57428
rect 0 57204 112 57232
rect 3332 57204 3388 57372
rect 4844 57316 4900 57372
rect 4844 57260 6076 57316
rect 6132 57260 19516 57316
rect 19572 57260 19582 57316
rect 4454 57204 4464 57260
rect 4520 57204 4568 57260
rect 4624 57204 4672 57260
rect 4728 57204 4738 57260
rect 24454 57204 24464 57260
rect 24520 57204 24568 57260
rect 24624 57204 24672 57260
rect 24728 57204 24738 57260
rect 0 57148 3388 57204
rect 16706 57148 16716 57204
rect 16772 57148 21196 57204
rect 21252 57148 21262 57204
rect 0 57120 112 57148
rect 8978 56924 8988 56980
rect 9044 56924 9548 56980
rect 9604 56924 10108 56980
rect 10164 56924 10174 56980
rect 10994 56924 11004 56980
rect 11060 56924 20188 56980
rect 20244 56924 20254 56980
rect 6626 56812 6636 56868
rect 6692 56812 8092 56868
rect 8148 56812 8158 56868
rect 9650 56812 9660 56868
rect 9716 56812 10444 56868
rect 10500 56812 10510 56868
rect 12226 56812 12236 56868
rect 12292 56812 13132 56868
rect 13188 56812 13198 56868
rect 0 56756 112 56784
rect 31584 56756 31696 56784
rect 0 56700 1260 56756
rect 1316 56700 1326 56756
rect 2930 56700 2940 56756
rect 2996 56700 4396 56756
rect 4452 56700 4462 56756
rect 30594 56700 30604 56756
rect 30660 56700 31696 56756
rect 0 56672 112 56700
rect 31584 56672 31696 56700
rect 4834 56588 4844 56644
rect 4900 56588 7420 56644
rect 7476 56588 14140 56644
rect 14196 56588 29260 56644
rect 29316 56588 29326 56644
rect 3794 56420 3804 56476
rect 3860 56420 3908 56476
rect 3964 56420 4012 56476
rect 4068 56420 4078 56476
rect 23794 56420 23804 56476
rect 23860 56420 23908 56476
rect 23964 56420 24012 56476
rect 24068 56420 24078 56476
rect 11442 56364 11452 56420
rect 11508 56364 15148 56420
rect 0 56308 112 56336
rect 15092 56308 15148 56364
rect 0 56252 3500 56308
rect 3556 56252 6860 56308
rect 6916 56252 6926 56308
rect 15092 56252 28252 56308
rect 28308 56252 28318 56308
rect 0 56224 112 56252
rect 4386 56140 4396 56196
rect 4452 56140 5852 56196
rect 5908 56140 6636 56196
rect 6692 56140 6702 56196
rect 14438 56140 14476 56196
rect 14532 56140 14542 56196
rect 9874 56028 9884 56084
rect 9940 56028 10332 56084
rect 10388 56028 11004 56084
rect 11060 56028 11070 56084
rect 11218 56028 11228 56084
rect 11284 56028 11676 56084
rect 11732 56028 12348 56084
rect 12404 56028 12414 56084
rect 21298 56028 21308 56084
rect 21364 56028 30268 56084
rect 30324 56028 30334 56084
rect 0 55860 112 55888
rect 0 55804 2492 55860
rect 2548 55804 3276 55860
rect 3332 55804 3342 55860
rect 0 55776 112 55804
rect 4454 55636 4464 55692
rect 4520 55636 4568 55692
rect 4624 55636 4672 55692
rect 4728 55636 4738 55692
rect 24454 55636 24464 55692
rect 24520 55636 24568 55692
rect 24624 55636 24672 55692
rect 24728 55636 24738 55692
rect 31584 55636 31696 55664
rect 30594 55580 30604 55636
rect 30660 55580 31696 55636
rect 31584 55552 31696 55580
rect 19282 55468 19292 55524
rect 19348 55468 20300 55524
rect 20356 55468 20366 55524
rect 0 55412 112 55440
rect 0 55356 1932 55412
rect 1988 55356 1998 55412
rect 5058 55356 5068 55412
rect 5124 55356 5292 55412
rect 5348 55356 5740 55412
rect 5796 55356 5806 55412
rect 9538 55356 9548 55412
rect 9604 55356 12348 55412
rect 12404 55356 12414 55412
rect 13122 55356 13132 55412
rect 13188 55356 14476 55412
rect 14532 55356 14542 55412
rect 0 55328 112 55356
rect 4610 55244 4620 55300
rect 4676 55244 6524 55300
rect 6580 55244 6590 55300
rect 8306 55244 8316 55300
rect 8372 55244 11900 55300
rect 11956 55244 11966 55300
rect 27682 55244 27692 55300
rect 27748 55244 28364 55300
rect 28420 55244 28430 55300
rect 23650 55132 23660 55188
rect 23716 55132 24780 55188
rect 24836 55132 24846 55188
rect 2594 55020 2604 55076
rect 2660 55020 3388 55076
rect 14578 55020 14588 55076
rect 14644 55020 15260 55076
rect 15316 55020 15326 55076
rect 0 54964 112 54992
rect 0 54908 1820 54964
rect 1876 54908 1886 54964
rect 0 54880 112 54908
rect 3332 54628 3388 55020
rect 3794 54852 3804 54908
rect 3860 54852 3908 54908
rect 3964 54852 4012 54908
rect 4068 54852 4078 54908
rect 23794 54852 23804 54908
rect 23860 54852 23908 54908
rect 23964 54852 24012 54908
rect 24068 54852 24078 54908
rect 6626 54796 6636 54852
rect 6692 54796 18732 54852
rect 18788 54796 18798 54852
rect 3714 54684 3724 54740
rect 3780 54684 5404 54740
rect 5460 54684 5470 54740
rect 5618 54684 5628 54740
rect 5684 54684 14140 54740
rect 14196 54684 14206 54740
rect 2146 54572 2156 54628
rect 2212 54572 2940 54628
rect 2996 54572 3006 54628
rect 3332 54572 20412 54628
rect 20468 54572 20478 54628
rect 0 54516 112 54544
rect 31584 54516 31696 54544
rect 0 54460 3388 54516
rect 7970 54460 7980 54516
rect 8036 54460 8764 54516
rect 8820 54460 8830 54516
rect 14886 54460 14924 54516
rect 14980 54460 14990 54516
rect 16370 54460 16380 54516
rect 16436 54460 17164 54516
rect 17220 54460 17230 54516
rect 30594 54460 30604 54516
rect 30660 54460 31696 54516
rect 0 54432 112 54460
rect 3332 54292 3388 54460
rect 31584 54432 31696 54460
rect 6290 54348 6300 54404
rect 6356 54348 9548 54404
rect 9604 54348 10892 54404
rect 10948 54348 10958 54404
rect 14130 54348 14140 54404
rect 14196 54348 15596 54404
rect 15652 54348 15662 54404
rect 3332 54236 15148 54292
rect 15092 54180 15148 54236
rect 15092 54124 18172 54180
rect 18228 54124 20188 54180
rect 0 54068 112 54096
rect 4454 54068 4464 54124
rect 4520 54068 4568 54124
rect 4624 54068 4672 54124
rect 4728 54068 4738 54124
rect 0 54012 1316 54068
rect 0 53984 112 54012
rect 1260 53844 1316 54012
rect 20132 53956 20188 54124
rect 24454 54068 24464 54124
rect 24520 54068 24568 54124
rect 24624 54068 24672 54124
rect 24728 54068 24738 54124
rect 1474 53900 1484 53956
rect 1540 53900 6300 53956
rect 6356 53900 6366 53956
rect 20132 53900 20300 53956
rect 20356 53900 20366 53956
rect 1260 53788 6636 53844
rect 6692 53788 6702 53844
rect 8194 53788 8204 53844
rect 8260 53788 9884 53844
rect 9940 53788 9950 53844
rect 10882 53788 10892 53844
rect 10948 53788 14924 53844
rect 14980 53788 19292 53844
rect 19348 53788 19358 53844
rect 6738 53676 6748 53732
rect 6804 53676 6972 53732
rect 7028 53676 7038 53732
rect 17154 53676 17164 53732
rect 17220 53676 21420 53732
rect 21476 53676 21486 53732
rect 21746 53676 21756 53732
rect 21812 53676 29932 53732
rect 29988 53676 29998 53732
rect 0 53620 112 53648
rect 0 53564 3276 53620
rect 3332 53564 3342 53620
rect 7522 53564 7532 53620
rect 7588 53564 9772 53620
rect 9828 53564 9838 53620
rect 14018 53564 14028 53620
rect 14084 53564 16156 53620
rect 16212 53564 16222 53620
rect 0 53536 112 53564
rect 2482 53452 2492 53508
rect 2548 53452 3500 53508
rect 3556 53452 4452 53508
rect 4610 53452 4620 53508
rect 4676 53452 5292 53508
rect 5348 53452 5358 53508
rect 15586 53452 15596 53508
rect 15652 53452 30156 53508
rect 30212 53452 30222 53508
rect 4396 53396 4452 53452
rect 31584 53396 31696 53424
rect 4396 53340 16492 53396
rect 16548 53340 16558 53396
rect 30594 53340 30604 53396
rect 30660 53340 31696 53396
rect 3794 53284 3804 53340
rect 3860 53284 3908 53340
rect 3964 53284 4012 53340
rect 4068 53284 4078 53340
rect 23794 53284 23804 53340
rect 23860 53284 23908 53340
rect 23964 53284 24012 53340
rect 24068 53284 24078 53340
rect 31584 53312 31696 53340
rect 5506 53228 5516 53284
rect 5572 53228 10892 53284
rect 10948 53228 10958 53284
rect 0 53172 112 53200
rect 0 53116 6300 53172
rect 6356 53116 6366 53172
rect 0 53088 112 53116
rect 7858 53004 7868 53060
rect 7924 53004 25004 53060
rect 25060 53004 25070 53060
rect 6514 52892 6524 52948
rect 6580 52892 6972 52948
rect 7028 52892 7038 52948
rect 8082 52892 8092 52948
rect 8148 52892 8316 52948
rect 8372 52892 8382 52948
rect 9174 52892 9212 52948
rect 9268 52892 9278 52948
rect 12226 52892 12236 52948
rect 12292 52892 15260 52948
rect 15316 52892 15326 52948
rect 1586 52780 1596 52836
rect 1652 52780 10108 52836
rect 10164 52780 10174 52836
rect 13682 52780 13692 52836
rect 13748 52780 14476 52836
rect 14532 52780 14700 52836
rect 14756 52780 14766 52836
rect 0 52724 112 52752
rect 10108 52724 10164 52780
rect 0 52668 1484 52724
rect 1540 52668 1550 52724
rect 4274 52668 4284 52724
rect 4340 52668 6412 52724
rect 6468 52668 6478 52724
rect 10108 52668 15148 52724
rect 15204 52668 15214 52724
rect 16818 52668 16828 52724
rect 16884 52668 30380 52724
rect 30436 52668 30446 52724
rect 0 52640 112 52668
rect 6626 52556 6636 52612
rect 6692 52556 12236 52612
rect 12292 52556 12302 52612
rect 14018 52556 14028 52612
rect 14084 52556 14476 52612
rect 14532 52556 14542 52612
rect 4454 52500 4464 52556
rect 4520 52500 4568 52556
rect 4624 52500 4672 52556
rect 4728 52500 4738 52556
rect 24454 52500 24464 52556
rect 24520 52500 24568 52556
rect 24624 52500 24672 52556
rect 24728 52500 24738 52556
rect 9762 52444 9772 52500
rect 9828 52444 16828 52500
rect 16884 52444 16894 52500
rect 4498 52332 4508 52388
rect 4564 52332 9660 52388
rect 9716 52332 9726 52388
rect 10210 52332 10220 52388
rect 10276 52332 11788 52388
rect 11844 52332 11854 52388
rect 0 52276 112 52304
rect 31584 52276 31696 52304
rect 0 52220 4844 52276
rect 4900 52220 4910 52276
rect 9762 52220 9772 52276
rect 9828 52220 10780 52276
rect 10836 52220 13132 52276
rect 13188 52220 13198 52276
rect 17042 52220 17052 52276
rect 17108 52220 30268 52276
rect 30324 52220 30334 52276
rect 30594 52220 30604 52276
rect 30660 52220 31696 52276
rect 0 52192 112 52220
rect 31584 52192 31696 52220
rect 3042 52108 3052 52164
rect 3108 52108 6636 52164
rect 6692 52108 6702 52164
rect 6850 52108 6860 52164
rect 6916 52108 8316 52164
rect 8372 52108 8382 52164
rect 9090 52108 9100 52164
rect 9156 52108 10892 52164
rect 10948 52108 10958 52164
rect 3052 51996 4844 52052
rect 4900 51996 4910 52052
rect 5618 51996 5628 52052
rect 5684 51996 10108 52052
rect 10164 51996 10174 52052
rect 14578 51996 14588 52052
rect 14644 51996 15372 52052
rect 15428 51996 19292 52052
rect 19348 51996 19358 52052
rect 0 51828 112 51856
rect 3052 51828 3108 51996
rect 0 51772 3108 51828
rect 3164 51884 20300 51940
rect 20356 51884 29484 51940
rect 29540 51884 29550 51940
rect 0 51744 112 51772
rect 0 51380 112 51408
rect 0 51324 1708 51380
rect 1764 51324 2940 51380
rect 2996 51324 3006 51380
rect 0 51296 112 51324
rect 0 50932 112 50960
rect 3164 50932 3220 51884
rect 9874 51772 9884 51828
rect 9940 51772 10668 51828
rect 10724 51772 10734 51828
rect 11442 51772 11452 51828
rect 11508 51772 20972 51828
rect 21028 51772 21038 51828
rect 3794 51716 3804 51772
rect 3860 51716 3908 51772
rect 3964 51716 4012 51772
rect 4068 51716 4078 51772
rect 23794 51716 23804 51772
rect 23860 51716 23908 51772
rect 23964 51716 24012 51772
rect 24068 51716 24078 51772
rect 3378 51548 3388 51604
rect 3444 51548 17948 51604
rect 18004 51548 18014 51604
rect 8530 51436 8540 51492
rect 8596 51436 9324 51492
rect 9380 51436 10444 51492
rect 10500 51436 10510 51492
rect 10322 51324 10332 51380
rect 10388 51324 11116 51380
rect 11172 51324 11182 51380
rect 11890 51324 11900 51380
rect 11956 51324 14812 51380
rect 14868 51324 14878 51380
rect 3378 51212 3388 51268
rect 3444 51212 6860 51268
rect 6916 51212 6926 51268
rect 10658 51212 10668 51268
rect 10724 51212 11564 51268
rect 11620 51212 11630 51268
rect 31584 51156 31696 51184
rect 4274 51100 4284 51156
rect 4340 51100 5516 51156
rect 5572 51100 5582 51156
rect 17266 51100 17276 51156
rect 17332 51100 30268 51156
rect 30324 51100 30334 51156
rect 30594 51100 30604 51156
rect 30660 51100 31696 51156
rect 31584 51072 31696 51100
rect 8754 50988 8764 51044
rect 8820 50988 9884 51044
rect 9940 50988 9950 51044
rect 10770 50988 10780 51044
rect 10836 50988 13244 51044
rect 13300 50988 13310 51044
rect 14914 50988 14924 51044
rect 14980 50988 15092 51044
rect 4454 50932 4464 50988
rect 4520 50932 4568 50988
rect 4624 50932 4672 50988
rect 4728 50932 4738 50988
rect 10780 50932 10836 50988
rect 0 50876 3220 50932
rect 6850 50876 6860 50932
rect 6916 50876 10836 50932
rect 10994 50876 11004 50932
rect 11060 50876 14588 50932
rect 14644 50876 14654 50932
rect 0 50848 112 50876
rect 1138 50764 1148 50820
rect 1204 50764 5068 50820
rect 5124 50764 5134 50820
rect 11218 50764 11228 50820
rect 11284 50764 13804 50820
rect 13860 50764 13870 50820
rect 802 50652 812 50708
rect 868 50652 1484 50708
rect 1540 50652 1550 50708
rect 2454 50652 2492 50708
rect 2548 50652 2558 50708
rect 3332 50652 11452 50708
rect 11508 50652 11518 50708
rect 12226 50652 12236 50708
rect 12292 50652 12796 50708
rect 12852 50652 12862 50708
rect 13570 50652 13580 50708
rect 13636 50652 14364 50708
rect 14420 50652 14430 50708
rect 2034 50540 2044 50596
rect 2100 50540 2828 50596
rect 2884 50540 2894 50596
rect 0 50484 112 50512
rect 3332 50484 3388 50652
rect 15036 50596 15092 50988
rect 24454 50932 24464 50988
rect 24520 50932 24568 50988
rect 24624 50932 24672 50988
rect 24728 50932 24738 50988
rect 15222 50876 15260 50932
rect 15316 50876 15326 50932
rect 17938 50652 17948 50708
rect 18004 50652 29372 50708
rect 29428 50652 29438 50708
rect 4946 50540 4956 50596
rect 5012 50540 5908 50596
rect 6066 50540 6076 50596
rect 6132 50540 6860 50596
rect 6916 50540 6926 50596
rect 7074 50540 7084 50596
rect 7140 50540 7644 50596
rect 7700 50540 8204 50596
rect 8260 50540 8270 50596
rect 10994 50540 11004 50596
rect 11060 50540 11228 50596
rect 11284 50540 11294 50596
rect 12562 50540 12572 50596
rect 12628 50540 13692 50596
rect 13748 50540 13758 50596
rect 14802 50540 14812 50596
rect 14868 50540 14878 50596
rect 15026 50540 15036 50596
rect 15092 50540 15102 50596
rect 5852 50484 5908 50540
rect 14812 50484 14868 50540
rect 0 50428 3388 50484
rect 4050 50428 4060 50484
rect 4116 50428 5628 50484
rect 5684 50428 5694 50484
rect 5852 50428 10332 50484
rect 10388 50428 11788 50484
rect 11844 50428 11854 50484
rect 12002 50428 12012 50484
rect 12068 50428 15820 50484
rect 15876 50428 15886 50484
rect 17938 50428 17948 50484
rect 18004 50428 18396 50484
rect 18452 50428 18462 50484
rect 0 50400 112 50428
rect 12572 50372 12628 50428
rect 12572 50316 12796 50372
rect 12852 50316 12862 50372
rect 8866 50204 8876 50260
rect 8932 50204 15316 50260
rect 15474 50204 15484 50260
rect 15540 50204 16380 50260
rect 16436 50204 16446 50260
rect 3794 50148 3804 50204
rect 3860 50148 3908 50204
rect 3964 50148 4012 50204
rect 4068 50148 4078 50204
rect 15260 50148 15316 50204
rect 23794 50148 23804 50204
rect 23860 50148 23908 50204
rect 23964 50148 24012 50204
rect 24068 50148 24078 50204
rect 15250 50092 15260 50148
rect 15316 50092 18396 50148
rect 18452 50092 18462 50148
rect 0 50036 112 50064
rect 31584 50036 31696 50064
rect 0 49980 1036 50036
rect 1092 49980 1102 50036
rect 2594 49980 2604 50036
rect 2660 49980 3276 50036
rect 3332 49980 3342 50036
rect 10658 49980 10668 50036
rect 10724 49980 11004 50036
rect 11060 49980 11070 50036
rect 14466 49980 14476 50036
rect 14532 49980 19516 50036
rect 19572 49980 19582 50036
rect 30594 49980 30604 50036
rect 30660 49980 31696 50036
rect 0 49952 112 49980
rect 31584 49952 31696 49980
rect 1250 49868 1260 49924
rect 1316 49868 3388 49924
rect 4946 49868 4956 49924
rect 5012 49868 15148 49924
rect 15204 49868 15214 49924
rect 3332 49812 3388 49868
rect 3332 49756 11004 49812
rect 11060 49756 11070 49812
rect 15810 49756 15820 49812
rect 15876 49756 16156 49812
rect 16212 49756 16222 49812
rect 6962 49644 6972 49700
rect 7028 49644 8988 49700
rect 9044 49644 10220 49700
rect 10276 49644 10556 49700
rect 10612 49644 14812 49700
rect 14868 49644 14878 49700
rect 15362 49644 15372 49700
rect 15428 49644 16268 49700
rect 16324 49644 16334 49700
rect 17154 49644 17164 49700
rect 17220 49644 30492 49700
rect 30548 49644 30558 49700
rect 0 49588 112 49616
rect 0 49532 1148 49588
rect 1204 49532 1214 49588
rect 2930 49532 2940 49588
rect 2996 49532 5292 49588
rect 5348 49532 6636 49588
rect 6692 49532 6702 49588
rect 7382 49532 7420 49588
rect 7476 49532 7486 49588
rect 16146 49532 16156 49588
rect 16212 49532 16380 49588
rect 16436 49532 16446 49588
rect 0 49504 112 49532
rect 11778 49420 11788 49476
rect 11844 49420 12684 49476
rect 12740 49420 12750 49476
rect 4454 49364 4464 49420
rect 4520 49364 4568 49420
rect 4624 49364 4672 49420
rect 4728 49364 4738 49420
rect 24454 49364 24464 49420
rect 24520 49364 24568 49420
rect 24624 49364 24672 49420
rect 24728 49364 24738 49420
rect 4834 49308 4844 49364
rect 4900 49308 10444 49364
rect 10500 49308 11340 49364
rect 11396 49308 11406 49364
rect 2258 49196 2268 49252
rect 2324 49196 9268 49252
rect 12674 49196 12684 49252
rect 12740 49196 14364 49252
rect 14420 49196 14430 49252
rect 0 49140 112 49168
rect 0 49084 3276 49140
rect 3332 49084 3342 49140
rect 3490 49084 3500 49140
rect 3556 49084 4844 49140
rect 4900 49084 4910 49140
rect 0 49056 112 49084
rect 9212 49028 9268 49196
rect 14364 49140 14420 49196
rect 14364 49084 17836 49140
rect 17892 49084 17902 49140
rect 19730 49084 19740 49140
rect 19796 49084 30380 49140
rect 30436 49084 30446 49140
rect 1922 48972 1932 49028
rect 1988 48972 3724 49028
rect 3780 48972 3790 49028
rect 5842 48972 5852 49028
rect 5908 48972 6748 49028
rect 6804 48972 7756 49028
rect 7812 48972 7822 49028
rect 9212 48972 20188 49028
rect 20244 48972 20254 49028
rect 31584 48916 31696 48944
rect 2706 48860 2716 48916
rect 2772 48860 5068 48916
rect 5124 48860 6188 48916
rect 6244 48860 6254 48916
rect 9986 48860 9996 48916
rect 10052 48860 10220 48916
rect 10276 48860 10286 48916
rect 12338 48860 12348 48916
rect 12404 48860 12908 48916
rect 12964 48860 12974 48916
rect 15250 48860 15260 48916
rect 15316 48860 17388 48916
rect 17444 48860 17454 48916
rect 30594 48860 30604 48916
rect 30660 48860 31696 48916
rect 31584 48832 31696 48860
rect 2716 48748 3612 48804
rect 3668 48748 4956 48804
rect 5012 48748 5022 48804
rect 9650 48748 9660 48804
rect 9716 48748 10668 48804
rect 10724 48748 10734 48804
rect 0 48692 112 48720
rect 2716 48692 2772 48748
rect 0 48636 2492 48692
rect 2548 48636 2558 48692
rect 2706 48636 2716 48692
rect 2772 48636 2782 48692
rect 7074 48636 7084 48692
rect 7140 48636 7532 48692
rect 7588 48636 7598 48692
rect 10098 48636 10108 48692
rect 10164 48636 12908 48692
rect 12964 48636 12974 48692
rect 0 48608 112 48636
rect 3794 48580 3804 48636
rect 3860 48580 3908 48636
rect 3964 48580 4012 48636
rect 4068 48580 4078 48636
rect 23794 48580 23804 48636
rect 23860 48580 23908 48636
rect 23964 48580 24012 48636
rect 24068 48580 24078 48636
rect 1362 48524 1372 48580
rect 1428 48524 3276 48580
rect 3332 48524 3342 48580
rect 9538 48524 9548 48580
rect 9604 48524 11340 48580
rect 11396 48524 11406 48580
rect 12226 48524 12236 48580
rect 12292 48524 12572 48580
rect 12628 48524 12638 48580
rect 14578 48524 14588 48580
rect 14644 48524 15036 48580
rect 15092 48524 15102 48580
rect 16594 48524 16604 48580
rect 16660 48524 17948 48580
rect 18004 48524 18014 48580
rect 1586 48412 1596 48468
rect 1652 48412 2156 48468
rect 2212 48412 2222 48468
rect 2380 48412 9156 48468
rect 9314 48412 9324 48468
rect 9380 48412 10108 48468
rect 10164 48412 10174 48468
rect 10994 48412 11004 48468
rect 11060 48412 11676 48468
rect 11732 48412 11742 48468
rect 2380 48356 2436 48412
rect 9100 48356 9156 48412
rect 1026 48300 1036 48356
rect 1092 48300 1708 48356
rect 1764 48300 2436 48356
rect 2818 48300 2828 48356
rect 2884 48300 3612 48356
rect 3668 48300 3678 48356
rect 3948 48300 7196 48356
rect 7252 48300 7262 48356
rect 9100 48300 13860 48356
rect 15026 48300 15036 48356
rect 15092 48300 16940 48356
rect 16996 48300 17006 48356
rect 18732 48300 30044 48356
rect 30100 48300 30110 48356
rect 0 48244 112 48272
rect 0 48188 1764 48244
rect 3490 48188 3500 48244
rect 3556 48188 3724 48244
rect 3780 48188 3790 48244
rect 0 48160 112 48188
rect 1708 47908 1764 48188
rect 3948 48132 4004 48300
rect 13804 48244 13860 48300
rect 18732 48244 18788 48300
rect 2258 48076 2268 48132
rect 2324 48076 2604 48132
rect 2660 48076 4004 48132
rect 4172 48188 5964 48244
rect 6020 48188 6030 48244
rect 6626 48188 6636 48244
rect 6692 48188 7868 48244
rect 7924 48188 7934 48244
rect 10770 48188 10780 48244
rect 10836 48188 11228 48244
rect 11284 48188 11294 48244
rect 11452 48188 11900 48244
rect 11956 48188 11966 48244
rect 12226 48188 12236 48244
rect 12292 48188 13580 48244
rect 13636 48188 13646 48244
rect 13804 48188 14924 48244
rect 14980 48188 16828 48244
rect 16884 48188 18788 48244
rect 18946 48188 18956 48244
rect 19012 48188 30268 48244
rect 30324 48188 30334 48244
rect 4172 48020 4228 48188
rect 11452 48132 11508 48188
rect 2034 47964 2044 48020
rect 2100 47964 2492 48020
rect 2548 47964 2558 48020
rect 3042 47964 3052 48020
rect 3108 47964 4060 48020
rect 4116 47964 4228 48020
rect 4284 48076 7084 48132
rect 7140 48076 7150 48132
rect 9874 48076 9884 48132
rect 9940 48076 11452 48132
rect 11508 48076 11518 48132
rect 11666 48076 11676 48132
rect 11732 48076 13020 48132
rect 13076 48076 13086 48132
rect 15092 48076 28812 48132
rect 28868 48076 28878 48132
rect 4284 47908 4340 48076
rect 15092 48020 15148 48076
rect 6402 47964 6412 48020
rect 6468 47964 6478 48020
rect 10210 47964 10220 48020
rect 10276 47964 10444 48020
rect 10500 47964 10510 48020
rect 14802 47964 14812 48020
rect 14868 47964 14924 48020
rect 14980 47964 15148 48020
rect 23538 47964 23548 48020
rect 23604 47964 30268 48020
rect 30324 47964 30334 48020
rect 1708 47852 4340 47908
rect 6412 47908 6468 47964
rect 14812 47908 14868 47964
rect 6412 47852 14868 47908
rect 14924 47852 16604 47908
rect 16660 47852 16670 47908
rect 0 47796 112 47824
rect 4454 47796 4464 47852
rect 4520 47796 4568 47852
rect 4624 47796 4672 47852
rect 4728 47796 4738 47852
rect 14924 47796 14980 47852
rect 24454 47796 24464 47852
rect 24520 47796 24568 47852
rect 24624 47796 24672 47852
rect 24728 47796 24738 47852
rect 31584 47796 31696 47824
rect 0 47740 2268 47796
rect 2324 47740 2334 47796
rect 14354 47740 14364 47796
rect 14420 47740 14980 47796
rect 15092 47740 19404 47796
rect 19460 47740 19470 47796
rect 30594 47740 30604 47796
rect 30660 47740 31696 47796
rect 0 47712 112 47740
rect 2268 47628 9212 47684
rect 9268 47628 9278 47684
rect 2268 47572 2324 47628
rect 1894 47516 1932 47572
rect 1988 47516 1998 47572
rect 2258 47516 2268 47572
rect 2324 47516 2334 47572
rect 2930 47516 2940 47572
rect 2996 47516 3724 47572
rect 3780 47516 3790 47572
rect 6514 47516 6524 47572
rect 6580 47516 7196 47572
rect 7252 47516 14980 47572
rect 14924 47460 14980 47516
rect 2706 47404 2716 47460
rect 2772 47404 4172 47460
rect 4228 47404 4238 47460
rect 5394 47404 5404 47460
rect 5460 47404 12236 47460
rect 12292 47404 12684 47460
rect 12740 47404 12750 47460
rect 14914 47404 14924 47460
rect 14980 47404 14990 47460
rect 0 47348 112 47376
rect 15092 47348 15148 47740
rect 31584 47712 31696 47740
rect 17490 47516 17500 47572
rect 17556 47516 19292 47572
rect 19348 47516 19358 47572
rect 15922 47404 15932 47460
rect 15988 47404 17052 47460
rect 17108 47404 17118 47460
rect 18694 47404 18732 47460
rect 18788 47404 18798 47460
rect 22642 47404 22652 47460
rect 22708 47404 30268 47460
rect 30324 47404 30334 47460
rect 0 47292 3388 47348
rect 3602 47292 3612 47348
rect 3668 47292 6076 47348
rect 6132 47292 6636 47348
rect 6692 47292 6702 47348
rect 6962 47292 6972 47348
rect 7028 47292 7084 47348
rect 7140 47292 7150 47348
rect 7420 47292 9212 47348
rect 9268 47292 15148 47348
rect 16566 47292 16604 47348
rect 16660 47292 19740 47348
rect 19796 47292 19806 47348
rect 0 47264 112 47292
rect 3332 47236 3388 47292
rect 7420 47236 7476 47292
rect 2706 47180 2716 47236
rect 2772 47180 3164 47236
rect 3220 47180 3230 47236
rect 3332 47180 7476 47236
rect 7858 47180 7868 47236
rect 7924 47180 8876 47236
rect 8932 47180 8942 47236
rect 2482 47068 2492 47124
rect 2548 47068 3052 47124
rect 3108 47068 3118 47124
rect 4834 47068 4844 47124
rect 4900 47068 6972 47124
rect 7028 47068 11228 47124
rect 11284 47068 11294 47124
rect 3794 47012 3804 47068
rect 3860 47012 3908 47068
rect 3964 47012 4012 47068
rect 4068 47012 4078 47068
rect 7532 47012 7588 47068
rect 23794 47012 23804 47068
rect 23860 47012 23908 47068
rect 23964 47012 24012 47068
rect 24068 47012 24078 47068
rect 5058 46956 5068 47012
rect 5124 46956 6748 47012
rect 6804 46956 6814 47012
rect 7522 46956 7532 47012
rect 7588 46956 7598 47012
rect 12450 46956 12460 47012
rect 12516 46956 13356 47012
rect 13412 46956 13422 47012
rect 20178 46956 20188 47012
rect 20244 46956 23548 47012
rect 23604 46956 23614 47012
rect 0 46900 112 46928
rect 0 46844 10892 46900
rect 10948 46844 18620 46900
rect 18676 46844 18686 46900
rect 0 46816 112 46844
rect 1474 46732 1484 46788
rect 1540 46732 3500 46788
rect 3556 46732 4956 46788
rect 5012 46732 5022 46788
rect 7074 46732 7084 46788
rect 7140 46732 10220 46788
rect 10276 46732 10444 46788
rect 10500 46732 10510 46788
rect 31584 46676 31696 46704
rect 2930 46620 2940 46676
rect 2996 46620 5852 46676
rect 5908 46620 5918 46676
rect 8978 46620 8988 46676
rect 9044 46620 11116 46676
rect 11172 46620 11182 46676
rect 30594 46620 30604 46676
rect 30660 46620 31696 46676
rect 31584 46592 31696 46620
rect 1698 46508 1708 46564
rect 1764 46508 7756 46564
rect 7812 46508 7822 46564
rect 9874 46508 9884 46564
rect 9940 46508 10108 46564
rect 10164 46508 11004 46564
rect 11060 46508 11070 46564
rect 11974 46508 12012 46564
rect 12068 46508 14364 46564
rect 14420 46508 14430 46564
rect 16370 46508 16380 46564
rect 16436 46508 16716 46564
rect 16772 46508 16782 46564
rect 0 46452 112 46480
rect 0 46396 11788 46452
rect 11844 46396 14812 46452
rect 14868 46396 23212 46452
rect 23268 46396 23278 46452
rect 0 46368 112 46396
rect 5404 46284 14028 46340
rect 14084 46284 14588 46340
rect 14644 46284 17276 46340
rect 17332 46284 17342 46340
rect 4454 46228 4464 46284
rect 4520 46228 4568 46284
rect 4624 46228 4672 46284
rect 4728 46228 4738 46284
rect 5404 46116 5460 46284
rect 24454 46228 24464 46284
rect 24520 46228 24568 46284
rect 24624 46228 24672 46284
rect 24728 46228 24738 46284
rect 10210 46172 10220 46228
rect 10276 46172 22764 46228
rect 22820 46172 22830 46228
rect 1810 46060 1820 46116
rect 1876 46060 5404 46116
rect 5460 46060 5470 46116
rect 9650 46060 9660 46116
rect 9716 46060 10108 46116
rect 10164 46060 10174 46116
rect 16034 46060 16044 46116
rect 16100 46060 17836 46116
rect 17892 46060 17902 46116
rect 0 46004 112 46032
rect 0 45948 5964 46004
rect 6020 45948 6030 46004
rect 7046 45948 7084 46004
rect 7140 45948 7150 46004
rect 10546 45948 10556 46004
rect 10612 45948 11004 46004
rect 11060 45948 15148 46004
rect 16370 45948 16380 46004
rect 16436 45948 16604 46004
rect 16660 45948 16670 46004
rect 0 45920 112 45948
rect 15092 45892 15148 45948
rect 690 45836 700 45892
rect 756 45836 1596 45892
rect 1652 45836 1662 45892
rect 4834 45836 4844 45892
rect 4900 45836 4956 45892
rect 5012 45836 5022 45892
rect 5282 45836 5292 45892
rect 5348 45836 6524 45892
rect 6580 45836 6590 45892
rect 8194 45836 8204 45892
rect 8260 45836 9100 45892
rect 9156 45836 9166 45892
rect 10332 45836 11228 45892
rect 11284 45836 11294 45892
rect 15092 45836 20076 45892
rect 20132 45836 22652 45892
rect 22708 45836 22718 45892
rect 4844 45780 4900 45836
rect 10332 45780 10388 45836
rect 1708 45724 4900 45780
rect 8978 45724 8988 45780
rect 9044 45724 10332 45780
rect 10388 45724 10398 45780
rect 0 45556 112 45584
rect 1708 45556 1764 45724
rect 2146 45612 2156 45668
rect 2212 45612 5068 45668
rect 5124 45612 5134 45668
rect 6626 45612 6636 45668
rect 6692 45612 9884 45668
rect 9940 45612 9950 45668
rect 10098 45612 10108 45668
rect 10164 45612 12348 45668
rect 12404 45612 12414 45668
rect 20850 45612 20860 45668
rect 20916 45612 21308 45668
rect 21364 45612 21374 45668
rect 31584 45556 31696 45584
rect 0 45500 1764 45556
rect 4386 45500 4396 45556
rect 4452 45500 5292 45556
rect 5348 45500 5358 45556
rect 6178 45500 6188 45556
rect 6244 45500 16604 45556
rect 16660 45500 16670 45556
rect 30594 45500 30604 45556
rect 30660 45500 31696 45556
rect 0 45472 112 45500
rect 3794 45444 3804 45500
rect 3860 45444 3908 45500
rect 3964 45444 4012 45500
rect 4068 45444 4078 45500
rect 23794 45444 23804 45500
rect 23860 45444 23908 45500
rect 23964 45444 24012 45500
rect 24068 45444 24078 45500
rect 31584 45472 31696 45500
rect 1138 45388 1148 45444
rect 1204 45388 1708 45444
rect 1764 45388 1774 45444
rect 4946 45388 4956 45444
rect 5012 45388 5460 45444
rect 5842 45388 5852 45444
rect 5908 45388 8876 45444
rect 8932 45388 8942 45444
rect 9874 45388 9884 45444
rect 9940 45388 10444 45444
rect 10500 45388 11228 45444
rect 11284 45388 12012 45444
rect 12068 45388 12078 45444
rect 5404 45332 5460 45388
rect 5404 45276 8596 45332
rect 9314 45276 9324 45332
rect 9380 45276 15260 45332
rect 15316 45276 15326 45332
rect 24882 45276 24892 45332
rect 24948 45276 29708 45332
rect 29764 45276 29774 45332
rect 8540 45220 8596 45276
rect 5954 45164 5964 45220
rect 6020 45164 7532 45220
rect 7588 45164 7598 45220
rect 8540 45164 13468 45220
rect 13524 45164 14364 45220
rect 14420 45164 14430 45220
rect 19730 45164 19740 45220
rect 19796 45164 23212 45220
rect 23268 45164 23278 45220
rect 0 45108 112 45136
rect 0 45052 2044 45108
rect 2100 45052 2110 45108
rect 6822 45052 6860 45108
rect 6916 45052 6926 45108
rect 8166 45052 8204 45108
rect 8260 45052 8270 45108
rect 10182 45052 10220 45108
rect 10276 45052 11340 45108
rect 11396 45052 11406 45108
rect 11666 45052 11676 45108
rect 11732 45052 18060 45108
rect 18116 45052 18126 45108
rect 0 45024 112 45052
rect 5170 44940 5180 44996
rect 5236 44940 5516 44996
rect 5572 44940 6076 44996
rect 6132 44940 6142 44996
rect 1586 44828 1596 44884
rect 1652 44828 2828 44884
rect 2884 44828 3388 44884
rect 3444 44828 3454 44884
rect 5618 44828 5628 44884
rect 5684 44828 8092 44884
rect 8148 44828 9660 44884
rect 9716 44828 9726 44884
rect 9874 44828 9884 44884
rect 9940 44828 9950 44884
rect 21858 44828 21868 44884
rect 21924 44828 29484 44884
rect 29540 44828 29550 44884
rect 9884 44772 9940 44828
rect 1698 44716 1708 44772
rect 1764 44716 2492 44772
rect 2548 44716 2558 44772
rect 9772 44716 9940 44772
rect 0 44660 112 44688
rect 4454 44660 4464 44716
rect 4520 44660 4568 44716
rect 4624 44660 4672 44716
rect 4728 44660 4738 44716
rect 0 44604 1484 44660
rect 1540 44604 1550 44660
rect 0 44576 112 44604
rect 7970 44492 7980 44548
rect 8036 44492 8092 44548
rect 8148 44492 8158 44548
rect 9772 44436 9828 44716
rect 24454 44660 24464 44716
rect 24520 44660 24568 44716
rect 24624 44660 24672 44716
rect 24728 44660 24738 44716
rect 10882 44492 10892 44548
rect 10948 44492 11340 44548
rect 11396 44492 11406 44548
rect 19506 44492 19516 44548
rect 19572 44492 19852 44548
rect 19908 44492 20524 44548
rect 20580 44492 20590 44548
rect 22194 44492 22204 44548
rect 22260 44492 22540 44548
rect 22596 44492 22606 44548
rect 31584 44436 31696 44464
rect 7074 44380 7084 44436
rect 7140 44380 8092 44436
rect 8148 44380 8158 44436
rect 9762 44380 9772 44436
rect 9828 44380 9838 44436
rect 11442 44380 11452 44436
rect 11508 44380 20412 44436
rect 20468 44380 20478 44436
rect 30594 44380 30604 44436
rect 30660 44380 31696 44436
rect 31584 44352 31696 44380
rect 8306 44268 8316 44324
rect 8372 44268 9100 44324
rect 9156 44268 9166 44324
rect 9874 44268 9884 44324
rect 9940 44268 14252 44324
rect 14308 44268 14318 44324
rect 0 44212 112 44240
rect 0 44156 1260 44212
rect 1316 44156 1326 44212
rect 19366 44156 19404 44212
rect 19460 44156 23100 44212
rect 23156 44156 23166 44212
rect 0 44128 112 44156
rect 1474 44044 1484 44100
rect 1540 44044 6748 44100
rect 6804 44044 7924 44100
rect 8082 44044 8092 44100
rect 8148 44044 9324 44100
rect 9380 44044 9390 44100
rect 14354 44044 14364 44100
rect 14420 44044 19740 44100
rect 19796 44044 19806 44100
rect 7868 43988 7924 44044
rect 7868 43932 10332 43988
rect 10388 43932 11004 43988
rect 11060 43932 11070 43988
rect 15474 43932 15484 43988
rect 15540 43932 16828 43988
rect 16884 43932 16894 43988
rect 18162 43932 18172 43988
rect 18228 43932 18844 43988
rect 18900 43932 18910 43988
rect 3794 43876 3804 43932
rect 3860 43876 3908 43932
rect 3964 43876 4012 43932
rect 4068 43876 4078 43932
rect 23794 43876 23804 43932
rect 23860 43876 23908 43932
rect 23964 43876 24012 43932
rect 24068 43876 24078 43932
rect 9314 43820 9324 43876
rect 9380 43820 10220 43876
rect 10276 43820 10286 43876
rect 0 43764 112 43792
rect 0 43708 4284 43764
rect 4340 43708 4350 43764
rect 4946 43708 4956 43764
rect 5012 43708 9772 43764
rect 9828 43708 9838 43764
rect 11442 43708 11452 43764
rect 11508 43708 11518 43764
rect 0 43680 112 43708
rect 1250 43596 1260 43652
rect 1316 43596 8260 43652
rect 9650 43596 9660 43652
rect 9716 43596 10892 43652
rect 10948 43596 10958 43652
rect 8204 43540 8260 43596
rect 11452 43540 11508 43708
rect 13010 43596 13020 43652
rect 13076 43596 17220 43652
rect 17378 43596 17388 43652
rect 17444 43596 17612 43652
rect 17668 43596 17678 43652
rect 17164 43540 17220 43596
rect 2034 43484 2044 43540
rect 2100 43484 4284 43540
rect 4340 43484 4350 43540
rect 8194 43484 8204 43540
rect 8260 43484 11508 43540
rect 14466 43484 14476 43540
rect 14532 43484 15036 43540
rect 15092 43484 15102 43540
rect 17154 43484 17164 43540
rect 17220 43484 18844 43540
rect 18900 43484 18910 43540
rect 21522 43484 21532 43540
rect 21588 43484 22092 43540
rect 22148 43484 22158 43540
rect 1810 43372 1820 43428
rect 1876 43372 14028 43428
rect 14084 43372 14094 43428
rect 17826 43372 17836 43428
rect 17892 43372 18620 43428
rect 18676 43372 18686 43428
rect 0 43316 112 43344
rect 31584 43316 31696 43344
rect 0 43260 6188 43316
rect 6244 43260 6254 43316
rect 7746 43260 7756 43316
rect 7812 43260 8652 43316
rect 8708 43260 9996 43316
rect 10052 43260 10062 43316
rect 14354 43260 14364 43316
rect 14420 43260 15036 43316
rect 15092 43260 15102 43316
rect 30594 43260 30604 43316
rect 30660 43260 31696 43316
rect 0 43232 112 43260
rect 4454 43092 4464 43148
rect 4520 43092 4568 43148
rect 4624 43092 4672 43148
rect 4728 43092 4738 43148
rect 7756 43092 7812 43260
rect 31584 43232 31696 43260
rect 11890 43148 11900 43204
rect 11956 43148 16044 43204
rect 16100 43148 16110 43204
rect 24454 43092 24464 43148
rect 24520 43092 24568 43148
rect 24624 43092 24672 43148
rect 24728 43092 24738 43148
rect 5730 43036 5740 43092
rect 5796 43036 6860 43092
rect 6916 43036 7812 43092
rect 10882 43036 10892 43092
rect 10948 43036 14812 43092
rect 14868 43036 14878 43092
rect 2034 42924 2044 42980
rect 2100 42924 5628 42980
rect 5684 42924 5852 42980
rect 5908 42924 5918 42980
rect 7186 42924 7196 42980
rect 7252 42924 9324 42980
rect 9380 42924 9390 42980
rect 12338 42924 12348 42980
rect 12404 42924 12684 42980
rect 12740 42924 12750 42980
rect 14242 42924 14252 42980
rect 14308 42924 15036 42980
rect 15092 42924 15102 42980
rect 16594 42924 16604 42980
rect 16660 42924 26908 42980
rect 0 42868 112 42896
rect 26852 42868 26908 42924
rect 0 42812 16772 42868
rect 26852 42812 30380 42868
rect 30436 42812 30446 42868
rect 0 42784 112 42812
rect 16716 42756 16772 42812
rect 7186 42700 7196 42756
rect 7252 42700 11452 42756
rect 11508 42700 12908 42756
rect 12964 42700 12974 42756
rect 14578 42700 14588 42756
rect 14644 42700 15708 42756
rect 15764 42700 15774 42756
rect 16716 42700 20188 42756
rect 20244 42700 20254 42756
rect 1138 42588 1148 42644
rect 1204 42588 1932 42644
rect 1988 42588 1998 42644
rect 4274 42588 4284 42644
rect 4340 42588 5852 42644
rect 5908 42588 11340 42644
rect 11396 42588 11406 42644
rect 3332 42476 7196 42532
rect 7252 42476 7262 42532
rect 9650 42476 9660 42532
rect 9716 42476 12012 42532
rect 12068 42476 13916 42532
rect 13972 42476 13982 42532
rect 0 42420 112 42448
rect 3332 42420 3388 42476
rect 0 42364 3388 42420
rect 9314 42364 9324 42420
rect 9380 42364 11900 42420
rect 11956 42364 11966 42420
rect 0 42336 112 42364
rect 3794 42308 3804 42364
rect 3860 42308 3908 42364
rect 3964 42308 4012 42364
rect 4068 42308 4078 42364
rect 23794 42308 23804 42364
rect 23860 42308 23908 42364
rect 23964 42308 24012 42364
rect 24068 42308 24078 42364
rect 31584 42196 31696 42224
rect 3332 42140 6076 42196
rect 6132 42140 6142 42196
rect 7746 42140 7756 42196
rect 7812 42140 7980 42196
rect 8036 42140 12348 42196
rect 12404 42140 12414 42196
rect 30594 42140 30604 42196
rect 30660 42140 31696 42196
rect 3332 42084 3388 42140
rect 31584 42112 31696 42140
rect 2930 42028 2940 42084
rect 2996 42028 3388 42084
rect 5842 42028 5852 42084
rect 5908 42028 8988 42084
rect 9044 42028 9054 42084
rect 10556 42028 11900 42084
rect 11956 42028 13468 42084
rect 13524 42028 13534 42084
rect 19730 42028 19740 42084
rect 19796 42028 22652 42084
rect 22708 42028 22718 42084
rect 0 41972 112 42000
rect 10556 41972 10612 42028
rect 0 41916 1820 41972
rect 1876 41916 1886 41972
rect 4162 41916 4172 41972
rect 4228 41916 4396 41972
rect 4452 41916 4956 41972
rect 5012 41916 5022 41972
rect 5730 41916 5740 41972
rect 5796 41916 5806 41972
rect 6402 41916 6412 41972
rect 6468 41916 8652 41972
rect 8708 41916 8718 41972
rect 10546 41916 10556 41972
rect 10612 41916 10622 41972
rect 10994 41916 11004 41972
rect 11060 41916 11788 41972
rect 11844 41916 11854 41972
rect 14466 41916 14476 41972
rect 14532 41916 15372 41972
rect 15428 41916 16492 41972
rect 16548 41916 16828 41972
rect 16884 41916 17612 41972
rect 17668 41916 17678 41972
rect 17826 41916 17836 41972
rect 17892 41916 17902 41972
rect 18274 41916 18284 41972
rect 18340 41916 18732 41972
rect 18788 41916 18798 41972
rect 19068 41916 20636 41972
rect 20692 41916 20702 41972
rect 20962 41916 20972 41972
rect 21028 41916 21308 41972
rect 21364 41916 21374 41972
rect 21522 41916 21532 41972
rect 21588 41916 22092 41972
rect 22148 41916 22158 41972
rect 0 41888 112 41916
rect 5740 41860 5796 41916
rect 17836 41860 17892 41916
rect 19068 41860 19124 41916
rect 1474 41804 1484 41860
rect 1540 41804 3164 41860
rect 3220 41804 3230 41860
rect 4274 41804 4284 41860
rect 4340 41804 5796 41860
rect 7298 41804 7308 41860
rect 7364 41804 9212 41860
rect 9268 41804 9278 41860
rect 9986 41804 9996 41860
rect 10052 41804 12572 41860
rect 12628 41804 12638 41860
rect 16258 41804 16268 41860
rect 16324 41804 17164 41860
rect 17220 41804 17230 41860
rect 17836 41804 19124 41860
rect 19282 41804 19292 41860
rect 19348 41804 19358 41860
rect 19618 41804 19628 41860
rect 19684 41804 21644 41860
rect 21700 41804 21710 41860
rect 19292 41748 19348 41804
rect 2146 41692 2156 41748
rect 2212 41692 5068 41748
rect 5124 41692 5134 41748
rect 5954 41692 5964 41748
rect 6020 41692 9548 41748
rect 9604 41692 9614 41748
rect 19292 41692 21756 41748
rect 21812 41692 21822 41748
rect 1586 41580 1596 41636
rect 1652 41580 2604 41636
rect 2660 41580 3388 41636
rect 3444 41580 3454 41636
rect 20850 41580 20860 41636
rect 20916 41580 23660 41636
rect 23716 41580 23726 41636
rect 0 41524 112 41552
rect 4454 41524 4464 41580
rect 4520 41524 4568 41580
rect 4624 41524 4672 41580
rect 4728 41524 4738 41580
rect 24454 41524 24464 41580
rect 24520 41524 24568 41580
rect 24624 41524 24672 41580
rect 24728 41524 24738 41580
rect 0 41468 2604 41524
rect 2660 41468 2670 41524
rect 3238 41468 3276 41524
rect 3332 41468 3342 41524
rect 15810 41468 15820 41524
rect 15876 41468 21420 41524
rect 21476 41468 21486 41524
rect 0 41440 112 41468
rect 242 41356 252 41412
rect 308 41356 4172 41412
rect 4228 41356 4238 41412
rect 4386 41356 4396 41412
rect 4452 41356 5292 41412
rect 5348 41356 5358 41412
rect 10994 41356 11004 41412
rect 11060 41356 11564 41412
rect 11620 41356 11630 41412
rect 20402 41356 20412 41412
rect 20468 41356 21420 41412
rect 21476 41356 22876 41412
rect 22932 41356 22942 41412
rect 4844 41244 6412 41300
rect 6468 41244 6478 41300
rect 4844 41188 4900 41244
rect 3378 41132 3388 41188
rect 3444 41132 4844 41188
rect 4900 41132 4910 41188
rect 5618 41132 5628 41188
rect 5684 41132 10780 41188
rect 10836 41132 10846 41188
rect 12674 41132 12684 41188
rect 12740 41132 13020 41188
rect 13076 41132 13086 41188
rect 21074 41132 21084 41188
rect 21140 41132 23772 41188
rect 23828 41132 23838 41188
rect 0 41076 112 41104
rect 31584 41076 31696 41104
rect 0 41020 1764 41076
rect 2930 41020 2940 41076
rect 2996 41020 3500 41076
rect 3556 41020 7868 41076
rect 7924 41020 7934 41076
rect 9986 41020 9996 41076
rect 10052 41020 10892 41076
rect 10948 41020 10958 41076
rect 30594 41020 30604 41076
rect 30660 41020 31696 41076
rect 0 40992 112 41020
rect 690 40908 700 40964
rect 756 40908 766 40964
rect 700 40852 756 40908
rect 1708 40852 1764 41020
rect 31584 40992 31696 41020
rect 2482 40908 2492 40964
rect 2548 40908 11116 40964
rect 11172 40908 14812 40964
rect 14868 40908 17052 40964
rect 17108 40908 17118 40964
rect 22418 40908 22428 40964
rect 22484 40908 28252 40964
rect 28308 40908 28318 40964
rect 700 40796 924 40852
rect 980 40796 990 40852
rect 1708 40796 2212 40852
rect 7756 40796 10668 40852
rect 10724 40796 10734 40852
rect 18834 40796 18844 40852
rect 18900 40796 21532 40852
rect 21588 40796 22988 40852
rect 23044 40796 23054 40852
rect 0 40628 112 40656
rect 0 40572 1148 40628
rect 1204 40572 1214 40628
rect 0 40544 112 40572
rect 2156 40516 2212 40796
rect 3794 40740 3804 40796
rect 3860 40740 3908 40796
rect 3964 40740 4012 40796
rect 4068 40740 4078 40796
rect 7756 40628 7812 40796
rect 23794 40740 23804 40796
rect 23860 40740 23908 40796
rect 23964 40740 24012 40796
rect 24068 40740 24078 40796
rect 7970 40684 7980 40740
rect 8036 40684 20636 40740
rect 20692 40684 20702 40740
rect 21298 40684 21308 40740
rect 21364 40684 22204 40740
rect 22260 40684 22270 40740
rect 2370 40572 2380 40628
rect 2436 40572 7812 40628
rect 8418 40572 8428 40628
rect 8484 40572 10332 40628
rect 10388 40572 10398 40628
rect 11330 40572 11340 40628
rect 11396 40572 26908 40628
rect 26852 40516 26908 40572
rect 2156 40460 7980 40516
rect 8036 40460 8046 40516
rect 8866 40460 8876 40516
rect 8932 40460 10220 40516
rect 10276 40460 10286 40516
rect 10658 40460 10668 40516
rect 10724 40460 11228 40516
rect 11284 40460 11294 40516
rect 13010 40460 13020 40516
rect 13076 40460 13804 40516
rect 13860 40460 14476 40516
rect 14532 40460 14542 40516
rect 16258 40460 16268 40516
rect 16324 40460 16716 40516
rect 16772 40460 16782 40516
rect 17154 40460 17164 40516
rect 17220 40460 18396 40516
rect 18452 40460 18462 40516
rect 18946 40460 18956 40516
rect 19012 40460 21644 40516
rect 21700 40460 21710 40516
rect 22082 40460 22092 40516
rect 22148 40460 22158 40516
rect 26852 40460 29484 40516
rect 29540 40460 29550 40516
rect 22092 40404 22148 40460
rect 3266 40348 3276 40404
rect 3332 40348 5180 40404
rect 5236 40348 5246 40404
rect 6178 40348 6188 40404
rect 6244 40348 10108 40404
rect 10164 40348 10174 40404
rect 10770 40348 10780 40404
rect 10836 40348 11564 40404
rect 11620 40348 11630 40404
rect 15810 40348 15820 40404
rect 15876 40348 16940 40404
rect 16996 40348 17006 40404
rect 18134 40348 18172 40404
rect 18228 40348 18238 40404
rect 19842 40348 19852 40404
rect 19908 40348 19964 40404
rect 20020 40348 20030 40404
rect 20962 40348 20972 40404
rect 21028 40348 22148 40404
rect 23090 40348 23100 40404
rect 23156 40348 23660 40404
rect 23716 40348 23726 40404
rect 2006 40236 2044 40292
rect 2100 40236 2110 40292
rect 2818 40236 2828 40292
rect 2884 40236 4956 40292
rect 5012 40236 5022 40292
rect 6066 40236 6076 40292
rect 6132 40236 6636 40292
rect 6692 40236 6702 40292
rect 11778 40236 11788 40292
rect 11844 40236 12572 40292
rect 12628 40236 13468 40292
rect 13524 40236 13534 40292
rect 15922 40236 15932 40292
rect 15988 40236 17388 40292
rect 17444 40236 17454 40292
rect 18610 40236 18620 40292
rect 18676 40236 19404 40292
rect 19460 40236 19470 40292
rect 20850 40236 20860 40292
rect 20916 40236 21308 40292
rect 21364 40236 21374 40292
rect 0 40180 112 40208
rect 0 40124 6412 40180
rect 6468 40124 6478 40180
rect 10098 40124 10108 40180
rect 10164 40124 18060 40180
rect 18116 40124 18126 40180
rect 0 40096 112 40124
rect 4946 40012 4956 40068
rect 5012 40012 5740 40068
rect 5796 40012 7308 40068
rect 7364 40012 15148 40068
rect 4454 39956 4464 40012
rect 4520 39956 4568 40012
rect 4624 39956 4672 40012
rect 4728 39956 4738 40012
rect 15092 39956 15148 40012
rect 24454 39956 24464 40012
rect 24520 39956 24568 40012
rect 24624 39956 24672 40012
rect 24728 39956 24738 40012
rect 31584 39956 31696 39984
rect 10210 39900 10220 39956
rect 10276 39900 11676 39956
rect 11732 39900 11742 39956
rect 15092 39900 17500 39956
rect 17556 39900 17566 39956
rect 30594 39900 30604 39956
rect 30660 39900 31696 39956
rect 31584 39872 31696 39900
rect 6178 39788 6188 39844
rect 6244 39788 26012 39844
rect 26068 39788 26078 39844
rect 0 39732 112 39760
rect 0 39676 14252 39732
rect 14308 39676 14318 39732
rect 0 39648 112 39676
rect 4946 39564 4956 39620
rect 5012 39564 6860 39620
rect 6916 39564 6926 39620
rect 7980 39564 12684 39620
rect 12740 39564 13916 39620
rect 13972 39564 13982 39620
rect 1250 39452 1260 39508
rect 1316 39452 1708 39508
rect 1764 39452 6076 39508
rect 6132 39452 6142 39508
rect 7980 39396 8036 39564
rect 10434 39452 10444 39508
rect 10500 39452 11564 39508
rect 11620 39452 11676 39508
rect 11732 39452 11742 39508
rect 18050 39452 18060 39508
rect 18116 39452 29484 39508
rect 29540 39452 29550 39508
rect 1138 39340 1148 39396
rect 1204 39340 1596 39396
rect 1652 39340 1662 39396
rect 4834 39340 4844 39396
rect 4900 39340 8036 39396
rect 8194 39340 8204 39396
rect 8260 39340 20524 39396
rect 20580 39340 20590 39396
rect 0 39284 112 39312
rect 0 39228 3388 39284
rect 5394 39228 5404 39284
rect 5460 39228 14924 39284
rect 14980 39228 14990 39284
rect 0 39200 112 39228
rect 3332 39060 3388 39228
rect 3794 39172 3804 39228
rect 3860 39172 3908 39228
rect 3964 39172 4012 39228
rect 4068 39172 4078 39228
rect 23794 39172 23804 39228
rect 23860 39172 23908 39228
rect 23964 39172 24012 39228
rect 24068 39172 24078 39228
rect 6514 39116 6524 39172
rect 6580 39116 7084 39172
rect 7140 39116 7150 39172
rect 8306 39116 8316 39172
rect 8372 39116 10108 39172
rect 10164 39116 10556 39172
rect 10612 39116 13468 39172
rect 13524 39116 13534 39172
rect 3332 39004 5068 39060
rect 5124 39004 5134 39060
rect 9874 39004 9884 39060
rect 9940 39004 11228 39060
rect 11284 39004 11294 39060
rect 11554 39004 11564 39060
rect 11620 39004 20860 39060
rect 20916 39004 20926 39060
rect 10770 38892 10780 38948
rect 10836 38892 11564 38948
rect 11620 38892 11630 38948
rect 0 38836 112 38864
rect 0 38780 4844 38836
rect 4900 38780 4910 38836
rect 6178 38780 6188 38836
rect 6244 38780 11564 38836
rect 11620 38780 11630 38836
rect 13234 38780 13244 38836
rect 13300 38780 14028 38836
rect 14084 38780 14094 38836
rect 14242 38780 14252 38836
rect 14308 38780 15260 38836
rect 15316 38780 15708 38836
rect 15764 38780 15774 38836
rect 0 38752 112 38780
rect 2818 38668 2828 38724
rect 2884 38668 4284 38724
rect 4340 38668 4350 38724
rect 6066 38668 6076 38724
rect 6132 38668 6636 38724
rect 6692 38668 6702 38724
rect 6850 38668 6860 38724
rect 6916 38668 8428 38724
rect 14662 38668 14700 38724
rect 14756 38668 14766 38724
rect 17490 38668 17500 38724
rect 17556 38668 21420 38724
rect 21476 38668 21486 38724
rect 8372 38612 8428 38668
rect 5506 38556 5516 38612
rect 5572 38556 5582 38612
rect 8372 38556 9436 38612
rect 9492 38556 9502 38612
rect 5516 38500 5572 38556
rect 5516 38444 5740 38500
rect 5796 38444 5806 38500
rect 6066 38444 6076 38500
rect 6132 38444 6188 38500
rect 6244 38444 6254 38500
rect 8866 38444 8876 38500
rect 8932 38444 10556 38500
rect 10612 38444 10622 38500
rect 15474 38444 15484 38500
rect 15540 38444 16044 38500
rect 16100 38444 16110 38500
rect 0 38388 112 38416
rect 4454 38388 4464 38444
rect 4520 38388 4568 38444
rect 4624 38388 4672 38444
rect 4728 38388 4738 38444
rect 24454 38388 24464 38444
rect 24520 38388 24568 38444
rect 24624 38388 24672 38444
rect 24728 38388 24738 38444
rect 0 38332 3388 38388
rect 5954 38332 5964 38388
rect 6020 38332 13580 38388
rect 13636 38332 14252 38388
rect 14308 38332 15148 38388
rect 16258 38332 16268 38388
rect 16324 38332 20188 38388
rect 20244 38332 22204 38388
rect 22260 38332 22270 38388
rect 0 38304 112 38332
rect 3332 38276 3388 38332
rect 15092 38276 15148 38332
rect 3332 38220 5180 38276
rect 5236 38220 5246 38276
rect 5618 38220 5628 38276
rect 5684 38220 9884 38276
rect 9940 38220 9950 38276
rect 11778 38220 11788 38276
rect 11844 38220 12124 38276
rect 12180 38220 12190 38276
rect 15092 38220 18396 38276
rect 18452 38220 18462 38276
rect 19842 38220 19852 38276
rect 19908 38220 24332 38276
rect 24388 38220 24398 38276
rect 1922 38108 1932 38164
rect 1988 38108 10220 38164
rect 10276 38108 10286 38164
rect 21074 38108 21084 38164
rect 21140 38108 27692 38164
rect 27748 38108 27758 38164
rect 3154 37996 3164 38052
rect 3220 37996 15036 38052
rect 15092 37996 15102 38052
rect 17826 37996 17836 38052
rect 17892 37996 19852 38052
rect 19908 37996 19918 38052
rect 22418 37996 22428 38052
rect 22484 37996 29484 38052
rect 29540 37996 29550 38052
rect 0 37940 112 37968
rect 14364 37940 14420 37996
rect 0 37884 8596 37940
rect 8754 37884 8764 37940
rect 8820 37884 9436 37940
rect 9492 37884 11676 37940
rect 11732 37884 13916 37940
rect 13972 37884 13982 37940
rect 14354 37884 14364 37940
rect 14420 37884 14430 37940
rect 18386 37884 18396 37940
rect 18452 37884 21308 37940
rect 21364 37884 21980 37940
rect 22036 37884 22046 37940
rect 0 37856 112 37884
rect 8540 37828 8596 37884
rect 3042 37772 3052 37828
rect 3108 37772 5292 37828
rect 5348 37772 5358 37828
rect 5618 37772 5628 37828
rect 5684 37772 6188 37828
rect 6244 37772 6254 37828
rect 6850 37772 6860 37828
rect 6916 37772 7196 37828
rect 7252 37772 7262 37828
rect 8540 37772 12236 37828
rect 12292 37772 12302 37828
rect 19394 37772 19404 37828
rect 19460 37772 31276 37828
rect 31332 37772 31342 37828
rect 5842 37660 5852 37716
rect 5908 37660 6076 37716
rect 6132 37660 6142 37716
rect 6290 37660 6300 37716
rect 6356 37660 10556 37716
rect 10612 37660 10622 37716
rect 3794 37604 3804 37660
rect 3860 37604 3908 37660
rect 3964 37604 4012 37660
rect 4068 37604 4078 37660
rect 23794 37604 23804 37660
rect 23860 37604 23908 37660
rect 23964 37604 24012 37660
rect 24068 37604 24078 37660
rect 5842 37548 5852 37604
rect 5908 37548 5964 37604
rect 6020 37548 6030 37604
rect 7410 37548 7420 37604
rect 7476 37548 7868 37604
rect 7924 37548 7934 37604
rect 18050 37548 18060 37604
rect 18116 37548 18620 37604
rect 18676 37548 18686 37604
rect 0 37492 112 37520
rect 0 37436 21308 37492
rect 21364 37436 22764 37492
rect 22820 37436 22830 37492
rect 0 37408 112 37436
rect 1474 37324 1484 37380
rect 1540 37324 2716 37380
rect 2772 37324 5628 37380
rect 5684 37324 5694 37380
rect 7494 37324 7532 37380
rect 7588 37324 7598 37380
rect 12226 37324 12236 37380
rect 12292 37324 12572 37380
rect 12628 37324 16156 37380
rect 16212 37324 16222 37380
rect 1922 37212 1932 37268
rect 1988 37212 2492 37268
rect 2548 37212 2558 37268
rect 5170 37212 5180 37268
rect 5236 37212 9436 37268
rect 9492 37212 9502 37268
rect 14466 37212 14476 37268
rect 14532 37212 15036 37268
rect 15092 37212 15102 37268
rect 16706 37212 16716 37268
rect 16772 37212 17276 37268
rect 17332 37212 17342 37268
rect 17910 37212 17948 37268
rect 18004 37212 18014 37268
rect 15036 37156 15092 37212
rect 5730 37100 5740 37156
rect 5796 37100 7308 37156
rect 7364 37100 7868 37156
rect 7924 37100 7934 37156
rect 9986 37100 9996 37156
rect 10052 37100 10062 37156
rect 15036 37100 19740 37156
rect 19796 37100 19806 37156
rect 0 37044 112 37072
rect 9996 37044 10052 37100
rect 0 36988 1820 37044
rect 1876 36988 1886 37044
rect 3126 36988 3164 37044
rect 3220 36988 3230 37044
rect 5506 36988 5516 37044
rect 5572 36988 5964 37044
rect 6020 36988 6030 37044
rect 7186 36988 7196 37044
rect 7252 36988 7532 37044
rect 7588 36988 9212 37044
rect 9268 36988 10052 37044
rect 10658 36988 10668 37044
rect 10724 36988 14812 37044
rect 14868 36988 14878 37044
rect 15250 36988 15260 37044
rect 15316 36988 15372 37044
rect 15428 36988 15438 37044
rect 21410 36988 21420 37044
rect 21476 36988 21486 37044
rect 0 36960 112 36988
rect 21420 36932 21476 36988
rect 10434 36876 10444 36932
rect 10500 36876 11004 36932
rect 11060 36876 11070 36932
rect 20178 36876 20188 36932
rect 20244 36876 21476 36932
rect 4454 36820 4464 36876
rect 4520 36820 4568 36876
rect 4624 36820 4672 36876
rect 4728 36820 4738 36876
rect 24454 36820 24464 36876
rect 24520 36820 24568 36876
rect 24624 36820 24672 36876
rect 24728 36820 24738 36876
rect 10770 36764 10780 36820
rect 10836 36764 11116 36820
rect 11172 36764 11182 36820
rect 11554 36764 11564 36820
rect 11620 36764 15036 36820
rect 15092 36764 15102 36820
rect 17490 36764 17500 36820
rect 17556 36764 18060 36820
rect 18116 36764 18126 36820
rect 4274 36652 4284 36708
rect 4340 36652 6636 36708
rect 6692 36652 7868 36708
rect 7924 36652 7934 36708
rect 9986 36652 9996 36708
rect 10052 36652 17948 36708
rect 18004 36652 29596 36708
rect 29652 36652 29662 36708
rect 0 36596 112 36624
rect 0 36540 6188 36596
rect 6244 36540 6254 36596
rect 7298 36540 7308 36596
rect 7364 36540 9772 36596
rect 9828 36540 9838 36596
rect 10658 36540 10668 36596
rect 10724 36540 11116 36596
rect 11172 36540 11182 36596
rect 11330 36540 11340 36596
rect 11396 36540 12684 36596
rect 12740 36540 12750 36596
rect 19170 36540 19180 36596
rect 19236 36540 19628 36596
rect 19684 36540 19694 36596
rect 23986 36540 23996 36596
rect 24052 36540 30268 36596
rect 30324 36540 30334 36596
rect 0 36512 112 36540
rect 1474 36428 1484 36484
rect 1540 36428 3388 36484
rect 3444 36428 3454 36484
rect 6402 36428 6412 36484
rect 6468 36428 8316 36484
rect 8372 36428 10332 36484
rect 10388 36428 12012 36484
rect 12068 36428 12078 36484
rect 13570 36428 13580 36484
rect 13636 36428 14364 36484
rect 14420 36428 14430 36484
rect 2258 36316 2268 36372
rect 2324 36316 2604 36372
rect 2660 36316 2670 36372
rect 8642 36316 8652 36372
rect 8708 36316 11116 36372
rect 11172 36316 11182 36372
rect 14578 36316 14588 36372
rect 14644 36316 15708 36372
rect 15764 36316 15774 36372
rect 16156 36316 20524 36372
rect 20580 36316 21308 36372
rect 21364 36316 21374 36372
rect 16156 36260 16212 36316
rect 11554 36204 11564 36260
rect 11620 36204 16212 36260
rect 18498 36204 18508 36260
rect 18564 36204 19292 36260
rect 19348 36204 19404 36260
rect 19460 36204 19470 36260
rect 0 36148 112 36176
rect 0 36092 3388 36148
rect 14242 36092 14252 36148
rect 14308 36092 17724 36148
rect 17780 36092 19964 36148
rect 20020 36092 20030 36148
rect 0 36064 112 36092
rect 3332 35924 3388 36092
rect 3794 36036 3804 36092
rect 3860 36036 3908 36092
rect 3964 36036 4012 36092
rect 4068 36036 4078 36092
rect 23794 36036 23804 36092
rect 23860 36036 23908 36092
rect 23964 36036 24012 36092
rect 24068 36036 24078 36092
rect 7522 35980 7532 36036
rect 7588 35980 13916 36036
rect 13972 35980 13982 36036
rect 14690 35980 14700 36036
rect 14756 35980 15036 36036
rect 15092 35980 15102 36036
rect 16930 35980 16940 36036
rect 16996 35980 17276 36036
rect 17332 35980 18284 36036
rect 18340 35980 19292 36036
rect 19348 35980 19358 36036
rect 3332 35868 7196 35924
rect 7252 35868 7262 35924
rect 10658 35868 10668 35924
rect 10724 35868 11228 35924
rect 11284 35868 11294 35924
rect 17490 35868 17500 35924
rect 17556 35868 17724 35924
rect 17780 35868 17790 35924
rect 20738 35868 20748 35924
rect 20804 35868 20814 35924
rect 20748 35812 20804 35868
rect 1138 35756 1148 35812
rect 1204 35756 3500 35812
rect 3556 35756 4508 35812
rect 4564 35756 4574 35812
rect 5170 35756 5180 35812
rect 5236 35756 12236 35812
rect 12292 35756 12302 35812
rect 17042 35756 17052 35812
rect 17108 35756 17612 35812
rect 17668 35756 17678 35812
rect 17826 35756 17836 35812
rect 17892 35756 18396 35812
rect 18452 35756 18462 35812
rect 20748 35756 20972 35812
rect 21028 35756 21038 35812
rect 0 35700 112 35728
rect 0 35644 3388 35700
rect 6178 35644 6188 35700
rect 6244 35644 12348 35700
rect 12404 35644 12414 35700
rect 16370 35644 16380 35700
rect 16436 35644 16828 35700
rect 16884 35644 16894 35700
rect 17154 35644 17164 35700
rect 17220 35644 19180 35700
rect 19236 35644 19246 35700
rect 21410 35644 21420 35700
rect 21476 35644 22428 35700
rect 22484 35644 22494 35700
rect 0 35616 112 35644
rect 3332 35588 3388 35644
rect 3332 35532 18228 35588
rect 18386 35532 18396 35588
rect 18452 35532 19740 35588
rect 19796 35532 19806 35588
rect 18172 35476 18228 35532
rect 6066 35420 6076 35476
rect 6132 35420 7420 35476
rect 7476 35420 8652 35476
rect 8708 35420 8718 35476
rect 9202 35420 9212 35476
rect 9268 35420 9436 35476
rect 9492 35420 9502 35476
rect 10182 35420 10220 35476
rect 10276 35420 10286 35476
rect 15026 35420 15036 35476
rect 15092 35420 15932 35476
rect 15988 35420 15998 35476
rect 16818 35420 16828 35476
rect 16884 35420 17500 35476
rect 17556 35420 17566 35476
rect 18172 35420 20748 35476
rect 20804 35420 20814 35476
rect 21970 35420 21980 35476
rect 22036 35420 25452 35476
rect 25508 35420 25518 35476
rect 2492 35308 3780 35364
rect 9650 35308 9660 35364
rect 9716 35308 11340 35364
rect 11396 35308 11406 35364
rect 11554 35308 11564 35364
rect 11620 35308 11788 35364
rect 11844 35308 11854 35364
rect 16034 35308 16044 35364
rect 16100 35308 17948 35364
rect 18004 35308 18732 35364
rect 18788 35308 18798 35364
rect 20178 35308 20188 35364
rect 20244 35308 20524 35364
rect 20580 35308 20590 35364
rect 0 35252 112 35280
rect 2492 35252 2548 35308
rect 0 35196 1036 35252
rect 1092 35196 1102 35252
rect 1362 35196 1372 35252
rect 1428 35196 2548 35252
rect 2706 35196 2716 35252
rect 2772 35196 3164 35252
rect 3220 35196 3230 35252
rect 0 35168 112 35196
rect 3724 35140 3780 35308
rect 4454 35252 4464 35308
rect 4520 35252 4568 35308
rect 4624 35252 4672 35308
rect 4728 35252 4738 35308
rect 24454 35252 24464 35308
rect 24520 35252 24568 35308
rect 24624 35252 24672 35308
rect 24728 35252 24738 35308
rect 31584 35252 31696 35280
rect 3938 35196 3948 35252
rect 4004 35196 4172 35252
rect 4228 35196 4238 35252
rect 4844 35196 16660 35252
rect 16818 35196 16828 35252
rect 16884 35196 17388 35252
rect 17444 35196 17454 35252
rect 18732 35196 20860 35252
rect 20916 35196 20926 35252
rect 30594 35196 30604 35252
rect 30660 35196 31696 35252
rect 4844 35140 4900 35196
rect 3724 35084 4900 35140
rect 5842 35084 5852 35140
rect 5908 35084 6188 35140
rect 6244 35084 6254 35140
rect 11106 35084 11116 35140
rect 11172 35084 13916 35140
rect 13972 35084 13982 35140
rect 14130 35084 14140 35140
rect 14196 35084 14700 35140
rect 14756 35084 15932 35140
rect 15988 35084 15998 35140
rect 16604 35028 16660 35196
rect 18732 35140 18788 35196
rect 31584 35168 31696 35196
rect 17714 35084 17724 35140
rect 17780 35084 18732 35140
rect 18788 35084 18798 35140
rect 20178 35084 20188 35140
rect 20244 35084 21196 35140
rect 21252 35084 21262 35140
rect 28018 35084 28028 35140
rect 28084 35084 30268 35140
rect 30324 35084 30334 35140
rect 1810 34972 1820 35028
rect 1876 34972 3388 35028
rect 3444 34972 3668 35028
rect 3938 34972 3948 35028
rect 4004 34972 4284 35028
rect 4340 34972 4350 35028
rect 6066 34972 6076 35028
rect 6132 34972 9100 35028
rect 9156 34972 9166 35028
rect 12450 34972 12460 35028
rect 12516 34972 13244 35028
rect 13300 34972 13310 35028
rect 13580 34972 14812 35028
rect 14868 34972 14878 35028
rect 16604 34972 17108 35028
rect 17826 34972 17836 35028
rect 17892 34972 18620 35028
rect 18676 34972 19404 35028
rect 19460 34972 19470 35028
rect 21858 34972 21868 35028
rect 21924 34972 24780 35028
rect 24836 34972 24846 35028
rect 3612 34916 3668 34972
rect 13580 34916 13636 34972
rect 3612 34860 4732 34916
rect 4788 34860 4798 34916
rect 5506 34860 5516 34916
rect 5572 34860 6188 34916
rect 6244 34860 6636 34916
rect 6692 34860 6702 34916
rect 7522 34860 7532 34916
rect 7588 34860 8092 34916
rect 8148 34860 8428 34916
rect 8484 34860 8494 34916
rect 9538 34860 9548 34916
rect 9604 34860 13636 34916
rect 13766 34860 13804 34916
rect 13860 34860 13870 34916
rect 0 34804 112 34832
rect 17052 34804 17108 34972
rect 17266 34860 17276 34916
rect 17332 34860 19068 34916
rect 19124 34860 19134 34916
rect 21186 34860 21196 34916
rect 21252 34860 22540 34916
rect 22596 34860 22606 34916
rect 23426 34860 23436 34916
rect 23492 34860 24668 34916
rect 24724 34860 24734 34916
rect 0 34748 1092 34804
rect 1698 34748 1708 34804
rect 1764 34748 3444 34804
rect 3602 34748 3612 34804
rect 3668 34748 3836 34804
rect 3892 34748 4900 34804
rect 5058 34748 5068 34804
rect 5124 34748 5292 34804
rect 5348 34748 5358 34804
rect 12450 34748 12460 34804
rect 12516 34748 12908 34804
rect 12964 34748 16604 34804
rect 16660 34748 16670 34804
rect 17052 34748 17612 34804
rect 17668 34748 18060 34804
rect 18116 34748 18126 34804
rect 0 34720 112 34748
rect 1036 34468 1092 34748
rect 3388 34692 3444 34748
rect 3388 34636 4172 34692
rect 4228 34636 4238 34692
rect 4844 34580 4900 34748
rect 5394 34636 5404 34692
rect 5460 34636 5852 34692
rect 5908 34636 5918 34692
rect 8530 34636 8540 34692
rect 8596 34636 9772 34692
rect 9828 34636 9838 34692
rect 16818 34636 16828 34692
rect 16884 34636 18956 34692
rect 19012 34636 19022 34692
rect 2034 34524 2044 34580
rect 2100 34524 3612 34580
rect 3668 34524 3678 34580
rect 4844 34524 11116 34580
rect 11172 34524 11182 34580
rect 12114 34524 12124 34580
rect 12180 34524 19068 34580
rect 19124 34524 22092 34580
rect 22148 34524 22158 34580
rect 3794 34468 3804 34524
rect 3860 34468 3908 34524
rect 3964 34468 4012 34524
rect 4068 34468 4078 34524
rect 23794 34468 23804 34524
rect 23860 34468 23908 34524
rect 23964 34468 24012 34524
rect 24068 34468 24078 34524
rect 1036 34412 3612 34468
rect 3668 34412 3678 34468
rect 7410 34412 7420 34468
rect 7476 34412 7532 34468
rect 7588 34412 7598 34468
rect 13794 34412 13804 34468
rect 13860 34412 16716 34468
rect 16772 34412 16782 34468
rect 20402 34412 20412 34468
rect 20468 34412 21476 34468
rect 0 34356 112 34384
rect 21420 34356 21476 34412
rect 31584 34356 31696 34384
rect 0 34300 6972 34356
rect 7028 34300 7038 34356
rect 7634 34300 7644 34356
rect 7700 34300 7868 34356
rect 7924 34300 7934 34356
rect 8978 34300 8988 34356
rect 9044 34300 9996 34356
rect 10052 34300 10062 34356
rect 10658 34300 10668 34356
rect 10724 34300 10780 34356
rect 10836 34300 10846 34356
rect 19842 34300 19852 34356
rect 19908 34300 21196 34356
rect 21252 34300 21262 34356
rect 21420 34300 30268 34356
rect 30324 34300 30334 34356
rect 30594 34300 30604 34356
rect 30660 34300 31696 34356
rect 0 34272 112 34300
rect 31584 34272 31696 34300
rect 2370 34188 2380 34244
rect 2436 34188 2940 34244
rect 2996 34188 3006 34244
rect 3164 34188 14924 34244
rect 14980 34188 14990 34244
rect 16790 34188 16828 34244
rect 16884 34188 16894 34244
rect 21410 34188 21420 34244
rect 21476 34188 22316 34244
rect 22372 34188 22382 34244
rect 3164 34132 3220 34188
rect 1250 34076 1260 34132
rect 1316 34076 3220 34132
rect 3332 34076 3500 34132
rect 3556 34076 3566 34132
rect 3714 34076 3724 34132
rect 3780 34076 5068 34132
rect 5124 34076 5134 34132
rect 5618 34076 5628 34132
rect 5684 34076 6412 34132
rect 6468 34076 6478 34132
rect 9874 34076 9884 34132
rect 9940 34076 10780 34132
rect 10836 34076 10846 34132
rect 11778 34076 11788 34132
rect 11844 34076 11900 34132
rect 11956 34076 11966 34132
rect 14130 34076 14140 34132
rect 14196 34076 14700 34132
rect 14756 34076 14766 34132
rect 16258 34076 16268 34132
rect 16324 34076 16492 34132
rect 16548 34076 16558 34132
rect 17154 34076 17164 34132
rect 17220 34076 17612 34132
rect 17668 34076 17678 34132
rect 17826 34076 17836 34132
rect 17892 34076 18172 34132
rect 18228 34076 18238 34132
rect 18806 34076 18844 34132
rect 18900 34076 18910 34132
rect 21970 34076 21980 34132
rect 22036 34076 25452 34132
rect 25508 34076 25518 34132
rect 3332 34020 3388 34076
rect 2258 33964 2268 34020
rect 2324 33964 3388 34020
rect 3612 33964 21700 34020
rect 21858 33964 21868 34020
rect 21924 33964 24668 34020
rect 24724 33964 24734 34020
rect 0 33908 112 33936
rect 3612 33908 3668 33964
rect 21644 33908 21700 33964
rect 0 33852 3668 33908
rect 4162 33852 4172 33908
rect 4228 33852 4956 33908
rect 5012 33852 5628 33908
rect 5684 33852 5694 33908
rect 9202 33852 9212 33908
rect 9268 33852 12796 33908
rect 12852 33852 14140 33908
rect 14196 33852 14206 33908
rect 15092 33852 15260 33908
rect 15316 33852 15326 33908
rect 19590 33852 19628 33908
rect 19684 33852 19694 33908
rect 21644 33852 22764 33908
rect 22820 33852 22830 33908
rect 0 33824 112 33852
rect 15092 33796 15148 33852
rect 1698 33740 1708 33796
rect 1764 33740 2044 33796
rect 2100 33740 2380 33796
rect 2436 33740 2446 33796
rect 2818 33740 2828 33796
rect 2884 33740 3948 33796
rect 4004 33740 4172 33796
rect 4228 33740 4238 33796
rect 9986 33740 9996 33796
rect 10052 33740 15148 33796
rect 18722 33740 18732 33796
rect 18788 33740 19740 33796
rect 19796 33740 19806 33796
rect 4454 33684 4464 33740
rect 4520 33684 4568 33740
rect 4624 33684 4672 33740
rect 4728 33684 4738 33740
rect 24454 33684 24464 33740
rect 24520 33684 24568 33740
rect 24624 33684 24672 33740
rect 24728 33684 24738 33740
rect 1362 33628 1372 33684
rect 1428 33628 2156 33684
rect 2212 33628 2222 33684
rect 11218 33628 11228 33684
rect 11284 33628 13692 33684
rect 13748 33628 13758 33684
rect 18050 33628 18060 33684
rect 18116 33628 18284 33684
rect 18340 33628 18350 33684
rect 19730 33628 19740 33684
rect 19796 33628 19806 33684
rect 21074 33628 21084 33684
rect 21140 33628 22652 33684
rect 22708 33628 22718 33684
rect 19740 33572 19796 33628
rect 4274 33516 4284 33572
rect 4340 33516 5516 33572
rect 5572 33516 5582 33572
rect 7970 33516 7980 33572
rect 8036 33516 8316 33572
rect 8372 33516 8382 33572
rect 19058 33516 19068 33572
rect 19124 33516 19292 33572
rect 19348 33516 19358 33572
rect 19740 33516 19852 33572
rect 19908 33516 19918 33572
rect 0 33460 112 33488
rect 31584 33460 31696 33488
rect 0 33404 1484 33460
rect 1540 33404 1550 33460
rect 2146 33404 2156 33460
rect 2212 33404 3612 33460
rect 3668 33404 3678 33460
rect 4060 33404 9660 33460
rect 9716 33404 9726 33460
rect 15698 33404 15708 33460
rect 15764 33404 18284 33460
rect 18340 33404 18350 33460
rect 18610 33404 18620 33460
rect 18676 33404 23772 33460
rect 23828 33404 23838 33460
rect 30706 33404 30716 33460
rect 30772 33404 31696 33460
rect 0 33376 112 33404
rect 4060 33348 4116 33404
rect 31584 33376 31696 33404
rect 3378 33292 3388 33348
rect 3444 33292 4116 33348
rect 4274 33292 4284 33348
rect 4340 33292 5068 33348
rect 5124 33292 5134 33348
rect 8082 33292 8092 33348
rect 8148 33292 8428 33348
rect 8484 33292 8494 33348
rect 10098 33292 10108 33348
rect 10164 33292 17052 33348
rect 17108 33292 17118 33348
rect 17714 33292 17724 33348
rect 17780 33292 18508 33348
rect 18564 33292 18574 33348
rect 19282 33292 19292 33348
rect 19348 33292 19516 33348
rect 19572 33292 19582 33348
rect 6402 33180 6412 33236
rect 6468 33180 7868 33236
rect 7924 33180 7934 33236
rect 16818 33180 16828 33236
rect 16884 33180 17500 33236
rect 17556 33180 17566 33236
rect 18050 33180 18060 33236
rect 18116 33180 19852 33236
rect 19908 33180 19918 33236
rect 3332 33068 7084 33124
rect 7140 33068 7150 33124
rect 8418 33068 8428 33124
rect 8484 33068 15148 33124
rect 15204 33068 16716 33124
rect 16772 33068 16782 33124
rect 17686 33068 17724 33124
rect 17780 33068 17790 33124
rect 18722 33068 18732 33124
rect 18788 33068 19180 33124
rect 19236 33068 20076 33124
rect 20132 33068 20142 33124
rect 0 33012 112 33040
rect 3332 33012 3388 33068
rect 0 32956 3388 33012
rect 8194 32956 8204 33012
rect 8260 32956 10332 33012
rect 10388 32956 10398 33012
rect 18946 32956 18956 33012
rect 19012 32956 21644 33012
rect 21700 32956 21710 33012
rect 0 32928 112 32956
rect 3794 32900 3804 32956
rect 3860 32900 3908 32956
rect 3964 32900 4012 32956
rect 4068 32900 4078 32956
rect 23794 32900 23804 32956
rect 23860 32900 23908 32956
rect 23964 32900 24012 32956
rect 24068 32900 24078 32956
rect 17490 32844 17500 32900
rect 17556 32844 20748 32900
rect 20804 32844 20814 32900
rect 25778 32844 25788 32900
rect 25844 32844 30380 32900
rect 30436 32844 30446 32900
rect 1138 32732 1148 32788
rect 1204 32732 1708 32788
rect 1764 32732 1774 32788
rect 6374 32732 6412 32788
rect 6468 32732 6478 32788
rect 7970 32732 7980 32788
rect 8036 32732 9212 32788
rect 9268 32732 9278 32788
rect 9874 32732 9884 32788
rect 9940 32732 10332 32788
rect 10388 32732 10398 32788
rect 10770 32732 10780 32788
rect 10836 32732 11452 32788
rect 11508 32732 13356 32788
rect 13412 32732 13422 32788
rect 14466 32732 14476 32788
rect 14532 32732 14700 32788
rect 14756 32732 14766 32788
rect 15138 32732 15148 32788
rect 15204 32732 23660 32788
rect 23716 32732 23726 32788
rect 3266 32620 3276 32676
rect 3332 32620 11004 32676
rect 11060 32620 11070 32676
rect 17276 32620 19292 32676
rect 19348 32620 19358 32676
rect 21074 32620 21084 32676
rect 21140 32620 29596 32676
rect 29652 32620 29662 32676
rect 0 32564 112 32592
rect 17276 32564 17332 32620
rect 31584 32564 31696 32592
rect 0 32508 11116 32564
rect 11172 32508 11182 32564
rect 14242 32508 14252 32564
rect 14308 32508 14924 32564
rect 14980 32508 14990 32564
rect 16370 32508 16380 32564
rect 16436 32508 16604 32564
rect 16660 32508 16670 32564
rect 17238 32508 17276 32564
rect 17332 32508 17342 32564
rect 18162 32508 18172 32564
rect 18228 32508 19852 32564
rect 19908 32508 19918 32564
rect 20290 32508 20300 32564
rect 20356 32508 20972 32564
rect 21028 32508 21038 32564
rect 30594 32508 30604 32564
rect 30660 32508 31696 32564
rect 0 32480 112 32508
rect 31584 32480 31696 32508
rect 2790 32396 2828 32452
rect 2884 32396 2894 32452
rect 5058 32396 5068 32452
rect 5124 32396 15148 32452
rect 15204 32396 15214 32452
rect 19702 32396 19740 32452
rect 19796 32396 21868 32452
rect 21924 32396 21934 32452
rect 3332 32284 5460 32340
rect 6850 32284 6860 32340
rect 6916 32284 6972 32340
rect 7028 32284 10780 32340
rect 10836 32284 10846 32340
rect 10994 32284 11004 32340
rect 11060 32284 11340 32340
rect 11396 32284 11406 32340
rect 14018 32284 14028 32340
rect 14084 32284 15596 32340
rect 15652 32284 15662 32340
rect 22306 32284 22316 32340
rect 22372 32284 22988 32340
rect 23044 32284 23054 32340
rect 1362 32172 1372 32228
rect 1428 32172 1820 32228
rect 1876 32172 1886 32228
rect 0 32116 112 32144
rect 3332 32116 3388 32284
rect 5404 32228 5460 32284
rect 5404 32172 18620 32228
rect 18676 32172 18686 32228
rect 4454 32116 4464 32172
rect 4520 32116 4568 32172
rect 4624 32116 4672 32172
rect 4728 32116 4738 32172
rect 24454 32116 24464 32172
rect 24520 32116 24568 32172
rect 24624 32116 24672 32172
rect 24728 32116 24738 32172
rect 0 32060 3388 32116
rect 7410 32060 7420 32116
rect 7476 32060 7868 32116
rect 7924 32060 7934 32116
rect 11666 32060 11676 32116
rect 11732 32060 16716 32116
rect 16772 32060 17948 32116
rect 18004 32060 18014 32116
rect 0 32032 112 32060
rect 6626 31948 6636 32004
rect 6692 31948 6748 32004
rect 6804 31948 6814 32004
rect 7186 31948 7196 32004
rect 7252 31948 9884 32004
rect 9940 31948 9950 32004
rect 10994 31948 11004 32004
rect 11060 31948 11564 32004
rect 11620 31948 11630 32004
rect 15596 31948 20188 32004
rect 20244 31948 20254 32004
rect 1698 31836 1708 31892
rect 1764 31836 2492 31892
rect 2548 31836 2558 31892
rect 2902 31836 2940 31892
rect 2996 31836 3006 31892
rect 4834 31836 4844 31892
rect 4900 31836 10220 31892
rect 10276 31836 10286 31892
rect 11330 31836 11340 31892
rect 11396 31836 11788 31892
rect 11844 31836 11854 31892
rect 13458 31836 13468 31892
rect 13524 31836 14812 31892
rect 14868 31836 14878 31892
rect 15596 31780 15652 31948
rect 19058 31836 19068 31892
rect 19124 31836 20860 31892
rect 20916 31836 20926 31892
rect 23202 31836 23212 31892
rect 23268 31836 24892 31892
rect 24948 31836 24958 31892
rect 2258 31724 2268 31780
rect 2324 31724 2716 31780
rect 2772 31724 3052 31780
rect 3108 31724 3118 31780
rect 4946 31724 4956 31780
rect 5012 31724 11900 31780
rect 11956 31724 15652 31780
rect 16146 31724 16156 31780
rect 16212 31724 17052 31780
rect 17108 31724 17118 31780
rect 17938 31724 17948 31780
rect 18004 31724 19292 31780
rect 19348 31724 19358 31780
rect 0 31668 112 31696
rect 31584 31668 31696 31696
rect 0 31612 252 31668
rect 308 31612 318 31668
rect 1810 31612 1820 31668
rect 1876 31612 1932 31668
rect 1988 31612 1998 31668
rect 2146 31612 2156 31668
rect 2212 31612 2940 31668
rect 2996 31612 3006 31668
rect 6738 31612 6748 31668
rect 6804 31612 8204 31668
rect 8260 31612 8270 31668
rect 9538 31612 9548 31668
rect 9604 31612 9996 31668
rect 10052 31612 10062 31668
rect 11218 31612 11228 31668
rect 11284 31612 15372 31668
rect 15428 31612 15932 31668
rect 15988 31612 15998 31668
rect 19618 31612 19628 31668
rect 19684 31612 20524 31668
rect 20580 31612 20590 31668
rect 30594 31612 30604 31668
rect 30660 31612 31696 31668
rect 0 31584 112 31612
rect 1932 31556 1988 31612
rect 31584 31584 31696 31612
rect 1932 31500 2716 31556
rect 2772 31500 2782 31556
rect 12002 31500 12012 31556
rect 12068 31500 12124 31556
rect 12180 31500 12190 31556
rect 13122 31500 13132 31556
rect 13188 31500 15708 31556
rect 15764 31500 15774 31556
rect 17042 31500 17052 31556
rect 17108 31500 19404 31556
rect 19460 31500 19470 31556
rect 11554 31388 11564 31444
rect 11620 31388 13692 31444
rect 13748 31388 13758 31444
rect 16146 31388 16156 31444
rect 16212 31388 18172 31444
rect 18228 31388 18844 31444
rect 18900 31388 18910 31444
rect 3794 31332 3804 31388
rect 3860 31332 3908 31388
rect 3964 31332 4012 31388
rect 4068 31332 4078 31388
rect 23794 31332 23804 31388
rect 23860 31332 23908 31388
rect 23964 31332 24012 31388
rect 24068 31332 24078 31388
rect 8754 31276 8764 31332
rect 8820 31276 16044 31332
rect 16100 31276 16110 31332
rect 0 31220 112 31248
rect 0 31164 7532 31220
rect 7588 31164 7598 31220
rect 15138 31164 15148 31220
rect 15204 31164 16940 31220
rect 16996 31164 17006 31220
rect 18470 31164 18508 31220
rect 18564 31164 18574 31220
rect 0 31136 112 31164
rect 2034 31052 2044 31108
rect 2100 31052 4956 31108
rect 5012 31052 5022 31108
rect 5394 31052 5404 31108
rect 5460 31052 6188 31108
rect 6244 31052 6254 31108
rect 7410 31052 7420 31108
rect 7476 31052 8652 31108
rect 8708 31052 9100 31108
rect 9156 31052 9166 31108
rect 17154 31052 17164 31108
rect 17220 31052 18620 31108
rect 18676 31052 18686 31108
rect 1698 30940 1708 30996
rect 1764 30940 2828 30996
rect 2884 30940 6748 30996
rect 6804 30940 7196 30996
rect 7252 30940 7262 30996
rect 10434 30940 10444 30996
rect 10500 30940 11564 30996
rect 11620 30940 11630 30996
rect 17042 30940 17052 30996
rect 17108 30940 17500 30996
rect 17556 30940 20076 30996
rect 20132 30940 20972 30996
rect 21028 30940 21038 30996
rect 3332 30828 11676 30884
rect 11732 30828 11742 30884
rect 12786 30828 12796 30884
rect 12852 30828 16044 30884
rect 16100 30828 16110 30884
rect 20514 30828 20524 30884
rect 20580 30828 30156 30884
rect 30212 30828 30222 30884
rect 0 30772 112 30800
rect 3332 30772 3388 30828
rect 31584 30772 31696 30800
rect 0 30716 3388 30772
rect 4284 30716 6076 30772
rect 6132 30716 6142 30772
rect 10658 30716 10668 30772
rect 10724 30716 11004 30772
rect 11060 30716 11070 30772
rect 15922 30716 15932 30772
rect 15988 30716 16380 30772
rect 16436 30716 16446 30772
rect 18834 30716 18844 30772
rect 18900 30716 20636 30772
rect 20692 30716 20702 30772
rect 21196 30716 29372 30772
rect 29428 30716 29438 30772
rect 30594 30716 30604 30772
rect 30660 30716 31696 30772
rect 0 30688 112 30716
rect 4284 30660 4340 30716
rect 21196 30660 21252 30716
rect 31584 30688 31696 30716
rect 3332 30604 4340 30660
rect 18844 30604 18956 30660
rect 19012 30604 21252 30660
rect 1586 30380 1596 30436
rect 1652 30380 2492 30436
rect 2548 30380 2558 30436
rect 0 30324 112 30352
rect 3332 30324 3388 30604
rect 4454 30548 4464 30604
rect 4520 30548 4568 30604
rect 4624 30548 4672 30604
rect 4728 30548 4738 30604
rect 18844 30548 18900 30604
rect 24454 30548 24464 30604
rect 24520 30548 24568 30604
rect 24624 30548 24672 30604
rect 24728 30548 24738 30604
rect 18834 30492 18844 30548
rect 18900 30492 18910 30548
rect 20066 30492 20076 30548
rect 20132 30492 21868 30548
rect 21924 30492 21934 30548
rect 3602 30380 3612 30436
rect 3668 30380 5068 30436
rect 5124 30380 5134 30436
rect 7074 30380 7084 30436
rect 7140 30380 10780 30436
rect 10836 30380 13468 30436
rect 13524 30380 13534 30436
rect 16258 30380 16268 30436
rect 16324 30380 16604 30436
rect 16660 30380 16670 30436
rect 17826 30380 17836 30436
rect 17892 30380 20300 30436
rect 20356 30380 20366 30436
rect 0 30268 3388 30324
rect 3500 30268 6524 30324
rect 6580 30268 6590 30324
rect 7298 30268 7308 30324
rect 7364 30268 7980 30324
rect 8036 30268 8046 30324
rect 8978 30268 8988 30324
rect 9044 30268 9772 30324
rect 9828 30268 10444 30324
rect 10500 30268 10510 30324
rect 15026 30268 15036 30324
rect 15092 30268 15708 30324
rect 15764 30268 15774 30324
rect 16034 30268 16044 30324
rect 16100 30268 17052 30324
rect 17108 30268 17118 30324
rect 0 30240 112 30268
rect 3500 30100 3556 30268
rect 4162 30156 4172 30212
rect 4228 30156 4956 30212
rect 5012 30156 5740 30212
rect 5796 30156 5806 30212
rect 6626 30156 6636 30212
rect 6692 30156 7532 30212
rect 7588 30156 7598 30212
rect 14242 30156 14252 30212
rect 14308 30156 14812 30212
rect 14868 30156 14878 30212
rect 15092 30156 17276 30212
rect 17332 30156 17342 30212
rect 17826 30156 17836 30212
rect 17892 30156 18060 30212
rect 18116 30156 21420 30212
rect 21476 30156 21486 30212
rect 26002 30156 26012 30212
rect 26068 30156 30268 30212
rect 30324 30156 30334 30212
rect 15092 30100 15148 30156
rect 2482 30044 2492 30100
rect 2548 30044 3556 30100
rect 3612 30044 9324 30100
rect 9380 30044 9390 30100
rect 12450 30044 12460 30100
rect 12516 30044 15148 30100
rect 18386 30044 18396 30100
rect 18452 30044 19068 30100
rect 19124 30044 19628 30100
rect 19684 30044 19694 30100
rect 2034 29932 2044 29988
rect 2100 29932 3388 29988
rect 3444 29932 3454 29988
rect 0 29876 112 29904
rect 3612 29876 3668 30044
rect 19852 29988 19908 30156
rect 8194 29932 8204 29988
rect 8260 29932 8652 29988
rect 8708 29932 8718 29988
rect 11330 29932 11340 29988
rect 11396 29932 13468 29988
rect 13524 29932 13534 29988
rect 17266 29932 17276 29988
rect 17332 29932 17388 29988
rect 17444 29932 17454 29988
rect 17602 29932 17612 29988
rect 17668 29932 18284 29988
rect 18340 29932 19516 29988
rect 19572 29932 19582 29988
rect 19852 29932 19964 29988
rect 20020 29932 20030 29988
rect 31584 29876 31696 29904
rect 0 29820 3668 29876
rect 30594 29820 30604 29876
rect 30660 29820 31696 29876
rect 0 29792 112 29820
rect 3794 29764 3804 29820
rect 3860 29764 3908 29820
rect 3964 29764 4012 29820
rect 4068 29764 4078 29820
rect 23794 29764 23804 29820
rect 23860 29764 23908 29820
rect 23964 29764 24012 29820
rect 24068 29764 24078 29820
rect 31584 29792 31696 29820
rect 10546 29708 10556 29764
rect 10612 29708 11116 29764
rect 11172 29708 11182 29764
rect 15092 29708 18844 29764
rect 18900 29708 18910 29764
rect 15092 29652 15148 29708
rect 354 29596 364 29652
rect 420 29596 15148 29652
rect 16604 29596 17388 29652
rect 17444 29596 17454 29652
rect 2482 29484 2492 29540
rect 2548 29484 2716 29540
rect 2772 29484 2782 29540
rect 10332 29484 11340 29540
rect 11396 29484 11406 29540
rect 0 29428 112 29456
rect 10332 29428 10388 29484
rect 0 29372 10388 29428
rect 10546 29372 10556 29428
rect 10612 29372 11452 29428
rect 11508 29372 13020 29428
rect 13076 29372 13580 29428
rect 13636 29372 14028 29428
rect 14084 29372 14364 29428
rect 14420 29372 14430 29428
rect 0 29344 112 29372
rect 16604 29316 16660 29596
rect 16790 29484 16828 29540
rect 16884 29484 16894 29540
rect 18722 29484 18732 29540
rect 18788 29484 21308 29540
rect 21364 29484 21374 29540
rect 16930 29372 16940 29428
rect 16996 29372 17388 29428
rect 17444 29372 17612 29428
rect 17668 29372 17678 29428
rect 18806 29372 18844 29428
rect 18900 29372 18910 29428
rect 19506 29372 19516 29428
rect 19572 29372 20636 29428
rect 20692 29372 20702 29428
rect 21634 29372 21644 29428
rect 21700 29372 22204 29428
rect 22260 29372 22270 29428
rect 2230 29260 2268 29316
rect 2324 29260 2334 29316
rect 3332 29260 5404 29316
rect 5460 29260 5470 29316
rect 5842 29260 5852 29316
rect 5908 29260 6188 29316
rect 6244 29260 6254 29316
rect 7634 29260 7644 29316
rect 7700 29260 8428 29316
rect 8484 29260 8494 29316
rect 9538 29260 9548 29316
rect 9604 29260 11004 29316
rect 11060 29260 11116 29316
rect 11172 29260 11182 29316
rect 15092 29260 16660 29316
rect 17714 29260 17724 29316
rect 17780 29260 21532 29316
rect 21588 29260 21598 29316
rect 3332 29204 3388 29260
rect 15092 29204 15148 29260
rect 1810 29148 1820 29204
rect 1876 29148 3388 29204
rect 4284 29148 15148 29204
rect 23212 29148 29148 29204
rect 29204 29148 29214 29204
rect 0 28980 112 29008
rect 4284 28980 4340 29148
rect 23212 29092 23268 29148
rect 8194 29036 8204 29092
rect 8260 29036 21308 29092
rect 21364 29036 23212 29092
rect 23268 29036 23278 29092
rect 4454 28980 4464 29036
rect 4520 28980 4568 29036
rect 4624 28980 4672 29036
rect 4728 28980 4738 29036
rect 24454 28980 24464 29036
rect 24520 28980 24568 29036
rect 24624 28980 24672 29036
rect 24728 28980 24738 29036
rect 31584 28980 31696 29008
rect 0 28924 4340 28980
rect 30594 28924 30604 28980
rect 30660 28924 31696 28980
rect 0 28896 112 28924
rect 31584 28896 31696 28924
rect 1474 28812 1484 28868
rect 1540 28812 2156 28868
rect 2212 28812 2268 28868
rect 2324 28812 2334 28868
rect 6290 28812 6300 28868
rect 6356 28812 7532 28868
rect 7588 28812 7598 28868
rect 13794 28812 13804 28868
rect 13860 28812 14364 28868
rect 14420 28812 14924 28868
rect 14980 28812 15708 28868
rect 15764 28812 15774 28868
rect 17826 28812 17836 28868
rect 17892 28812 18060 28868
rect 18116 28812 18620 28868
rect 18676 28812 18686 28868
rect 19842 28812 19852 28868
rect 19908 28812 20300 28868
rect 20356 28812 20366 28868
rect 6962 28700 6972 28756
rect 7028 28700 8428 28756
rect 8484 28700 8988 28756
rect 9044 28700 9054 28756
rect 9874 28700 9884 28756
rect 9940 28700 10108 28756
rect 10164 28700 10174 28756
rect 13906 28700 13916 28756
rect 13972 28700 17612 28756
rect 17668 28700 17678 28756
rect 18834 28700 18844 28756
rect 18900 28700 30268 28756
rect 30324 28700 30334 28756
rect 1250 28588 1260 28644
rect 1316 28588 1708 28644
rect 1764 28588 1774 28644
rect 8642 28588 8652 28644
rect 8708 28588 10220 28644
rect 10276 28588 10286 28644
rect 12114 28588 12124 28644
rect 12180 28588 13244 28644
rect 13300 28588 14700 28644
rect 14756 28588 14766 28644
rect 18386 28588 18396 28644
rect 18452 28588 19012 28644
rect 19842 28588 19852 28644
rect 19908 28588 20076 28644
rect 20132 28588 20142 28644
rect 0 28532 112 28560
rect 18956 28532 19012 28588
rect 0 28476 3388 28532
rect 11330 28476 11340 28532
rect 11396 28476 15036 28532
rect 15092 28476 18508 28532
rect 18564 28476 18574 28532
rect 18956 28476 19068 28532
rect 19124 28476 20860 28532
rect 20916 28476 20926 28532
rect 0 28448 112 28476
rect 3332 28420 3388 28476
rect 3332 28364 16156 28420
rect 16212 28364 17276 28420
rect 17332 28364 20076 28420
rect 20132 28364 20142 28420
rect 5618 28252 5628 28308
rect 5684 28252 7868 28308
rect 7924 28252 7934 28308
rect 9090 28252 9100 28308
rect 9156 28252 9772 28308
rect 9828 28252 13916 28308
rect 13972 28252 13982 28308
rect 3794 28196 3804 28252
rect 3860 28196 3908 28252
rect 3964 28196 4012 28252
rect 4068 28196 4078 28252
rect 23794 28196 23804 28252
rect 23860 28196 23908 28252
rect 23964 28196 24012 28252
rect 24068 28196 24078 28252
rect 9090 28140 9100 28196
rect 9156 28140 18172 28196
rect 18228 28140 18238 28196
rect 0 28084 112 28112
rect 31584 28084 31696 28112
rect 0 28028 3388 28084
rect 10322 28028 10332 28084
rect 10388 28028 11228 28084
rect 11284 28028 11294 28084
rect 11554 28028 11564 28084
rect 11620 28028 16828 28084
rect 16884 28028 16894 28084
rect 19170 28028 19180 28084
rect 19236 28028 19516 28084
rect 19572 28028 19964 28084
rect 20020 28028 20030 28084
rect 20626 28028 20636 28084
rect 20692 28028 21868 28084
rect 21924 28028 22540 28084
rect 22596 28028 22606 28084
rect 30594 28028 30604 28084
rect 30660 28028 31696 28084
rect 0 28000 112 28028
rect 3332 27972 3388 28028
rect 31584 28000 31696 28028
rect 1138 27916 1148 27972
rect 1204 27916 1484 27972
rect 1540 27916 1820 27972
rect 1876 27916 1886 27972
rect 3332 27916 8540 27972
rect 8596 27916 17388 27972
rect 17444 27916 17454 27972
rect 21970 27916 21980 27972
rect 22036 27916 22428 27972
rect 22484 27916 22494 27972
rect 28130 27916 28140 27972
rect 28196 27916 30268 27972
rect 30324 27916 30334 27972
rect 3266 27804 3276 27860
rect 3332 27804 3612 27860
rect 3668 27804 3678 27860
rect 3938 27804 3948 27860
rect 4004 27804 8372 27860
rect 10546 27804 10556 27860
rect 10612 27804 10892 27860
rect 10948 27804 10958 27860
rect 11890 27804 11900 27860
rect 11956 27804 12684 27860
rect 12740 27804 12750 27860
rect 21074 27804 21084 27860
rect 21140 27804 29596 27860
rect 29652 27804 29662 27860
rect 8316 27748 8372 27804
rect 1922 27692 1932 27748
rect 1988 27692 2492 27748
rect 2548 27692 2558 27748
rect 6626 27692 6636 27748
rect 6692 27692 7084 27748
rect 7140 27692 7150 27748
rect 8306 27692 8316 27748
rect 8372 27692 13580 27748
rect 13636 27692 13646 27748
rect 18694 27692 18732 27748
rect 18788 27692 18798 27748
rect 19814 27692 19852 27748
rect 19908 27692 19918 27748
rect 29698 27692 29708 27748
rect 29764 27692 31500 27748
rect 31556 27692 31566 27748
rect 0 27636 112 27664
rect 0 27580 8932 27636
rect 9202 27580 9212 27636
rect 9268 27580 10332 27636
rect 10388 27580 10398 27636
rect 15250 27580 15260 27636
rect 15316 27580 16156 27636
rect 16212 27580 16222 27636
rect 18732 27580 19292 27636
rect 19348 27580 19358 27636
rect 0 27552 112 27580
rect 8876 27524 8932 27580
rect 18732 27524 18788 27580
rect 8876 27468 11452 27524
rect 11508 27468 11518 27524
rect 18722 27468 18732 27524
rect 18788 27468 18798 27524
rect 4454 27412 4464 27468
rect 4520 27412 4568 27468
rect 4624 27412 4672 27468
rect 4728 27412 4738 27468
rect 24454 27412 24464 27468
rect 24520 27412 24568 27468
rect 24624 27412 24672 27468
rect 24728 27412 24738 27468
rect 2146 27356 2156 27412
rect 2212 27356 2380 27412
rect 2436 27356 2446 27412
rect 14130 27356 14140 27412
rect 14196 27356 20300 27412
rect 20356 27356 20524 27412
rect 20580 27356 20590 27412
rect 3714 27244 3724 27300
rect 3780 27244 6748 27300
rect 6804 27244 6814 27300
rect 9090 27244 9100 27300
rect 9156 27244 9772 27300
rect 9828 27244 9838 27300
rect 13010 27244 13020 27300
rect 13076 27244 13132 27300
rect 13188 27244 14252 27300
rect 14308 27244 17052 27300
rect 17108 27244 17118 27300
rect 18610 27244 18620 27300
rect 18676 27244 19292 27300
rect 19348 27244 19358 27300
rect 20066 27244 20076 27300
rect 20132 27244 21084 27300
rect 21140 27244 21150 27300
rect 0 27188 112 27216
rect 31584 27188 31696 27216
rect 0 27132 9100 27188
rect 9156 27132 9166 27188
rect 9874 27132 9884 27188
rect 9940 27132 11676 27188
rect 11732 27132 11742 27188
rect 15138 27132 15148 27188
rect 15204 27132 16940 27188
rect 16996 27132 17006 27188
rect 30706 27132 30716 27188
rect 30772 27132 31696 27188
rect 0 27104 112 27132
rect 31584 27104 31696 27132
rect 2594 27020 2604 27076
rect 2660 27020 3948 27076
rect 4004 27020 4014 27076
rect 4162 27020 4172 27076
rect 4228 27020 4508 27076
rect 4564 27020 4574 27076
rect 7746 27020 7756 27076
rect 7812 27020 9212 27076
rect 9268 27020 10444 27076
rect 10500 27020 10510 27076
rect 10882 27020 10892 27076
rect 10948 27020 12572 27076
rect 12628 27020 15260 27076
rect 15316 27020 15326 27076
rect 16258 27020 16268 27076
rect 16324 27020 16828 27076
rect 16884 27020 16894 27076
rect 18834 27020 18844 27076
rect 18900 27020 19180 27076
rect 19236 27020 19246 27076
rect 2482 26908 2492 26964
rect 2548 26908 6860 26964
rect 6916 26908 6926 26964
rect 7522 26908 7532 26964
rect 7588 26908 12684 26964
rect 12740 26908 12750 26964
rect 14690 26908 14700 26964
rect 14756 26908 15708 26964
rect 15764 26908 15774 26964
rect 18162 26908 18172 26964
rect 18228 26908 19124 26964
rect 19506 26908 19516 26964
rect 19572 26908 19628 26964
rect 19684 26908 19694 26964
rect 21298 26908 21308 26964
rect 21364 26908 21756 26964
rect 21812 26908 22204 26964
rect 22260 26908 22270 26964
rect 19068 26852 19124 26908
rect 3332 26796 5180 26852
rect 5236 26796 5246 26852
rect 8866 26796 8876 26852
rect 8932 26796 13916 26852
rect 13972 26796 16156 26852
rect 16212 26796 16222 26852
rect 17938 26796 17948 26852
rect 18004 26796 18620 26852
rect 18676 26796 18686 26852
rect 19058 26796 19068 26852
rect 19124 26796 19134 26852
rect 20738 26796 20748 26852
rect 20804 26796 28028 26852
rect 28084 26796 28094 26852
rect 0 26740 112 26768
rect 3332 26740 3388 26796
rect 0 26684 3388 26740
rect 9538 26684 9548 26740
rect 9604 26684 16716 26740
rect 16772 26684 16782 26740
rect 0 26656 112 26684
rect 3794 26628 3804 26684
rect 3860 26628 3908 26684
rect 3964 26628 4012 26684
rect 4068 26628 4078 26684
rect 23794 26628 23804 26684
rect 23860 26628 23908 26684
rect 23964 26628 24012 26684
rect 24068 26628 24078 26684
rect 6962 26572 6972 26628
rect 7028 26572 7420 26628
rect 7476 26572 7486 26628
rect 10210 26572 10220 26628
rect 10276 26572 11228 26628
rect 11284 26572 11294 26628
rect 1698 26460 1708 26516
rect 1764 26460 1932 26516
rect 1988 26460 1998 26516
rect 3602 26460 3612 26516
rect 3668 26460 4844 26516
rect 4900 26460 4910 26516
rect 6178 26460 6188 26516
rect 6244 26460 18732 26516
rect 18788 26460 18798 26516
rect 20738 26460 20748 26516
rect 20804 26460 21644 26516
rect 21700 26460 21710 26516
rect 4162 26348 4172 26404
rect 4228 26348 12124 26404
rect 12180 26348 12190 26404
rect 18274 26348 18284 26404
rect 18340 26348 20188 26404
rect 20244 26348 20254 26404
rect 0 26292 112 26320
rect 31584 26292 31696 26320
rect 0 26236 364 26292
rect 420 26236 430 26292
rect 1922 26236 1932 26292
rect 1988 26236 6972 26292
rect 7028 26236 7038 26292
rect 8306 26236 8316 26292
rect 8372 26236 9100 26292
rect 9156 26236 9166 26292
rect 9538 26236 9548 26292
rect 9604 26236 9884 26292
rect 9940 26236 11564 26292
rect 11620 26236 11630 26292
rect 11890 26236 11900 26292
rect 11956 26236 12460 26292
rect 12516 26236 12526 26292
rect 14018 26236 14028 26292
rect 14084 26236 14476 26292
rect 14532 26236 14542 26292
rect 15250 26236 15260 26292
rect 15316 26236 15820 26292
rect 15876 26236 15886 26292
rect 16342 26236 16380 26292
rect 16436 26236 16446 26292
rect 17154 26236 17164 26292
rect 17220 26236 17724 26292
rect 17780 26236 17790 26292
rect 20290 26236 20300 26292
rect 20356 26236 22316 26292
rect 22372 26236 22382 26292
rect 30594 26236 30604 26292
rect 30660 26236 31696 26292
rect 0 26208 112 26236
rect 31584 26208 31696 26236
rect 1586 26124 1596 26180
rect 1652 26124 17500 26180
rect 17556 26124 20748 26180
rect 20804 26124 20814 26180
rect 3154 26012 3164 26068
rect 3220 26012 3500 26068
rect 3556 26012 3566 26068
rect 8082 26012 8092 26068
rect 8148 26012 9772 26068
rect 9828 26012 9838 26068
rect 14998 26012 15036 26068
rect 15092 26012 15102 26068
rect 15810 26012 15820 26068
rect 15876 26012 16604 26068
rect 16660 26012 18060 26068
rect 18116 26012 18126 26068
rect 3332 25900 3612 25956
rect 3668 25900 3678 25956
rect 6514 25900 6524 25956
rect 6580 25900 6748 25956
rect 6804 25900 6814 25956
rect 7186 25900 7196 25956
rect 7252 25900 9660 25956
rect 9716 25900 9726 25956
rect 9986 25900 9996 25956
rect 10052 25900 21868 25956
rect 21924 25900 21934 25956
rect 0 25844 112 25872
rect 3332 25844 3388 25900
rect 4454 25844 4464 25900
rect 4520 25844 4568 25900
rect 4624 25844 4672 25900
rect 4728 25844 4738 25900
rect 24454 25844 24464 25900
rect 24520 25844 24568 25900
rect 24624 25844 24672 25900
rect 24728 25844 24738 25900
rect 0 25788 3388 25844
rect 11890 25788 11900 25844
rect 11956 25788 12908 25844
rect 12964 25788 12974 25844
rect 13906 25788 13916 25844
rect 13972 25788 14924 25844
rect 14980 25788 15596 25844
rect 15652 25788 15662 25844
rect 0 25760 112 25788
rect 3714 25676 3724 25732
rect 3780 25676 4508 25732
rect 4564 25676 4574 25732
rect 5282 25676 5292 25732
rect 5348 25676 5628 25732
rect 5684 25676 5694 25732
rect 5842 25676 5852 25732
rect 5908 25676 9996 25732
rect 10052 25676 10062 25732
rect 14018 25676 14028 25732
rect 14084 25676 17948 25732
rect 18004 25676 18014 25732
rect 20066 25676 20076 25732
rect 20132 25676 30268 25732
rect 30324 25676 30334 25732
rect 4172 25564 4956 25620
rect 5012 25564 5022 25620
rect 5170 25564 5180 25620
rect 5236 25564 5404 25620
rect 5460 25564 5470 25620
rect 5730 25564 5740 25620
rect 5796 25564 8988 25620
rect 9044 25564 9884 25620
rect 9940 25564 9950 25620
rect 12898 25564 12908 25620
rect 12964 25564 15484 25620
rect 15540 25564 15550 25620
rect 4172 25508 4228 25564
rect 2146 25452 2156 25508
rect 2212 25452 4172 25508
rect 4228 25452 4238 25508
rect 4498 25452 4508 25508
rect 4564 25452 5628 25508
rect 5684 25452 5694 25508
rect 6626 25452 6636 25508
rect 6692 25452 9100 25508
rect 9156 25452 10612 25508
rect 11554 25452 11564 25508
rect 11620 25452 14924 25508
rect 14980 25452 14990 25508
rect 15698 25452 15708 25508
rect 15764 25452 17388 25508
rect 17444 25452 17454 25508
rect 21858 25452 21868 25508
rect 21924 25452 22092 25508
rect 22148 25452 22540 25508
rect 22596 25452 22606 25508
rect 0 25396 112 25424
rect 10556 25396 10612 25452
rect 31584 25396 31696 25424
rect 0 25340 9548 25396
rect 9604 25340 9614 25396
rect 10546 25340 10556 25396
rect 10612 25340 18620 25396
rect 18676 25340 20300 25396
rect 20356 25340 20366 25396
rect 30594 25340 30604 25396
rect 30660 25340 31696 25396
rect 0 25312 112 25340
rect 31584 25312 31696 25340
rect 1138 25228 1148 25284
rect 1204 25228 1820 25284
rect 1876 25228 1886 25284
rect 3154 25228 3164 25284
rect 3220 25228 3444 25284
rect 3602 25228 3612 25284
rect 3668 25228 5292 25284
rect 5348 25228 5358 25284
rect 5516 25228 5852 25284
rect 5908 25228 5918 25284
rect 8530 25228 8540 25284
rect 8596 25228 12572 25284
rect 12628 25228 12638 25284
rect 14914 25228 14924 25284
rect 14980 25228 15932 25284
rect 15988 25228 15998 25284
rect 16342 25228 16380 25284
rect 16436 25228 16446 25284
rect 18946 25228 18956 25284
rect 19012 25228 19516 25284
rect 19572 25228 22764 25284
rect 22820 25228 22830 25284
rect 3388 25172 3444 25228
rect 5516 25172 5572 25228
rect 3388 25116 3668 25172
rect 4274 25116 4284 25172
rect 4340 25116 4350 25172
rect 5170 25116 5180 25172
rect 5236 25116 5572 25172
rect 5628 25116 8316 25172
rect 8372 25116 8382 25172
rect 8642 25116 8652 25172
rect 8708 25116 9548 25172
rect 9604 25116 9614 25172
rect 12002 25116 12012 25172
rect 12068 25116 12236 25172
rect 12292 25116 12302 25172
rect 16230 25116 16268 25172
rect 16324 25116 16334 25172
rect 3612 25060 3668 25116
rect 3794 25060 3804 25116
rect 3860 25060 3908 25116
rect 3964 25060 4012 25116
rect 4068 25060 4078 25116
rect 4284 25060 4340 25116
rect 5628 25060 5684 25116
rect 23794 25060 23804 25116
rect 23860 25060 23908 25116
rect 23964 25060 24012 25116
rect 24068 25060 24078 25116
rect 3602 25004 3612 25060
rect 3668 25004 3678 25060
rect 4162 25004 4172 25060
rect 4228 25004 5684 25060
rect 6524 25004 14252 25060
rect 14308 25004 14318 25060
rect 29474 25004 29484 25060
rect 29540 25004 30492 25060
rect 30548 25004 30558 25060
rect 0 24948 112 24976
rect 6524 24948 6580 25004
rect 0 24892 6580 24948
rect 6738 24892 6748 24948
rect 6804 24892 7980 24948
rect 8036 24892 8046 24948
rect 10098 24892 10108 24948
rect 10164 24892 10892 24948
rect 10948 24892 10958 24948
rect 16146 24892 16156 24948
rect 16212 24892 17164 24948
rect 17220 24892 17230 24948
rect 0 24864 112 24892
rect 13010 24780 13020 24836
rect 13076 24780 14140 24836
rect 14196 24780 14206 24836
rect 20850 24780 20860 24836
rect 20916 24780 21644 24836
rect 21700 24780 21710 24836
rect 1250 24668 1260 24724
rect 1316 24668 1708 24724
rect 1764 24668 1774 24724
rect 7522 24668 7532 24724
rect 7588 24668 9324 24724
rect 9380 24668 9390 24724
rect 14466 24668 14476 24724
rect 14532 24668 17276 24724
rect 17332 24668 17724 24724
rect 17780 24668 17790 24724
rect 28354 24668 28364 24724
rect 28420 24668 30268 24724
rect 30324 24668 30334 24724
rect 3490 24556 3500 24612
rect 3556 24556 3612 24612
rect 3668 24556 3678 24612
rect 7298 24556 7308 24612
rect 7364 24556 8988 24612
rect 9044 24556 9054 24612
rect 10658 24556 10668 24612
rect 10724 24556 10780 24612
rect 10836 24556 10846 24612
rect 16678 24556 16716 24612
rect 16772 24556 17948 24612
rect 18004 24556 18014 24612
rect 0 24500 112 24528
rect 31584 24500 31696 24528
rect 0 24444 11788 24500
rect 11844 24444 12684 24500
rect 12740 24444 12750 24500
rect 30594 24444 30604 24500
rect 30660 24444 31696 24500
rect 0 24416 112 24444
rect 31584 24416 31696 24444
rect 7410 24332 7420 24388
rect 7476 24332 13356 24388
rect 13412 24332 18060 24388
rect 18116 24332 18126 24388
rect 4454 24276 4464 24332
rect 4520 24276 4568 24332
rect 4624 24276 4672 24332
rect 4728 24276 4738 24332
rect 24454 24276 24464 24332
rect 24520 24276 24568 24332
rect 24624 24276 24672 24332
rect 24728 24276 24738 24332
rect 2370 24220 2380 24276
rect 2436 24220 2716 24276
rect 2772 24220 4172 24276
rect 4228 24220 4238 24276
rect 9538 24220 9548 24276
rect 9604 24220 15148 24276
rect 21634 24220 21644 24276
rect 21700 24220 21710 24276
rect 15092 24164 15148 24220
rect 21644 24164 21700 24220
rect 2258 24108 2268 24164
rect 2324 24108 3388 24164
rect 3444 24108 3454 24164
rect 6850 24108 6860 24164
rect 6916 24108 7420 24164
rect 7476 24108 7486 24164
rect 12114 24108 12124 24164
rect 12180 24108 12572 24164
rect 12628 24108 12638 24164
rect 15092 24108 21700 24164
rect 0 24052 112 24080
rect 0 23996 140 24052
rect 196 23996 206 24052
rect 2930 23996 2940 24052
rect 2996 23996 3052 24052
rect 3108 23996 3118 24052
rect 3388 23996 11900 24052
rect 11956 23996 12908 24052
rect 12964 23996 12974 24052
rect 14774 23996 14812 24052
rect 14868 23996 14878 24052
rect 15362 23996 15372 24052
rect 15428 23996 30268 24052
rect 30324 23996 30334 24052
rect 0 23968 112 23996
rect 3388 23940 3444 23996
rect 242 23884 252 23940
rect 308 23884 3444 23940
rect 4162 23884 4172 23940
rect 4228 23884 4956 23940
rect 5012 23884 5022 23940
rect 5730 23884 5740 23940
rect 5796 23884 6188 23940
rect 6244 23884 6254 23940
rect 10444 23884 14140 23940
rect 14196 23884 18396 23940
rect 18452 23884 18462 23940
rect 10444 23828 10500 23884
rect 1810 23772 1820 23828
rect 1876 23772 1932 23828
rect 1988 23772 1998 23828
rect 4050 23772 4060 23828
rect 4116 23772 4396 23828
rect 4452 23772 4462 23828
rect 5170 23772 5180 23828
rect 5236 23772 5852 23828
rect 5908 23772 10444 23828
rect 10500 23772 10510 23828
rect 20402 23772 20412 23828
rect 20468 23772 21756 23828
rect 21812 23772 21822 23828
rect 1250 23660 1260 23716
rect 1316 23660 2716 23716
rect 2772 23660 2782 23716
rect 3332 23660 17164 23716
rect 17220 23660 18172 23716
rect 18228 23660 20300 23716
rect 20356 23660 20366 23716
rect 0 23604 112 23632
rect 3332 23604 3388 23660
rect 31584 23604 31696 23632
rect 0 23548 3388 23604
rect 4162 23548 4172 23604
rect 4228 23548 7420 23604
rect 7476 23548 7486 23604
rect 7634 23548 7644 23604
rect 7700 23548 7980 23604
rect 8036 23548 8046 23604
rect 17714 23548 17724 23604
rect 17780 23548 19404 23604
rect 19460 23548 21644 23604
rect 21700 23548 21710 23604
rect 23202 23548 23212 23604
rect 23268 23548 23278 23604
rect 30594 23548 30604 23604
rect 30660 23548 31696 23604
rect 0 23520 112 23548
rect 3794 23492 3804 23548
rect 3860 23492 3908 23548
rect 3964 23492 4012 23548
rect 4068 23492 4078 23548
rect 23212 23492 23268 23548
rect 23794 23492 23804 23548
rect 23860 23492 23908 23548
rect 23964 23492 24012 23548
rect 24068 23492 24078 23548
rect 31584 23520 31696 23548
rect 12674 23436 12684 23492
rect 12740 23436 12796 23492
rect 12852 23436 14756 23492
rect 14886 23436 14924 23492
rect 14980 23436 14990 23492
rect 15250 23436 15260 23492
rect 15316 23436 18732 23492
rect 18788 23436 18798 23492
rect 20066 23436 20076 23492
rect 20132 23436 20524 23492
rect 20580 23436 20590 23492
rect 23090 23436 23100 23492
rect 23156 23436 23268 23492
rect 14700 23380 14756 23436
rect 802 23324 812 23380
rect 868 23324 4956 23380
rect 5012 23324 5022 23380
rect 6738 23324 6748 23380
rect 6804 23324 7756 23380
rect 7812 23324 7822 23380
rect 9212 23324 13580 23380
rect 13636 23324 13646 23380
rect 14018 23324 14028 23380
rect 14084 23324 14364 23380
rect 14420 23324 14430 23380
rect 14700 23324 15092 23380
rect 21858 23324 21868 23380
rect 21924 23324 30268 23380
rect 30324 23324 30334 23380
rect 2258 23212 2268 23268
rect 2324 23212 8988 23268
rect 9044 23212 9054 23268
rect 0 23156 112 23184
rect 9212 23156 9268 23324
rect 15036 23268 15092 23324
rect 13234 23212 13244 23268
rect 13300 23212 14868 23268
rect 15036 23212 19404 23268
rect 19460 23212 19470 23268
rect 14812 23156 14868 23212
rect 0 23100 9268 23156
rect 10658 23100 10668 23156
rect 10724 23100 11004 23156
rect 11060 23100 11070 23156
rect 13906 23100 13916 23156
rect 13972 23100 14588 23156
rect 14644 23100 14654 23156
rect 14802 23100 14812 23156
rect 14868 23100 15484 23156
rect 15540 23100 15550 23156
rect 17042 23100 17052 23156
rect 17108 23100 17500 23156
rect 17556 23100 17566 23156
rect 18386 23100 18396 23156
rect 18452 23100 22428 23156
rect 22484 23100 22494 23156
rect 23202 23100 23212 23156
rect 23268 23100 23436 23156
rect 23492 23100 23502 23156
rect 0 23072 112 23100
rect 802 22988 812 23044
rect 868 22988 1596 23044
rect 1652 22988 1662 23044
rect 4386 22988 4396 23044
rect 4452 22988 4844 23044
rect 4900 22988 4910 23044
rect 5170 22988 5180 23044
rect 5236 22988 5404 23044
rect 5460 22988 10220 23044
rect 10276 22988 10286 23044
rect 12002 22988 12012 23044
rect 12068 22988 13972 23044
rect 14326 22988 14364 23044
rect 14420 22988 14430 23044
rect 15026 22988 15036 23044
rect 15092 22988 16492 23044
rect 16548 22988 16558 23044
rect 18022 22988 18060 23044
rect 18116 22988 18126 23044
rect 18834 22988 18844 23044
rect 18900 22988 18956 23044
rect 19012 22988 19022 23044
rect 21858 22988 21868 23044
rect 21924 22988 22988 23044
rect 23044 22988 23054 23044
rect 13916 22932 13972 22988
rect 2146 22876 2156 22932
rect 2212 22876 3164 22932
rect 3220 22876 3230 22932
rect 5590 22876 5628 22932
rect 5684 22876 6412 22932
rect 6468 22876 6478 22932
rect 13916 22876 18844 22932
rect 18900 22876 18910 22932
rect 23062 22876 23100 22932
rect 23156 22876 24108 22932
rect 24164 22876 24174 22932
rect 7980 22764 13748 22820
rect 13906 22764 13916 22820
rect 13972 22764 14010 22820
rect 15092 22764 15596 22820
rect 15652 22764 15662 22820
rect 20514 22764 20524 22820
rect 20580 22764 23212 22820
rect 23268 22764 23278 22820
rect 0 22708 112 22736
rect 4454 22708 4464 22764
rect 4520 22708 4568 22764
rect 4624 22708 4672 22764
rect 4728 22708 4738 22764
rect 7980 22708 8036 22764
rect 13692 22708 13748 22764
rect 15092 22708 15148 22764
rect 24454 22708 24464 22764
rect 24520 22708 24568 22764
rect 24624 22708 24672 22764
rect 24728 22708 24738 22764
rect 31584 22708 31696 22736
rect 0 22652 4060 22708
rect 4116 22652 4126 22708
rect 4834 22652 4844 22708
rect 4900 22652 5740 22708
rect 5796 22652 8036 22708
rect 11340 22652 13020 22708
rect 13076 22652 13468 22708
rect 13524 22652 13534 22708
rect 13692 22652 15148 22708
rect 22754 22652 22764 22708
rect 22820 22652 23548 22708
rect 23604 22652 23614 22708
rect 30594 22652 30604 22708
rect 30660 22652 31696 22708
rect 0 22624 112 22652
rect 11340 22596 11396 22652
rect 31584 22624 31696 22652
rect 1708 22540 11396 22596
rect 11554 22540 11564 22596
rect 11620 22540 12628 22596
rect 13122 22540 13132 22596
rect 13188 22540 14924 22596
rect 14980 22540 15708 22596
rect 15764 22540 15774 22596
rect 17602 22540 17612 22596
rect 17668 22540 30268 22596
rect 30324 22540 30334 22596
rect 0 22260 112 22288
rect 1708 22260 1764 22540
rect 12572 22484 12628 22540
rect 2594 22428 2604 22484
rect 2660 22428 6860 22484
rect 6916 22428 9996 22484
rect 10052 22428 10062 22484
rect 12002 22428 12012 22484
rect 12068 22428 12348 22484
rect 12404 22428 12414 22484
rect 12572 22428 16940 22484
rect 16996 22428 17006 22484
rect 2482 22316 2492 22372
rect 2548 22316 7084 22372
rect 7140 22316 18060 22372
rect 18116 22316 22540 22372
rect 22596 22316 22606 22372
rect 0 22204 1764 22260
rect 4050 22204 4060 22260
rect 4116 22204 5124 22260
rect 6178 22204 6188 22260
rect 6244 22204 6636 22260
rect 6692 22204 6702 22260
rect 9314 22204 9324 22260
rect 9380 22204 15148 22260
rect 15362 22204 15372 22260
rect 15428 22204 16380 22260
rect 16436 22204 16446 22260
rect 16818 22204 16828 22260
rect 16884 22204 17276 22260
rect 17332 22204 17342 22260
rect 17602 22204 17612 22260
rect 17668 22204 18396 22260
rect 18452 22204 18462 22260
rect 23650 22204 23660 22260
rect 23716 22204 23772 22260
rect 23828 22204 23838 22260
rect 0 22176 112 22204
rect 1922 22092 1932 22148
rect 1988 22092 4844 22148
rect 4900 22092 4910 22148
rect 5068 22036 5124 22204
rect 15092 22148 15148 22204
rect 5842 22092 5852 22148
rect 5908 22092 7308 22148
rect 7364 22092 7374 22148
rect 7746 22092 7756 22148
rect 7812 22092 10444 22148
rect 10500 22092 10510 22148
rect 11666 22092 11676 22148
rect 11732 22092 13132 22148
rect 13188 22092 13198 22148
rect 13458 22092 13468 22148
rect 13524 22092 14364 22148
rect 14420 22092 14430 22148
rect 14690 22092 14700 22148
rect 14756 22092 14812 22148
rect 14868 22092 14878 22148
rect 15092 22092 18844 22148
rect 18900 22092 18910 22148
rect 20514 22092 20524 22148
rect 20580 22092 21756 22148
rect 21812 22092 24220 22148
rect 24276 22092 24286 22148
rect 5068 21980 7980 22036
rect 8036 21980 8046 22036
rect 10098 21980 10108 22036
rect 10164 21980 12348 22036
rect 12404 21980 22092 22036
rect 22148 21980 22158 22036
rect 3794 21924 3804 21980
rect 3860 21924 3908 21980
rect 3964 21924 4012 21980
rect 4068 21924 4078 21980
rect 23794 21924 23804 21980
rect 23860 21924 23908 21980
rect 23964 21924 24012 21980
rect 24068 21924 24078 21980
rect 7074 21868 7084 21924
rect 7140 21868 13244 21924
rect 13300 21868 13310 21924
rect 13570 21868 13580 21924
rect 13636 21868 14812 21924
rect 14868 21868 14878 21924
rect 19506 21868 19516 21924
rect 19572 21868 21196 21924
rect 21252 21868 21262 21924
rect 0 21812 112 21840
rect 31584 21812 31696 21840
rect 0 21756 10612 21812
rect 12786 21756 12796 21812
rect 12852 21756 13804 21812
rect 13860 21756 13870 21812
rect 15026 21756 15036 21812
rect 15092 21756 17388 21812
rect 17444 21756 17454 21812
rect 22530 21756 22540 21812
rect 22596 21756 23324 21812
rect 23380 21756 23390 21812
rect 30594 21756 30604 21812
rect 30660 21756 31696 21812
rect 0 21728 112 21756
rect 10556 21700 10612 21756
rect 31584 21728 31696 21756
rect 1362 21644 1372 21700
rect 1428 21644 2156 21700
rect 2212 21644 2222 21700
rect 2594 21644 2604 21700
rect 2660 21644 3388 21700
rect 3444 21644 3454 21700
rect 3602 21644 3612 21700
rect 3668 21644 5404 21700
rect 5460 21644 5470 21700
rect 10556 21644 13132 21700
rect 13188 21644 15820 21700
rect 15876 21644 15886 21700
rect 2156 21588 2212 21644
rect 2156 21532 2716 21588
rect 2772 21532 2782 21588
rect 13570 21532 13580 21588
rect 13636 21532 14140 21588
rect 14196 21532 14206 21588
rect 14354 21532 14364 21588
rect 14420 21532 14700 21588
rect 14756 21532 14766 21588
rect 17826 21532 17836 21588
rect 17892 21532 18172 21588
rect 18228 21532 18238 21588
rect 18386 21532 18396 21588
rect 18452 21532 19180 21588
rect 19236 21532 19246 21588
rect 19842 21532 19852 21588
rect 19908 21532 22764 21588
rect 22820 21532 22830 21588
rect 2034 21420 2044 21476
rect 2100 21420 7868 21476
rect 7924 21420 7934 21476
rect 12450 21420 12460 21476
rect 12516 21420 14700 21476
rect 14756 21420 14766 21476
rect 21382 21420 21420 21476
rect 21476 21420 21486 21476
rect 0 21364 112 21392
rect 0 21308 1036 21364
rect 1092 21308 1102 21364
rect 4050 21308 4060 21364
rect 4116 21308 15148 21364
rect 0 21280 112 21308
rect 15092 21252 15148 21308
rect 19068 21308 19852 21364
rect 19908 21308 19918 21364
rect 7298 21196 7308 21252
rect 7364 21196 7868 21252
rect 7924 21196 7934 21252
rect 12786 21196 12796 21252
rect 12852 21196 13468 21252
rect 13524 21196 13534 21252
rect 13794 21196 13804 21252
rect 13860 21196 14364 21252
rect 14420 21196 14430 21252
rect 15092 21196 16604 21252
rect 16660 21196 16670 21252
rect 4454 21140 4464 21196
rect 4520 21140 4568 21196
rect 4624 21140 4672 21196
rect 4728 21140 4738 21196
rect 19068 21140 19124 21308
rect 19282 21196 19292 21252
rect 19348 21196 20748 21252
rect 20804 21196 20814 21252
rect 24454 21140 24464 21196
rect 24520 21140 24568 21196
rect 24624 21140 24672 21196
rect 24728 21140 24738 21196
rect 4946 21084 4956 21140
rect 5012 21084 9212 21140
rect 9268 21084 9996 21140
rect 10052 21084 10062 21140
rect 12674 21084 12684 21140
rect 12740 21084 13916 21140
rect 13972 21084 13982 21140
rect 14130 21084 14140 21140
rect 14196 21084 19124 21140
rect 19618 21084 19628 21140
rect 19684 21084 19852 21140
rect 19908 21084 21308 21140
rect 21364 21084 21374 21140
rect 1698 20972 1708 21028
rect 1764 20972 4172 21028
rect 4228 20972 4396 21028
rect 4452 20972 4462 21028
rect 6178 20972 6188 21028
rect 6244 20972 12012 21028
rect 12068 20972 12078 21028
rect 13906 20972 13916 21028
rect 13972 20972 14812 21028
rect 14868 20972 14878 21028
rect 16454 20972 16492 21028
rect 16548 20972 16558 21028
rect 0 20916 112 20944
rect 31584 20916 31696 20944
rect 0 20860 1596 20916
rect 1652 20860 1662 20916
rect 6962 20860 6972 20916
rect 7028 20860 15708 20916
rect 15764 20860 15774 20916
rect 16034 20860 16044 20916
rect 16100 20860 17612 20916
rect 17668 20860 17678 20916
rect 18050 20860 18060 20916
rect 18116 20860 19516 20916
rect 19572 20860 19582 20916
rect 30706 20860 30716 20916
rect 30772 20860 31696 20916
rect 0 20832 112 20860
rect 31584 20832 31696 20860
rect 7298 20748 7308 20804
rect 7364 20748 9436 20804
rect 9492 20748 9502 20804
rect 11218 20748 11228 20804
rect 11284 20748 13132 20804
rect 13188 20748 13198 20804
rect 13906 20748 13916 20804
rect 13972 20748 17052 20804
rect 17108 20748 17118 20804
rect 21522 20748 21532 20804
rect 21588 20748 30268 20804
rect 30324 20748 30334 20804
rect 2594 20636 2604 20692
rect 2660 20636 3164 20692
rect 3220 20636 5964 20692
rect 6020 20636 15708 20692
rect 15764 20636 15774 20692
rect 16034 20636 16044 20692
rect 16100 20636 30156 20692
rect 30212 20636 30222 20692
rect 4722 20524 4732 20580
rect 4788 20524 4844 20580
rect 4900 20524 4910 20580
rect 5058 20524 5068 20580
rect 5124 20524 5162 20580
rect 7522 20524 7532 20580
rect 7588 20524 12124 20580
rect 12180 20524 12190 20580
rect 15586 20524 15596 20580
rect 15652 20524 18060 20580
rect 18116 20524 18126 20580
rect 0 20468 112 20496
rect 0 20412 924 20468
rect 980 20412 990 20468
rect 1698 20412 1708 20468
rect 1764 20412 2156 20468
rect 2212 20412 2222 20468
rect 7970 20412 7980 20468
rect 8036 20412 14476 20468
rect 14532 20412 14542 20468
rect 0 20384 112 20412
rect 3794 20356 3804 20412
rect 3860 20356 3908 20412
rect 3964 20356 4012 20412
rect 4068 20356 4078 20412
rect 23794 20356 23804 20412
rect 23860 20356 23908 20412
rect 23964 20356 24012 20412
rect 24068 20356 24078 20412
rect 1250 20300 1260 20356
rect 1316 20300 1596 20356
rect 1652 20300 1662 20356
rect 9538 20300 9548 20356
rect 9604 20300 9884 20356
rect 9940 20300 9950 20356
rect 19954 20300 19964 20356
rect 20020 20300 20636 20356
rect 20692 20300 20702 20356
rect 3332 20188 3612 20244
rect 3668 20188 3678 20244
rect 4172 20188 4396 20244
rect 4452 20188 4956 20244
rect 5012 20188 8092 20244
rect 8148 20188 8158 20244
rect 8540 20188 10780 20244
rect 10836 20188 11676 20244
rect 11732 20188 11742 20244
rect 12002 20188 12012 20244
rect 12068 20188 26012 20244
rect 26068 20188 26078 20244
rect 1138 20076 1148 20132
rect 1204 20076 1932 20132
rect 1988 20076 1998 20132
rect 0 20020 112 20048
rect 3332 20020 3388 20188
rect 4172 20020 4228 20188
rect 8540 20132 8596 20188
rect 7410 20076 7420 20132
rect 7476 20076 8540 20132
rect 8596 20076 8606 20132
rect 8754 20076 8764 20132
rect 8820 20076 9436 20132
rect 9492 20076 9502 20132
rect 9650 20076 9660 20132
rect 9716 20076 10556 20132
rect 10612 20076 10622 20132
rect 31584 20020 31696 20048
rect 0 19964 3388 20020
rect 4162 19964 4172 20020
rect 4228 19964 4238 20020
rect 5366 19964 5404 20020
rect 5460 19964 5470 20020
rect 6738 19964 6748 20020
rect 6804 19964 7196 20020
rect 7252 19964 7262 20020
rect 8194 19964 8204 20020
rect 8260 19964 10108 20020
rect 10164 19964 10174 20020
rect 13122 19964 13132 20020
rect 13188 19964 15260 20020
rect 15316 19964 20860 20020
rect 20916 19964 20926 20020
rect 30594 19964 30604 20020
rect 30660 19964 31696 20020
rect 0 19936 112 19964
rect 31584 19936 31696 19964
rect 354 19852 364 19908
rect 420 19852 8652 19908
rect 8708 19852 9548 19908
rect 9604 19852 9614 19908
rect 13682 19852 13692 19908
rect 13748 19852 15484 19908
rect 15540 19852 16044 19908
rect 16100 19852 17948 19908
rect 18004 19852 18014 19908
rect 18386 19852 18396 19908
rect 18452 19852 18620 19908
rect 18676 19852 19180 19908
rect 19236 19852 23212 19908
rect 23268 19852 23278 19908
rect 18396 19796 18452 19852
rect 578 19740 588 19796
rect 644 19740 2156 19796
rect 2212 19740 2222 19796
rect 2706 19740 2716 19796
rect 2772 19740 3500 19796
rect 3556 19740 5852 19796
rect 5908 19740 9660 19796
rect 9716 19740 12460 19796
rect 12516 19740 12526 19796
rect 15586 19740 15596 19796
rect 15652 19740 16940 19796
rect 16996 19740 18452 19796
rect 4834 19628 4844 19684
rect 4900 19628 5068 19684
rect 5124 19628 5134 19684
rect 0 19572 112 19600
rect 4454 19572 4464 19628
rect 4520 19572 4568 19628
rect 4624 19572 4672 19628
rect 4728 19572 4738 19628
rect 24454 19572 24464 19628
rect 24520 19572 24568 19628
rect 24624 19572 24672 19628
rect 24728 19572 24738 19628
rect 0 19516 3276 19572
rect 3332 19516 3342 19572
rect 7522 19516 7532 19572
rect 7588 19516 7980 19572
rect 8036 19516 12348 19572
rect 12404 19516 12414 19572
rect 13570 19516 13580 19572
rect 13636 19516 14252 19572
rect 14308 19516 14318 19572
rect 19058 19516 19068 19572
rect 19124 19516 19852 19572
rect 19908 19516 19918 19572
rect 0 19488 112 19516
rect 1922 19404 1932 19460
rect 1988 19404 4844 19460
rect 4900 19404 4910 19460
rect 6850 19404 6860 19460
rect 6916 19404 7756 19460
rect 7812 19404 7822 19460
rect 8194 19404 8204 19460
rect 8260 19404 8988 19460
rect 9044 19404 9054 19460
rect 11890 19404 11900 19460
rect 11956 19404 13580 19460
rect 13636 19404 13646 19460
rect 17714 19404 17724 19460
rect 17780 19404 18284 19460
rect 18340 19404 18508 19460
rect 18564 19404 18574 19460
rect 19954 19404 19964 19460
rect 20020 19404 21980 19460
rect 22036 19404 22046 19460
rect 27906 19404 27916 19460
rect 27972 19404 30268 19460
rect 30324 19404 30334 19460
rect 1250 19292 1260 19348
rect 1316 19292 5964 19348
rect 6020 19292 6030 19348
rect 6738 19292 6748 19348
rect 6804 19292 9100 19348
rect 9156 19292 9166 19348
rect 9986 19292 9996 19348
rect 10052 19292 10220 19348
rect 10276 19292 11228 19348
rect 11284 19292 11294 19348
rect 12562 19292 12572 19348
rect 12628 19292 13244 19348
rect 13300 19292 13310 19348
rect 15922 19292 15932 19348
rect 15988 19292 17164 19348
rect 17220 19292 17230 19348
rect 2034 19180 2044 19236
rect 2100 19180 2716 19236
rect 2772 19180 2782 19236
rect 3378 19180 3388 19236
rect 3444 19180 3948 19236
rect 4004 19180 4014 19236
rect 11106 19180 11116 19236
rect 11172 19180 11900 19236
rect 11956 19180 11966 19236
rect 13570 19180 13580 19236
rect 13636 19180 15148 19236
rect 17378 19180 17388 19236
rect 17444 19180 17724 19236
rect 17780 19180 17790 19236
rect 0 19124 112 19152
rect 15092 19124 15148 19180
rect 31584 19124 31696 19152
rect 0 19068 3612 19124
rect 3668 19068 3678 19124
rect 6178 19068 6188 19124
rect 6244 19068 6636 19124
rect 6692 19068 13020 19124
rect 13076 19068 13086 19124
rect 15092 19068 17948 19124
rect 18004 19068 18014 19124
rect 30594 19068 30604 19124
rect 30660 19068 31696 19124
rect 0 19040 112 19068
rect 31584 19040 31696 19068
rect 4050 18956 4060 19012
rect 4116 18956 5740 19012
rect 5796 18956 5806 19012
rect 9650 18956 9660 19012
rect 9716 18956 9884 19012
rect 9940 18956 9950 19012
rect 10546 18956 10556 19012
rect 10612 18956 11340 19012
rect 11396 18956 11406 19012
rect 15138 18956 15148 19012
rect 15204 18956 15596 19012
rect 15652 18956 15662 19012
rect 8866 18844 8876 18900
rect 8932 18844 19180 18900
rect 19236 18844 19246 18900
rect 3794 18788 3804 18844
rect 3860 18788 3908 18844
rect 3964 18788 4012 18844
rect 4068 18788 4078 18844
rect 23794 18788 23804 18844
rect 23860 18788 23908 18844
rect 23964 18788 24012 18844
rect 24068 18788 24078 18844
rect 6066 18732 6076 18788
rect 6132 18732 10948 18788
rect 13906 18732 13916 18788
rect 13972 18732 14588 18788
rect 14644 18732 15260 18788
rect 15316 18732 15326 18788
rect 0 18676 112 18704
rect 10892 18676 10948 18732
rect 0 18620 5516 18676
rect 5572 18620 5582 18676
rect 9762 18620 9772 18676
rect 9828 18620 10668 18676
rect 10724 18620 10734 18676
rect 10892 18620 23660 18676
rect 23716 18620 23726 18676
rect 0 18592 112 18620
rect 3378 18508 3388 18564
rect 3444 18508 4956 18564
rect 5012 18508 7084 18564
rect 7140 18508 7150 18564
rect 10322 18508 10332 18564
rect 10388 18508 11900 18564
rect 11956 18508 11966 18564
rect 13010 18508 13020 18564
rect 13076 18508 13132 18564
rect 13188 18508 13198 18564
rect 14466 18508 14476 18564
rect 14532 18508 15148 18564
rect 15204 18508 15214 18564
rect 15362 18508 15372 18564
rect 15428 18508 16996 18564
rect 16940 18452 16996 18508
rect 1586 18396 1596 18452
rect 1652 18396 4172 18452
rect 4228 18396 4238 18452
rect 8950 18396 8988 18452
rect 9044 18396 9054 18452
rect 12002 18396 12012 18452
rect 12068 18396 12460 18452
rect 12516 18396 12526 18452
rect 16930 18396 16940 18452
rect 16996 18396 17006 18452
rect 24994 18396 25004 18452
rect 25060 18396 30268 18452
rect 30324 18396 30334 18452
rect 2118 18284 2156 18340
rect 2212 18284 2222 18340
rect 2706 18284 2716 18340
rect 2772 18284 7868 18340
rect 7924 18284 7934 18340
rect 11666 18284 11676 18340
rect 11732 18284 12908 18340
rect 12964 18284 12974 18340
rect 13458 18284 13468 18340
rect 13524 18284 14812 18340
rect 14868 18284 15596 18340
rect 15652 18284 16940 18340
rect 16996 18284 17006 18340
rect 0 18228 112 18256
rect 31584 18228 31696 18256
rect 0 18172 4956 18228
rect 5012 18172 5022 18228
rect 5590 18172 5628 18228
rect 5684 18172 5694 18228
rect 16146 18172 16156 18228
rect 16212 18172 17836 18228
rect 17892 18172 17902 18228
rect 30594 18172 30604 18228
rect 30660 18172 31696 18228
rect 0 18144 112 18172
rect 31584 18144 31696 18172
rect 1698 18060 1708 18116
rect 1764 18060 2716 18116
rect 2772 18060 2782 18116
rect 5954 18060 5964 18116
rect 6020 18060 15596 18116
rect 15652 18060 15662 18116
rect 4454 18004 4464 18060
rect 4520 18004 4568 18060
rect 4624 18004 4672 18060
rect 4728 18004 4738 18060
rect 24454 18004 24464 18060
rect 24520 18004 24568 18060
rect 24624 18004 24672 18060
rect 24728 18004 24738 18060
rect 6178 17948 6188 18004
rect 6244 17948 6636 18004
rect 6692 17948 6702 18004
rect 11218 17948 11228 18004
rect 11284 17948 18508 18004
rect 18564 17948 18574 18004
rect 1810 17836 1820 17892
rect 1876 17836 3276 17892
rect 3332 17836 5460 17892
rect 11554 17836 11564 17892
rect 11620 17836 16716 17892
rect 16772 17836 16782 17892
rect 18946 17836 18956 17892
rect 19012 17836 20188 17892
rect 20244 17836 20254 17892
rect 27794 17836 27804 17892
rect 27860 17836 30268 17892
rect 30324 17836 30334 17892
rect 0 17780 112 17808
rect 0 17724 3612 17780
rect 3668 17724 3678 17780
rect 4162 17724 4172 17780
rect 4228 17724 4284 17780
rect 4340 17724 4350 17780
rect 0 17696 112 17724
rect 5404 17668 5460 17836
rect 6738 17724 6748 17780
rect 6804 17724 7084 17780
rect 7140 17724 7150 17780
rect 11442 17724 11452 17780
rect 11508 17724 14924 17780
rect 14980 17724 14990 17780
rect 18610 17724 18620 17780
rect 18676 17724 19964 17780
rect 20020 17724 20030 17780
rect 21634 17724 21644 17780
rect 21700 17724 27020 17780
rect 27076 17724 27086 17780
rect 2258 17612 2268 17668
rect 2324 17612 3612 17668
rect 3668 17612 3678 17668
rect 5394 17612 5404 17668
rect 5460 17612 5470 17668
rect 5730 17612 5740 17668
rect 5796 17612 6860 17668
rect 6916 17612 6926 17668
rect 7858 17612 7868 17668
rect 7924 17612 9100 17668
rect 9156 17612 14700 17668
rect 14756 17612 14766 17668
rect 25778 17612 25788 17668
rect 25844 17612 26796 17668
rect 26852 17612 26862 17668
rect 2146 17500 2156 17556
rect 2212 17500 3780 17556
rect 3938 17500 3948 17556
rect 4004 17500 5516 17556
rect 5572 17500 6188 17556
rect 6244 17500 6254 17556
rect 3724 17444 3780 17500
rect 690 17388 700 17444
rect 756 17388 3388 17444
rect 3444 17388 3454 17444
rect 3724 17388 5124 17444
rect 5282 17388 5292 17444
rect 5348 17388 18284 17444
rect 18340 17388 18350 17444
rect 0 17332 112 17360
rect 5068 17332 5124 17388
rect 31584 17332 31696 17360
rect 0 17276 3164 17332
rect 3220 17276 3230 17332
rect 5068 17276 5852 17332
rect 5908 17276 5918 17332
rect 6626 17276 6636 17332
rect 6692 17276 11340 17332
rect 11396 17276 11564 17332
rect 11620 17276 11630 17332
rect 30594 17276 30604 17332
rect 30660 17276 31696 17332
rect 0 17248 112 17276
rect 3794 17220 3804 17276
rect 3860 17220 3908 17276
rect 3964 17220 4012 17276
rect 4068 17220 4078 17276
rect 23794 17220 23804 17276
rect 23860 17220 23908 17276
rect 23964 17220 24012 17276
rect 24068 17220 24078 17276
rect 31584 17248 31696 17276
rect 2706 17164 2716 17220
rect 2772 17164 3276 17220
rect 3332 17164 3342 17220
rect 4274 17164 4284 17220
rect 4340 17164 15036 17220
rect 15092 17164 15102 17220
rect 5394 17052 5404 17108
rect 5460 17052 6636 17108
rect 6692 17052 6702 17108
rect 6962 17052 6972 17108
rect 7028 17052 7196 17108
rect 7252 17052 7262 17108
rect 9202 17052 9212 17108
rect 9268 17052 12908 17108
rect 12964 17052 12974 17108
rect 14914 17052 14924 17108
rect 14980 17052 20188 17108
rect 20244 17052 21644 17108
rect 21700 17052 21710 17108
rect 3238 16940 3276 16996
rect 3332 16940 3342 16996
rect 13346 16940 13356 16996
rect 13412 16940 13804 16996
rect 13860 16940 13870 16996
rect 0 16884 112 16912
rect 0 16828 4844 16884
rect 4900 16828 4910 16884
rect 6290 16828 6300 16884
rect 6356 16828 9996 16884
rect 10052 16828 10062 16884
rect 18498 16828 18508 16884
rect 18564 16828 20076 16884
rect 20132 16828 20142 16884
rect 0 16800 112 16828
rect 1474 16716 1484 16772
rect 1540 16716 7980 16772
rect 8036 16716 8046 16772
rect 8194 16716 8204 16772
rect 8260 16716 8298 16772
rect 15092 16716 18844 16772
rect 18900 16716 20636 16772
rect 20692 16716 20702 16772
rect 22306 16716 22316 16772
rect 22372 16716 24892 16772
rect 24948 16716 24958 16772
rect 3332 16604 5628 16660
rect 5684 16604 5694 16660
rect 11078 16604 11116 16660
rect 11172 16604 11182 16660
rect 14326 16604 14364 16660
rect 14420 16604 14430 16660
rect 0 16436 112 16464
rect 3332 16436 3388 16604
rect 11116 16548 11172 16604
rect 15092 16548 15148 16716
rect 17826 16604 17836 16660
rect 17892 16604 17948 16660
rect 18004 16604 18014 16660
rect 22642 16604 22652 16660
rect 22708 16604 30268 16660
rect 30324 16604 30334 16660
rect 5954 16492 5964 16548
rect 6020 16492 15148 16548
rect 20962 16492 20972 16548
rect 21028 16492 21196 16548
rect 21252 16492 21262 16548
rect 4454 16436 4464 16492
rect 4520 16436 4568 16492
rect 4624 16436 4672 16492
rect 4728 16436 4738 16492
rect 24454 16436 24464 16492
rect 24520 16436 24568 16492
rect 24624 16436 24672 16492
rect 24728 16436 24738 16492
rect 31584 16436 31696 16464
rect 0 16380 3388 16436
rect 5730 16380 5740 16436
rect 5796 16380 5852 16436
rect 5908 16380 5918 16436
rect 30594 16380 30604 16436
rect 30660 16380 31696 16436
rect 0 16352 112 16380
rect 31584 16352 31696 16380
rect 2482 16268 2492 16324
rect 2548 16268 3276 16324
rect 3332 16268 3342 16324
rect 6514 16268 6524 16324
rect 6580 16268 7084 16324
rect 7140 16268 7150 16324
rect 11890 16268 11900 16324
rect 11956 16268 15932 16324
rect 15988 16268 19852 16324
rect 19908 16268 19918 16324
rect 25890 16268 25900 16324
rect 25956 16268 30268 16324
rect 30324 16268 30334 16324
rect 3602 16156 3612 16212
rect 3668 16156 11228 16212
rect 11284 16156 11294 16212
rect 11554 16156 11564 16212
rect 11620 16156 12908 16212
rect 12964 16156 12974 16212
rect 2380 16044 4116 16100
rect 4246 16044 4284 16100
rect 4340 16044 4350 16100
rect 5506 16044 5516 16100
rect 5572 16044 8988 16100
rect 9044 16044 9054 16100
rect 12002 16044 12012 16100
rect 12068 16044 12236 16100
rect 12292 16044 12302 16100
rect 14018 16044 14028 16100
rect 14084 16044 14924 16100
rect 14980 16044 14990 16100
rect 21186 16044 21196 16100
rect 21252 16044 23100 16100
rect 23156 16044 23166 16100
rect 0 15988 112 16016
rect 2380 15988 2436 16044
rect 0 15932 2436 15988
rect 4060 15988 4116 16044
rect 4060 15932 4844 15988
rect 4900 15932 4910 15988
rect 9874 15932 9884 15988
rect 9940 15932 11564 15988
rect 11620 15932 11630 15988
rect 18050 15932 18060 15988
rect 18116 15932 19404 15988
rect 19460 15932 19470 15988
rect 26534 15932 26572 15988
rect 26628 15932 26638 15988
rect 0 15904 112 15932
rect 10098 15820 10108 15876
rect 10164 15820 10668 15876
rect 10724 15820 10734 15876
rect 11778 15820 11788 15876
rect 11844 15820 12460 15876
rect 12516 15820 12526 15876
rect 12786 15820 12796 15876
rect 12852 15820 18956 15876
rect 19012 15820 19022 15876
rect 5618 15708 5628 15764
rect 5684 15708 9324 15764
rect 9380 15708 18172 15764
rect 18228 15708 18238 15764
rect 3794 15652 3804 15708
rect 3860 15652 3908 15708
rect 3964 15652 4012 15708
rect 4068 15652 4078 15708
rect 23794 15652 23804 15708
rect 23860 15652 23908 15708
rect 23964 15652 24012 15708
rect 24068 15652 24078 15708
rect 5058 15596 5068 15652
rect 5124 15596 5404 15652
rect 5460 15596 5470 15652
rect 11106 15596 11116 15652
rect 11172 15596 14476 15652
rect 14532 15596 14542 15652
rect 17042 15596 17052 15652
rect 17108 15596 17724 15652
rect 17780 15596 17790 15652
rect 0 15540 112 15568
rect 31584 15540 31696 15568
rect 0 15484 1036 15540
rect 1092 15484 1102 15540
rect 2706 15484 2716 15540
rect 2772 15484 5068 15540
rect 5124 15484 5134 15540
rect 7532 15484 17388 15540
rect 17444 15484 17454 15540
rect 30594 15484 30604 15540
rect 30660 15484 31696 15540
rect 0 15456 112 15484
rect 1250 15372 1260 15428
rect 1316 15372 1932 15428
rect 1988 15372 1998 15428
rect 4162 15372 4172 15428
rect 4228 15372 4396 15428
rect 4452 15372 4462 15428
rect 7532 15316 7588 15484
rect 31584 15456 31696 15484
rect 11778 15372 11788 15428
rect 11844 15372 12124 15428
rect 12180 15372 12190 15428
rect 12422 15372 12460 15428
rect 12516 15372 12526 15428
rect 14018 15372 14028 15428
rect 14084 15372 17948 15428
rect 18004 15372 18014 15428
rect 1362 15260 1372 15316
rect 1428 15260 4060 15316
rect 4116 15260 4126 15316
rect 4284 15260 7588 15316
rect 7858 15260 7868 15316
rect 7924 15260 8764 15316
rect 8820 15260 8830 15316
rect 10658 15260 10668 15316
rect 10724 15260 12572 15316
rect 12628 15260 13916 15316
rect 13972 15260 13982 15316
rect 15922 15260 15932 15316
rect 15988 15260 18060 15316
rect 18116 15260 18126 15316
rect 23426 15260 23436 15316
rect 23492 15260 31388 15316
rect 31444 15260 31454 15316
rect 4284 15204 4340 15260
rect 802 15148 812 15204
rect 868 15148 1596 15204
rect 1652 15148 1662 15204
rect 1932 15148 4340 15204
rect 4610 15148 4620 15204
rect 4676 15148 6076 15204
rect 6132 15148 6142 15204
rect 8306 15148 8316 15204
rect 8372 15148 9436 15204
rect 9492 15148 9502 15204
rect 9650 15148 9660 15204
rect 9716 15148 12908 15204
rect 12964 15148 12974 15204
rect 14130 15148 14140 15204
rect 14196 15148 15484 15204
rect 15540 15148 16268 15204
rect 16324 15148 16334 15204
rect 26450 15148 26460 15204
rect 26516 15148 27804 15204
rect 27860 15148 27870 15204
rect 0 15092 112 15120
rect 1932 15092 1988 15148
rect 0 15036 1092 15092
rect 1474 15036 1484 15092
rect 1540 15036 1988 15092
rect 4284 15036 6188 15092
rect 6244 15036 6748 15092
rect 6804 15036 6814 15092
rect 8082 15036 8092 15092
rect 8148 15036 9324 15092
rect 9380 15036 9390 15092
rect 26338 15036 26348 15092
rect 26404 15036 26516 15092
rect 0 15008 112 15036
rect 1036 14980 1092 15036
rect 1036 14924 1820 14980
rect 1876 14924 1886 14980
rect 4284 14868 4340 15036
rect 5170 14924 5180 14980
rect 5236 14924 5628 14980
rect 5684 14924 5694 14980
rect 11890 14924 11900 14980
rect 11956 14924 12460 14980
rect 12516 14924 12908 14980
rect 12964 14924 12974 14980
rect 17042 14924 17052 14980
rect 17108 14924 22484 14980
rect 4454 14868 4464 14924
rect 4520 14868 4568 14924
rect 4624 14868 4672 14924
rect 4728 14868 4738 14924
rect 1474 14812 1484 14868
rect 1540 14812 4340 14868
rect 8418 14812 8428 14868
rect 8484 14812 10892 14868
rect 10948 14812 14028 14868
rect 14084 14812 14094 14868
rect 18722 14812 18732 14868
rect 18788 14812 19068 14868
rect 19124 14812 19134 14868
rect 22428 14756 22484 14924
rect 24454 14868 24464 14924
rect 24520 14868 24568 14924
rect 24624 14868 24672 14924
rect 24728 14868 24738 14924
rect 26460 14868 26516 15036
rect 24882 14812 24892 14868
rect 24948 14812 26236 14868
rect 26292 14812 26302 14868
rect 26450 14812 26460 14868
rect 26516 14812 26526 14868
rect 1250 14700 1260 14756
rect 1316 14700 1708 14756
rect 1764 14700 8036 14756
rect 8978 14700 8988 14756
rect 9044 14700 10444 14756
rect 10500 14700 10510 14756
rect 12450 14700 12460 14756
rect 12516 14700 13468 14756
rect 13524 14700 13534 14756
rect 13906 14700 13916 14756
rect 13972 14700 15372 14756
rect 15428 14700 15438 14756
rect 21522 14700 21532 14756
rect 21588 14700 22204 14756
rect 22260 14700 22270 14756
rect 22428 14700 30268 14756
rect 30324 14700 30334 14756
rect 0 14644 112 14672
rect 7980 14644 8036 14700
rect 31584 14644 31696 14672
rect 0 14588 924 14644
rect 980 14588 990 14644
rect 2034 14588 2044 14644
rect 2100 14588 3724 14644
rect 3780 14588 3790 14644
rect 4946 14588 4956 14644
rect 5012 14588 5068 14644
rect 5124 14588 5134 14644
rect 7970 14588 7980 14644
rect 8036 14588 11004 14644
rect 11060 14588 20412 14644
rect 20468 14588 20478 14644
rect 25974 14588 26012 14644
rect 26068 14588 26078 14644
rect 26534 14588 26572 14644
rect 26628 14588 26638 14644
rect 30706 14588 30716 14644
rect 30772 14588 31696 14644
rect 0 14560 112 14588
rect 31584 14560 31696 14588
rect 2258 14476 2268 14532
rect 2324 14476 3836 14532
rect 3892 14476 3902 14532
rect 4386 14476 4396 14532
rect 4452 14476 6300 14532
rect 6356 14476 6366 14532
rect 9874 14476 9884 14532
rect 9940 14476 12684 14532
rect 12740 14476 12750 14532
rect 13122 14476 13132 14532
rect 13188 14476 13580 14532
rect 13636 14476 13646 14532
rect 14018 14476 14028 14532
rect 14084 14476 17500 14532
rect 17556 14476 17566 14532
rect 18386 14476 18396 14532
rect 18452 14476 18732 14532
rect 18788 14476 21196 14532
rect 21252 14476 21756 14532
rect 21812 14476 21822 14532
rect 3836 14420 3892 14476
rect 3836 14364 5852 14420
rect 5908 14364 5918 14420
rect 10658 14364 10668 14420
rect 10724 14364 11116 14420
rect 11172 14364 11182 14420
rect 11330 14364 11340 14420
rect 11396 14364 13804 14420
rect 13860 14364 14812 14420
rect 14868 14364 14878 14420
rect 15026 14364 15036 14420
rect 15092 14364 19516 14420
rect 19572 14364 21532 14420
rect 21588 14364 21598 14420
rect 14812 14308 14868 14364
rect 2706 14252 2716 14308
rect 2772 14252 11900 14308
rect 11956 14252 11966 14308
rect 14812 14252 19740 14308
rect 19796 14252 19806 14308
rect 0 14196 112 14224
rect 0 14140 3612 14196
rect 3668 14140 3678 14196
rect 4386 14140 4396 14196
rect 4452 14140 4732 14196
rect 4788 14140 4956 14196
rect 5012 14140 5022 14196
rect 9090 14140 9100 14196
rect 9156 14140 12460 14196
rect 12516 14140 12684 14196
rect 12740 14140 12750 14196
rect 0 14112 112 14140
rect 3794 14084 3804 14140
rect 3860 14084 3908 14140
rect 3964 14084 4012 14140
rect 4068 14084 4078 14140
rect 23794 14084 23804 14140
rect 23860 14084 23908 14140
rect 23964 14084 24012 14140
rect 24068 14084 24078 14140
rect 4274 14028 4284 14084
rect 4340 14028 4844 14084
rect 4900 14028 4910 14084
rect 5068 14028 9548 14084
rect 9604 14028 9614 14084
rect 14578 14028 14588 14084
rect 14644 14028 15036 14084
rect 15092 14028 15102 14084
rect 5068 13972 5124 14028
rect 3154 13916 3164 13972
rect 3220 13916 5124 13972
rect 5282 13916 5292 13972
rect 5348 13916 7756 13972
rect 7812 13916 7822 13972
rect 10434 13916 10444 13972
rect 10500 13916 13916 13972
rect 13972 13916 22316 13972
rect 22372 13916 22382 13972
rect 1708 13804 3164 13860
rect 3220 13804 3230 13860
rect 4050 13804 4060 13860
rect 4116 13804 18284 13860
rect 18340 13804 18350 13860
rect 0 13748 112 13776
rect 1708 13748 1764 13804
rect 31584 13748 31696 13776
rect 0 13692 1764 13748
rect 2258 13692 2268 13748
rect 2324 13692 2492 13748
rect 2548 13692 2558 13748
rect 3490 13692 3500 13748
rect 3556 13692 3948 13748
rect 4004 13692 7532 13748
rect 7588 13692 7598 13748
rect 7858 13692 7868 13748
rect 7924 13692 8652 13748
rect 8708 13692 8718 13748
rect 9762 13692 9772 13748
rect 9828 13692 11228 13748
rect 11284 13692 11294 13748
rect 14018 13692 14028 13748
rect 14084 13692 14700 13748
rect 14756 13692 14766 13748
rect 16818 13692 16828 13748
rect 16884 13692 17724 13748
rect 17780 13692 21812 13748
rect 30594 13692 30604 13748
rect 30660 13692 31696 13748
rect 0 13664 112 13692
rect 21756 13636 21812 13692
rect 31584 13664 31696 13692
rect 2930 13580 2940 13636
rect 2996 13580 4844 13636
rect 4900 13580 4910 13636
rect 5394 13580 5404 13636
rect 5460 13580 6300 13636
rect 6356 13580 6366 13636
rect 6626 13580 6636 13636
rect 6692 13580 6748 13636
rect 6804 13580 8540 13636
rect 8596 13580 8606 13636
rect 10658 13580 10668 13636
rect 10724 13580 12236 13636
rect 12292 13580 12302 13636
rect 13010 13580 13020 13636
rect 13076 13580 14588 13636
rect 14644 13580 14654 13636
rect 16902 13580 16940 13636
rect 16996 13580 17276 13636
rect 17332 13580 17342 13636
rect 20290 13580 20300 13636
rect 20356 13580 20748 13636
rect 20804 13580 20814 13636
rect 21746 13580 21756 13636
rect 21812 13580 22092 13636
rect 22148 13580 22158 13636
rect 3266 13468 3276 13524
rect 3332 13468 3388 13524
rect 3444 13468 3454 13524
rect 4274 13468 4284 13524
rect 4340 13468 5964 13524
rect 6020 13468 6030 13524
rect 6290 13468 6300 13524
rect 6356 13468 8876 13524
rect 8932 13468 8942 13524
rect 9986 13468 9996 13524
rect 10052 13468 10332 13524
rect 10388 13468 10398 13524
rect 10546 13468 10556 13524
rect 10612 13468 12348 13524
rect 12404 13468 12414 13524
rect 13794 13468 13804 13524
rect 13860 13468 16604 13524
rect 16660 13468 16670 13524
rect 17826 13468 17836 13524
rect 17892 13468 18732 13524
rect 18788 13468 18798 13524
rect 20402 13468 20412 13524
rect 20468 13468 21308 13524
rect 21364 13468 21374 13524
rect 3042 13356 3052 13412
rect 3108 13356 3500 13412
rect 3556 13356 3566 13412
rect 13458 13356 13468 13412
rect 13524 13356 16044 13412
rect 16100 13356 16716 13412
rect 16772 13356 16782 13412
rect 0 13300 112 13328
rect 4454 13300 4464 13356
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4728 13300 4738 13356
rect 24454 13300 24464 13356
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24728 13300 24738 13356
rect 0 13244 700 13300
rect 756 13244 766 13300
rect 6962 13244 6972 13300
rect 7028 13244 10780 13300
rect 10836 13244 13020 13300
rect 13076 13244 13086 13300
rect 13766 13244 13804 13300
rect 13860 13244 13870 13300
rect 19730 13244 19740 13300
rect 19796 13244 20748 13300
rect 20804 13244 21196 13300
rect 21252 13244 21262 13300
rect 0 13216 112 13244
rect 2370 13132 2380 13188
rect 2436 13132 8876 13188
rect 8932 13132 8942 13188
rect 13346 13132 13356 13188
rect 13412 13132 14140 13188
rect 14196 13132 14206 13188
rect 19170 13132 19180 13188
rect 19236 13132 30268 13188
rect 30324 13132 30334 13188
rect 5058 13020 5068 13076
rect 5124 13020 5180 13076
rect 5236 13020 5246 13076
rect 13010 13020 13020 13076
rect 13076 13020 22540 13076
rect 22596 13020 22606 13076
rect 2258 12908 2268 12964
rect 2324 12908 5740 12964
rect 5796 12908 5806 12964
rect 6738 12908 6748 12964
rect 6804 12908 7196 12964
rect 7252 12908 7262 12964
rect 8054 12908 8092 12964
rect 8148 12908 8158 12964
rect 9426 12908 9436 12964
rect 9492 12908 13916 12964
rect 13972 12908 13982 12964
rect 18722 12908 18732 12964
rect 18788 12908 18956 12964
rect 19012 12908 19022 12964
rect 19954 12908 19964 12964
rect 20020 12908 20412 12964
rect 20468 12908 21868 12964
rect 21924 12908 21934 12964
rect 0 12852 112 12880
rect 31584 12852 31696 12880
rect 0 12796 476 12852
rect 532 12796 542 12852
rect 2818 12796 2828 12852
rect 2884 12796 5068 12852
rect 5124 12796 5134 12852
rect 8418 12796 8428 12852
rect 8484 12796 10332 12852
rect 10388 12796 10892 12852
rect 10948 12796 12572 12852
rect 12628 12796 13468 12852
rect 13524 12796 13534 12852
rect 18274 12796 18284 12852
rect 18340 12796 25116 12852
rect 25172 12796 25182 12852
rect 30594 12796 30604 12852
rect 30660 12796 31696 12852
rect 0 12768 112 12796
rect 31584 12768 31696 12796
rect 12002 12684 12012 12740
rect 12068 12684 17724 12740
rect 17780 12684 17790 12740
rect 4722 12572 4732 12628
rect 4788 12572 4956 12628
rect 5012 12572 5852 12628
rect 5908 12572 11900 12628
rect 11956 12572 11966 12628
rect 16818 12572 16828 12628
rect 16884 12572 19964 12628
rect 20020 12572 20030 12628
rect 3794 12516 3804 12572
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 4068 12516 4078 12572
rect 23794 12516 23804 12572
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 24068 12516 24078 12572
rect 2268 12460 2492 12516
rect 2548 12460 2558 12516
rect 4386 12460 4396 12516
rect 4452 12460 15708 12516
rect 15764 12460 15774 12516
rect 0 12404 112 12432
rect 2268 12404 2324 12460
rect 0 12348 2324 12404
rect 2380 12348 17052 12404
rect 17108 12348 17118 12404
rect 26852 12348 27692 12404
rect 27748 12348 27758 12404
rect 0 12320 112 12348
rect 2380 12292 2436 12348
rect 26852 12292 26908 12348
rect 1250 12236 1260 12292
rect 1316 12236 2436 12292
rect 3602 12236 3612 12292
rect 3668 12236 4956 12292
rect 5012 12236 5022 12292
rect 6178 12236 6188 12292
rect 6244 12236 11228 12292
rect 11284 12236 11294 12292
rect 11890 12236 11900 12292
rect 11956 12236 12796 12292
rect 12852 12236 26908 12292
rect 802 12124 812 12180
rect 868 12124 3388 12180
rect 3490 12124 3500 12180
rect 3556 12124 4172 12180
rect 4228 12124 4238 12180
rect 6290 12124 6300 12180
rect 6356 12124 8428 12180
rect 8484 12124 8494 12180
rect 9202 12124 9212 12180
rect 9268 12124 12124 12180
rect 12180 12124 12190 12180
rect 16370 12124 16380 12180
rect 16436 12124 16716 12180
rect 16772 12124 16782 12180
rect 22418 12124 22428 12180
rect 22484 12124 22988 12180
rect 23044 12124 23054 12180
rect 3332 12068 3388 12124
rect 3332 12012 10892 12068
rect 10948 12012 10958 12068
rect 14018 12012 14028 12068
rect 14084 12012 18452 12068
rect 18610 12012 18620 12068
rect 18676 12012 20188 12068
rect 20244 12012 20254 12068
rect 0 11956 112 11984
rect 18396 11956 18452 12012
rect 31584 11956 31696 11984
rect 0 11900 364 11956
rect 420 11900 430 11956
rect 2370 11900 2380 11956
rect 2436 11900 5292 11956
rect 5348 11900 5358 11956
rect 6066 11900 6076 11956
rect 6132 11900 6748 11956
rect 6804 11900 8764 11956
rect 8820 11900 8830 11956
rect 8978 11900 8988 11956
rect 9044 11900 12012 11956
rect 12068 11900 12078 11956
rect 18396 11900 19516 11956
rect 19572 11900 19582 11956
rect 30594 11900 30604 11956
rect 30660 11900 31696 11956
rect 0 11872 112 11900
rect 31584 11872 31696 11900
rect 5730 11788 5740 11844
rect 5796 11788 9436 11844
rect 9492 11788 9502 11844
rect 10770 11788 10780 11844
rect 10836 11788 17612 11844
rect 17668 11788 21868 11844
rect 21924 11788 21934 11844
rect 4454 11732 4464 11788
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4728 11732 4738 11788
rect 24454 11732 24464 11788
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24728 11732 24738 11788
rect 5394 11676 5404 11732
rect 5460 11676 10556 11732
rect 10612 11676 10622 11732
rect 13916 11676 17164 11732
rect 17220 11676 17948 11732
rect 18004 11676 18014 11732
rect 1586 11564 1596 11620
rect 1652 11564 3388 11620
rect 3444 11564 3454 11620
rect 4274 11564 4284 11620
rect 4340 11564 5404 11620
rect 5460 11564 5470 11620
rect 6066 11564 6076 11620
rect 6132 11564 6412 11620
rect 6468 11564 6478 11620
rect 6626 11564 6636 11620
rect 6692 11564 7308 11620
rect 7364 11564 7374 11620
rect 10434 11564 10444 11620
rect 10500 11564 11228 11620
rect 11284 11564 11294 11620
rect 0 11508 112 11536
rect 13916 11508 13972 11676
rect 17378 11564 17388 11620
rect 17444 11564 19180 11620
rect 19236 11564 19246 11620
rect 28018 11564 28028 11620
rect 28084 11564 30268 11620
rect 30324 11564 30334 11620
rect 0 11452 7756 11508
rect 7812 11452 7822 11508
rect 9874 11452 9884 11508
rect 9940 11452 13916 11508
rect 13972 11452 13982 11508
rect 15092 11452 19404 11508
rect 19460 11452 19470 11508
rect 0 11424 112 11452
rect 4946 11340 4956 11396
rect 5012 11340 6524 11396
rect 6580 11340 6590 11396
rect 10434 11340 10444 11396
rect 10500 11340 12012 11396
rect 12068 11340 12078 11396
rect 15092 11284 15148 11452
rect 15698 11340 15708 11396
rect 15764 11340 23660 11396
rect 23716 11340 23726 11396
rect 2370 11228 2380 11284
rect 2436 11228 2828 11284
rect 2884 11228 2894 11284
rect 5730 11228 5740 11284
rect 5796 11228 6076 11284
rect 6132 11228 6300 11284
rect 6356 11228 6366 11284
rect 8754 11228 8764 11284
rect 8820 11228 15148 11284
rect 21186 11228 21196 11284
rect 21252 11228 21644 11284
rect 21700 11228 21710 11284
rect 2034 11116 2044 11172
rect 2100 11116 4844 11172
rect 4900 11116 4910 11172
rect 5842 11116 5852 11172
rect 5908 11116 15708 11172
rect 15764 11116 15774 11172
rect 0 11060 112 11088
rect 31584 11060 31696 11088
rect 0 11004 1820 11060
rect 1876 11004 1886 11060
rect 4610 11004 4620 11060
rect 4676 11004 8204 11060
rect 8260 11004 8270 11060
rect 10994 11004 11004 11060
rect 11060 11004 12348 11060
rect 12404 11004 14700 11060
rect 14756 11004 14766 11060
rect 30594 11004 30604 11060
rect 30660 11004 31696 11060
rect 0 10976 112 11004
rect 3794 10948 3804 11004
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 4068 10948 4078 11004
rect 23794 10948 23804 11004
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 24068 10948 24078 11004
rect 31584 10976 31696 11004
rect 1922 10892 1932 10948
rect 1988 10892 1998 10948
rect 3266 10892 3276 10948
rect 3332 10892 3388 10948
rect 3444 10892 3454 10948
rect 4946 10892 4956 10948
rect 5012 10892 11900 10948
rect 11956 10892 11966 10948
rect 12226 10892 12236 10948
rect 12292 10892 12796 10948
rect 12852 10892 12862 10948
rect 13906 10892 13916 10948
rect 13972 10892 14140 10948
rect 14196 10892 14206 10948
rect 1932 10836 1988 10892
rect 1250 10780 1260 10836
rect 1316 10780 2716 10836
rect 2772 10780 2782 10836
rect 2930 10780 2940 10836
rect 2996 10780 3500 10836
rect 3556 10780 3566 10836
rect 7298 10780 7308 10836
rect 7364 10780 11004 10836
rect 11060 10780 11070 10836
rect 11554 10780 11564 10836
rect 11620 10780 14924 10836
rect 14980 10780 14990 10836
rect 1922 10668 1932 10724
rect 1988 10668 3612 10724
rect 3668 10668 3678 10724
rect 7074 10668 7084 10724
rect 7140 10668 8764 10724
rect 8820 10668 9436 10724
rect 9492 10668 9502 10724
rect 9650 10668 9660 10724
rect 9716 10668 22092 10724
rect 22148 10668 22158 10724
rect 0 10612 112 10640
rect 0 10556 7644 10612
rect 7700 10556 7710 10612
rect 8418 10556 8428 10612
rect 8484 10556 9660 10612
rect 9716 10556 9996 10612
rect 10052 10556 10062 10612
rect 11554 10556 11564 10612
rect 11620 10556 12908 10612
rect 12964 10556 12974 10612
rect 13458 10556 13468 10612
rect 13524 10556 14364 10612
rect 14420 10556 14430 10612
rect 20514 10556 20524 10612
rect 20580 10556 21196 10612
rect 21252 10556 21262 10612
rect 0 10528 112 10556
rect 3154 10444 3164 10500
rect 3220 10444 3948 10500
rect 4004 10444 4014 10500
rect 4274 10444 4284 10500
rect 4340 10444 5628 10500
rect 5684 10444 5694 10500
rect 5926 10444 5964 10500
rect 6020 10444 6030 10500
rect 7084 10444 10892 10500
rect 10948 10444 10958 10500
rect 11778 10444 11788 10500
rect 11844 10444 20748 10500
rect 20804 10444 20814 10500
rect 7084 10388 7140 10444
rect 802 10332 812 10388
rect 868 10332 1260 10388
rect 1316 10332 1326 10388
rect 2146 10332 2156 10388
rect 2212 10332 7140 10388
rect 7970 10332 7980 10388
rect 8036 10332 10332 10388
rect 10388 10332 10398 10388
rect 11890 10332 11900 10388
rect 11956 10332 12460 10388
rect 12516 10332 12526 10388
rect 14242 10332 14252 10388
rect 14308 10332 18508 10388
rect 18564 10332 18574 10388
rect 20626 10332 20636 10388
rect 20692 10332 20702 10388
rect 22978 10332 22988 10388
rect 23044 10332 25004 10388
rect 25060 10332 25070 10388
rect 2706 10220 2716 10276
rect 2772 10220 4284 10276
rect 4340 10220 4350 10276
rect 7522 10220 7532 10276
rect 7588 10220 16044 10276
rect 16100 10220 16110 10276
rect 0 10164 112 10192
rect 4454 10164 4464 10220
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4728 10164 4738 10220
rect 0 10108 812 10164
rect 868 10108 878 10164
rect 1810 10108 1820 10164
rect 1876 10108 2604 10164
rect 2660 10108 2670 10164
rect 6626 10108 6636 10164
rect 6692 10108 10668 10164
rect 10724 10108 10734 10164
rect 12450 10108 12460 10164
rect 12516 10108 15708 10164
rect 15764 10108 15774 10164
rect 0 10080 112 10108
rect 20636 10052 20692 10332
rect 24454 10164 24464 10220
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24728 10164 24738 10220
rect 31584 10164 31696 10192
rect 31490 10108 31500 10164
rect 31556 10108 31696 10164
rect 31584 10080 31696 10108
rect 2258 9996 2268 10052
rect 2324 9996 2492 10052
rect 2548 9996 2558 10052
rect 3154 9996 3164 10052
rect 3220 9996 4732 10052
rect 4788 9996 4798 10052
rect 5506 9996 5516 10052
rect 5572 9996 5964 10052
rect 6020 9996 6030 10052
rect 6178 9996 6188 10052
rect 6244 9996 9100 10052
rect 9156 9996 9166 10052
rect 9314 9996 9324 10052
rect 9380 9996 16716 10052
rect 16772 9996 16782 10052
rect 20636 9996 20804 10052
rect 21634 9996 21644 10052
rect 21700 9996 22428 10052
rect 22484 9996 22494 10052
rect 25106 9996 25116 10052
rect 25172 9996 25676 10052
rect 25732 9996 25742 10052
rect 20748 9940 20804 9996
rect 242 9884 252 9940
rect 308 9884 8876 9940
rect 8932 9884 8942 9940
rect 13570 9884 13580 9940
rect 13636 9884 18396 9940
rect 18452 9884 18462 9940
rect 20748 9884 26124 9940
rect 26180 9884 26190 9940
rect 690 9772 700 9828
rect 756 9772 8148 9828
rect 8306 9772 8316 9828
rect 8372 9772 9772 9828
rect 9828 9772 9838 9828
rect 9986 9772 9996 9828
rect 10052 9772 11788 9828
rect 11844 9772 12124 9828
rect 12180 9772 12190 9828
rect 13990 9772 14028 9828
rect 14084 9772 14094 9828
rect 16930 9772 16940 9828
rect 16996 9772 18060 9828
rect 18116 9772 18126 9828
rect 0 9716 112 9744
rect 8092 9716 8148 9772
rect 0 9660 4844 9716
rect 4900 9660 4910 9716
rect 8092 9660 15260 9716
rect 15316 9660 15326 9716
rect 21074 9660 21084 9716
rect 21140 9660 21308 9716
rect 21364 9660 21532 9716
rect 21588 9660 21598 9716
rect 0 9632 112 9660
rect 2034 9548 2044 9604
rect 2100 9548 6804 9604
rect 8194 9548 8204 9604
rect 8260 9548 11900 9604
rect 11956 9548 11966 9604
rect 6748 9492 6804 9548
rect 4722 9436 4732 9492
rect 4788 9436 6188 9492
rect 6244 9436 6254 9492
rect 6748 9436 10108 9492
rect 10164 9436 10174 9492
rect 10434 9436 10444 9492
rect 10500 9436 10668 9492
rect 10724 9436 10734 9492
rect 13682 9436 13692 9492
rect 13748 9436 14700 9492
rect 14756 9436 19180 9492
rect 19236 9436 19246 9492
rect 3794 9380 3804 9436
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 4068 9380 4078 9436
rect 23794 9380 23804 9436
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 24068 9380 24078 9436
rect 5618 9324 5628 9380
rect 5684 9324 15148 9380
rect 21970 9324 21980 9380
rect 22036 9324 22764 9380
rect 22820 9324 22830 9380
rect 0 9268 112 9296
rect 0 9212 1820 9268
rect 1876 9212 1886 9268
rect 3332 9212 14588 9268
rect 14644 9212 14654 9268
rect 0 9184 112 9212
rect 3332 9156 3388 9212
rect 15092 9156 15148 9324
rect 31584 9268 31696 9296
rect 21858 9212 21868 9268
rect 21924 9212 22428 9268
rect 22484 9212 22494 9268
rect 28242 9212 28252 9268
rect 28308 9212 31696 9268
rect 31584 9184 31696 9212
rect 2930 9100 2940 9156
rect 2996 9100 3388 9156
rect 4386 9100 4396 9156
rect 4452 9100 6076 9156
rect 6132 9100 6142 9156
rect 7074 9100 7084 9156
rect 7140 9100 9324 9156
rect 9380 9100 9390 9156
rect 10658 9100 10668 9156
rect 10724 9100 12572 9156
rect 12628 9100 12638 9156
rect 13542 9100 13580 9156
rect 13636 9100 14476 9156
rect 14532 9100 14542 9156
rect 15092 9100 17276 9156
rect 17332 9100 17342 9156
rect 18834 9100 18844 9156
rect 18900 9100 22316 9156
rect 22372 9100 24556 9156
rect 24612 9100 24892 9156
rect 24948 9100 24958 9156
rect 2706 8988 2716 9044
rect 2772 8988 2828 9044
rect 2884 8988 2894 9044
rect 3938 8988 3948 9044
rect 4004 8988 4284 9044
rect 4340 8988 5068 9044
rect 5124 8988 5134 9044
rect 5254 8988 5292 9044
rect 5348 8988 5358 9044
rect 5954 8988 5964 9044
rect 6020 8988 6860 9044
rect 6916 8988 6926 9044
rect 10994 8988 11004 9044
rect 11060 8988 11070 9044
rect 12114 8988 12124 9044
rect 12180 8988 13916 9044
rect 13972 8988 13982 9044
rect 14354 8988 14364 9044
rect 14420 8988 15484 9044
rect 15540 8988 16828 9044
rect 16884 8988 16894 9044
rect 19170 8988 19180 9044
rect 19236 8988 20860 9044
rect 20916 8988 21644 9044
rect 21700 8988 21868 9044
rect 21924 8988 21934 9044
rect 11004 8932 11060 8988
rect 4274 8876 4284 8932
rect 4340 8876 7868 8932
rect 7924 8876 7934 8932
rect 11004 8876 13020 8932
rect 13076 8876 14588 8932
rect 14644 8876 14654 8932
rect 17378 8876 17388 8932
rect 17444 8876 24108 8932
rect 24164 8876 24174 8932
rect 0 8820 112 8848
rect 0 8764 3612 8820
rect 3668 8764 3678 8820
rect 4284 8764 7420 8820
rect 7476 8764 7486 8820
rect 13122 8764 13132 8820
rect 13188 8764 15484 8820
rect 15540 8764 15550 8820
rect 20066 8764 20076 8820
rect 20132 8764 21644 8820
rect 21700 8764 21710 8820
rect 0 8736 112 8764
rect 4284 8708 4340 8764
rect 2930 8652 2940 8708
rect 2996 8652 4340 8708
rect 8642 8652 8652 8708
rect 8708 8652 15148 8708
rect 18498 8652 18508 8708
rect 18564 8652 18956 8708
rect 19012 8652 19022 8708
rect 4454 8596 4464 8652
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4728 8596 4738 8652
rect 15092 8596 15148 8652
rect 24454 8596 24464 8652
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24728 8596 24738 8652
rect 1250 8540 1260 8596
rect 1316 8540 3276 8596
rect 3332 8540 3342 8596
rect 8418 8540 8428 8596
rect 8484 8540 8764 8596
rect 8820 8540 8830 8596
rect 9398 8540 9436 8596
rect 9492 8540 9502 8596
rect 11106 8540 11116 8596
rect 11172 8540 11340 8596
rect 11396 8540 11406 8596
rect 15092 8540 21196 8596
rect 21252 8540 21262 8596
rect 21746 8540 21756 8596
rect 21812 8540 21822 8596
rect 1474 8428 1484 8484
rect 1540 8428 4956 8484
rect 5012 8428 5022 8484
rect 8082 8428 8092 8484
rect 8148 8428 10220 8484
rect 10276 8428 10286 8484
rect 10994 8428 11004 8484
rect 11060 8428 17388 8484
rect 17444 8428 17454 8484
rect 0 8372 112 8400
rect 0 8316 7308 8372
rect 7364 8316 7374 8372
rect 7522 8316 7532 8372
rect 7588 8316 7644 8372
rect 7700 8316 7710 8372
rect 8418 8316 8428 8372
rect 8484 8316 9772 8372
rect 9828 8316 9838 8372
rect 9986 8316 9996 8372
rect 10052 8316 10780 8372
rect 10836 8316 10846 8372
rect 12114 8316 12124 8372
rect 12180 8316 13020 8372
rect 13076 8316 13086 8372
rect 17938 8316 17948 8372
rect 18004 8316 19068 8372
rect 19124 8316 19134 8372
rect 19478 8316 19516 8372
rect 19572 8316 19582 8372
rect 0 8288 112 8316
rect 690 8204 700 8260
rect 756 8204 1092 8260
rect 1362 8204 1372 8260
rect 1428 8204 1484 8260
rect 1540 8204 1550 8260
rect 3490 8204 3500 8260
rect 3556 8204 4956 8260
rect 5012 8204 5022 8260
rect 5954 8204 5964 8260
rect 6020 8204 8204 8260
rect 8260 8204 8270 8260
rect 9314 8204 9324 8260
rect 9380 8204 12796 8260
rect 12852 8204 12862 8260
rect 13346 8204 13356 8260
rect 13412 8204 14028 8260
rect 14084 8204 14588 8260
rect 14644 8204 14654 8260
rect 19730 8204 19740 8260
rect 19796 8204 19964 8260
rect 20020 8204 20030 8260
rect 1036 8148 1092 8204
rect 21756 8148 21812 8540
rect 31584 8372 31696 8400
rect 31378 8316 31388 8372
rect 31444 8316 31696 8372
rect 31584 8288 31696 8316
rect 1026 8092 1036 8148
rect 1092 8092 1102 8148
rect 3602 8092 3612 8148
rect 3668 8092 6636 8148
rect 6692 8092 6702 8148
rect 9212 8092 17556 8148
rect 18386 8092 18396 8148
rect 18452 8092 21084 8148
rect 21140 8092 21420 8148
rect 21476 8092 21486 8148
rect 21756 8092 23548 8148
rect 23604 8092 23614 8148
rect 3332 7980 7980 8036
rect 8036 7980 8046 8036
rect 8614 7980 8652 8036
rect 8708 7980 8718 8036
rect 0 7924 112 7952
rect 3332 7924 3388 7980
rect 9212 7924 9268 8092
rect 9762 7980 9772 8036
rect 9828 7980 12908 8036
rect 12964 7980 13580 8036
rect 13636 7980 13646 8036
rect 16258 7980 16268 8036
rect 16324 7980 16828 8036
rect 16884 7980 16894 8036
rect 17500 7924 17556 8092
rect 17714 7980 17724 8036
rect 17780 7980 21756 8036
rect 21812 7980 21822 8036
rect 22194 7980 22204 8036
rect 22260 7980 25452 8036
rect 25508 7980 25518 8036
rect 0 7868 3388 7924
rect 4946 7868 4956 7924
rect 5012 7868 9268 7924
rect 11554 7868 11564 7924
rect 11620 7868 13804 7924
rect 13860 7868 15596 7924
rect 15652 7868 15662 7924
rect 17500 7868 22876 7924
rect 22932 7868 22942 7924
rect 0 7840 112 7868
rect 3794 7812 3804 7868
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 4068 7812 4078 7868
rect 23794 7812 23804 7868
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 24068 7812 24078 7868
rect 4722 7756 4732 7812
rect 4788 7756 9212 7812
rect 9268 7756 9278 7812
rect 10994 7756 11004 7812
rect 11060 7756 16604 7812
rect 16660 7756 16940 7812
rect 16996 7756 17006 7812
rect 20066 7756 20076 7812
rect 20132 7756 20748 7812
rect 20804 7756 20814 7812
rect 21634 7756 21644 7812
rect 21700 7756 23660 7812
rect 23716 7756 23726 7812
rect 2818 7644 2828 7700
rect 2884 7644 3388 7700
rect 3444 7644 3454 7700
rect 6402 7644 6412 7700
rect 6468 7644 6748 7700
rect 6804 7644 10220 7700
rect 10276 7644 18732 7700
rect 18788 7644 21140 7700
rect 21298 7644 21308 7700
rect 21364 7644 25004 7700
rect 25060 7644 25070 7700
rect 21084 7588 21140 7644
rect 6066 7532 6076 7588
rect 6132 7532 9380 7588
rect 9538 7532 9548 7588
rect 9604 7532 10556 7588
rect 10612 7532 11004 7588
rect 11060 7532 11070 7588
rect 13570 7532 13580 7588
rect 13636 7532 20412 7588
rect 20468 7532 20478 7588
rect 21084 7532 21420 7588
rect 21476 7532 21486 7588
rect 23650 7532 23660 7588
rect 23716 7532 28588 7588
rect 28644 7532 28654 7588
rect 0 7476 112 7504
rect 9324 7476 9380 7532
rect 31584 7476 31696 7504
rect 0 7420 6636 7476
rect 6692 7420 6702 7476
rect 7410 7420 7420 7476
rect 7476 7420 7644 7476
rect 7700 7420 9100 7476
rect 9156 7420 9166 7476
rect 9324 7420 9436 7476
rect 9492 7420 9772 7476
rect 9828 7420 13356 7476
rect 13412 7420 13422 7476
rect 13682 7420 13692 7476
rect 13748 7420 15372 7476
rect 15428 7420 15484 7476
rect 15540 7420 15550 7476
rect 18834 7420 18844 7476
rect 18900 7420 19404 7476
rect 19460 7420 20580 7476
rect 31266 7420 31276 7476
rect 31332 7420 31696 7476
rect 0 7392 112 7420
rect 20524 7364 20580 7420
rect 31584 7392 31696 7420
rect 2230 7308 2268 7364
rect 2324 7308 2334 7364
rect 3378 7308 3388 7364
rect 3444 7308 11788 7364
rect 11844 7308 11854 7364
rect 13234 7308 13244 7364
rect 13300 7308 18956 7364
rect 19012 7308 19022 7364
rect 20514 7308 20524 7364
rect 20580 7308 20590 7364
rect 24882 7308 24892 7364
rect 24948 7308 26572 7364
rect 26628 7308 26638 7364
rect 7970 7196 7980 7252
rect 8036 7196 11004 7252
rect 11060 7196 11070 7252
rect 12226 7196 12236 7252
rect 12292 7196 13916 7252
rect 13972 7196 13982 7252
rect 14140 7196 17836 7252
rect 17892 7196 17902 7252
rect 14140 7140 14196 7196
rect 10770 7084 10780 7140
rect 10836 7084 14196 7140
rect 15092 7084 17500 7140
rect 17556 7084 17566 7140
rect 20066 7084 20076 7140
rect 20132 7084 20636 7140
rect 20692 7084 20702 7140
rect 0 7028 112 7056
rect 4454 7028 4464 7084
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4728 7028 4738 7084
rect 0 6972 2492 7028
rect 2548 6972 2558 7028
rect 5954 6972 5964 7028
rect 6020 6972 6972 7028
rect 7028 6972 7038 7028
rect 13570 6972 13580 7028
rect 13636 6972 14140 7028
rect 14196 6972 14206 7028
rect 0 6944 112 6972
rect 15092 6916 15148 7084
rect 24454 7028 24464 7084
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 24728 7028 24738 7084
rect 20290 6972 20300 7028
rect 20356 6972 22876 7028
rect 22932 6972 22942 7028
rect 25750 6972 25788 7028
rect 25844 6972 25854 7028
rect 4722 6860 4732 6916
rect 4788 6860 5628 6916
rect 5684 6860 5694 6916
rect 5842 6860 5852 6916
rect 5908 6860 9436 6916
rect 9492 6860 9502 6916
rect 11442 6860 11452 6916
rect 11508 6860 15148 6916
rect 19730 6860 19740 6916
rect 19796 6860 19964 6916
rect 20020 6860 20030 6916
rect 23650 6860 23660 6916
rect 23716 6860 27356 6916
rect 27412 6860 27422 6916
rect 3938 6748 3948 6804
rect 4004 6748 4284 6804
rect 4340 6748 5740 6804
rect 5796 6748 5806 6804
rect 6962 6748 6972 6804
rect 7028 6748 7308 6804
rect 7364 6748 7374 6804
rect 8316 6748 8428 6804
rect 8484 6748 8652 6804
rect 8708 6748 8718 6804
rect 9202 6748 9212 6804
rect 9268 6748 15148 6804
rect 15204 6748 15214 6804
rect 15474 6748 15484 6804
rect 15540 6748 18060 6804
rect 18116 6748 18126 6804
rect 20514 6748 20524 6804
rect 20580 6748 25788 6804
rect 25844 6748 25854 6804
rect 8316 6692 8372 6748
rect 1334 6636 1372 6692
rect 1428 6636 1438 6692
rect 2118 6636 2156 6692
rect 2212 6636 2222 6692
rect 2370 6636 2380 6692
rect 2436 6636 2474 6692
rect 3378 6636 3388 6692
rect 3444 6636 3482 6692
rect 4050 6636 4060 6692
rect 4116 6636 7980 6692
rect 8036 6636 8046 6692
rect 8306 6636 8316 6692
rect 8372 6636 8382 6692
rect 9538 6636 9548 6692
rect 9604 6636 10108 6692
rect 10164 6636 10174 6692
rect 12450 6636 12460 6692
rect 12516 6636 14364 6692
rect 14420 6636 14430 6692
rect 16146 6636 16156 6692
rect 16212 6636 19068 6692
rect 19124 6636 19134 6692
rect 19618 6636 19628 6692
rect 19684 6636 21420 6692
rect 21476 6636 21486 6692
rect 22082 6636 22092 6692
rect 22148 6636 22988 6692
rect 23044 6636 23054 6692
rect 0 6580 112 6608
rect 19628 6580 19684 6636
rect 31584 6580 31696 6608
rect 0 6524 6412 6580
rect 6468 6524 6478 6580
rect 6626 6524 6636 6580
rect 6692 6524 8092 6580
rect 8148 6524 8158 6580
rect 9762 6524 9772 6580
rect 9828 6524 9996 6580
rect 10052 6524 10062 6580
rect 10882 6524 10892 6580
rect 10948 6524 13580 6580
rect 13636 6524 13646 6580
rect 14242 6524 14252 6580
rect 14308 6524 15932 6580
rect 15988 6524 16604 6580
rect 16660 6524 17612 6580
rect 17668 6524 17678 6580
rect 18274 6524 18284 6580
rect 18340 6524 19180 6580
rect 19236 6524 19684 6580
rect 20178 6524 20188 6580
rect 20244 6524 20412 6580
rect 20468 6524 20478 6580
rect 22866 6524 22876 6580
rect 22932 6524 25564 6580
rect 25620 6524 25630 6580
rect 27682 6524 27692 6580
rect 27748 6524 31696 6580
rect 0 6496 112 6524
rect 31584 6496 31696 6524
rect 1698 6412 1708 6468
rect 1764 6412 7868 6468
rect 7924 6412 7934 6468
rect 12898 6412 12908 6468
rect 12964 6412 14476 6468
rect 14532 6412 14812 6468
rect 14868 6412 14878 6468
rect 22194 6412 22204 6468
rect 22260 6412 23212 6468
rect 23268 6412 23278 6468
rect 23436 6412 27468 6468
rect 27524 6412 27534 6468
rect 23436 6356 23492 6412
rect 1810 6300 1820 6356
rect 1876 6300 1886 6356
rect 13570 6300 13580 6356
rect 13636 6300 14700 6356
rect 14756 6300 14766 6356
rect 16930 6300 16940 6356
rect 16996 6300 23492 6356
rect 1820 6244 1876 6300
rect 3794 6244 3804 6300
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 4068 6244 4078 6300
rect 23794 6244 23804 6300
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 24068 6244 24078 6300
rect 1820 6188 2268 6244
rect 2324 6188 2334 6244
rect 4946 6188 4956 6244
rect 5012 6188 22988 6244
rect 23044 6188 23054 6244
rect 0 6132 112 6160
rect 0 6076 8876 6132
rect 8932 6076 8942 6132
rect 21746 6076 21756 6132
rect 21812 6076 24108 6132
rect 24164 6076 24174 6132
rect 0 6048 112 6076
rect 3378 5964 3388 6020
rect 3444 5964 6132 6020
rect 10322 5964 10332 6020
rect 10388 5964 23212 6020
rect 23268 5964 23278 6020
rect 6076 5908 6132 5964
rect 3490 5852 3500 5908
rect 3556 5852 3836 5908
rect 3892 5852 3902 5908
rect 5030 5852 5068 5908
rect 5124 5852 5134 5908
rect 6066 5852 6076 5908
rect 6132 5852 6972 5908
rect 7028 5852 7038 5908
rect 7858 5852 7868 5908
rect 7924 5852 8316 5908
rect 8372 5852 8382 5908
rect 15474 5852 15484 5908
rect 15540 5852 15596 5908
rect 15652 5852 15662 5908
rect 18834 5852 18844 5908
rect 18900 5852 19964 5908
rect 20020 5852 21868 5908
rect 21924 5852 21934 5908
rect 22306 5852 22316 5908
rect 22372 5852 24556 5908
rect 24612 5852 25340 5908
rect 25396 5852 25406 5908
rect 25554 5852 25564 5908
rect 25620 5852 29540 5908
rect 2716 5740 4172 5796
rect 4228 5740 4238 5796
rect 7634 5740 7644 5796
rect 7700 5740 9100 5796
rect 9156 5740 9166 5796
rect 10332 5740 26908 5796
rect 26964 5740 26974 5796
rect 0 5684 112 5712
rect 2716 5684 2772 5740
rect 10332 5684 10388 5740
rect 29484 5684 29540 5852
rect 31584 5684 31696 5712
rect 0 5628 252 5684
rect 308 5628 318 5684
rect 2146 5628 2156 5684
rect 2212 5628 2716 5684
rect 2772 5628 2782 5684
rect 3042 5628 3052 5684
rect 3108 5628 5908 5684
rect 6066 5628 6076 5684
rect 6132 5628 10388 5684
rect 10546 5628 10556 5684
rect 10612 5628 11900 5684
rect 11956 5628 11966 5684
rect 14690 5628 14700 5684
rect 14756 5628 18844 5684
rect 18900 5628 18910 5684
rect 19058 5628 19068 5684
rect 19124 5628 29260 5684
rect 29316 5628 29326 5684
rect 29484 5628 31696 5684
rect 0 5600 112 5628
rect 5852 5572 5908 5628
rect 31584 5600 31696 5628
rect 5852 5516 6412 5572
rect 6468 5516 9660 5572
rect 9716 5516 9726 5572
rect 9986 5516 9996 5572
rect 10052 5516 14924 5572
rect 14980 5516 15484 5572
rect 15540 5516 16828 5572
rect 16884 5516 16894 5572
rect 19394 5516 19404 5572
rect 19460 5516 20412 5572
rect 20468 5516 20478 5572
rect 20738 5516 20748 5572
rect 20804 5516 21644 5572
rect 21700 5516 21710 5572
rect 4454 5460 4464 5516
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4728 5460 4738 5516
rect 24454 5460 24464 5516
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24728 5460 24738 5516
rect 5068 5404 7532 5460
rect 7588 5404 7598 5460
rect 9090 5404 9100 5460
rect 9156 5404 9548 5460
rect 9604 5404 9614 5460
rect 10630 5404 10668 5460
rect 10724 5404 10734 5460
rect 10882 5404 10892 5460
rect 10948 5404 13468 5460
rect 13524 5404 13534 5460
rect 17826 5404 17836 5460
rect 17892 5404 19740 5460
rect 19796 5404 19806 5460
rect 20850 5404 20860 5460
rect 20916 5404 22316 5460
rect 22372 5404 22382 5460
rect 25106 5404 25116 5460
rect 25172 5404 25228 5460
rect 25284 5404 25294 5460
rect 5068 5348 5124 5404
rect 466 5292 476 5348
rect 532 5292 1036 5348
rect 1092 5292 1102 5348
rect 1250 5292 1260 5348
rect 1316 5292 1372 5348
rect 1428 5292 1438 5348
rect 2006 5292 2044 5348
rect 2100 5292 2110 5348
rect 2706 5292 2716 5348
rect 2772 5292 5124 5348
rect 5282 5292 5292 5348
rect 5348 5292 7084 5348
rect 7140 5292 7150 5348
rect 8082 5292 8092 5348
rect 8148 5292 13244 5348
rect 13300 5292 13310 5348
rect 13570 5292 13580 5348
rect 13636 5292 14028 5348
rect 14084 5292 14094 5348
rect 15334 5292 15372 5348
rect 15428 5292 15438 5348
rect 15698 5292 15708 5348
rect 15764 5292 22428 5348
rect 22484 5292 22494 5348
rect 23286 5292 23324 5348
rect 23380 5292 23390 5348
rect 23986 5292 23996 5348
rect 24052 5292 25116 5348
rect 25172 5292 25182 5348
rect 0 5236 112 5264
rect 0 5180 5852 5236
rect 5908 5180 5918 5236
rect 6402 5180 6412 5236
rect 6468 5180 6748 5236
rect 6804 5180 6814 5236
rect 7298 5180 7308 5236
rect 7364 5180 12236 5236
rect 12292 5180 12302 5236
rect 15922 5180 15932 5236
rect 15988 5180 26348 5236
rect 26404 5180 26414 5236
rect 0 5152 112 5180
rect 1698 5068 1708 5124
rect 1764 5068 2492 5124
rect 2548 5068 2558 5124
rect 4162 5068 4172 5124
rect 4228 5068 4844 5124
rect 4900 5068 7868 5124
rect 7924 5068 7934 5124
rect 8092 5068 8652 5124
rect 8708 5068 9548 5124
rect 9604 5068 9614 5124
rect 11218 5068 11228 5124
rect 11284 5068 12908 5124
rect 12964 5068 12974 5124
rect 13346 5068 13356 5124
rect 13412 5068 13916 5124
rect 13972 5068 13982 5124
rect 14214 5068 14252 5124
rect 14308 5068 14318 5124
rect 15362 5068 15372 5124
rect 15428 5068 16492 5124
rect 16548 5068 16558 5124
rect 17714 5068 17724 5124
rect 17780 5068 18284 5124
rect 18340 5068 18350 5124
rect 22418 5068 22428 5124
rect 22484 5068 23436 5124
rect 23492 5068 23502 5124
rect 24210 5068 24220 5124
rect 24276 5068 27244 5124
rect 27300 5068 27310 5124
rect 8092 5012 8148 5068
rect 3154 4956 3164 5012
rect 3220 4956 8148 5012
rect 8306 4956 8316 5012
rect 8372 4956 17052 5012
rect 17108 4956 17118 5012
rect 19842 4956 19852 5012
rect 19908 4956 22988 5012
rect 23044 4956 23054 5012
rect 3332 4844 8428 4900
rect 8484 4844 8494 4900
rect 15138 4844 15148 4900
rect 15204 4844 18956 4900
rect 19012 4844 19022 4900
rect 19954 4844 19964 4900
rect 20020 4844 27356 4900
rect 27412 4844 27422 4900
rect 0 4788 112 4816
rect 3332 4788 3388 4844
rect 31584 4788 31696 4816
rect 0 4732 3388 4788
rect 9762 4732 9772 4788
rect 9828 4732 22988 4788
rect 23044 4732 23054 4788
rect 25106 4732 25116 4788
rect 25172 4732 25564 4788
rect 25620 4732 25630 4788
rect 27682 4732 27692 4788
rect 27748 4732 31696 4788
rect 0 4704 112 4732
rect 3794 4676 3804 4732
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 4068 4676 4078 4732
rect 23794 4676 23804 4732
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 24068 4676 24078 4732
rect 31584 4704 31696 4732
rect 2706 4620 2716 4676
rect 2772 4620 2828 4676
rect 2884 4620 2894 4676
rect 9090 4620 9100 4676
rect 9156 4620 9324 4676
rect 9380 4620 9390 4676
rect 11526 4620 11564 4676
rect 11620 4620 11630 4676
rect 15092 4620 20076 4676
rect 20132 4620 20142 4676
rect 20290 4620 20300 4676
rect 20356 4620 20804 4676
rect 22754 4620 22764 4676
rect 22820 4620 23436 4676
rect 23492 4620 23502 4676
rect 1148 4508 5404 4564
rect 5460 4508 5470 4564
rect 9202 4508 9212 4564
rect 9268 4508 13580 4564
rect 13636 4508 13646 4564
rect 0 4340 112 4368
rect 1148 4340 1204 4508
rect 15092 4452 15148 4620
rect 15586 4508 15596 4564
rect 15652 4508 16268 4564
rect 16324 4508 16334 4564
rect 17154 4508 17164 4564
rect 17220 4508 20692 4564
rect 2034 4396 2044 4452
rect 2100 4396 15148 4452
rect 17164 4340 17220 4508
rect 18722 4396 18732 4452
rect 18788 4396 19628 4452
rect 19684 4396 19694 4452
rect 20636 4340 20692 4508
rect 20748 4452 20804 4620
rect 21522 4508 21532 4564
rect 21588 4508 26908 4564
rect 26852 4452 26908 4508
rect 20748 4396 23660 4452
rect 23716 4396 23726 4452
rect 26450 4396 26460 4452
rect 26516 4396 26526 4452
rect 26852 4396 31668 4452
rect 0 4284 1204 4340
rect 1362 4284 1372 4340
rect 1428 4284 1932 4340
rect 1988 4284 1998 4340
rect 8866 4284 8876 4340
rect 8932 4284 10556 4340
rect 10612 4284 10622 4340
rect 11330 4284 11340 4340
rect 11396 4284 11564 4340
rect 11620 4284 11630 4340
rect 12198 4284 12236 4340
rect 12292 4284 12302 4340
rect 13318 4284 13356 4340
rect 13412 4284 13422 4340
rect 16258 4284 16268 4340
rect 16324 4284 17220 4340
rect 18246 4284 18284 4340
rect 18340 4284 18350 4340
rect 19282 4284 19292 4340
rect 19348 4284 20412 4340
rect 20468 4284 20478 4340
rect 20636 4284 22428 4340
rect 22484 4284 22494 4340
rect 23762 4284 23772 4340
rect 23828 4284 25116 4340
rect 25172 4284 25182 4340
rect 0 4256 112 4284
rect 26460 4228 26516 4396
rect 354 4172 364 4228
rect 420 4172 1036 4228
rect 1092 4172 1102 4228
rect 1698 4172 1708 4228
rect 1764 4172 2604 4228
rect 2660 4172 2670 4228
rect 5394 4172 5404 4228
rect 5460 4172 6524 4228
rect 6580 4172 6590 4228
rect 8642 4172 8652 4228
rect 8708 4172 21476 4228
rect 21858 4172 21868 4228
rect 21924 4172 24108 4228
rect 24164 4172 24174 4228
rect 24658 4172 24668 4228
rect 24724 4172 25004 4228
rect 25060 4172 25070 4228
rect 26338 4172 26348 4228
rect 26404 4172 26516 4228
rect 21420 4116 21476 4172
rect 31612 4116 31668 4396
rect 3266 4060 3276 4116
rect 3332 4060 5740 4116
rect 5796 4060 5806 4116
rect 6962 4060 6972 4116
rect 7028 4060 7980 4116
rect 8036 4060 8046 4116
rect 9538 4060 9548 4116
rect 9604 4060 11228 4116
rect 11284 4060 11294 4116
rect 15932 4060 21196 4116
rect 21252 4060 21262 4116
rect 21410 4060 21420 4116
rect 21476 4060 21486 4116
rect 21644 4060 26572 4116
rect 26628 4060 26638 4116
rect 31388 4060 31668 4116
rect 15932 4004 15988 4060
rect 21644 4004 21700 4060
rect 4946 3948 4956 4004
rect 5012 3948 9660 4004
rect 9716 3948 9726 4004
rect 10658 3948 10668 4004
rect 10724 3948 14476 4004
rect 14532 3948 15932 4004
rect 15988 3948 15998 4004
rect 18834 3948 18844 4004
rect 18900 3948 21700 4004
rect 24892 3948 25452 4004
rect 25508 3948 25518 4004
rect 0 3892 112 3920
rect 4454 3892 4464 3948
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4728 3892 4738 3948
rect 24454 3892 24464 3948
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24728 3892 24738 3948
rect 0 3836 1764 3892
rect 6066 3836 6076 3892
rect 6132 3836 12964 3892
rect 21186 3836 21196 3892
rect 21252 3836 22540 3892
rect 22596 3836 22606 3892
rect 0 3808 112 3836
rect 1708 3668 1764 3836
rect 12908 3780 12964 3836
rect 24892 3780 24948 3948
rect 31388 3892 31444 4060
rect 31584 3892 31696 3920
rect 26646 3836 26684 3892
rect 26740 3836 26750 3892
rect 31388 3836 31696 3892
rect 31584 3808 31696 3836
rect 2034 3724 2044 3780
rect 2100 3724 3556 3780
rect 5394 3724 5404 3780
rect 5460 3724 6300 3780
rect 6356 3724 6366 3780
rect 9090 3724 9100 3780
rect 9156 3724 9772 3780
rect 9828 3724 9838 3780
rect 10882 3724 10892 3780
rect 10948 3724 12684 3780
rect 12740 3724 12750 3780
rect 12908 3724 22876 3780
rect 22932 3724 22942 3780
rect 23510 3724 23548 3780
rect 23604 3724 23614 3780
rect 24882 3724 24892 3780
rect 24948 3724 24958 3780
rect 25218 3724 25228 3780
rect 25284 3724 25294 3780
rect 3500 3668 3556 3724
rect 25228 3668 25284 3724
rect 1708 3612 3388 3668
rect 3500 3612 18396 3668
rect 18452 3612 18462 3668
rect 20514 3612 20524 3668
rect 20580 3612 25284 3668
rect 3332 3556 3388 3612
rect 2258 3500 2268 3556
rect 2324 3500 3164 3556
rect 3220 3500 3230 3556
rect 3332 3500 9212 3556
rect 9268 3500 9278 3556
rect 10994 3500 11004 3556
rect 11060 3500 11228 3556
rect 11284 3500 11452 3556
rect 11508 3500 11518 3556
rect 11778 3500 11788 3556
rect 11844 3500 13692 3556
rect 13748 3500 13758 3556
rect 14466 3500 14476 3556
rect 14532 3500 14588 3556
rect 14644 3500 14654 3556
rect 16818 3500 16828 3556
rect 16884 3500 17164 3556
rect 17220 3500 17230 3556
rect 21074 3500 21084 3556
rect 21140 3500 23772 3556
rect 23828 3500 23838 3556
rect 25890 3500 25900 3556
rect 25956 3500 25966 3556
rect 26758 3500 26796 3556
rect 26852 3500 26862 3556
rect 0 3444 112 3472
rect 25900 3444 25956 3500
rect 0 3388 6300 3444
rect 6356 3388 6366 3444
rect 8306 3388 8316 3444
rect 8372 3388 13356 3444
rect 13412 3388 13422 3444
rect 13580 3388 15148 3444
rect 15204 3388 17724 3444
rect 17780 3388 17790 3444
rect 19394 3388 19404 3444
rect 19460 3388 25956 3444
rect 0 3360 112 3388
rect 13580 3332 13636 3388
rect 1586 3276 1596 3332
rect 1652 3276 5852 3332
rect 5908 3276 5918 3332
rect 6066 3276 6076 3332
rect 6132 3276 7196 3332
rect 7252 3276 7262 3332
rect 9314 3276 9324 3332
rect 9380 3276 10220 3332
rect 10276 3276 10286 3332
rect 10882 3276 10892 3332
rect 10948 3276 13636 3332
rect 23874 3276 23884 3332
rect 23940 3276 28476 3332
rect 28532 3276 28542 3332
rect 9426 3164 9436 3220
rect 9492 3164 20748 3220
rect 20804 3164 20814 3220
rect 22978 3164 22988 3220
rect 23044 3164 23548 3220
rect 25218 3164 25228 3220
rect 25284 3164 26012 3220
rect 26068 3164 26078 3220
rect 3794 3108 3804 3164
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 4068 3108 4078 3164
rect 4162 3052 4172 3108
rect 4228 3052 8988 3108
rect 9044 3052 9054 3108
rect 13458 3052 13468 3108
rect 13524 3052 16716 3108
rect 16772 3052 16782 3108
rect 17612 3052 20860 3108
rect 20916 3052 23100 3108
rect 23156 3052 23166 3108
rect 0 2996 112 3024
rect 17612 2996 17668 3052
rect 23492 2996 23548 3164
rect 23794 3108 23804 3164
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 24068 3108 24078 3164
rect 31584 2996 31696 3024
rect 0 2940 2548 2996
rect 3378 2940 3388 2996
rect 3444 2940 4844 2996
rect 4900 2940 4910 2996
rect 5180 2940 9212 2996
rect 9268 2940 9278 2996
rect 10098 2940 10108 2996
rect 10164 2940 11340 2996
rect 11396 2940 11406 2996
rect 13234 2940 13244 2996
rect 13300 2940 13692 2996
rect 13748 2940 14028 2996
rect 14084 2940 14094 2996
rect 16566 2940 16604 2996
rect 16660 2940 17612 2996
rect 17668 2940 17678 2996
rect 18610 2940 18620 2996
rect 18676 2940 19628 2996
rect 19684 2940 19694 2996
rect 23492 2940 23660 2996
rect 23716 2940 24556 2996
rect 24612 2940 25004 2996
rect 25060 2940 25900 2996
rect 25956 2940 25966 2996
rect 28578 2940 28588 2996
rect 28644 2940 31696 2996
rect 0 2912 112 2940
rect 2492 2884 2548 2940
rect 2492 2828 4956 2884
rect 5012 2828 5022 2884
rect 3602 2716 3612 2772
rect 3668 2716 3836 2772
rect 3892 2716 3902 2772
rect 5180 2660 5236 2940
rect 31584 2912 31696 2940
rect 7970 2828 7980 2884
rect 8036 2828 15036 2884
rect 15092 2828 15102 2884
rect 16706 2828 16716 2884
rect 16772 2828 17052 2884
rect 17108 2828 21420 2884
rect 21476 2828 21486 2884
rect 7718 2716 7756 2772
rect 7812 2716 7822 2772
rect 8082 2716 8092 2772
rect 8148 2716 8652 2772
rect 8708 2716 8718 2772
rect 9202 2716 9212 2772
rect 9268 2716 14140 2772
rect 14196 2716 14206 2772
rect 15586 2716 15596 2772
rect 15652 2716 15708 2772
rect 15764 2716 15774 2772
rect 18582 2716 18620 2772
rect 18676 2716 18686 2772
rect 20962 2716 20972 2772
rect 21028 2716 21756 2772
rect 21812 2716 22316 2772
rect 22372 2716 22382 2772
rect 25414 2716 25452 2772
rect 25508 2716 25518 2772
rect 26086 2716 26124 2772
rect 26180 2716 26190 2772
rect 1596 2604 3164 2660
rect 3220 2604 3230 2660
rect 3378 2604 3388 2660
rect 3444 2604 5236 2660
rect 5702 2604 5740 2660
rect 5796 2604 5806 2660
rect 11554 2604 11564 2660
rect 11620 2604 11676 2660
rect 11732 2604 11742 2660
rect 14018 2604 14028 2660
rect 14084 2604 14700 2660
rect 14756 2604 14766 2660
rect 18274 2604 18284 2660
rect 18340 2604 25844 2660
rect 0 2548 112 2576
rect 1596 2548 1652 2604
rect 25788 2548 25844 2604
rect 0 2492 1652 2548
rect 1810 2492 1820 2548
rect 1876 2492 7532 2548
rect 7588 2492 7598 2548
rect 11554 2492 11564 2548
rect 11620 2492 11788 2548
rect 11844 2492 11854 2548
rect 14102 2492 14140 2548
rect 14196 2492 14206 2548
rect 16930 2492 16940 2548
rect 16996 2492 19292 2548
rect 19348 2492 19358 2548
rect 19842 2492 19852 2548
rect 19908 2492 21252 2548
rect 21410 2492 21420 2548
rect 21476 2492 24108 2548
rect 24164 2492 24174 2548
rect 25778 2492 25788 2548
rect 25844 2492 25854 2548
rect 0 2464 112 2492
rect 21196 2436 21252 2492
rect 5282 2380 5292 2436
rect 5348 2380 5628 2436
rect 5684 2380 6412 2436
rect 6468 2380 10220 2436
rect 10276 2380 10286 2436
rect 10546 2380 10556 2436
rect 10612 2380 20188 2436
rect 20244 2380 20254 2436
rect 21196 2380 22876 2436
rect 22932 2380 23660 2436
rect 23716 2380 23726 2436
rect 4454 2324 4464 2380
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4728 2324 4738 2380
rect 24454 2324 24464 2380
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24728 2324 24738 2380
rect 2454 2268 2492 2324
rect 2548 2268 2558 2324
rect 8306 2268 8316 2324
rect 8372 2268 15260 2324
rect 15316 2268 15326 2324
rect 18610 2268 18620 2324
rect 18676 2268 23548 2324
rect 23604 2268 23614 2324
rect 24882 2268 24892 2324
rect 24948 2268 25228 2324
rect 25284 2268 25294 2324
rect 25778 2268 25788 2324
rect 25844 2268 26684 2324
rect 26740 2268 26750 2324
rect 1698 2156 1708 2212
rect 1764 2156 2828 2212
rect 2884 2156 3444 2212
rect 4946 2156 4956 2212
rect 5012 2156 8428 2212
rect 8484 2156 8494 2212
rect 11778 2156 11788 2212
rect 11844 2156 12908 2212
rect 12964 2156 12974 2212
rect 15670 2156 15708 2212
rect 15764 2156 15774 2212
rect 17490 2156 17500 2212
rect 17556 2156 18172 2212
rect 18228 2156 21868 2212
rect 21924 2156 21934 2212
rect 22054 2156 22092 2212
rect 22148 2156 22158 2212
rect 22642 2156 22652 2212
rect 22708 2156 23100 2212
rect 23156 2156 25452 2212
rect 25508 2156 25518 2212
rect 26310 2156 26348 2212
rect 26404 2156 26414 2212
rect 0 2100 112 2128
rect 3388 2100 3444 2156
rect 21868 2100 21924 2156
rect 0 2044 2940 2100
rect 2996 2044 3006 2100
rect 3388 2044 5628 2100
rect 5684 2044 5694 2100
rect 7634 2044 7644 2100
rect 7700 2044 10220 2100
rect 10276 2044 10286 2100
rect 12786 2044 12796 2100
rect 12852 2044 13468 2100
rect 13524 2044 13534 2100
rect 16034 2044 16044 2100
rect 16100 2044 17164 2100
rect 17220 2044 17230 2100
rect 21868 2044 23212 2100
rect 23268 2044 23278 2100
rect 23538 2044 23548 2100
rect 23604 2044 26796 2100
rect 26852 2044 26862 2100
rect 0 2016 112 2044
rect 2146 1932 2156 1988
rect 2212 1932 8540 1988
rect 8596 1932 8606 1988
rect 9884 1932 10444 1988
rect 10500 1932 10510 1988
rect 12338 1932 12348 1988
rect 12404 1932 13244 1988
rect 13300 1932 13310 1988
rect 14354 1932 14364 1988
rect 14420 1932 14476 1988
rect 14532 1932 14542 1988
rect 20850 1932 20860 1988
rect 20916 1932 27132 1988
rect 27188 1932 27198 1988
rect 9884 1876 9940 1932
rect 914 1820 924 1876
rect 980 1820 3668 1876
rect 3826 1820 3836 1876
rect 3892 1820 9940 1876
rect 10098 1820 10108 1876
rect 10164 1820 10220 1876
rect 10276 1820 17836 1876
rect 17892 1820 17902 1876
rect 19954 1820 19964 1876
rect 20020 1820 25116 1876
rect 25172 1820 25182 1876
rect 25890 1820 25900 1876
rect 25956 1820 26236 1876
rect 26292 1820 26302 1876
rect 3612 1764 3668 1820
rect 17836 1764 17892 1820
rect 1810 1708 1820 1764
rect 1876 1708 3388 1764
rect 3444 1708 3454 1764
rect 3612 1708 7084 1764
rect 7140 1708 7150 1764
rect 9538 1708 9548 1764
rect 9604 1708 15372 1764
rect 15428 1708 15438 1764
rect 17836 1708 19852 1764
rect 19908 1708 19918 1764
rect 20962 1708 20972 1764
rect 21028 1708 28140 1764
rect 28196 1708 28206 1764
rect 0 1652 112 1680
rect 0 1596 700 1652
rect 756 1596 766 1652
rect 6038 1596 6076 1652
rect 6132 1596 6142 1652
rect 6486 1596 6524 1652
rect 6580 1596 6590 1652
rect 6738 1596 6748 1652
rect 6804 1596 6842 1652
rect 6962 1596 6972 1652
rect 7028 1596 7066 1652
rect 7382 1596 7420 1652
rect 7476 1596 7486 1652
rect 7634 1596 7644 1652
rect 7700 1596 7738 1652
rect 7830 1596 7868 1652
rect 7924 1596 7934 1652
rect 8278 1596 8316 1652
rect 8372 1596 8382 1652
rect 8530 1596 8540 1652
rect 8596 1596 8634 1652
rect 8754 1596 8764 1652
rect 8820 1596 8858 1652
rect 9314 1596 9324 1652
rect 9380 1596 9660 1652
rect 9716 1596 9726 1652
rect 10070 1596 10108 1652
rect 10164 1596 10174 1652
rect 10294 1596 10332 1652
rect 10388 1596 10398 1652
rect 11190 1596 11228 1652
rect 11284 1596 11294 1652
rect 11414 1596 11452 1652
rect 11508 1596 11518 1652
rect 11862 1596 11900 1652
rect 11956 1596 11966 1652
rect 12086 1596 12124 1652
rect 12180 1596 12190 1652
rect 12338 1596 12348 1652
rect 12404 1596 12442 1652
rect 12534 1596 12572 1652
rect 12628 1596 12638 1652
rect 12786 1596 12796 1652
rect 12852 1596 12890 1652
rect 12982 1596 13020 1652
rect 13076 1596 13086 1652
rect 13234 1596 13244 1652
rect 13300 1596 13338 1652
rect 14690 1596 14700 1652
rect 14756 1596 22540 1652
rect 22596 1596 22606 1652
rect 24994 1596 25004 1652
rect 25060 1596 25116 1652
rect 25172 1596 25182 1652
rect 26002 1596 26012 1652
rect 26068 1596 28364 1652
rect 28420 1596 28430 1652
rect 0 1568 112 1596
rect 3794 1540 3804 1596
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 4068 1540 4078 1596
rect 23794 1540 23804 1596
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 24068 1540 24078 1596
rect 6290 1484 6300 1540
rect 6356 1484 7756 1540
rect 7812 1484 7822 1540
rect 9202 1484 9212 1540
rect 9268 1484 10556 1540
rect 10612 1484 10622 1540
rect 10882 1484 10892 1540
rect 10948 1484 11676 1540
rect 11732 1484 11742 1540
rect 21494 1484 21532 1540
rect 21588 1484 21598 1540
rect 24322 1484 24332 1540
rect 24388 1484 27020 1540
rect 27076 1484 27086 1540
rect 2258 1372 2268 1428
rect 2324 1372 5964 1428
rect 6020 1372 6030 1428
rect 8978 1372 8988 1428
rect 9044 1372 12012 1428
rect 12068 1372 12078 1428
rect 23650 1372 23660 1428
rect 23716 1372 23772 1428
rect 23828 1372 23838 1428
rect 26226 1372 26236 1428
rect 26292 1372 28588 1428
rect 28644 1372 28654 1428
rect 5618 1260 5628 1316
rect 5684 1260 11340 1316
rect 11396 1260 11406 1316
rect 11554 1260 11564 1316
rect 11620 1260 13916 1316
rect 13972 1260 13982 1316
rect 19282 1260 19292 1316
rect 19348 1260 19964 1316
rect 20020 1260 20030 1316
rect 23426 1260 23436 1316
rect 23492 1260 24892 1316
rect 24948 1260 24958 1316
rect 25106 1260 25116 1316
rect 25172 1260 27692 1316
rect 27748 1260 27758 1316
rect 0 1204 112 1232
rect 0 1148 2716 1204
rect 2772 1148 2782 1204
rect 4162 1148 4172 1204
rect 4228 1148 8652 1204
rect 8708 1148 8718 1204
rect 9548 1148 13132 1204
rect 13188 1148 13198 1204
rect 14802 1148 14812 1204
rect 14868 1148 15148 1204
rect 15204 1148 15214 1204
rect 17276 1148 21756 1204
rect 21812 1148 21822 1204
rect 23986 1148 23996 1204
rect 24052 1148 27244 1204
rect 27300 1148 27310 1204
rect 27990 1148 28028 1204
rect 28084 1148 28094 1204
rect 0 1120 112 1148
rect 9548 1092 9604 1148
rect 17276 1092 17332 1148
rect 4834 1036 4844 1092
rect 4900 1036 9604 1092
rect 10210 1036 10220 1092
rect 10276 1036 12684 1092
rect 12740 1036 17332 1092
rect 17490 1036 17500 1092
rect 17556 1036 26124 1092
rect 26180 1036 26190 1092
rect 26852 1036 28364 1092
rect 28420 1036 28430 1092
rect 26852 980 26908 1036
rect 5618 924 5628 980
rect 5684 924 9212 980
rect 9268 924 9278 980
rect 9426 924 9436 980
rect 9492 924 9884 980
rect 9940 924 9950 980
rect 10994 924 11004 980
rect 11060 924 11116 980
rect 11172 924 11182 980
rect 11330 924 11340 980
rect 11396 924 14812 980
rect 14868 924 14878 980
rect 15026 924 15036 980
rect 15092 924 16940 980
rect 16996 924 17006 980
rect 17266 924 17276 980
rect 17332 924 22988 980
rect 23044 924 23054 980
rect 23212 924 26908 980
rect 23212 868 23268 924
rect 5842 812 5852 868
rect 5908 812 15092 868
rect 15698 812 15708 868
rect 15764 812 16156 868
rect 16212 812 16222 868
rect 18386 812 18396 868
rect 18452 812 23268 868
rect 25554 812 25564 868
rect 25620 812 25788 868
rect 25844 812 25854 868
rect 0 756 112 784
rect 4454 756 4464 812
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4728 756 4738 812
rect 15036 756 15092 812
rect 24454 756 24464 812
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24728 756 24738 812
rect 0 700 924 756
rect 980 700 990 756
rect 5170 700 5180 756
rect 5236 700 14588 756
rect 14644 700 14654 756
rect 15026 700 15036 756
rect 15092 700 15102 756
rect 0 672 112 700
rect 10770 588 10780 644
rect 10836 588 11676 644
rect 11732 588 11742 644
rect 12226 588 12236 644
rect 12292 588 15708 644
rect 15764 588 15774 644
rect 17938 588 17948 644
rect 18004 588 22596 644
rect 24210 588 24220 644
rect 24276 588 24444 644
rect 24500 588 24510 644
rect 24658 588 24668 644
rect 24724 588 24892 644
rect 24948 588 24958 644
rect 22540 532 22596 588
rect 10546 476 10556 532
rect 10612 476 15596 532
rect 15652 476 15662 532
rect 17042 476 17052 532
rect 17108 476 22316 532
rect 22372 476 22382 532
rect 22540 476 25116 532
rect 25172 476 25182 532
rect 26852 476 27468 532
rect 27524 476 27534 532
rect 26852 420 26908 476
rect 5394 364 5404 420
rect 5460 364 9324 420
rect 9380 364 9390 420
rect 9538 364 9548 420
rect 9604 364 14812 420
rect 14868 364 14878 420
rect 19730 364 19740 420
rect 19796 364 26908 420
rect 0 308 112 336
rect 0 252 1596 308
rect 1652 252 1662 308
rect 7186 252 7196 308
rect 7252 252 11116 308
rect 11172 252 11182 308
rect 13122 252 13132 308
rect 13188 252 14028 308
rect 14084 252 14094 308
rect 19926 252 19964 308
rect 20020 252 20030 308
rect 20626 252 20636 308
rect 20692 252 29036 308
rect 29092 252 29102 308
rect 0 224 112 252
rect 17714 140 17724 196
rect 17780 140 26796 196
rect 26852 140 26862 196
rect 9314 28 9324 84
rect 9380 28 14252 84
rect 14308 28 14318 84
rect 19954 28 19964 84
rect 20020 28 26460 84
rect 26516 28 26526 84
<< via3 >>
rect 6636 114604 6692 114660
rect 4284 114492 4340 114548
rect 19964 113932 20020 113988
rect 5404 113820 5460 113876
rect 11900 113820 11956 113876
rect 4464 113652 4520 113708
rect 4568 113652 4624 113708
rect 4672 113652 4728 113708
rect 24464 113652 24520 113708
rect 24568 113652 24624 113708
rect 24672 113652 24728 113708
rect 27356 113596 27412 113652
rect 15036 113484 15092 113540
rect 19516 113484 19572 113540
rect 5292 113372 5348 113428
rect 8764 113372 8820 113428
rect 9884 113372 9940 113428
rect 13692 113372 13748 113428
rect 14140 113372 14196 113428
rect 14588 113372 14644 113428
rect 7308 113260 7364 113316
rect 7532 113260 7588 113316
rect 9324 113036 9380 113092
rect 10668 113036 10724 113092
rect 4956 112924 5012 112980
rect 11676 112924 11732 112980
rect 3804 112868 3860 112924
rect 3908 112868 3964 112924
rect 4012 112868 4068 112924
rect 23804 112868 23860 112924
rect 23908 112868 23964 112924
rect 24012 112868 24068 112924
rect 5180 112700 5236 112756
rect 7532 112700 7588 112756
rect 12684 112700 12740 112756
rect 5740 112588 5796 112644
rect 14364 112588 14420 112644
rect 14812 112588 14868 112644
rect 15148 112588 15204 112644
rect 16044 112588 16100 112644
rect 17052 112588 17108 112644
rect 6300 112476 6356 112532
rect 6860 112476 6916 112532
rect 10668 112476 10724 112532
rect 11228 112364 11284 112420
rect 11900 112364 11956 112420
rect 1820 112252 1876 112308
rect 5068 112252 5124 112308
rect 6412 112252 6468 112308
rect 7980 112252 8036 112308
rect 14700 112252 14756 112308
rect 16156 112252 16212 112308
rect 17388 112252 17444 112308
rect 6636 112140 6692 112196
rect 12684 112140 12740 112196
rect 4464 112084 4520 112140
rect 4568 112084 4624 112140
rect 4672 112084 4728 112140
rect 24464 112084 24520 112140
rect 24568 112084 24624 112140
rect 24672 112084 24728 112140
rect 15260 112028 15316 112084
rect 16156 112028 16212 112084
rect 25340 112028 25396 112084
rect 17948 111804 18004 111860
rect 21644 111804 21700 111860
rect 22204 111804 22260 111860
rect 3500 111692 3556 111748
rect 7084 111692 7140 111748
rect 10556 111692 10612 111748
rect 11228 111580 11284 111636
rect 11452 111580 11508 111636
rect 14476 111580 14532 111636
rect 16828 111468 16884 111524
rect 17724 111468 17780 111524
rect 3804 111300 3860 111356
rect 3908 111300 3964 111356
rect 4012 111300 4068 111356
rect 8988 111356 9044 111412
rect 13468 111356 13524 111412
rect 23804 111300 23860 111356
rect 23908 111300 23964 111356
rect 24012 111300 24068 111356
rect 7084 111132 7140 111188
rect 11452 111132 11508 111188
rect 17724 111132 17780 111188
rect 3500 111020 3556 111076
rect 5516 110908 5572 110964
rect 11116 110908 11172 110964
rect 12796 110908 12852 110964
rect 17836 110908 17892 110964
rect 18620 110908 18676 110964
rect 22316 110908 22372 110964
rect 23212 110908 23268 110964
rect 6748 110796 6804 110852
rect 27020 110796 27076 110852
rect 11676 110684 11732 110740
rect 26908 110684 26964 110740
rect 11340 110572 11396 110628
rect 14588 110572 14644 110628
rect 15820 110572 15876 110628
rect 25340 110572 25396 110628
rect 4464 110516 4520 110572
rect 4568 110516 4624 110572
rect 4672 110516 4728 110572
rect 24464 110516 24520 110572
rect 24568 110516 24624 110572
rect 24672 110516 24728 110572
rect 6188 110460 6244 110516
rect 13916 110460 13972 110516
rect 27132 110348 27188 110404
rect 27356 110348 27412 110404
rect 4956 110236 5012 110292
rect 5628 110236 5684 110292
rect 25228 110236 25284 110292
rect 10332 110124 10388 110180
rect 14252 110124 14308 110180
rect 14924 110124 14980 110180
rect 12908 110012 12964 110068
rect 14028 110012 14084 110068
rect 5628 109788 5684 109844
rect 3804 109732 3860 109788
rect 3908 109732 3964 109788
rect 4012 109732 4068 109788
rect 23804 109732 23860 109788
rect 23908 109732 23964 109788
rect 24012 109732 24068 109788
rect 4844 109676 4900 109732
rect 7980 109676 8036 109732
rect 3388 109564 3444 109620
rect 5404 109564 5460 109620
rect 14924 109564 14980 109620
rect 7980 109452 8036 109508
rect 13580 109452 13636 109508
rect 15820 109452 15876 109508
rect 18620 109452 18676 109508
rect 3612 109340 3668 109396
rect 8092 109340 8148 109396
rect 9996 109340 10052 109396
rect 1596 109228 1652 109284
rect 4172 109228 4228 109284
rect 4844 109228 4900 109284
rect 5852 109228 5908 109284
rect 9548 109116 9604 109172
rect 10220 109116 10276 109172
rect 19404 109116 19460 109172
rect 28028 109116 28084 109172
rect 3500 109004 3556 109060
rect 5068 109004 5124 109060
rect 10444 109004 10500 109060
rect 25340 109004 25396 109060
rect 27132 109004 27188 109060
rect 4464 108948 4520 109004
rect 4568 108948 4624 109004
rect 4672 108948 4728 109004
rect 24464 108948 24520 109004
rect 24568 108948 24624 109004
rect 24672 108948 24728 109004
rect 4284 108892 4340 108948
rect 13468 108892 13524 108948
rect 15260 108892 15316 108948
rect 3388 108668 3444 108724
rect 26908 108780 26964 108836
rect 8092 108668 8148 108724
rect 8540 108668 8596 108724
rect 8876 108556 8932 108612
rect 9548 108556 9604 108612
rect 19404 108556 19460 108612
rect 26236 108556 26292 108612
rect 4956 108444 5012 108500
rect 15260 108444 15316 108500
rect 23436 108444 23492 108500
rect 3276 108220 3332 108276
rect 11564 108332 11620 108388
rect 10444 108220 10500 108276
rect 3804 108164 3860 108220
rect 3908 108164 3964 108220
rect 4012 108164 4068 108220
rect 23804 108164 23860 108220
rect 23908 108164 23964 108220
rect 24012 108164 24068 108220
rect 6300 107884 6356 107940
rect 9884 107884 9940 107940
rect 14028 107884 14084 107940
rect 25228 107884 25284 107940
rect 1708 107772 1764 107828
rect 3276 107772 3332 107828
rect 5292 107772 5348 107828
rect 9324 107772 9380 107828
rect 10668 107772 10724 107828
rect 11340 107772 11396 107828
rect 13468 107772 13524 107828
rect 13916 107772 13972 107828
rect 14588 107772 14644 107828
rect 4284 107548 4340 107604
rect 8764 107548 8820 107604
rect 11340 107548 11396 107604
rect 14028 107548 14084 107604
rect 14812 107548 14868 107604
rect 15036 107548 15092 107604
rect 26796 107548 26852 107604
rect 14700 107436 14756 107492
rect 3612 107324 3668 107380
rect 4464 107380 4520 107436
rect 4568 107380 4624 107436
rect 4672 107380 4728 107436
rect 24464 107380 24520 107436
rect 24568 107380 24624 107436
rect 24672 107380 24728 107436
rect 5180 107324 5236 107380
rect 2380 106988 2436 107044
rect 3276 106988 3332 107044
rect 8316 106876 8372 106932
rect 8764 106876 8820 106932
rect 9548 106876 9604 106932
rect 10780 106876 10836 106932
rect 14588 106876 14644 106932
rect 21308 106876 21364 106932
rect 14476 106764 14532 106820
rect 20188 106652 20244 106708
rect 3804 106596 3860 106652
rect 3908 106596 3964 106652
rect 4012 106596 4068 106652
rect 23804 106596 23860 106652
rect 23908 106596 23964 106652
rect 24012 106596 24068 106652
rect 2156 106428 2212 106484
rect 2044 106204 2100 106260
rect 3052 106204 3108 106260
rect 1484 106092 1540 106148
rect 1932 105980 1988 106036
rect 3500 105868 3556 105924
rect 5964 105868 6020 105924
rect 4464 105812 4520 105868
rect 4568 105812 4624 105868
rect 4672 105812 4728 105868
rect 26124 106204 26180 106260
rect 7196 106092 7252 106148
rect 11228 105868 11284 105924
rect 13244 105868 13300 105924
rect 24464 105812 24520 105868
rect 24568 105812 24624 105868
rect 24672 105812 24728 105868
rect 2268 105644 2324 105700
rect 9212 105644 9268 105700
rect 2716 105532 2772 105588
rect 17948 105532 18004 105588
rect 19068 105532 19124 105588
rect 3612 105420 3668 105476
rect 6972 105420 7028 105476
rect 5068 105196 5124 105252
rect 13580 105196 13636 105252
rect 7980 105084 8036 105140
rect 3804 105028 3860 105084
rect 3908 105028 3964 105084
rect 4012 105028 4068 105084
rect 23804 105028 23860 105084
rect 23908 105028 23964 105084
rect 24012 105028 24068 105084
rect 16156 104524 16212 104580
rect 4844 104412 4900 104468
rect 8092 104412 8148 104468
rect 9324 104412 9380 104468
rect 9660 104412 9716 104468
rect 11452 104412 11508 104468
rect 11676 104412 11732 104468
rect 2268 104300 2324 104356
rect 4464 104244 4520 104300
rect 4568 104244 4624 104300
rect 4672 104244 4728 104300
rect 24464 104244 24520 104300
rect 24568 104244 24624 104300
rect 24672 104244 24728 104300
rect 2604 104188 2660 104244
rect 6076 104188 6132 104244
rect 6748 104188 6804 104244
rect 7420 104188 7476 104244
rect 17724 104188 17780 104244
rect 19068 104188 19124 104244
rect 6188 104076 6244 104132
rect 11900 104076 11956 104132
rect 13468 104076 13524 104132
rect 14700 104076 14756 104132
rect 1596 103964 1652 104020
rect 2716 103964 2772 104020
rect 5404 103964 5460 104020
rect 8092 103964 8148 104020
rect 11676 103964 11732 104020
rect 2604 103740 2660 103796
rect 5068 103740 5124 103796
rect 20300 103740 20356 103796
rect 5404 103628 5460 103684
rect 3804 103460 3860 103516
rect 3908 103460 3964 103516
rect 4012 103460 4068 103516
rect 10444 103516 10500 103572
rect 13580 103516 13636 103572
rect 23804 103460 23860 103516
rect 23908 103460 23964 103516
rect 24012 103460 24068 103516
rect 3500 103180 3556 103236
rect 2156 103068 2212 103124
rect 9324 103068 9380 103124
rect 5740 102956 5796 103012
rect 10444 102844 10500 102900
rect 16604 102844 16660 102900
rect 1484 102732 1540 102788
rect 8092 102732 8148 102788
rect 4464 102676 4520 102732
rect 4568 102676 4624 102732
rect 4672 102676 4728 102732
rect 24464 102676 24520 102732
rect 24568 102676 24624 102732
rect 24672 102676 24728 102732
rect 1372 102396 1428 102452
rect 5404 102172 5460 102228
rect 7644 102060 7700 102116
rect 3804 101892 3860 101948
rect 3908 101892 3964 101948
rect 4012 101892 4068 101948
rect 23804 101892 23860 101948
rect 23908 101892 23964 101948
rect 24012 101892 24068 101948
rect 5404 101500 5460 101556
rect 3612 101388 3668 101444
rect 13468 101388 13524 101444
rect 3612 101164 3668 101220
rect 17388 101164 17444 101220
rect 4464 101108 4520 101164
rect 4568 101108 4624 101164
rect 4672 101108 4728 101164
rect 24464 101108 24520 101164
rect 24568 101108 24624 101164
rect 24672 101108 24728 101164
rect 2380 100940 2436 100996
rect 3500 100716 3556 100772
rect 7308 100716 7364 100772
rect 2716 100604 2772 100660
rect 7196 100380 7252 100436
rect 16828 100380 16884 100436
rect 3804 100324 3860 100380
rect 3908 100324 3964 100380
rect 4012 100324 4068 100380
rect 5068 100268 5124 100324
rect 5404 100268 5460 100324
rect 23804 100324 23860 100380
rect 23908 100324 23964 100380
rect 24012 100324 24068 100380
rect 17836 100156 17892 100212
rect 5180 99932 5236 99988
rect 17724 99820 17780 99876
rect 10108 99708 10164 99764
rect 140 99596 196 99652
rect 4464 99540 4520 99596
rect 4568 99540 4624 99596
rect 4672 99540 4728 99596
rect 24464 99540 24520 99596
rect 24568 99540 24624 99596
rect 24672 99540 24728 99596
rect 7196 99484 7252 99540
rect 13916 99484 13972 99540
rect 2268 99260 2324 99316
rect 3612 99260 3668 99316
rect 3388 99148 3444 99204
rect 5292 99148 5348 99204
rect 2380 99036 2436 99092
rect 6188 99036 6244 99092
rect 3276 98924 3332 98980
rect 20076 98924 20132 98980
rect 3804 98756 3860 98812
rect 3908 98756 3964 98812
rect 4012 98756 4068 98812
rect 6076 98700 6132 98756
rect 10332 98812 10388 98868
rect 13020 98812 13076 98868
rect 18396 98812 18452 98868
rect 23804 98756 23860 98812
rect 23908 98756 23964 98812
rect 24012 98756 24068 98812
rect 252 98476 308 98532
rect 12572 98476 12628 98532
rect 14364 98476 14420 98532
rect 18172 98364 18228 98420
rect 5068 98252 5124 98308
rect 5740 98252 5796 98308
rect 6860 98252 6916 98308
rect 7980 98252 8036 98308
rect 16156 98252 16212 98308
rect 14364 98028 14420 98084
rect 14812 98028 14868 98084
rect 4464 97972 4520 98028
rect 4568 97972 4624 98028
rect 4672 97972 4728 98028
rect 24464 97972 24520 98028
rect 24568 97972 24624 98028
rect 24672 97972 24728 98028
rect 13692 97916 13748 97972
rect 17836 97916 17892 97972
rect 20076 97804 20132 97860
rect 4956 97692 5012 97748
rect 14364 97692 14420 97748
rect 7756 97580 7812 97636
rect 11116 97580 11172 97636
rect 16940 97580 16996 97636
rect 7756 97356 7812 97412
rect 3804 97188 3860 97244
rect 3908 97188 3964 97244
rect 4012 97188 4068 97244
rect 23804 97188 23860 97244
rect 23908 97188 23964 97244
rect 24012 97188 24068 97244
rect 14364 97132 14420 97188
rect 3276 97020 3332 97076
rect 5404 96908 5460 96964
rect 14140 96908 14196 96964
rect 9884 96796 9940 96852
rect 3612 96684 3668 96740
rect 6188 96684 6244 96740
rect 14140 96684 14196 96740
rect 17836 96684 17892 96740
rect 15708 96572 15764 96628
rect 4464 96404 4520 96460
rect 4568 96404 4624 96460
rect 4672 96404 4728 96460
rect 24464 96404 24520 96460
rect 24568 96404 24624 96460
rect 24672 96404 24728 96460
rect 2604 96236 2660 96292
rect 1708 96124 1764 96180
rect 17836 96124 17892 96180
rect 3500 96012 3556 96068
rect 7532 96012 7588 96068
rect 18172 96012 18228 96068
rect 1372 95900 1428 95956
rect 5068 95900 5124 95956
rect 14364 95900 14420 95956
rect 476 95788 532 95844
rect 2380 95788 2436 95844
rect 3612 95788 3668 95844
rect 11788 95788 11844 95844
rect 8652 95676 8708 95732
rect 14028 95676 14084 95732
rect 3804 95620 3860 95676
rect 3908 95620 3964 95676
rect 4012 95620 4068 95676
rect 23804 95620 23860 95676
rect 23908 95620 23964 95676
rect 24012 95620 24068 95676
rect 5180 95452 5236 95508
rect 3612 95340 3668 95396
rect 10444 95340 10500 95396
rect 4284 95228 4340 95284
rect 3500 95116 3556 95172
rect 6972 95116 7028 95172
rect 14812 95116 14868 95172
rect 4464 94836 4520 94892
rect 4568 94836 4624 94892
rect 4672 94836 4728 94892
rect 24464 94836 24520 94892
rect 24568 94836 24624 94892
rect 24672 94836 24728 94892
rect 3500 94780 3556 94836
rect 4284 94780 4340 94836
rect 8652 94668 8708 94724
rect 8988 94668 9044 94724
rect 6972 94556 7028 94612
rect 11900 94556 11956 94612
rect 2492 94444 2548 94500
rect 5404 94444 5460 94500
rect 5516 94332 5572 94388
rect 8428 94332 8484 94388
rect 13916 94332 13972 94388
rect 17164 94220 17220 94276
rect 2492 94108 2548 94164
rect 13580 94108 13636 94164
rect 3804 94052 3860 94108
rect 3908 94052 3964 94108
rect 4012 94052 4068 94108
rect 23804 94052 23860 94108
rect 23908 94052 23964 94108
rect 24012 94052 24068 94108
rect 3500 93996 3556 94052
rect 10892 93996 10948 94052
rect 3164 93772 3220 93828
rect 4284 93772 4340 93828
rect 17836 93660 17892 93716
rect 476 93436 532 93492
rect 17948 93436 18004 93492
rect 5068 93324 5124 93380
rect 4464 93268 4520 93324
rect 4568 93268 4624 93324
rect 4672 93268 4728 93324
rect 24464 93268 24520 93324
rect 24568 93268 24624 93324
rect 24672 93268 24728 93324
rect 7084 93212 7140 93268
rect 15596 92988 15652 93044
rect 11004 92876 11060 92932
rect 6300 92540 6356 92596
rect 15596 92540 15652 92596
rect 3804 92484 3860 92540
rect 3908 92484 3964 92540
rect 4012 92484 4068 92540
rect 23804 92484 23860 92540
rect 23908 92484 23964 92540
rect 24012 92484 24068 92540
rect 17836 92316 17892 92372
rect 20076 92316 20132 92372
rect 5068 92092 5124 92148
rect 17276 92092 17332 92148
rect 1484 91980 1540 92036
rect 6524 91868 6580 91924
rect 4464 91700 4520 91756
rect 4568 91700 4624 91756
rect 4672 91700 4728 91756
rect 7420 91532 7476 91588
rect 24464 91700 24520 91756
rect 24568 91700 24624 91756
rect 24672 91700 24728 91756
rect 21980 91644 22036 91700
rect 7084 91420 7140 91476
rect 7980 91420 8036 91476
rect 6524 91084 6580 91140
rect 3804 90916 3860 90972
rect 3908 90916 3964 90972
rect 4012 90916 4068 90972
rect 23804 90916 23860 90972
rect 23908 90916 23964 90972
rect 24012 90916 24068 90972
rect 5964 90748 6020 90804
rect 3612 90524 3668 90580
rect 2380 90300 2436 90356
rect 11228 90300 11284 90356
rect 11676 90188 11732 90244
rect 4464 90132 4520 90188
rect 4568 90132 4624 90188
rect 4672 90132 4728 90188
rect 24464 90132 24520 90188
rect 24568 90132 24624 90188
rect 24672 90132 24728 90188
rect 9884 90076 9940 90132
rect 17836 89964 17892 90020
rect 252 89852 308 89908
rect 7644 89852 7700 89908
rect 7868 89852 7924 89908
rect 3388 89740 3444 89796
rect 2604 89516 2660 89572
rect 7868 89516 7924 89572
rect 3804 89348 3860 89404
rect 3908 89348 3964 89404
rect 4012 89348 4068 89404
rect 23804 89348 23860 89404
rect 23908 89348 23964 89404
rect 24012 89348 24068 89404
rect 8204 89292 8260 89348
rect 5068 89068 5124 89124
rect 1708 88956 1764 89012
rect 6972 88956 7028 89012
rect 8764 88956 8820 89012
rect 4844 88844 4900 88900
rect 5852 88732 5908 88788
rect 4464 88564 4520 88620
rect 4568 88564 4624 88620
rect 4672 88564 4728 88620
rect 24464 88564 24520 88620
rect 24568 88564 24624 88620
rect 24672 88564 24728 88620
rect 5740 88508 5796 88564
rect 6636 88508 6692 88564
rect 9884 88284 9940 88340
rect 11228 88284 11284 88340
rect 3500 88172 3556 88228
rect 3276 88060 3332 88116
rect 3804 87780 3860 87836
rect 3908 87780 3964 87836
rect 4012 87780 4068 87836
rect 23804 87780 23860 87836
rect 23908 87780 23964 87836
rect 24012 87780 24068 87836
rect 10556 87724 10612 87780
rect 3388 87612 3444 87668
rect 1708 87500 1764 87556
rect 22652 87500 22708 87556
rect 1372 87388 1428 87444
rect 8428 87388 8484 87444
rect 11788 87388 11844 87444
rect 140 87276 196 87332
rect 14364 87276 14420 87332
rect 18844 87164 18900 87220
rect 4464 86996 4520 87052
rect 4568 86996 4624 87052
rect 4672 86996 4728 87052
rect 24464 86996 24520 87052
rect 24568 86996 24624 87052
rect 24672 86996 24728 87052
rect 6300 86940 6356 86996
rect 2044 86828 2100 86884
rect 11004 86716 11060 86772
rect 18732 86716 18788 86772
rect 23100 86716 23156 86772
rect 13468 86604 13524 86660
rect 13468 86268 13524 86324
rect 3804 86212 3860 86268
rect 3908 86212 3964 86268
rect 4012 86212 4068 86268
rect 23804 86212 23860 86268
rect 23908 86212 23964 86268
rect 24012 86212 24068 86268
rect 2380 86156 2436 86212
rect 1596 86044 1652 86100
rect 23548 86044 23604 86100
rect 1820 85820 1876 85876
rect 5628 85820 5684 85876
rect 14812 85820 14868 85876
rect 1484 85708 1540 85764
rect 3388 85708 3444 85764
rect 14140 85708 14196 85764
rect 17052 85596 17108 85652
rect 21980 85596 22036 85652
rect 14140 85484 14196 85540
rect 23548 85484 23604 85540
rect 1484 85372 1540 85428
rect 4464 85428 4520 85484
rect 4568 85428 4624 85484
rect 4672 85428 4728 85484
rect 24464 85428 24520 85484
rect 24568 85428 24624 85484
rect 24672 85428 24728 85484
rect 17276 85372 17332 85428
rect 13356 85260 13412 85316
rect 23100 85260 23156 85316
rect 2940 85148 2996 85204
rect 15148 85036 15204 85092
rect 16828 85036 16884 85092
rect 8204 84924 8260 84980
rect 11228 84924 11284 84980
rect 13356 84924 13412 84980
rect 14364 84812 14420 84868
rect 6188 84700 6244 84756
rect 3804 84644 3860 84700
rect 3908 84644 3964 84700
rect 4012 84644 4068 84700
rect 23804 84644 23860 84700
rect 23908 84644 23964 84700
rect 24012 84644 24068 84700
rect 4956 84588 5012 84644
rect 9884 84588 9940 84644
rect 10892 84588 10948 84644
rect 3164 84476 3220 84532
rect 11004 84364 11060 84420
rect 6188 84252 6244 84308
rect 13692 84140 13748 84196
rect 2044 84028 2100 84084
rect 3052 84028 3108 84084
rect 8204 83916 8260 83972
rect 4464 83860 4520 83916
rect 4568 83860 4624 83916
rect 4672 83860 4728 83916
rect 24464 83860 24520 83916
rect 24568 83860 24624 83916
rect 24672 83860 24728 83916
rect 5404 83692 5460 83748
rect 5628 83692 5684 83748
rect 2716 83580 2772 83636
rect 8988 83580 9044 83636
rect 700 83468 756 83524
rect 14364 83356 14420 83412
rect 18844 83244 18900 83300
rect 5404 83132 5460 83188
rect 11676 83132 11732 83188
rect 3804 83076 3860 83132
rect 3908 83076 3964 83132
rect 4012 83076 4068 83132
rect 23804 83076 23860 83132
rect 23908 83076 23964 83132
rect 24012 83076 24068 83132
rect 1820 82684 1876 82740
rect 16716 82572 16772 82628
rect 8092 82460 8148 82516
rect 17388 82348 17444 82404
rect 4464 82292 4520 82348
rect 4568 82292 4624 82348
rect 4672 82292 4728 82348
rect 24464 82292 24520 82348
rect 24568 82292 24624 82348
rect 24672 82292 24728 82348
rect 2380 82236 2436 82292
rect 6748 82124 6804 82180
rect 8428 82012 8484 82068
rect 2156 81788 2212 81844
rect 2492 81788 2548 81844
rect 3804 81508 3860 81564
rect 3908 81508 3964 81564
rect 4012 81508 4068 81564
rect 9100 81452 9156 81508
rect 14364 81452 14420 81508
rect 23804 81508 23860 81564
rect 23908 81508 23964 81564
rect 24012 81508 24068 81564
rect 13132 81340 13188 81396
rect 15148 81228 15204 81284
rect 9884 81116 9940 81172
rect 14812 81116 14868 81172
rect 7756 81004 7812 81060
rect 4844 80892 4900 80948
rect 15036 81004 15092 81060
rect 22428 80892 22484 80948
rect 8204 80780 8260 80836
rect 4464 80724 4520 80780
rect 4568 80724 4624 80780
rect 4672 80724 4728 80780
rect 24464 80724 24520 80780
rect 24568 80724 24624 80780
rect 24672 80724 24728 80780
rect 15036 80668 15092 80724
rect 3612 80444 3668 80500
rect 2828 80332 2884 80388
rect 3276 80332 3332 80388
rect 6748 80220 6804 80276
rect 1708 80108 1764 80164
rect 10332 79996 10388 80052
rect 26572 79996 26628 80052
rect 3804 79940 3860 79996
rect 3908 79940 3964 79996
rect 4012 79940 4068 79996
rect 23804 79940 23860 79996
rect 23908 79940 23964 79996
rect 24012 79940 24068 79996
rect 9100 79884 9156 79940
rect 10556 79884 10612 79940
rect 1708 79548 1764 79604
rect 7532 79548 7588 79604
rect 10332 79548 10388 79604
rect 22428 79548 22484 79604
rect 6860 79436 6916 79492
rect 3388 79324 3444 79380
rect 9100 79324 9156 79380
rect 10556 79324 10612 79380
rect 11228 79324 11284 79380
rect 17948 79324 18004 79380
rect 4464 79156 4520 79212
rect 4568 79156 4624 79212
rect 4672 79156 4728 79212
rect 24464 79156 24520 79212
rect 24568 79156 24624 79212
rect 24672 79156 24728 79212
rect 6860 79100 6916 79156
rect 1708 78988 1764 79044
rect 2716 78988 2772 79044
rect 11676 78988 11732 79044
rect 17612 78876 17668 78932
rect 3804 78372 3860 78428
rect 3908 78372 3964 78428
rect 4012 78372 4068 78428
rect 23804 78372 23860 78428
rect 23908 78372 23964 78428
rect 24012 78372 24068 78428
rect 1820 78316 1876 78372
rect 5628 77868 5684 77924
rect 3164 77756 3220 77812
rect 15148 77980 15204 78036
rect 10332 77868 10388 77924
rect 10892 77756 10948 77812
rect 22988 77644 23044 77700
rect 4464 77588 4520 77644
rect 4568 77588 4624 77644
rect 4672 77588 4728 77644
rect 24464 77588 24520 77644
rect 24568 77588 24624 77644
rect 24672 77588 24728 77644
rect 6636 77420 6692 77476
rect 1596 77308 1652 77364
rect 8092 77196 8148 77252
rect 11452 77196 11508 77252
rect 12124 77196 12180 77252
rect 4284 77084 4340 77140
rect 9212 76972 9268 77028
rect 10668 76972 10724 77028
rect 3804 76804 3860 76860
rect 3908 76804 3964 76860
rect 4012 76804 4068 76860
rect 23804 76804 23860 76860
rect 23908 76804 23964 76860
rect 24012 76804 24068 76860
rect 3612 76748 3668 76804
rect 1708 76524 1764 76580
rect 12684 76524 12740 76580
rect 3388 76412 3444 76468
rect 3612 76412 3668 76468
rect 26572 76412 26628 76468
rect 2716 76300 2772 76356
rect 1260 76188 1316 76244
rect 6300 76076 6356 76132
rect 4464 76020 4520 76076
rect 4568 76020 4624 76076
rect 4672 76020 4728 76076
rect 24464 76020 24520 76076
rect 24568 76020 24624 76076
rect 24672 76020 24728 76076
rect 7084 75852 7140 75908
rect 7980 75852 8036 75908
rect 3804 75236 3860 75292
rect 3908 75236 3964 75292
rect 4012 75236 4068 75292
rect 23804 75236 23860 75292
rect 23908 75236 23964 75292
rect 24012 75236 24068 75292
rect 8428 75180 8484 75236
rect 4284 74844 4340 74900
rect 700 74732 756 74788
rect 4956 74732 5012 74788
rect 14364 74732 14420 74788
rect 17612 74732 17668 74788
rect 924 74508 980 74564
rect 4464 74452 4520 74508
rect 4568 74452 4624 74508
rect 4672 74452 4728 74508
rect 24464 74452 24520 74508
rect 24568 74452 24624 74508
rect 24672 74452 24728 74508
rect 3164 74396 3220 74452
rect 12908 74396 12964 74452
rect 3500 74172 3556 74228
rect 1372 74060 1428 74116
rect 17612 73948 17668 74004
rect 7532 73724 7588 73780
rect 3804 73668 3860 73724
rect 3908 73668 3964 73724
rect 4012 73668 4068 73724
rect 23804 73668 23860 73724
rect 23908 73668 23964 73724
rect 24012 73668 24068 73724
rect 2716 73500 2772 73556
rect 12684 73388 12740 73444
rect 2828 73276 2884 73332
rect 11676 73164 11732 73220
rect 20076 73164 20132 73220
rect 5628 72940 5684 72996
rect 4464 72884 4520 72940
rect 4568 72884 4624 72940
rect 4672 72884 4728 72940
rect 24464 72884 24520 72940
rect 24568 72884 24624 72940
rect 24672 72884 24728 72940
rect 1820 72828 1876 72884
rect 17388 72716 17444 72772
rect 6300 72604 6356 72660
rect 1596 72492 1652 72548
rect 11228 72492 11284 72548
rect 16044 72380 16100 72436
rect 3804 72100 3860 72156
rect 3908 72100 3964 72156
rect 4012 72100 4068 72156
rect 23804 72100 23860 72156
rect 23908 72100 23964 72156
rect 24012 72100 24068 72156
rect 924 72044 980 72100
rect 4844 71932 4900 71988
rect 6076 71820 6132 71876
rect 10892 71596 10948 71652
rect 4464 71316 4520 71372
rect 4568 71316 4624 71372
rect 4672 71316 4728 71372
rect 24464 71316 24520 71372
rect 24568 71316 24624 71372
rect 24672 71316 24728 71372
rect 3500 70924 3556 70980
rect 8876 70588 8932 70644
rect 3804 70532 3860 70588
rect 3908 70532 3964 70588
rect 4012 70532 4068 70588
rect 23804 70532 23860 70588
rect 23908 70532 23964 70588
rect 24012 70532 24068 70588
rect 1820 70364 1876 70420
rect 2940 70028 2996 70084
rect 4464 69748 4520 69804
rect 4568 69748 4624 69804
rect 4672 69748 4728 69804
rect 24464 69748 24520 69804
rect 24568 69748 24624 69804
rect 24672 69748 24728 69804
rect 3276 69356 3332 69412
rect 3804 68964 3860 69020
rect 3908 68964 3964 69020
rect 4012 68964 4068 69020
rect 23804 68964 23860 69020
rect 23908 68964 23964 69020
rect 24012 68964 24068 69020
rect 7084 68908 7140 68964
rect 7756 68796 7812 68852
rect 1372 68684 1428 68740
rect 1036 68572 1092 68628
rect 7756 68460 7812 68516
rect 9324 68460 9380 68516
rect 11228 68460 11284 68516
rect 8204 68348 8260 68404
rect 1036 67788 1092 67844
rect 4464 68180 4520 68236
rect 4568 68180 4624 68236
rect 4672 68180 4728 68236
rect 24464 68180 24520 68236
rect 24568 68180 24624 68236
rect 24672 68180 24728 68236
rect 4956 67900 5012 67956
rect 3500 67676 3556 67732
rect 20748 67564 20804 67620
rect 9436 67452 9492 67508
rect 10220 67452 10276 67508
rect 3804 67396 3860 67452
rect 3908 67396 3964 67452
rect 4012 67396 4068 67452
rect 23804 67396 23860 67452
rect 23908 67396 23964 67452
rect 24012 67396 24068 67452
rect 4172 67340 4228 67396
rect 3388 67228 3444 67284
rect 6636 67004 6692 67060
rect 4464 66612 4520 66668
rect 4568 66612 4624 66668
rect 4672 66612 4728 66668
rect 24464 66612 24520 66668
rect 24568 66612 24624 66668
rect 24672 66612 24728 66668
rect 20748 66444 20804 66500
rect 5180 66220 5236 66276
rect 3388 66108 3444 66164
rect 9100 65996 9156 66052
rect 3804 65828 3860 65884
rect 3908 65828 3964 65884
rect 4012 65828 4068 65884
rect 23804 65828 23860 65884
rect 23908 65828 23964 65884
rect 24012 65828 24068 65884
rect 1260 65660 1316 65716
rect 16268 65660 16324 65716
rect 8204 65436 8260 65492
rect 3500 65324 3556 65380
rect 4464 65044 4520 65100
rect 4568 65044 4624 65100
rect 4672 65044 4728 65100
rect 24464 65044 24520 65100
rect 24568 65044 24624 65100
rect 24672 65044 24728 65100
rect 3612 64764 3668 64820
rect 3804 64260 3860 64316
rect 3908 64260 3964 64316
rect 4012 64260 4068 64316
rect 23804 64260 23860 64316
rect 23908 64260 23964 64316
rect 24012 64260 24068 64316
rect 12572 63980 12628 64036
rect 2492 63756 2548 63812
rect 7980 63756 8036 63812
rect 4464 63476 4520 63532
rect 4568 63476 4624 63532
rect 4672 63476 4728 63532
rect 24464 63476 24520 63532
rect 24568 63476 24624 63532
rect 24672 63476 24728 63532
rect 5180 63196 5236 63252
rect 7980 63084 8036 63140
rect 12572 62860 12628 62916
rect 12908 62860 12964 62916
rect 3804 62692 3860 62748
rect 3908 62692 3964 62748
rect 4012 62692 4068 62748
rect 23804 62692 23860 62748
rect 23908 62692 23964 62748
rect 24012 62692 24068 62748
rect 9884 62636 9940 62692
rect 2492 62524 2548 62580
rect 3276 62412 3332 62468
rect 21196 62412 21252 62468
rect 21756 62188 21812 62244
rect 21196 62076 21252 62132
rect 4464 61908 4520 61964
rect 4568 61908 4624 61964
rect 4672 61908 4728 61964
rect 24464 61908 24520 61964
rect 24568 61908 24624 61964
rect 24672 61908 24728 61964
rect 2044 61740 2100 61796
rect 21532 61180 21588 61236
rect 3804 61124 3860 61180
rect 3908 61124 3964 61180
rect 4012 61124 4068 61180
rect 23804 61124 23860 61180
rect 23908 61124 23964 61180
rect 24012 61124 24068 61180
rect 16268 60844 16324 60900
rect 7756 60620 7812 60676
rect 4464 60340 4520 60396
rect 4568 60340 4624 60396
rect 4672 60340 4728 60396
rect 24464 60340 24520 60396
rect 24568 60340 24624 60396
rect 24672 60340 24728 60396
rect 3804 59556 3860 59612
rect 3908 59556 3964 59612
rect 4012 59556 4068 59612
rect 23804 59556 23860 59612
rect 23908 59556 23964 59612
rect 24012 59556 24068 59612
rect 4464 58772 4520 58828
rect 4568 58772 4624 58828
rect 4672 58772 4728 58828
rect 24464 58772 24520 58828
rect 24568 58772 24624 58828
rect 24672 58772 24728 58828
rect 2268 58716 2324 58772
rect 1372 58156 1428 58212
rect 1932 58156 1988 58212
rect 3804 57988 3860 58044
rect 3908 57988 3964 58044
rect 4012 57988 4068 58044
rect 23804 57988 23860 58044
rect 23908 57988 23964 58044
rect 24012 57988 24068 58044
rect 3164 57708 3220 57764
rect 6076 57260 6132 57316
rect 4464 57204 4520 57260
rect 4568 57204 4624 57260
rect 4672 57204 4728 57260
rect 24464 57204 24520 57260
rect 24568 57204 24624 57260
rect 24672 57204 24728 57260
rect 10108 56924 10164 56980
rect 20188 56924 20244 56980
rect 7420 56588 7476 56644
rect 3804 56420 3860 56476
rect 3908 56420 3964 56476
rect 4012 56420 4068 56476
rect 23804 56420 23860 56476
rect 23908 56420 23964 56476
rect 24012 56420 24068 56476
rect 14476 56140 14532 56196
rect 4464 55636 4520 55692
rect 4568 55636 4624 55692
rect 4672 55636 4728 55692
rect 24464 55636 24520 55692
rect 24568 55636 24624 55692
rect 24672 55636 24728 55692
rect 19292 55468 19348 55524
rect 20300 55468 20356 55524
rect 5292 55356 5348 55412
rect 9548 55356 9604 55412
rect 12348 55356 12404 55412
rect 13132 55356 13188 55412
rect 14476 55356 14532 55412
rect 8316 55244 8372 55300
rect 11900 55244 11956 55300
rect 2604 55020 2660 55076
rect 3804 54852 3860 54908
rect 3908 54852 3964 54908
rect 4012 54852 4068 54908
rect 23804 54852 23860 54908
rect 23908 54852 23964 54908
rect 24012 54852 24068 54908
rect 20412 54572 20468 54628
rect 14924 54460 14980 54516
rect 9548 54348 9604 54404
rect 15596 54348 15652 54404
rect 4464 54068 4520 54124
rect 4568 54068 4624 54124
rect 4672 54068 4728 54124
rect 24464 54068 24520 54124
rect 24568 54068 24624 54124
rect 24672 54068 24728 54124
rect 6972 53676 7028 53732
rect 3276 53564 3332 53620
rect 3804 53284 3860 53340
rect 3908 53284 3964 53340
rect 4012 53284 4068 53340
rect 23804 53284 23860 53340
rect 23908 53284 23964 53340
rect 24012 53284 24068 53340
rect 7868 53004 7924 53060
rect 6524 52892 6580 52948
rect 8316 52892 8372 52948
rect 9212 52892 9268 52948
rect 15148 52668 15204 52724
rect 4464 52500 4520 52556
rect 4568 52500 4624 52556
rect 4672 52500 4728 52556
rect 24464 52500 24520 52556
rect 24568 52500 24624 52556
rect 24672 52500 24728 52556
rect 8316 52108 8372 52164
rect 4844 51996 4900 52052
rect 1708 51324 1764 51380
rect 2940 51324 2996 51380
rect 3804 51716 3860 51772
rect 3908 51716 3964 51772
rect 4012 51716 4068 51772
rect 23804 51716 23860 51772
rect 23908 51716 23964 51772
rect 24012 51716 24068 51772
rect 3388 51548 3444 51604
rect 4464 50932 4520 50988
rect 4568 50932 4624 50988
rect 4672 50932 4728 50988
rect 2492 50652 2548 50708
rect 12236 50652 12292 50708
rect 24464 50932 24520 50988
rect 24568 50932 24624 50988
rect 24672 50932 24728 50988
rect 15260 50876 15316 50932
rect 6860 50540 6916 50596
rect 8204 50540 8260 50596
rect 3804 50148 3860 50204
rect 3908 50148 3964 50204
rect 4012 50148 4068 50204
rect 23804 50148 23860 50204
rect 23908 50148 23964 50204
rect 24012 50148 24068 50204
rect 10668 49980 10724 50036
rect 11004 49980 11060 50036
rect 11004 49756 11060 49812
rect 15820 49756 15876 49812
rect 17164 49644 17220 49700
rect 7420 49532 7476 49588
rect 4464 49364 4520 49420
rect 4568 49364 4624 49420
rect 4672 49364 4728 49420
rect 24464 49364 24520 49420
rect 24568 49364 24624 49420
rect 24672 49364 24728 49420
rect 4844 49308 4900 49364
rect 3500 49084 3556 49140
rect 4844 49084 4900 49140
rect 2492 48636 2548 48692
rect 3804 48580 3860 48636
rect 3908 48580 3964 48636
rect 4012 48580 4068 48636
rect 23804 48580 23860 48636
rect 23908 48580 23964 48636
rect 24012 48580 24068 48636
rect 14924 47964 14980 48020
rect 4464 47796 4520 47852
rect 4568 47796 4624 47852
rect 4672 47796 4728 47852
rect 24464 47796 24520 47852
rect 24568 47796 24624 47852
rect 24672 47796 24728 47852
rect 1932 47516 1988 47572
rect 19292 47516 19348 47572
rect 18732 47404 18788 47460
rect 7084 47292 7140 47348
rect 16604 47292 16660 47348
rect 7868 47180 7924 47236
rect 2492 47068 2548 47124
rect 3052 47068 3108 47124
rect 3804 47012 3860 47068
rect 3908 47012 3964 47068
rect 4012 47012 4068 47068
rect 23804 47012 23860 47068
rect 23908 47012 23964 47068
rect 24012 47012 24068 47068
rect 23548 46956 23604 47012
rect 7084 46732 7140 46788
rect 10108 46508 10164 46564
rect 12012 46508 12068 46564
rect 16716 46508 16772 46564
rect 11788 46396 11844 46452
rect 4464 46228 4520 46284
rect 4568 46228 4624 46284
rect 4672 46228 4728 46284
rect 24464 46228 24520 46284
rect 24568 46228 24624 46284
rect 24672 46228 24728 46284
rect 5404 46060 5460 46116
rect 5964 45948 6020 46004
rect 7084 45948 7140 46004
rect 10556 45948 10612 46004
rect 11004 45948 11060 46004
rect 4956 45836 5012 45892
rect 8988 45724 9044 45780
rect 9884 45612 9940 45668
rect 10108 45612 10164 45668
rect 3804 45444 3860 45500
rect 3908 45444 3964 45500
rect 4012 45444 4068 45500
rect 23804 45444 23860 45500
rect 23908 45444 23964 45500
rect 24012 45444 24068 45500
rect 9884 45388 9940 45444
rect 12012 45388 12068 45444
rect 9324 45276 9380 45332
rect 2044 45052 2100 45108
rect 6860 45052 6916 45108
rect 8204 45052 8260 45108
rect 10220 45052 10276 45108
rect 11676 45052 11732 45108
rect 5180 44940 5236 44996
rect 2492 44716 2548 44772
rect 4464 44660 4520 44716
rect 4568 44660 4624 44716
rect 4672 44660 4728 44716
rect 8092 44492 8148 44548
rect 24464 44660 24520 44716
rect 24568 44660 24624 44716
rect 24672 44660 24728 44716
rect 11340 44492 11396 44548
rect 11452 44380 11508 44436
rect 9884 44268 9940 44324
rect 19404 44156 19460 44212
rect 6748 44044 6804 44100
rect 8092 44044 8148 44100
rect 16828 43932 16884 43988
rect 3804 43876 3860 43932
rect 3908 43876 3964 43932
rect 4012 43876 4068 43932
rect 23804 43876 23860 43932
rect 23908 43876 23964 43932
rect 24012 43876 24068 43932
rect 4284 43708 4340 43764
rect 9660 43596 9716 43652
rect 10892 43596 10948 43652
rect 17388 43596 17444 43652
rect 18844 43484 18900 43540
rect 1820 43372 1876 43428
rect 6188 43260 6244 43316
rect 14364 43260 14420 43316
rect 4464 43092 4520 43148
rect 4568 43092 4624 43148
rect 4672 43092 4728 43148
rect 24464 43092 24520 43148
rect 24568 43092 24624 43148
rect 24672 43092 24728 43148
rect 2044 42924 2100 42980
rect 5628 42924 5684 42980
rect 14252 42924 14308 42980
rect 1148 42588 1204 42644
rect 4284 42588 4340 42644
rect 5852 42588 5908 42644
rect 3804 42308 3860 42364
rect 3908 42308 3964 42364
rect 4012 42308 4068 42364
rect 23804 42308 23860 42364
rect 23908 42308 23964 42364
rect 24012 42308 24068 42364
rect 1820 41916 1876 41972
rect 6412 41916 6468 41972
rect 11004 41916 11060 41972
rect 18284 41916 18340 41972
rect 1484 41804 1540 41860
rect 9996 41804 10052 41860
rect 12572 41804 12628 41860
rect 17164 41804 17220 41860
rect 4464 41524 4520 41580
rect 4568 41524 4624 41580
rect 4672 41524 4728 41580
rect 24464 41524 24520 41580
rect 24568 41524 24624 41580
rect 24672 41524 24728 41580
rect 2604 41468 2660 41524
rect 3276 41468 3332 41524
rect 11564 41356 11620 41412
rect 21420 41356 21476 41412
rect 2492 40908 2548 40964
rect 11116 40908 11172 40964
rect 1148 40572 1204 40628
rect 3804 40740 3860 40796
rect 3908 40740 3964 40796
rect 4012 40740 4068 40796
rect 23804 40740 23860 40796
rect 23908 40740 23964 40796
rect 24012 40740 24068 40796
rect 8876 40460 8932 40516
rect 18396 40460 18452 40516
rect 6188 40348 6244 40404
rect 11564 40348 11620 40404
rect 18172 40348 18228 40404
rect 19852 40348 19908 40404
rect 2044 40236 2100 40292
rect 6076 40236 6132 40292
rect 6636 40236 6692 40292
rect 18060 40124 18116 40180
rect 4956 40012 5012 40068
rect 5740 40012 5796 40068
rect 4464 39956 4520 40012
rect 4568 39956 4624 40012
rect 4672 39956 4728 40012
rect 24464 39956 24520 40012
rect 24568 39956 24624 40012
rect 24672 39956 24728 40012
rect 14252 39676 14308 39732
rect 11564 39452 11620 39508
rect 18060 39452 18116 39508
rect 4844 39340 4900 39396
rect 20524 39340 20580 39396
rect 14924 39228 14980 39284
rect 3804 39172 3860 39228
rect 3908 39172 3964 39228
rect 4012 39172 4068 39228
rect 23804 39172 23860 39228
rect 23908 39172 23964 39228
rect 24012 39172 24068 39228
rect 5068 39004 5124 39060
rect 11564 39004 11620 39060
rect 11564 38780 11620 38836
rect 14252 38780 14308 38836
rect 6636 38668 6692 38724
rect 14700 38668 14756 38724
rect 6188 38444 6244 38500
rect 10556 38444 10612 38500
rect 4464 38388 4520 38444
rect 4568 38388 4624 38444
rect 4672 38388 4728 38444
rect 24464 38388 24520 38444
rect 24568 38388 24624 38444
rect 24672 38388 24728 38444
rect 5964 38332 6020 38388
rect 5628 38220 5684 38276
rect 11788 38220 11844 38276
rect 19852 38220 19908 38276
rect 3164 37996 3220 38052
rect 3804 37604 3860 37660
rect 3908 37604 3964 37660
rect 4012 37604 4068 37660
rect 23804 37604 23860 37660
rect 23908 37604 23964 37660
rect 24012 37604 24068 37660
rect 5852 37548 5908 37604
rect 18620 37548 18676 37604
rect 7532 37324 7588 37380
rect 17948 37212 18004 37268
rect 3164 36988 3220 37044
rect 5964 36988 6020 37044
rect 14812 36988 14868 37044
rect 15372 36988 15428 37044
rect 20188 36876 20244 36932
rect 4464 36820 4520 36876
rect 4568 36820 4624 36876
rect 4672 36820 4728 36876
rect 24464 36820 24520 36876
rect 24568 36820 24624 36876
rect 24672 36820 24728 36876
rect 11116 36764 11172 36820
rect 15036 36764 15092 36820
rect 10668 36540 10724 36596
rect 11116 36540 11172 36596
rect 14588 36316 14644 36372
rect 15708 36316 15764 36372
rect 18508 36204 18564 36260
rect 19292 36204 19348 36260
rect 17724 36092 17780 36148
rect 3804 36036 3860 36092
rect 3908 36036 3964 36092
rect 4012 36036 4068 36092
rect 23804 36036 23860 36092
rect 23908 36036 23964 36092
rect 24012 36036 24068 36092
rect 7532 35980 7588 36036
rect 17500 35868 17556 35924
rect 10220 35420 10276 35476
rect 15036 35420 15092 35476
rect 1372 35196 1428 35252
rect 4464 35252 4520 35308
rect 4568 35252 4624 35308
rect 4672 35252 4728 35308
rect 24464 35252 24520 35308
rect 24568 35252 24624 35308
rect 24672 35252 24728 35308
rect 4172 35196 4228 35252
rect 16828 35196 16884 35252
rect 14140 35084 14196 35140
rect 14700 35084 14756 35140
rect 1820 34972 1876 35028
rect 4284 34972 4340 35028
rect 13804 34860 13860 34916
rect 3612 34748 3668 34804
rect 17612 34748 17668 34804
rect 8540 34636 8596 34692
rect 3612 34524 3668 34580
rect 3804 34468 3860 34524
rect 3908 34468 3964 34524
rect 4012 34468 4068 34524
rect 23804 34468 23860 34524
rect 23908 34468 23964 34524
rect 24012 34468 24068 34524
rect 7532 34412 7588 34468
rect 13804 34412 13860 34468
rect 20412 34412 20468 34468
rect 10668 34300 10724 34356
rect 16828 34188 16884 34244
rect 1260 34076 1316 34132
rect 3500 34076 3556 34132
rect 6412 34076 6468 34132
rect 11788 34076 11844 34132
rect 16268 34076 16324 34132
rect 18844 34076 18900 34132
rect 2268 33964 2324 34020
rect 9212 33852 9268 33908
rect 14140 33852 14196 33908
rect 19628 33852 19684 33908
rect 1708 33740 1764 33796
rect 2828 33740 2884 33796
rect 4172 33740 4228 33796
rect 19740 33740 19796 33796
rect 4464 33684 4520 33740
rect 4568 33684 4624 33740
rect 4672 33684 4728 33740
rect 24464 33684 24520 33740
rect 24568 33684 24624 33740
rect 24672 33684 24728 33740
rect 1372 33628 1428 33684
rect 19852 33516 19908 33572
rect 1484 33404 1540 33460
rect 18620 33404 18676 33460
rect 17052 33292 17108 33348
rect 19292 33292 19348 33348
rect 6412 33180 6468 33236
rect 17724 33068 17780 33124
rect 8204 32956 8260 33012
rect 10332 32956 10388 33012
rect 3804 32900 3860 32956
rect 3908 32900 3964 32956
rect 4012 32900 4068 32956
rect 23804 32900 23860 32956
rect 23908 32900 23964 32956
rect 24012 32900 24068 32956
rect 6412 32732 6468 32788
rect 14476 32732 14532 32788
rect 14700 32732 14756 32788
rect 3276 32620 3332 32676
rect 19292 32620 19348 32676
rect 17276 32508 17332 32564
rect 19852 32508 19908 32564
rect 2828 32396 2884 32452
rect 5068 32396 5124 32452
rect 19740 32396 19796 32452
rect 6972 32284 7028 32340
rect 18620 32172 18676 32228
rect 4464 32116 4520 32172
rect 4568 32116 4624 32172
rect 4672 32116 4728 32172
rect 24464 32116 24520 32172
rect 24568 32116 24624 32172
rect 24672 32116 24728 32172
rect 16716 32060 16772 32116
rect 17948 32060 18004 32116
rect 6748 31948 6804 32004
rect 20188 31948 20244 32004
rect 2940 31836 2996 31892
rect 10220 31836 10276 31892
rect 11340 31836 11396 31892
rect 13468 31836 13524 31892
rect 4956 31724 5012 31780
rect 1820 31612 1876 31668
rect 6748 31612 6804 31668
rect 8204 31612 8260 31668
rect 12012 31500 12068 31556
rect 3804 31332 3860 31388
rect 3908 31332 3964 31388
rect 4012 31332 4068 31388
rect 23804 31332 23860 31388
rect 23908 31332 23964 31388
rect 24012 31332 24068 31388
rect 8764 31276 8820 31332
rect 16940 31164 16996 31220
rect 18508 31164 18564 31220
rect 4956 31052 5012 31108
rect 5404 31052 5460 31108
rect 2828 30940 2884 30996
rect 6748 30940 6804 30996
rect 20524 30828 20580 30884
rect 18956 30604 19012 30660
rect 4464 30548 4520 30604
rect 4568 30548 4624 30604
rect 4672 30548 4728 30604
rect 24464 30548 24520 30604
rect 24568 30548 24624 30604
rect 24672 30548 24728 30604
rect 13468 30380 13524 30436
rect 7980 30268 8036 30324
rect 15708 30268 15764 30324
rect 17388 29932 17444 29988
rect 3804 29764 3860 29820
rect 3908 29764 3964 29820
rect 4012 29764 4068 29820
rect 23804 29764 23860 29820
rect 23908 29764 23964 29820
rect 24012 29764 24068 29820
rect 10556 29708 10612 29764
rect 11116 29708 11172 29764
rect 18844 29708 18900 29764
rect 16828 29484 16884 29540
rect 18844 29372 18900 29428
rect 2268 29260 2324 29316
rect 5852 29260 5908 29316
rect 7644 29260 7700 29316
rect 9548 29260 9604 29316
rect 11116 29260 11172 29316
rect 17724 29260 17780 29316
rect 8204 29036 8260 29092
rect 4464 28980 4520 29036
rect 4568 28980 4624 29036
rect 4672 28980 4728 29036
rect 24464 28980 24520 29036
rect 24568 28980 24624 29036
rect 24672 28980 24728 29036
rect 2268 28812 2324 28868
rect 17836 28812 17892 28868
rect 18060 28812 18116 28868
rect 18844 28700 18900 28756
rect 19852 28588 19908 28644
rect 15036 28476 15092 28532
rect 17276 28364 17332 28420
rect 3804 28196 3860 28252
rect 3908 28196 3964 28252
rect 4012 28196 4068 28252
rect 23804 28196 23860 28252
rect 23908 28196 23964 28252
rect 24012 28196 24068 28252
rect 9100 28140 9156 28196
rect 18172 28140 18228 28196
rect 16828 28028 16884 28084
rect 1820 27916 1876 27972
rect 3612 27804 3668 27860
rect 7084 27692 7140 27748
rect 18732 27692 18788 27748
rect 19852 27692 19908 27748
rect 4464 27412 4520 27468
rect 4568 27412 4624 27468
rect 4672 27412 4728 27468
rect 24464 27412 24520 27468
rect 24568 27412 24624 27468
rect 24672 27412 24728 27468
rect 2380 27356 2436 27412
rect 13132 27244 13188 27300
rect 9100 27132 9156 27188
rect 2604 27020 2660 27076
rect 4172 27020 4228 27076
rect 6860 26908 6916 26964
rect 18172 26908 18228 26964
rect 19628 26908 19684 26964
rect 18620 26796 18676 26852
rect 9548 26684 9604 26740
rect 3804 26628 3860 26684
rect 3908 26628 3964 26684
rect 4012 26628 4068 26684
rect 23804 26628 23860 26684
rect 23908 26628 23964 26684
rect 24012 26628 24068 26684
rect 3612 26460 3668 26516
rect 4844 26460 4900 26516
rect 18732 26460 18788 26516
rect 20188 26348 20244 26404
rect 6972 26236 7028 26292
rect 16380 26236 16436 26292
rect 17500 26124 17556 26180
rect 3500 26012 3556 26068
rect 15036 26012 15092 26068
rect 3612 25900 3668 25956
rect 6748 25900 6804 25956
rect 9996 25900 10052 25956
rect 4464 25844 4520 25900
rect 4568 25844 4624 25900
rect 4672 25844 4728 25900
rect 24464 25844 24520 25900
rect 24568 25844 24624 25900
rect 24672 25844 24728 25900
rect 5852 25676 5908 25732
rect 9996 25676 10052 25732
rect 20076 25676 20132 25732
rect 5404 25564 5460 25620
rect 4172 25452 4228 25508
rect 9548 25340 9604 25396
rect 5292 25228 5348 25284
rect 8540 25228 8596 25284
rect 16380 25228 16436 25284
rect 12012 25116 12068 25172
rect 16268 25116 16324 25172
rect 3804 25060 3860 25116
rect 3908 25060 3964 25116
rect 4012 25060 4068 25116
rect 23804 25060 23860 25116
rect 23908 25060 23964 25116
rect 24012 25060 24068 25116
rect 4172 25004 4228 25060
rect 3500 24556 3556 24612
rect 10668 24556 10724 24612
rect 16716 24556 16772 24612
rect 11788 24444 11844 24500
rect 7420 24332 7476 24388
rect 4464 24276 4520 24332
rect 4568 24276 4624 24332
rect 4672 24276 4728 24332
rect 24464 24276 24520 24332
rect 24568 24276 24624 24332
rect 24672 24276 24728 24332
rect 4172 24220 4228 24276
rect 140 23996 196 24052
rect 3052 23996 3108 24052
rect 14812 23996 14868 24052
rect 252 23884 308 23940
rect 5740 23884 5796 23940
rect 6188 23884 6244 23940
rect 1820 23772 1876 23828
rect 4172 23548 4228 23604
rect 7420 23548 7476 23604
rect 7980 23548 8036 23604
rect 19404 23548 19460 23604
rect 3804 23492 3860 23548
rect 3908 23492 3964 23548
rect 4012 23492 4068 23548
rect 23804 23492 23860 23548
rect 23908 23492 23964 23548
rect 24012 23492 24068 23548
rect 12684 23436 12740 23492
rect 14924 23436 14980 23492
rect 18732 23436 18788 23492
rect 23100 23436 23156 23492
rect 13580 23324 13636 23380
rect 14028 23324 14084 23380
rect 2268 23212 2324 23268
rect 4844 22988 4900 23044
rect 5404 22988 5460 23044
rect 14364 22988 14420 23044
rect 16492 22988 16548 23044
rect 18060 22988 18116 23044
rect 18956 22988 19012 23044
rect 2156 22876 2212 22932
rect 3164 22876 3220 22932
rect 5628 22876 5684 22932
rect 18844 22876 18900 22932
rect 23100 22876 23156 22932
rect 13916 22764 13972 22820
rect 4464 22708 4520 22764
rect 4568 22708 4624 22764
rect 4672 22708 4728 22764
rect 24464 22708 24520 22764
rect 24568 22708 24624 22764
rect 24672 22708 24728 22764
rect 4844 22652 4900 22708
rect 5740 22652 5796 22708
rect 2492 22316 2548 22372
rect 23660 22204 23716 22260
rect 1932 22092 1988 22148
rect 14700 22092 14756 22148
rect 21756 22092 21812 22148
rect 7980 21980 8036 22036
rect 3804 21924 3860 21980
rect 3908 21924 3964 21980
rect 4012 21924 4068 21980
rect 23804 21924 23860 21980
rect 23908 21924 23964 21980
rect 24012 21924 24068 21980
rect 7084 21868 7140 21924
rect 15036 21756 15092 21812
rect 3612 21644 3668 21700
rect 13132 21644 13188 21700
rect 13580 21532 13636 21588
rect 14700 21420 14756 21476
rect 21420 21420 21476 21476
rect 14364 21196 14420 21252
rect 4464 21140 4520 21196
rect 4568 21140 4624 21196
rect 4672 21140 4728 21196
rect 24464 21140 24520 21196
rect 24568 21140 24624 21196
rect 24672 21140 24728 21196
rect 6188 20972 6244 21028
rect 12012 20972 12068 21028
rect 13916 20972 13972 21028
rect 16492 20972 16548 21028
rect 6972 20860 7028 20916
rect 18060 20860 18116 20916
rect 4844 20524 4900 20580
rect 5068 20524 5124 20580
rect 7980 20412 8036 20468
rect 3804 20356 3860 20412
rect 3908 20356 3964 20412
rect 4012 20356 4068 20412
rect 23804 20356 23860 20412
rect 23908 20356 23964 20412
rect 24012 20356 24068 20412
rect 10780 20188 10836 20244
rect 12012 20188 12068 20244
rect 26012 20188 26068 20244
rect 7420 20076 7476 20132
rect 9436 20076 9492 20132
rect 5404 19964 5460 20020
rect 7196 19964 7252 20020
rect 9548 19852 9604 19908
rect 4844 19628 4900 19684
rect 4464 19572 4520 19628
rect 4568 19572 4624 19628
rect 4672 19572 4728 19628
rect 24464 19572 24520 19628
rect 24568 19572 24624 19628
rect 24672 19572 24728 19628
rect 3276 19516 3332 19572
rect 13580 19516 13636 19572
rect 14252 19516 14308 19572
rect 4844 19404 4900 19460
rect 6748 19292 6804 19348
rect 9100 19292 9156 19348
rect 3804 18788 3860 18844
rect 3908 18788 3964 18844
rect 4012 18788 4068 18844
rect 23804 18788 23860 18844
rect 23908 18788 23964 18844
rect 24012 18788 24068 18844
rect 6076 18732 6132 18788
rect 9772 18620 9828 18676
rect 23660 18620 23716 18676
rect 3388 18508 3444 18564
rect 4956 18508 5012 18564
rect 13132 18508 13188 18564
rect 8988 18396 9044 18452
rect 2156 18284 2212 18340
rect 12908 18284 12964 18340
rect 14812 18284 14868 18340
rect 16940 18284 16996 18340
rect 5628 18172 5684 18228
rect 4464 18004 4520 18060
rect 4568 18004 4624 18060
rect 4672 18004 4728 18060
rect 24464 18004 24520 18060
rect 24568 18004 24624 18060
rect 24672 18004 24728 18060
rect 4172 17724 4228 17780
rect 7084 17724 7140 17780
rect 21644 17724 21700 17780
rect 3612 17612 3668 17668
rect 5852 17276 5908 17332
rect 3804 17220 3860 17276
rect 3908 17220 3964 17276
rect 4012 17220 4068 17276
rect 23804 17220 23860 17276
rect 23908 17220 23964 17276
rect 24012 17220 24068 17276
rect 7196 17052 7252 17108
rect 3276 16940 3332 16996
rect 13356 16940 13412 16996
rect 13804 16940 13860 16996
rect 6300 16828 6356 16884
rect 8204 16716 8260 16772
rect 22316 16716 22372 16772
rect 5628 16604 5684 16660
rect 11116 16604 11172 16660
rect 14364 16604 14420 16660
rect 17836 16604 17892 16660
rect 22652 16604 22708 16660
rect 4464 16436 4520 16492
rect 4568 16436 4624 16492
rect 4672 16436 4728 16492
rect 24464 16436 24520 16492
rect 24568 16436 24624 16492
rect 24672 16436 24728 16492
rect 5740 16380 5796 16436
rect 15932 16268 15988 16324
rect 4284 16044 4340 16100
rect 14924 16044 14980 16100
rect 26572 15932 26628 15988
rect 12460 15820 12516 15876
rect 5628 15708 5684 15764
rect 3804 15652 3860 15708
rect 3908 15652 3964 15708
rect 4012 15652 4068 15708
rect 23804 15652 23860 15708
rect 23908 15652 23964 15708
rect 24012 15652 24068 15708
rect 5404 15596 5460 15652
rect 5068 15484 5124 15540
rect 12460 15372 12516 15428
rect 1484 15036 1540 15092
rect 5628 14924 5684 14980
rect 17052 14924 17108 14980
rect 4464 14868 4520 14924
rect 4568 14868 4624 14924
rect 4672 14868 4728 14924
rect 24464 14868 24520 14924
rect 24568 14868 24624 14924
rect 24672 14868 24728 14924
rect 4956 14588 5012 14644
rect 26012 14588 26068 14644
rect 26572 14588 26628 14644
rect 6300 14476 6356 14532
rect 13132 14476 13188 14532
rect 14028 14476 14084 14532
rect 10668 14364 10724 14420
rect 11116 14364 11172 14420
rect 13804 14364 13860 14420
rect 19516 14364 19572 14420
rect 2716 14252 2772 14308
rect 3612 14140 3668 14196
rect 4956 14140 5012 14196
rect 12684 14140 12740 14196
rect 3804 14084 3860 14140
rect 3908 14084 3964 14140
rect 4012 14084 4068 14140
rect 23804 14084 23860 14140
rect 23908 14084 23964 14140
rect 24012 14084 24068 14140
rect 3164 13916 3220 13972
rect 14028 13692 14084 13748
rect 4844 13580 4900 13636
rect 6636 13580 6692 13636
rect 16940 13580 16996 13636
rect 3276 13468 3332 13524
rect 6300 13468 6356 13524
rect 10556 13468 10612 13524
rect 3052 13356 3108 13412
rect 3500 13356 3556 13412
rect 4464 13300 4520 13356
rect 4568 13300 4624 13356
rect 4672 13300 4728 13356
rect 24464 13300 24520 13356
rect 24568 13300 24624 13356
rect 24672 13300 24728 13356
rect 13804 13244 13860 13300
rect 2380 13132 2436 13188
rect 5180 13020 5236 13076
rect 8092 12908 8148 12964
rect 5068 12796 5124 12852
rect 4956 12572 5012 12628
rect 19964 12572 20020 12628
rect 3804 12516 3860 12572
rect 3908 12516 3964 12572
rect 4012 12516 4068 12572
rect 23804 12516 23860 12572
rect 23908 12516 23964 12572
rect 24012 12516 24068 12572
rect 27692 12348 27748 12404
rect 1260 12236 1316 12292
rect 3612 12236 3668 12292
rect 2380 11900 2436 11956
rect 19516 11900 19572 11956
rect 5740 11788 5796 11844
rect 4464 11732 4520 11788
rect 4568 11732 4624 11788
rect 4672 11732 4728 11788
rect 24464 11732 24520 11788
rect 24568 11732 24624 11788
rect 24672 11732 24728 11788
rect 5404 11676 5460 11732
rect 3388 11564 3444 11620
rect 21644 11228 21700 11284
rect 5852 11116 5908 11172
rect 3804 10948 3860 11004
rect 3908 10948 3964 11004
rect 4012 10948 4068 11004
rect 23804 10948 23860 11004
rect 23908 10948 23964 11004
rect 24012 10948 24068 11004
rect 3388 10892 3444 10948
rect 4956 10892 5012 10948
rect 2940 10780 2996 10836
rect 9660 10668 9716 10724
rect 22092 10668 22148 10724
rect 4284 10444 4340 10500
rect 5964 10444 6020 10500
rect 11788 10444 11844 10500
rect 2156 10332 2212 10388
rect 22988 10332 23044 10388
rect 4284 10220 4340 10276
rect 4464 10164 4520 10220
rect 4568 10164 4624 10220
rect 4672 10164 4728 10220
rect 24464 10164 24520 10220
rect 24568 10164 24624 10220
rect 24672 10164 24728 10220
rect 2492 9996 2548 10052
rect 25116 9996 25172 10052
rect 700 9772 756 9828
rect 14028 9772 14084 9828
rect 2044 9548 2100 9604
rect 6188 9436 6244 9492
rect 10668 9436 10724 9492
rect 3804 9380 3860 9436
rect 3908 9380 3964 9436
rect 4012 9380 4068 9436
rect 23804 9380 23860 9436
rect 23908 9380 23964 9436
rect 24012 9380 24068 9436
rect 5628 9324 5684 9380
rect 2940 9100 2996 9156
rect 7084 9100 7140 9156
rect 13580 9100 13636 9156
rect 2828 8988 2884 9044
rect 4284 8988 4340 9044
rect 5292 8988 5348 9044
rect 6860 8988 6916 9044
rect 15484 8988 15540 9044
rect 3612 8764 3668 8820
rect 4464 8596 4520 8652
rect 4568 8596 4624 8652
rect 4672 8596 4728 8652
rect 24464 8596 24520 8652
rect 24568 8596 24624 8652
rect 24672 8596 24728 8652
rect 8428 8540 8484 8596
rect 9436 8540 9492 8596
rect 7532 8316 7588 8372
rect 19516 8316 19572 8372
rect 1484 8204 1540 8260
rect 14028 8204 14084 8260
rect 3612 8092 3668 8148
rect 8652 7980 8708 8036
rect 22204 7980 22260 8036
rect 25452 7980 25508 8036
rect 3804 7812 3860 7868
rect 3908 7812 3964 7868
rect 4012 7812 4068 7868
rect 23804 7812 23860 7868
rect 23908 7812 23964 7868
rect 24012 7812 24068 7868
rect 16604 7756 16660 7812
rect 21644 7756 21700 7812
rect 21308 7644 21364 7700
rect 25004 7644 25060 7700
rect 28588 7532 28644 7588
rect 9436 7420 9492 7476
rect 15484 7420 15540 7476
rect 2268 7308 2324 7364
rect 3388 7308 3444 7364
rect 11788 7308 11844 7364
rect 24892 7308 24948 7364
rect 7980 7196 8036 7252
rect 4464 7028 4520 7084
rect 4568 7028 4624 7084
rect 4672 7028 4728 7084
rect 2492 6972 2548 7028
rect 14140 6972 14196 7028
rect 24464 7028 24520 7084
rect 24568 7028 24624 7084
rect 24672 7028 24728 7084
rect 25788 6972 25844 7028
rect 5628 6860 5684 6916
rect 23660 6860 23716 6916
rect 4284 6748 4340 6804
rect 9212 6748 9268 6804
rect 15484 6748 15540 6804
rect 1372 6636 1428 6692
rect 2156 6636 2212 6692
rect 2380 6636 2436 6692
rect 3388 6636 3444 6692
rect 9548 6636 9604 6692
rect 6412 6524 6468 6580
rect 8092 6524 8148 6580
rect 14252 6524 14308 6580
rect 25564 6524 25620 6580
rect 3804 6244 3860 6300
rect 3908 6244 3964 6300
rect 4012 6244 4068 6300
rect 23804 6244 23860 6300
rect 23908 6244 23964 6300
rect 24012 6244 24068 6300
rect 3500 5852 3556 5908
rect 5068 5852 5124 5908
rect 15484 5852 15540 5908
rect 25564 5852 25620 5908
rect 4172 5740 4228 5796
rect 21644 5516 21700 5572
rect 4464 5460 4520 5516
rect 4568 5460 4624 5516
rect 4672 5460 4728 5516
rect 24464 5460 24520 5516
rect 24568 5460 24624 5516
rect 24672 5460 24728 5516
rect 7532 5404 7588 5460
rect 10668 5404 10724 5460
rect 25228 5404 25284 5460
rect 1260 5292 1316 5348
rect 2044 5292 2100 5348
rect 15372 5292 15428 5348
rect 23324 5292 23380 5348
rect 25116 5292 25172 5348
rect 6412 5180 6468 5236
rect 26348 5180 26404 5236
rect 8652 5068 8708 5124
rect 14252 5068 14308 5124
rect 24220 5068 24276 5124
rect 8428 4844 8484 4900
rect 27692 4732 27748 4788
rect 3804 4676 3860 4732
rect 3908 4676 3964 4732
rect 4012 4676 4068 4732
rect 23804 4676 23860 4732
rect 23908 4676 23964 4732
rect 24012 4676 24068 4732
rect 2828 4620 2884 4676
rect 11564 4620 11620 4676
rect 5404 4508 5460 4564
rect 18732 4396 18788 4452
rect 8876 4284 8932 4340
rect 11340 4284 11396 4340
rect 12236 4284 12292 4340
rect 13356 4284 13412 4340
rect 18284 4284 18340 4340
rect 3276 4060 3332 4116
rect 7980 4060 8036 4116
rect 9660 3948 9716 4004
rect 15932 3948 15988 4004
rect 4464 3892 4520 3948
rect 4568 3892 4624 3948
rect 4672 3892 4728 3948
rect 24464 3892 24520 3948
rect 24568 3892 24624 3948
rect 24672 3892 24728 3948
rect 26684 3836 26740 3892
rect 9772 3724 9828 3780
rect 23548 3724 23604 3780
rect 9212 3500 9268 3556
rect 11004 3500 11060 3556
rect 13692 3500 13748 3556
rect 14476 3500 14532 3556
rect 17164 3500 17220 3556
rect 26796 3500 26852 3556
rect 6300 3388 6356 3444
rect 17724 3388 17780 3444
rect 5852 3276 5908 3332
rect 10220 3276 10276 3332
rect 3804 3108 3860 3164
rect 3908 3108 3964 3164
rect 4012 3108 4068 3164
rect 13468 3052 13524 3108
rect 23100 3052 23156 3108
rect 23804 3108 23860 3164
rect 23908 3108 23964 3164
rect 24012 3108 24068 3164
rect 4844 2940 4900 2996
rect 16604 2940 16660 2996
rect 25900 2940 25956 2996
rect 28588 2940 28644 2996
rect 4956 2828 5012 2884
rect 3612 2716 3668 2772
rect 7756 2716 7812 2772
rect 15596 2716 15652 2772
rect 18620 2716 18676 2772
rect 25452 2716 25508 2772
rect 26124 2716 26180 2772
rect 3164 2604 3220 2660
rect 5740 2604 5796 2660
rect 11564 2604 11620 2660
rect 14140 2492 14196 2548
rect 10220 2380 10276 2436
rect 4464 2324 4520 2380
rect 4568 2324 4624 2380
rect 4672 2324 4728 2380
rect 24464 2324 24520 2380
rect 24568 2324 24624 2380
rect 24672 2324 24728 2380
rect 2492 2268 2548 2324
rect 23548 2268 23604 2324
rect 25228 2268 25284 2324
rect 26684 2268 26740 2324
rect 2828 2156 2884 2212
rect 15708 2156 15764 2212
rect 22092 2156 22148 2212
rect 23100 2156 23156 2212
rect 26348 2156 26404 2212
rect 2940 2044 2996 2100
rect 13468 2044 13524 2100
rect 23548 2044 23604 2100
rect 14476 1932 14532 1988
rect 10220 1820 10276 1876
rect 25900 1820 25956 1876
rect 7084 1708 7140 1764
rect 700 1596 756 1652
rect 6076 1596 6132 1652
rect 6524 1596 6580 1652
rect 6748 1596 6804 1652
rect 6972 1596 7028 1652
rect 7420 1596 7476 1652
rect 7644 1596 7700 1652
rect 7868 1596 7924 1652
rect 8316 1596 8372 1652
rect 8540 1596 8596 1652
rect 8764 1596 8820 1652
rect 9324 1596 9380 1652
rect 10108 1596 10164 1652
rect 10332 1596 10388 1652
rect 11228 1596 11284 1652
rect 11452 1596 11508 1652
rect 11900 1596 11956 1652
rect 12124 1596 12180 1652
rect 12348 1596 12404 1652
rect 12572 1596 12628 1652
rect 12796 1596 12852 1652
rect 13020 1596 13076 1652
rect 13244 1596 13300 1652
rect 25004 1596 25060 1652
rect 3804 1540 3860 1596
rect 3908 1540 3964 1596
rect 4012 1540 4068 1596
rect 23804 1540 23860 1596
rect 23908 1540 23964 1596
rect 24012 1540 24068 1596
rect 7756 1484 7812 1540
rect 9212 1484 9268 1540
rect 10556 1484 10612 1540
rect 10892 1484 10948 1540
rect 21532 1484 21588 1540
rect 27020 1484 27076 1540
rect 5964 1372 6020 1428
rect 23660 1372 23716 1428
rect 26236 1372 26292 1428
rect 11340 1260 11396 1316
rect 23436 1260 23492 1316
rect 25116 1260 25172 1316
rect 2716 1148 2772 1204
rect 15148 1148 15204 1204
rect 28028 1148 28084 1204
rect 9212 924 9268 980
rect 9884 924 9940 980
rect 11116 924 11172 980
rect 11340 924 11396 980
rect 25788 812 25844 868
rect 4464 756 4520 812
rect 4568 756 4624 812
rect 4672 756 4728 812
rect 24464 756 24520 812
rect 24568 756 24624 812
rect 24672 756 24728 812
rect 11676 588 11732 644
rect 24220 588 24276 644
rect 24892 588 24948 644
rect 25116 476 25172 532
rect 9324 364 9380 420
rect 19964 252 20020 308
rect 9324 28 9380 84
rect 14252 28 14308 84
rect 19964 28 20020 84
<< metal4 >>
rect 3776 112924 4096 114912
rect 3776 112868 3804 112924
rect 3860 112868 3908 112924
rect 3964 112868 4012 112924
rect 4068 112868 4096 112924
rect 1820 112308 1876 112318
rect 1596 109284 1652 109294
rect 1596 106318 1652 109228
rect 1484 106262 1652 106318
rect 1708 107828 1764 107838
rect 1484 106148 1540 106262
rect 1484 102788 1540 106092
rect 1372 102452 1428 102462
rect 140 99652 196 99662
rect 140 87332 196 99596
rect 252 98532 308 98542
rect 252 89908 308 98476
rect 1372 95956 1428 102396
rect 1372 95890 1428 95900
rect 476 95844 532 95854
rect 476 93492 532 95788
rect 476 93426 532 93436
rect 1484 92036 1540 102732
rect 1484 91970 1540 91980
rect 1596 104020 1652 104030
rect 252 89842 308 89852
rect 140 87266 196 87276
rect 1372 87444 1428 87454
rect 700 83524 756 83534
rect 700 74788 756 83468
rect 1372 79858 1428 87388
rect 1596 86100 1652 103964
rect 1708 96180 1764 107772
rect 1708 96114 1764 96124
rect 1708 89012 1764 89022
rect 1708 87556 1764 88956
rect 1708 87490 1764 87500
rect 1596 86034 1652 86044
rect 1820 85876 1876 112252
rect 3500 111748 3556 111758
rect 3500 111076 3556 111692
rect 3500 111010 3556 111020
rect 3776 111356 4096 112868
rect 3776 111300 3804 111356
rect 3860 111300 3908 111356
rect 3964 111300 4012 111356
rect 4068 111300 4096 111356
rect 3776 109788 4096 111300
rect 3776 109732 3804 109788
rect 3860 109732 3908 109788
rect 3964 109732 4012 109788
rect 4068 109732 4096 109788
rect 3388 109620 3444 109630
rect 3388 108724 3444 109564
rect 3612 109396 3668 109406
rect 3388 108658 3444 108668
rect 3500 109060 3556 109070
rect 3276 108276 3332 108286
rect 3276 107828 3332 108220
rect 2380 107044 2436 107054
rect 2156 106484 2212 106494
rect 2044 106260 2100 106270
rect 1820 85810 1876 85820
rect 1932 106036 1988 106046
rect 1484 85764 1540 85774
rect 1484 85428 1540 85708
rect 1484 85362 1540 85372
rect 1820 82740 1876 82750
rect 1708 80164 1764 80174
rect 1372 79802 1540 79858
rect 700 74722 756 74732
rect 1260 76244 1316 76254
rect 924 74564 980 74574
rect 924 72100 980 74508
rect 924 72034 980 72044
rect 1036 68628 1092 68638
rect 1036 67844 1092 68572
rect 1036 67778 1092 67788
rect 1260 65716 1316 76188
rect 1372 74116 1428 74126
rect 1372 68740 1428 74060
rect 1372 68674 1428 68684
rect 1260 65650 1316 65660
rect 1372 58212 1428 58222
rect 1372 44758 1428 58156
rect 1260 44702 1428 44758
rect 1148 42644 1204 42654
rect 1148 40628 1204 42588
rect 1148 40562 1204 40572
rect 1260 34132 1316 44702
rect 1484 44578 1540 79802
rect 1708 79604 1764 80108
rect 1708 79538 1764 79548
rect 1708 79044 1764 79054
rect 1596 77364 1652 77374
rect 1596 72548 1652 77308
rect 1708 76580 1764 78988
rect 1820 78372 1876 82684
rect 1820 78306 1876 78316
rect 1708 76514 1764 76524
rect 1596 72482 1652 72492
rect 1820 72884 1876 72894
rect 1820 70420 1876 72828
rect 1820 70354 1876 70364
rect 1932 58212 1988 105980
rect 2044 86884 2100 106204
rect 2156 103124 2212 106428
rect 2156 103058 2212 103068
rect 2268 105700 2324 105710
rect 2268 104356 2324 105644
rect 2268 102898 2324 104300
rect 2044 86818 2100 86828
rect 2156 102842 2324 102898
rect 2044 84084 2100 84094
rect 2044 61796 2100 84028
rect 2156 81844 2212 102842
rect 2380 100996 2436 106988
rect 3276 107044 3332 107772
rect 3276 106978 3332 106988
rect 3052 106260 3108 106270
rect 2716 105588 2772 105598
rect 2156 81778 2212 81788
rect 2268 99316 2324 99326
rect 2044 61730 2100 61740
rect 2268 58772 2324 99260
rect 2380 99092 2436 100940
rect 2380 99026 2436 99036
rect 2604 104244 2660 104254
rect 2604 103796 2660 104188
rect 2604 96292 2660 103740
rect 2604 96226 2660 96236
rect 2716 104020 2772 105532
rect 2716 100660 2772 103964
rect 2380 95844 2436 95854
rect 2380 90356 2436 95788
rect 2492 94500 2548 94510
rect 2492 94164 2548 94444
rect 2492 94098 2548 94108
rect 2380 90290 2436 90300
rect 2604 89572 2660 89582
rect 2380 86212 2436 86222
rect 2380 82292 2436 86156
rect 2380 82226 2436 82236
rect 2492 81844 2548 81854
rect 2492 63812 2548 81788
rect 2492 62580 2548 63756
rect 2492 62514 2548 62524
rect 2268 58706 2324 58716
rect 1932 58146 1988 58156
rect 2604 55076 2660 89516
rect 2716 83636 2772 100604
rect 2716 79044 2772 83580
rect 2940 85204 2996 85214
rect 2716 76356 2772 78988
rect 2716 73556 2772 76300
rect 2716 73490 2772 73500
rect 2828 80388 2884 80398
rect 2828 73332 2884 80332
rect 2828 73266 2884 73276
rect 2940 70084 2996 85148
rect 3052 84084 3108 106204
rect 3500 105924 3556 109004
rect 3612 107380 3668 109340
rect 3612 107314 3668 107324
rect 3776 108220 4096 109732
rect 4284 114548 4340 114558
rect 3776 108164 3804 108220
rect 3860 108164 3908 108220
rect 3964 108164 4012 108220
rect 4068 108164 4096 108220
rect 3500 105858 3556 105868
rect 3776 106652 4096 108164
rect 3776 106596 3804 106652
rect 3860 106596 3908 106652
rect 3964 106596 4012 106652
rect 4068 106596 4096 106652
rect 3612 105476 3668 105486
rect 3500 103236 3556 103246
rect 3500 100772 3556 103180
rect 3612 101444 3668 105420
rect 3612 101378 3668 101388
rect 3776 105084 4096 106596
rect 3776 105028 3804 105084
rect 3860 105028 3908 105084
rect 3964 105028 4012 105084
rect 4068 105028 4096 105084
rect 3776 103516 4096 105028
rect 3776 103460 3804 103516
rect 3860 103460 3908 103516
rect 3964 103460 4012 103516
rect 4068 103460 4096 103516
rect 3776 101948 4096 103460
rect 3776 101892 3804 101948
rect 3860 101892 3908 101948
rect 3964 101892 4012 101948
rect 4068 101892 4096 101948
rect 3388 99204 3444 99214
rect 3276 98980 3332 98990
rect 3276 97076 3332 98924
rect 3164 93828 3220 93838
rect 3164 84532 3220 93772
rect 3276 88116 3332 97020
rect 3388 89796 3444 99148
rect 3500 96068 3556 100716
rect 3612 101220 3668 101230
rect 3612 99316 3668 101164
rect 3612 99250 3668 99260
rect 3776 100380 4096 101892
rect 3776 100324 3804 100380
rect 3860 100324 3908 100380
rect 3964 100324 4012 100380
rect 4068 100324 4096 100380
rect 3776 98812 4096 100324
rect 3776 98756 3804 98812
rect 3860 98756 3908 98812
rect 3964 98756 4012 98812
rect 4068 98756 4096 98812
rect 3776 97244 4096 98756
rect 3776 97188 3804 97244
rect 3860 97188 3908 97244
rect 3964 97188 4012 97244
rect 4068 97188 4096 97244
rect 3500 96002 3556 96012
rect 3612 96740 3668 96750
rect 3612 95844 3668 96684
rect 3612 95778 3668 95788
rect 3776 95676 4096 97188
rect 3776 95620 3804 95676
rect 3860 95620 3908 95676
rect 3964 95620 4012 95676
rect 4068 95620 4096 95676
rect 3612 95396 3668 95406
rect 3500 95172 3556 95182
rect 3500 94836 3556 95116
rect 3500 94770 3556 94780
rect 3388 89730 3444 89740
rect 3500 94052 3556 94062
rect 3500 88228 3556 93996
rect 3612 90580 3668 95340
rect 3612 90514 3668 90524
rect 3776 94108 4096 95620
rect 3776 94052 3804 94108
rect 3860 94052 3908 94108
rect 3964 94052 4012 94108
rect 4068 94052 4096 94108
rect 3776 92540 4096 94052
rect 3776 92484 3804 92540
rect 3860 92484 3908 92540
rect 3964 92484 4012 92540
rect 4068 92484 4096 92540
rect 3776 90972 4096 92484
rect 3776 90916 3804 90972
rect 3860 90916 3908 90972
rect 3964 90916 4012 90972
rect 4068 90916 4096 90972
rect 3500 88162 3556 88172
rect 3776 89404 4096 90916
rect 3776 89348 3804 89404
rect 3860 89348 3908 89404
rect 3964 89348 4012 89404
rect 4068 89348 4096 89404
rect 3276 88050 3332 88060
rect 3776 87836 4096 89348
rect 3776 87780 3804 87836
rect 3860 87780 3908 87836
rect 3964 87780 4012 87836
rect 4068 87780 4096 87836
rect 3388 87668 3444 87678
rect 3388 85764 3444 87612
rect 3388 85698 3444 85708
rect 3776 86268 4096 87780
rect 3776 86212 3804 86268
rect 3860 86212 3908 86268
rect 3964 86212 4012 86268
rect 4068 86212 4096 86268
rect 3164 84466 3220 84476
rect 3776 84700 4096 86212
rect 3776 84644 3804 84700
rect 3860 84644 3908 84700
rect 3964 84644 4012 84700
rect 4068 84644 4096 84700
rect 3052 84018 3108 84028
rect 3776 83132 4096 84644
rect 3776 83076 3804 83132
rect 3860 83076 3908 83132
rect 3964 83076 4012 83132
rect 4068 83076 4096 83132
rect 3776 81564 4096 83076
rect 3776 81508 3804 81564
rect 3860 81508 3908 81564
rect 3964 81508 4012 81564
rect 4068 81508 4096 81564
rect 3612 80500 3668 80510
rect 3276 80388 3332 80398
rect 3164 77812 3220 77822
rect 3164 74452 3220 77756
rect 3276 76078 3332 80332
rect 3388 79380 3444 79390
rect 3388 76468 3444 79324
rect 3612 76978 3668 80444
rect 3388 76402 3444 76412
rect 3500 76922 3668 76978
rect 3776 79996 4096 81508
rect 3776 79940 3804 79996
rect 3860 79940 3908 79996
rect 3964 79940 4012 79996
rect 4068 79940 4096 79996
rect 3776 78428 4096 79940
rect 3776 78372 3804 78428
rect 3860 78372 3908 78428
rect 3964 78372 4012 78428
rect 4068 78372 4096 78428
rect 3500 76258 3556 76922
rect 3776 76860 4096 78372
rect 3612 76804 3668 76814
rect 3612 76468 3668 76748
rect 3612 76402 3668 76412
rect 3776 76804 3804 76860
rect 3860 76804 3908 76860
rect 3964 76804 4012 76860
rect 4068 76804 4096 76860
rect 3500 76202 3668 76258
rect 3276 76022 3556 76078
rect 3164 74386 3220 74396
rect 3500 74228 3556 76022
rect 3500 70980 3556 74172
rect 3500 70914 3556 70924
rect 2940 70018 2996 70028
rect 3276 69412 3332 69422
rect 3276 62468 3332 69356
rect 3500 67732 3556 67742
rect 3388 67284 3444 67294
rect 3388 66164 3444 67228
rect 3388 66098 3444 66108
rect 3500 65380 3556 67676
rect 3500 65314 3556 65324
rect 3612 64820 3668 76202
rect 3612 64754 3668 64764
rect 3776 75292 4096 76804
rect 3776 75236 3804 75292
rect 3860 75236 3908 75292
rect 3964 75236 4012 75292
rect 4068 75236 4096 75292
rect 3776 73724 4096 75236
rect 3776 73668 3804 73724
rect 3860 73668 3908 73724
rect 3964 73668 4012 73724
rect 4068 73668 4096 73724
rect 3776 72156 4096 73668
rect 3776 72100 3804 72156
rect 3860 72100 3908 72156
rect 3964 72100 4012 72156
rect 4068 72100 4096 72156
rect 3776 70588 4096 72100
rect 3776 70532 3804 70588
rect 3860 70532 3908 70588
rect 3964 70532 4012 70588
rect 4068 70532 4096 70588
rect 3776 69020 4096 70532
rect 3776 68964 3804 69020
rect 3860 68964 3908 69020
rect 3964 68964 4012 69020
rect 4068 68964 4096 69020
rect 3776 67452 4096 68964
rect 3776 67396 3804 67452
rect 3860 67396 3908 67452
rect 3964 67396 4012 67452
rect 4068 67396 4096 67452
rect 3776 65884 4096 67396
rect 4172 109284 4228 109294
rect 4172 67396 4228 109228
rect 4284 108948 4340 114492
rect 4284 108882 4340 108892
rect 4436 113708 4756 114912
rect 6636 114660 6692 114670
rect 4436 113652 4464 113708
rect 4520 113652 4568 113708
rect 4624 113652 4672 113708
rect 4728 113652 4756 113708
rect 4436 112140 4756 113652
rect 5404 113876 5460 113886
rect 5292 113428 5348 113438
rect 4436 112084 4464 112140
rect 4520 112084 4568 112140
rect 4624 112084 4672 112140
rect 4728 112084 4756 112140
rect 4436 110572 4756 112084
rect 4436 110516 4464 110572
rect 4520 110516 4568 110572
rect 4624 110516 4672 110572
rect 4728 110516 4756 110572
rect 4436 109004 4756 110516
rect 4956 112980 5012 112990
rect 4956 110292 5012 112924
rect 5180 112756 5236 112766
rect 4956 110226 5012 110236
rect 5068 112308 5124 112318
rect 4844 109732 4900 109742
rect 4844 109284 4900 109676
rect 4844 109218 4900 109228
rect 4436 108948 4464 109004
rect 4520 108948 4568 109004
rect 4624 108948 4672 109004
rect 4728 108948 4756 109004
rect 5068 109060 5124 112252
rect 5068 108994 5124 109004
rect 4284 107604 4340 107614
rect 4284 95284 4340 107548
rect 4284 95218 4340 95228
rect 4436 107436 4756 108948
rect 4436 107380 4464 107436
rect 4520 107380 4568 107436
rect 4624 107380 4672 107436
rect 4728 107380 4756 107436
rect 4436 105868 4756 107380
rect 4436 105812 4464 105868
rect 4520 105812 4568 105868
rect 4624 105812 4672 105868
rect 4728 105812 4756 105868
rect 4436 104300 4756 105812
rect 4956 108500 5012 108510
rect 4436 104244 4464 104300
rect 4520 104244 4568 104300
rect 4624 104244 4672 104300
rect 4728 104244 4756 104300
rect 4436 102732 4756 104244
rect 4436 102676 4464 102732
rect 4520 102676 4568 102732
rect 4624 102676 4672 102732
rect 4728 102676 4756 102732
rect 4436 101164 4756 102676
rect 4436 101108 4464 101164
rect 4520 101108 4568 101164
rect 4624 101108 4672 101164
rect 4728 101108 4756 101164
rect 4436 99596 4756 101108
rect 4436 99540 4464 99596
rect 4520 99540 4568 99596
rect 4624 99540 4672 99596
rect 4728 99540 4756 99596
rect 4436 98028 4756 99540
rect 4436 97972 4464 98028
rect 4520 97972 4568 98028
rect 4624 97972 4672 98028
rect 4728 97972 4756 98028
rect 4436 96460 4756 97972
rect 4436 96404 4464 96460
rect 4520 96404 4568 96460
rect 4624 96404 4672 96460
rect 4728 96404 4756 96460
rect 4436 94892 4756 96404
rect 4284 94836 4340 94846
rect 4284 93828 4340 94780
rect 4284 77140 4340 93772
rect 4284 74900 4340 77084
rect 4284 74834 4340 74844
rect 4436 94836 4464 94892
rect 4520 94836 4568 94892
rect 4624 94836 4672 94892
rect 4728 94836 4756 94892
rect 4436 93324 4756 94836
rect 4436 93268 4464 93324
rect 4520 93268 4568 93324
rect 4624 93268 4672 93324
rect 4728 93268 4756 93324
rect 4436 91756 4756 93268
rect 4436 91700 4464 91756
rect 4520 91700 4568 91756
rect 4624 91700 4672 91756
rect 4728 91700 4756 91756
rect 4436 90188 4756 91700
rect 4436 90132 4464 90188
rect 4520 90132 4568 90188
rect 4624 90132 4672 90188
rect 4728 90132 4756 90188
rect 4436 88620 4756 90132
rect 4844 104468 4900 104478
rect 4844 88900 4900 104412
rect 4844 88834 4900 88844
rect 4956 97748 5012 108444
rect 5180 107380 5236 112700
rect 5292 107828 5348 113372
rect 5404 109620 5460 113820
rect 5740 112644 5796 112654
rect 5404 109554 5460 109564
rect 5516 110964 5572 110974
rect 5292 107762 5348 107772
rect 5180 107314 5236 107324
rect 5068 105252 5124 105262
rect 5068 103796 5124 105196
rect 5068 100324 5124 103740
rect 5404 104020 5460 104030
rect 5404 103684 5460 103964
rect 5404 103618 5460 103628
rect 5404 102228 5460 102238
rect 5404 101556 5460 102172
rect 5404 101490 5460 101500
rect 5068 100258 5124 100268
rect 5404 100324 5460 100334
rect 5180 99988 5236 99998
rect 4436 88564 4464 88620
rect 4520 88564 4568 88620
rect 4624 88564 4672 88620
rect 4728 88564 4756 88620
rect 4436 87052 4756 88564
rect 4436 86996 4464 87052
rect 4520 86996 4568 87052
rect 4624 86996 4672 87052
rect 4728 86996 4756 87052
rect 4436 85484 4756 86996
rect 4436 85428 4464 85484
rect 4520 85428 4568 85484
rect 4624 85428 4672 85484
rect 4728 85428 4756 85484
rect 4436 83916 4756 85428
rect 4436 83860 4464 83916
rect 4520 83860 4568 83916
rect 4624 83860 4672 83916
rect 4728 83860 4756 83916
rect 4436 82348 4756 83860
rect 4436 82292 4464 82348
rect 4520 82292 4568 82348
rect 4624 82292 4672 82348
rect 4728 82292 4756 82348
rect 4436 80780 4756 82292
rect 4956 84644 5012 97692
rect 5068 98308 5124 98318
rect 5068 95956 5124 98252
rect 5068 95890 5124 95900
rect 5180 95508 5236 99932
rect 5180 95442 5236 95452
rect 5292 99204 5348 99214
rect 5068 93380 5124 93390
rect 5068 92148 5124 93324
rect 5068 89124 5124 92092
rect 5068 89058 5124 89068
rect 4436 80724 4464 80780
rect 4520 80724 4568 80780
rect 4624 80724 4672 80780
rect 4728 80724 4756 80780
rect 4436 79212 4756 80724
rect 4436 79156 4464 79212
rect 4520 79156 4568 79212
rect 4624 79156 4672 79212
rect 4728 79156 4756 79212
rect 4436 77644 4756 79156
rect 4436 77588 4464 77644
rect 4520 77588 4568 77644
rect 4624 77588 4672 77644
rect 4728 77588 4756 77644
rect 4436 76076 4756 77588
rect 4436 76020 4464 76076
rect 4520 76020 4568 76076
rect 4624 76020 4672 76076
rect 4728 76020 4756 76076
rect 4172 67330 4228 67340
rect 4436 74508 4756 76020
rect 4436 74452 4464 74508
rect 4520 74452 4568 74508
rect 4624 74452 4672 74508
rect 4728 74452 4756 74508
rect 4436 72940 4756 74452
rect 4436 72884 4464 72940
rect 4520 72884 4568 72940
rect 4624 72884 4672 72940
rect 4728 72884 4756 72940
rect 4436 71372 4756 72884
rect 4844 80948 4900 80958
rect 4844 71988 4900 80892
rect 4844 71922 4900 71932
rect 4956 74788 5012 84588
rect 4436 71316 4464 71372
rect 4520 71316 4568 71372
rect 4624 71316 4672 71372
rect 4728 71316 4756 71372
rect 4436 69804 4756 71316
rect 4436 69748 4464 69804
rect 4520 69748 4568 69804
rect 4624 69748 4672 69804
rect 4728 69748 4756 69804
rect 4436 68236 4756 69748
rect 4436 68180 4464 68236
rect 4520 68180 4568 68236
rect 4624 68180 4672 68236
rect 4728 68180 4756 68236
rect 3776 65828 3804 65884
rect 3860 65828 3908 65884
rect 3964 65828 4012 65884
rect 4068 65828 4096 65884
rect 3276 62402 3332 62412
rect 3776 64316 4096 65828
rect 3776 64260 3804 64316
rect 3860 64260 3908 64316
rect 3964 64260 4012 64316
rect 4068 64260 4096 64316
rect 3776 62748 4096 64260
rect 3776 62692 3804 62748
rect 3860 62692 3908 62748
rect 3964 62692 4012 62748
rect 4068 62692 4096 62748
rect 3776 61180 4096 62692
rect 3776 61124 3804 61180
rect 3860 61124 3908 61180
rect 3964 61124 4012 61180
rect 4068 61124 4096 61180
rect 3776 59612 4096 61124
rect 3776 59556 3804 59612
rect 3860 59556 3908 59612
rect 3964 59556 4012 59612
rect 4068 59556 4096 59612
rect 3776 58044 4096 59556
rect 3776 57988 3804 58044
rect 3860 57988 3908 58044
rect 3964 57988 4012 58044
rect 4068 57988 4096 58044
rect 2604 55010 2660 55020
rect 3164 57764 3220 57774
rect 3164 51418 3220 57708
rect 3776 56476 4096 57988
rect 3776 56420 3804 56476
rect 3860 56420 3908 56476
rect 3964 56420 4012 56476
rect 4068 56420 4096 56476
rect 3776 54908 4096 56420
rect 3776 54852 3804 54908
rect 3860 54852 3908 54908
rect 3964 54852 4012 54908
rect 4068 54852 4096 54908
rect 1372 44522 1540 44578
rect 1708 51380 1764 51390
rect 1372 35252 1428 44522
rect 1372 35186 1428 35196
rect 1484 41860 1540 41870
rect 1260 34066 1316 34076
rect 1372 33684 1428 33694
rect 140 24058 196 24062
rect 140 24052 308 24058
rect 196 24002 308 24052
rect 140 23986 196 23996
rect 252 23940 308 24002
rect 252 23874 308 23884
rect 1260 12292 1316 12302
rect 700 9828 756 9838
rect 700 1652 756 9772
rect 1260 5348 1316 12236
rect 1372 6692 1428 33628
rect 1484 33460 1540 41804
rect 1708 33796 1764 51324
rect 2940 51380 3220 51418
rect 2996 51362 3220 51380
rect 3276 53620 3332 53630
rect 3276 51598 3332 53564
rect 3776 53340 4096 54852
rect 3776 53284 3804 53340
rect 3860 53284 3908 53340
rect 3964 53284 4012 53340
rect 4068 53284 4096 53340
rect 3776 51772 4096 53284
rect 3776 51716 3804 51772
rect 3860 51716 3908 51772
rect 3964 51716 4012 51772
rect 4068 51716 4096 51772
rect 3388 51604 3444 51614
rect 3276 51548 3388 51598
rect 3276 51542 3444 51548
rect 2940 51314 2996 51324
rect 2492 50708 2548 50718
rect 2492 48692 2548 50652
rect 1932 47572 1988 47582
rect 1820 43428 1876 43438
rect 1820 41972 1876 43372
rect 1820 41906 1876 41916
rect 1708 33730 1764 33740
rect 1820 35028 1876 35038
rect 1484 33394 1540 33404
rect 1820 31668 1876 34972
rect 1820 27972 1876 31612
rect 1820 23828 1876 27916
rect 1820 23762 1876 23772
rect 1932 22148 1988 47516
rect 2492 47124 2548 48636
rect 2492 47058 2548 47068
rect 3052 47124 3108 47134
rect 2044 45108 2100 45118
rect 2044 42980 2100 45052
rect 2044 40292 2100 42924
rect 2492 44772 2548 44782
rect 2492 40964 2548 44716
rect 2492 40898 2548 40908
rect 2604 41524 2660 41534
rect 2044 40226 2100 40236
rect 2268 34020 2324 34030
rect 2268 29316 2324 33964
rect 2324 29260 2548 29278
rect 2268 29222 2548 29260
rect 2268 28868 2324 28878
rect 2268 23268 2324 28812
rect 1932 22082 1988 22092
rect 2156 22932 2212 22942
rect 2156 18340 2212 22876
rect 2156 18274 2212 18284
rect 1484 15092 1540 15102
rect 1484 8260 1540 15036
rect 2156 10388 2212 10398
rect 1484 8194 1540 8204
rect 2044 9604 2100 9614
rect 1372 6626 1428 6636
rect 1260 5282 1316 5292
rect 2044 5348 2100 9548
rect 2156 6692 2212 10332
rect 2268 7364 2324 23212
rect 2380 27412 2436 27422
rect 2380 13188 2436 27356
rect 2380 13122 2436 13132
rect 2492 22372 2548 29222
rect 2604 27076 2660 41468
rect 3052 38098 3108 47068
rect 3276 41524 3332 51542
rect 3388 51538 3444 51542
rect 3776 50204 4096 51716
rect 3776 50148 3804 50204
rect 3860 50148 3908 50204
rect 3964 50148 4012 50204
rect 4068 50148 4096 50204
rect 3052 38052 3220 38098
rect 3052 38042 3164 38052
rect 3164 37044 3220 37996
rect 2828 33796 2884 33806
rect 2828 32452 2884 33740
rect 2828 30996 2884 32396
rect 2828 30930 2884 30940
rect 2940 31892 2996 31902
rect 2604 27010 2660 27020
rect 2268 7298 2324 7308
rect 2380 11956 2436 11966
rect 2156 6626 2212 6636
rect 2380 6692 2436 11900
rect 2492 10052 2548 22316
rect 2492 9986 2548 9996
rect 2716 14308 2772 14318
rect 2380 6626 2436 6636
rect 2492 7028 2548 7038
rect 2044 5282 2100 5292
rect 2492 2324 2548 6972
rect 2492 2258 2548 2268
rect 700 1586 756 1596
rect 2716 1204 2772 14252
rect 2940 10836 2996 31836
rect 3052 24052 3108 24062
rect 3052 13412 3108 23996
rect 3164 22932 3220 36988
rect 3276 32676 3332 41468
rect 3500 49140 3556 49150
rect 3500 34132 3556 49084
rect 3776 48636 4096 50148
rect 3776 48580 3804 48636
rect 3860 48580 3908 48636
rect 3964 48580 4012 48636
rect 4068 48580 4096 48636
rect 3776 47068 4096 48580
rect 3776 47012 3804 47068
rect 3860 47012 3908 47068
rect 3964 47012 4012 47068
rect 4068 47012 4096 47068
rect 3776 45500 4096 47012
rect 3776 45444 3804 45500
rect 3860 45444 3908 45500
rect 3964 45444 4012 45500
rect 4068 45444 4096 45500
rect 3776 43932 4096 45444
rect 3776 43876 3804 43932
rect 3860 43876 3908 43932
rect 3964 43876 4012 43932
rect 4068 43876 4096 43932
rect 3776 42364 4096 43876
rect 4436 66668 4756 68180
rect 4956 67956 5012 74732
rect 4956 67890 5012 67900
rect 4436 66612 4464 66668
rect 4520 66612 4568 66668
rect 4624 66612 4672 66668
rect 4728 66612 4756 66668
rect 4436 65100 4756 66612
rect 4436 65044 4464 65100
rect 4520 65044 4568 65100
rect 4624 65044 4672 65100
rect 4728 65044 4756 65100
rect 4436 63532 4756 65044
rect 4436 63476 4464 63532
rect 4520 63476 4568 63532
rect 4624 63476 4672 63532
rect 4728 63476 4756 63532
rect 4436 61964 4756 63476
rect 5180 66276 5236 66286
rect 5180 63252 5236 66220
rect 5180 63186 5236 63196
rect 4436 61908 4464 61964
rect 4520 61908 4568 61964
rect 4624 61908 4672 61964
rect 4728 61908 4756 61964
rect 4436 60396 4756 61908
rect 4436 60340 4464 60396
rect 4520 60340 4568 60396
rect 4624 60340 4672 60396
rect 4728 60340 4756 60396
rect 4436 58828 4756 60340
rect 4436 58772 4464 58828
rect 4520 58772 4568 58828
rect 4624 58772 4672 58828
rect 4728 58772 4756 58828
rect 4436 57260 4756 58772
rect 4436 57204 4464 57260
rect 4520 57204 4568 57260
rect 4624 57204 4672 57260
rect 4728 57204 4756 57260
rect 4436 55692 4756 57204
rect 4436 55636 4464 55692
rect 4520 55636 4568 55692
rect 4624 55636 4672 55692
rect 4728 55636 4756 55692
rect 4436 54124 4756 55636
rect 5292 55412 5348 99148
rect 5404 96964 5460 100268
rect 5404 94500 5460 96908
rect 5404 94434 5460 94444
rect 5516 94388 5572 110908
rect 5628 110292 5684 110302
rect 5628 109844 5684 110236
rect 5628 101638 5684 109788
rect 5740 103012 5796 112588
rect 6300 112532 6356 112542
rect 6188 110516 6244 110526
rect 5740 102946 5796 102956
rect 5852 109284 5908 109294
rect 5628 101582 5796 101638
rect 5516 94322 5572 94332
rect 5740 98308 5796 101582
rect 5740 88564 5796 98252
rect 5852 88788 5908 109228
rect 5964 105924 6020 105934
rect 5964 90804 6020 105868
rect 5964 90738 6020 90748
rect 6076 104244 6132 104254
rect 6076 98756 6132 104188
rect 6188 104132 6244 110460
rect 6300 107940 6356 112476
rect 6300 107874 6356 107884
rect 6412 112308 6468 112318
rect 6188 104066 6244 104076
rect 5852 88722 5908 88732
rect 5740 88498 5796 88508
rect 5628 85876 5684 85886
rect 5404 83748 5460 83758
rect 5404 83188 5460 83692
rect 5628 83748 5684 85820
rect 5628 83682 5684 83692
rect 5404 83122 5460 83132
rect 5628 77924 5684 77934
rect 5628 72996 5684 77868
rect 5628 72930 5684 72940
rect 6076 71876 6132 98700
rect 6188 99092 6244 99102
rect 6188 96740 6244 99036
rect 6188 84756 6244 96684
rect 6300 92596 6356 92606
rect 6300 86996 6356 92540
rect 6300 86930 6356 86940
rect 6188 84308 6244 84700
rect 6188 84242 6244 84252
rect 6300 76132 6356 76142
rect 6300 72660 6356 76076
rect 6300 72594 6356 72604
rect 6076 71810 6132 71820
rect 5292 55346 5348 55356
rect 6076 57316 6132 57326
rect 4436 54068 4464 54124
rect 4520 54068 4568 54124
rect 4624 54068 4672 54124
rect 4728 54068 4756 54124
rect 4436 52556 4756 54068
rect 4436 52500 4464 52556
rect 4520 52500 4568 52556
rect 4624 52500 4672 52556
rect 4728 52500 4756 52556
rect 4436 50988 4756 52500
rect 4436 50932 4464 50988
rect 4520 50932 4568 50988
rect 4624 50932 4672 50988
rect 4728 50932 4756 50988
rect 4436 49420 4756 50932
rect 4436 49364 4464 49420
rect 4520 49364 4568 49420
rect 4624 49364 4672 49420
rect 4728 49364 4756 49420
rect 4436 47852 4756 49364
rect 4844 52052 4900 52062
rect 4844 49364 4900 51996
rect 4844 49140 4900 49308
rect 4844 49074 4900 49084
rect 4436 47796 4464 47852
rect 4520 47796 4568 47852
rect 4624 47796 4672 47852
rect 4728 47796 4756 47852
rect 4436 46284 4756 47796
rect 4436 46228 4464 46284
rect 4520 46228 4568 46284
rect 4624 46228 4672 46284
rect 4728 46228 4756 46284
rect 4436 44716 4756 46228
rect 5404 46116 5460 46126
rect 4436 44660 4464 44716
rect 4520 44660 4568 44716
rect 4624 44660 4672 44716
rect 4728 44660 4756 44716
rect 4284 43764 4340 43774
rect 4284 42644 4340 43708
rect 4284 42578 4340 42588
rect 4436 43148 4756 44660
rect 4436 43092 4464 43148
rect 4520 43092 4568 43148
rect 4624 43092 4672 43148
rect 4728 43092 4756 43148
rect 3776 42308 3804 42364
rect 3860 42308 3908 42364
rect 3964 42308 4012 42364
rect 4068 42308 4096 42364
rect 3776 40796 4096 42308
rect 3776 40740 3804 40796
rect 3860 40740 3908 40796
rect 3964 40740 4012 40796
rect 4068 40740 4096 40796
rect 3776 39228 4096 40740
rect 3776 39172 3804 39228
rect 3860 39172 3908 39228
rect 3964 39172 4012 39228
rect 4068 39172 4096 39228
rect 3776 37660 4096 39172
rect 3776 37604 3804 37660
rect 3860 37604 3908 37660
rect 3964 37604 4012 37660
rect 4068 37604 4096 37660
rect 3776 36092 4096 37604
rect 3776 36036 3804 36092
rect 3860 36036 3908 36092
rect 3964 36036 4012 36092
rect 4068 36036 4096 36092
rect 3500 34066 3556 34076
rect 3612 34804 3668 34814
rect 3612 34580 3668 34748
rect 3276 32610 3332 32620
rect 3612 27860 3668 34524
rect 3612 27794 3668 27804
rect 3776 34524 4096 36036
rect 4436 41580 4756 43092
rect 4436 41524 4464 41580
rect 4520 41524 4568 41580
rect 4624 41524 4672 41580
rect 4728 41524 4756 41580
rect 4436 40012 4756 41524
rect 4436 39956 4464 40012
rect 4520 39956 4568 40012
rect 4624 39956 4672 40012
rect 4728 39956 4756 40012
rect 4956 45892 5012 45902
rect 4956 40068 5012 45836
rect 4956 40002 5012 40012
rect 5180 44996 5236 45006
rect 4436 38444 4756 39956
rect 4436 38388 4464 38444
rect 4520 38388 4568 38444
rect 4624 38388 4672 38444
rect 4728 38388 4756 38444
rect 4436 36876 4756 38388
rect 4436 36820 4464 36876
rect 4520 36820 4568 36876
rect 4624 36820 4672 36876
rect 4728 36820 4756 36876
rect 4436 35308 4756 36820
rect 3776 34468 3804 34524
rect 3860 34468 3908 34524
rect 3964 34468 4012 34524
rect 4068 34468 4096 34524
rect 3776 32956 4096 34468
rect 4172 35252 4228 35262
rect 4172 33796 4228 35196
rect 4436 35252 4464 35308
rect 4520 35252 4568 35308
rect 4624 35252 4672 35308
rect 4728 35252 4756 35308
rect 4172 33730 4228 33740
rect 4284 35028 4340 35038
rect 3776 32900 3804 32956
rect 3860 32900 3908 32956
rect 3964 32900 4012 32956
rect 4068 32900 4096 32956
rect 3776 31388 4096 32900
rect 3776 31332 3804 31388
rect 3860 31332 3908 31388
rect 3964 31332 4012 31388
rect 4068 31332 4096 31388
rect 3776 29820 4096 31332
rect 3776 29764 3804 29820
rect 3860 29764 3908 29820
rect 3964 29764 4012 29820
rect 4068 29764 4096 29820
rect 3776 28252 4096 29764
rect 3776 28196 3804 28252
rect 3860 28196 3908 28252
rect 3964 28196 4012 28252
rect 4068 28196 4096 28252
rect 3776 26684 4096 28196
rect 3776 26628 3804 26684
rect 3860 26628 3908 26684
rect 3964 26628 4012 26684
rect 4068 26628 4096 26684
rect 3612 26516 3668 26526
rect 3500 26068 3556 26078
rect 3500 24612 3556 26012
rect 3612 25956 3668 26460
rect 3612 25890 3668 25900
rect 3500 24546 3556 24556
rect 3776 25116 4096 26628
rect 4172 27076 4228 27086
rect 4172 25508 4228 27020
rect 4172 25442 4228 25452
rect 3776 25060 3804 25116
rect 3860 25060 3908 25116
rect 3964 25060 4012 25116
rect 4068 25060 4096 25116
rect 3164 22866 3220 22876
rect 3776 23548 4096 25060
rect 4172 25060 4228 25070
rect 4172 24276 4228 25004
rect 4172 24210 4228 24220
rect 3776 23492 3804 23548
rect 3860 23492 3908 23548
rect 3964 23492 4012 23548
rect 4068 23492 4096 23548
rect 3776 21980 4096 23492
rect 3776 21924 3804 21980
rect 3860 21924 3908 21980
rect 3964 21924 4012 21980
rect 4068 21924 4096 21980
rect 3612 21700 3668 21710
rect 3276 19572 3332 19582
rect 3276 16996 3332 19516
rect 3276 16930 3332 16940
rect 3388 18564 3444 18574
rect 3052 13346 3108 13356
rect 3164 13972 3220 13982
rect 2940 10770 2996 10780
rect 2940 9156 2996 9166
rect 2828 9044 2884 9054
rect 2828 4676 2884 8988
rect 2828 2212 2884 4620
rect 2828 2146 2884 2156
rect 2940 2100 2996 9100
rect 3164 2660 3220 13916
rect 3276 13524 3332 13534
rect 3276 4116 3332 13468
rect 3388 11620 3444 18508
rect 3612 17668 3668 21644
rect 3612 17602 3668 17612
rect 3776 20412 4096 21924
rect 3776 20356 3804 20412
rect 3860 20356 3908 20412
rect 3964 20356 4012 20412
rect 4068 20356 4096 20412
rect 3776 18844 4096 20356
rect 3776 18788 3804 18844
rect 3860 18788 3908 18844
rect 3964 18788 4012 18844
rect 4068 18788 4096 18844
rect 3776 17276 4096 18788
rect 3776 17220 3804 17276
rect 3860 17220 3908 17276
rect 3964 17220 4012 17276
rect 4068 17220 4096 17276
rect 3776 15708 4096 17220
rect 3776 15652 3804 15708
rect 3860 15652 3908 15708
rect 3964 15652 4012 15708
rect 4068 15652 4096 15708
rect 3612 14196 3668 14206
rect 3388 11554 3444 11564
rect 3500 13412 3556 13422
rect 3388 10948 3444 10958
rect 3388 7498 3444 10892
rect 3500 7858 3556 13356
rect 3612 12292 3668 14140
rect 3612 12226 3668 12236
rect 3776 14140 4096 15652
rect 3776 14084 3804 14140
rect 3860 14084 3908 14140
rect 3964 14084 4012 14140
rect 4068 14084 4096 14140
rect 3776 12572 4096 14084
rect 3776 12516 3804 12572
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 4068 12516 4096 12572
rect 3776 11004 4096 12516
rect 3776 10948 3804 11004
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 4068 10948 4096 11004
rect 3776 9436 4096 10948
rect 3776 9380 3804 9436
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 4068 9380 4096 9436
rect 3612 8820 3668 8830
rect 3612 8148 3668 8764
rect 3612 8082 3668 8092
rect 3776 7868 4096 9380
rect 3500 7802 3668 7858
rect 3388 7442 3556 7498
rect 3388 7364 3444 7374
rect 3388 6692 3444 7308
rect 3388 6626 3444 6636
rect 3500 5908 3556 7442
rect 3500 5842 3556 5852
rect 3276 4050 3332 4060
rect 3612 2772 3668 7802
rect 3612 2706 3668 2716
rect 3776 7812 3804 7868
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 4068 7812 4096 7868
rect 3776 6300 4096 7812
rect 3776 6244 3804 6300
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 4068 6244 4096 6300
rect 3776 4732 4096 6244
rect 4172 23604 4228 23614
rect 4172 17780 4228 23548
rect 4172 5796 4228 17724
rect 4284 16100 4340 34972
rect 4284 16034 4340 16044
rect 4436 33740 4756 35252
rect 4436 33684 4464 33740
rect 4520 33684 4568 33740
rect 4624 33684 4672 33740
rect 4728 33684 4756 33740
rect 4436 32172 4756 33684
rect 4436 32116 4464 32172
rect 4520 32116 4568 32172
rect 4624 32116 4672 32172
rect 4728 32116 4756 32172
rect 4436 30604 4756 32116
rect 4436 30548 4464 30604
rect 4520 30548 4568 30604
rect 4624 30548 4672 30604
rect 4728 30548 4756 30604
rect 4436 29036 4756 30548
rect 4436 28980 4464 29036
rect 4520 28980 4568 29036
rect 4624 28980 4672 29036
rect 4728 28980 4756 29036
rect 4436 27468 4756 28980
rect 4436 27412 4464 27468
rect 4520 27412 4568 27468
rect 4624 27412 4672 27468
rect 4728 27412 4756 27468
rect 4436 25900 4756 27412
rect 4844 39396 4900 39406
rect 4844 26516 4900 39340
rect 5068 39060 5124 39070
rect 5068 32452 5124 39004
rect 5068 32386 5124 32396
rect 4844 26450 4900 26460
rect 4956 31780 5012 31790
rect 4956 31108 5012 31724
rect 4436 25844 4464 25900
rect 4520 25844 4568 25900
rect 4624 25844 4672 25900
rect 4728 25844 4756 25900
rect 4436 24332 4756 25844
rect 4436 24276 4464 24332
rect 4520 24276 4568 24332
rect 4624 24276 4672 24332
rect 4728 24276 4756 24332
rect 4436 22764 4756 24276
rect 4436 22708 4464 22764
rect 4520 22708 4568 22764
rect 4624 22708 4672 22764
rect 4728 22708 4756 22764
rect 4436 21196 4756 22708
rect 4844 23044 4900 23054
rect 4844 22708 4900 22988
rect 4844 22642 4900 22652
rect 4436 21140 4464 21196
rect 4520 21140 4568 21196
rect 4624 21140 4672 21196
rect 4728 21140 4756 21196
rect 4436 19628 4756 21140
rect 4436 19572 4464 19628
rect 4520 19572 4568 19628
rect 4624 19572 4672 19628
rect 4728 19572 4756 19628
rect 4436 18060 4756 19572
rect 4844 20580 4900 20590
rect 4844 19684 4900 20524
rect 4844 19460 4900 19628
rect 4844 18298 4900 19404
rect 4956 18564 5012 31052
rect 4956 18498 5012 18508
rect 5068 20580 5124 20590
rect 4844 18242 5012 18298
rect 4436 18004 4464 18060
rect 4520 18004 4568 18060
rect 4624 18004 4672 18060
rect 4728 18004 4756 18060
rect 4436 16492 4756 18004
rect 4436 16436 4464 16492
rect 4520 16436 4568 16492
rect 4624 16436 4672 16492
rect 4728 16436 4756 16492
rect 4436 14924 4756 16436
rect 4436 14868 4464 14924
rect 4520 14868 4568 14924
rect 4624 14868 4672 14924
rect 4728 14868 4756 14924
rect 4436 13356 4756 14868
rect 4956 14644 5012 18242
rect 5068 15540 5124 20524
rect 5068 15474 5124 15484
rect 4956 14196 5012 14588
rect 4436 13300 4464 13356
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4728 13300 4756 13356
rect 4436 11788 4756 13300
rect 4436 11732 4464 11788
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4728 11732 4756 11788
rect 4284 10500 4340 10510
rect 4284 10276 4340 10444
rect 4284 10210 4340 10220
rect 4436 10220 4756 11732
rect 4436 10164 4464 10220
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4728 10164 4756 10220
rect 4284 9044 4340 9054
rect 4284 6804 4340 8988
rect 4284 6738 4340 6748
rect 4436 8652 4756 10164
rect 4436 8596 4464 8652
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4728 8596 4756 8652
rect 4436 7084 4756 8596
rect 4436 7028 4464 7084
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4728 7028 4756 7084
rect 4172 5730 4228 5740
rect 3776 4676 3804 4732
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 4068 4676 4096 4732
rect 3776 3164 4096 4676
rect 3776 3108 3804 3164
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 4068 3108 4096 3164
rect 3164 2594 3220 2604
rect 2940 2034 2996 2044
rect 2716 1138 2772 1148
rect 3776 1596 4096 3108
rect 3776 1540 3804 1596
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 4068 1540 4096 1596
rect 3776 0 4096 1540
rect 4436 5516 4756 7028
rect 4436 5460 4464 5516
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4728 5460 4756 5516
rect 4436 3948 4756 5460
rect 4436 3892 4464 3948
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4728 3892 4756 3948
rect 4436 2380 4756 3892
rect 4844 13636 4900 13646
rect 4844 2996 4900 13580
rect 4956 12628 5012 14140
rect 5180 13076 5236 44940
rect 5404 31108 5460 46060
rect 5964 46004 6020 46014
rect 5404 31042 5460 31052
rect 5628 42980 5684 42990
rect 5628 38276 5684 42924
rect 5852 42644 5908 42654
rect 5404 25620 5460 25630
rect 5180 13010 5236 13020
rect 5292 25284 5348 25294
rect 4956 12562 5012 12572
rect 5068 12852 5124 12862
rect 4844 2930 4900 2940
rect 4956 10948 5012 10958
rect 4956 2884 5012 10892
rect 5068 5908 5124 12796
rect 5292 9044 5348 25228
rect 5404 23044 5460 25564
rect 5404 22978 5460 22988
rect 5628 22932 5684 38220
rect 5740 40068 5796 40078
rect 5740 23940 5796 40012
rect 5852 37604 5908 42588
rect 5852 37538 5908 37548
rect 5964 38388 6020 45948
rect 6076 40292 6132 57260
rect 6076 40226 6132 40236
rect 6188 43316 6244 43326
rect 6188 40404 6244 43260
rect 6412 41972 6468 112252
rect 6636 112196 6692 114604
rect 19964 113988 20020 113998
rect 11900 113876 11956 113886
rect 8764 113428 8820 113438
rect 7308 113316 7364 113326
rect 6636 112130 6692 112140
rect 6860 112532 6916 112542
rect 6748 110852 6804 110862
rect 6748 104244 6804 110796
rect 6860 108118 6916 112476
rect 7084 111748 7140 111758
rect 7084 111188 7140 111692
rect 6860 108062 7028 108118
rect 6748 104178 6804 104188
rect 6972 105476 7028 108062
rect 6860 98308 6916 98318
rect 6524 91924 6580 91934
rect 6524 91140 6580 91868
rect 6524 91074 6580 91084
rect 6636 88564 6692 88574
rect 6636 77476 6692 88508
rect 6748 82180 6804 82190
rect 6748 80276 6804 82124
rect 6748 80210 6804 80220
rect 6860 79492 6916 98252
rect 6972 95172 7028 105420
rect 6972 94612 7028 95116
rect 6972 94546 7028 94556
rect 7084 93268 7140 111132
rect 7196 106148 7252 106158
rect 7196 100436 7252 106092
rect 7308 100772 7364 113260
rect 7532 113316 7588 113326
rect 7532 112756 7588 113260
rect 7532 112690 7588 112700
rect 7980 112308 8036 112318
rect 7980 109732 8036 112252
rect 7980 109508 8036 109676
rect 7980 109442 8036 109452
rect 8092 109396 8148 109406
rect 8092 108724 8148 109340
rect 7980 105140 8036 105150
rect 7308 100706 7364 100716
rect 7420 104244 7476 104254
rect 7196 99540 7252 100380
rect 7196 99474 7252 99484
rect 7084 91476 7140 93212
rect 7420 91588 7476 104188
rect 7644 102116 7700 102126
rect 7420 91522 7476 91532
rect 7532 96068 7588 96078
rect 7084 91410 7140 91420
rect 6860 79156 6916 79436
rect 6860 79090 6916 79100
rect 6972 89012 7028 89022
rect 6636 67060 6692 77420
rect 6636 66994 6692 67004
rect 6972 53732 7028 88956
rect 7532 79604 7588 96012
rect 7644 89908 7700 102060
rect 7980 98308 8036 105084
rect 8092 104468 8148 108668
rect 8540 108724 8596 108734
rect 8092 104402 8148 104412
rect 8316 106932 8372 106942
rect 7980 98242 8036 98252
rect 8092 104020 8148 104030
rect 8092 102788 8148 103964
rect 7756 97636 7812 97646
rect 7756 97412 7812 97580
rect 7756 97346 7812 97356
rect 7980 91476 8036 91486
rect 7644 89842 7700 89852
rect 7868 89908 7924 89918
rect 7868 89758 7924 89852
rect 7084 75908 7140 75918
rect 7084 68964 7140 75852
rect 7532 73780 7588 79548
rect 7532 73714 7588 73724
rect 7756 89702 7924 89758
rect 7756 81060 7812 89702
rect 7084 68898 7140 68908
rect 7756 68852 7812 81004
rect 7756 68516 7812 68796
rect 7756 68450 7812 68460
rect 7868 89572 7924 89582
rect 7756 60676 7812 60686
rect 6972 53666 7028 53676
rect 7420 56644 7476 56654
rect 6412 41906 6468 41916
rect 6524 52948 6580 52958
rect 6188 38500 6244 40348
rect 6188 38434 6244 38444
rect 5964 37044 6020 38332
rect 5964 36978 6020 36988
rect 6412 34132 6468 34142
rect 6412 33236 6468 34076
rect 6412 32788 6468 33180
rect 6412 32722 6468 32732
rect 5740 23874 5796 23884
rect 5852 29316 5908 29326
rect 5852 25732 5908 29260
rect 5628 22866 5684 22876
rect 5740 22708 5796 22718
rect 5404 20020 5460 20030
rect 5404 15652 5460 19964
rect 5628 18228 5684 18238
rect 5628 16660 5684 18172
rect 5628 16594 5684 16604
rect 5740 16436 5796 22652
rect 5852 17332 5908 25676
rect 6188 23940 6244 23950
rect 6188 21028 6244 23884
rect 5852 17266 5908 17276
rect 6076 18788 6132 18798
rect 5740 16370 5796 16380
rect 5404 15586 5460 15596
rect 5628 15764 5684 15774
rect 5628 14980 5684 15708
rect 5628 14914 5684 14924
rect 5740 11844 5796 11854
rect 5292 8978 5348 8988
rect 5404 11732 5460 11742
rect 5068 5842 5124 5852
rect 5404 4564 5460 11676
rect 5628 9380 5684 9390
rect 5628 6916 5684 9324
rect 5628 6850 5684 6860
rect 5404 4498 5460 4508
rect 4956 2818 5012 2828
rect 5740 2660 5796 11788
rect 5852 11172 5908 11182
rect 5852 3332 5908 11116
rect 5852 3266 5908 3276
rect 5964 10500 6020 10510
rect 5740 2594 5796 2604
rect 4436 2324 4464 2380
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4728 2324 4756 2380
rect 4436 812 4756 2324
rect 5964 1428 6020 10444
rect 6076 1652 6132 18732
rect 6188 9492 6244 20972
rect 6300 16884 6356 16894
rect 6300 14532 6356 16828
rect 6300 14466 6356 14476
rect 6188 9426 6244 9436
rect 6300 13524 6356 13534
rect 6300 3444 6356 13468
rect 6412 6580 6468 6590
rect 6412 5236 6468 6524
rect 6412 5170 6468 5180
rect 6300 3378 6356 3388
rect 6076 1586 6132 1596
rect 6524 1652 6580 52892
rect 6860 50596 6916 50606
rect 6860 45108 6916 50540
rect 7420 49588 7476 56588
rect 6860 45042 6916 45052
rect 7084 47348 7140 47358
rect 7084 46788 7140 47292
rect 7084 46004 7140 46732
rect 6748 44100 6804 44110
rect 6636 40292 6692 40302
rect 6636 38724 6692 40236
rect 6636 13636 6692 38668
rect 6748 32004 6804 44044
rect 6748 31668 6804 31948
rect 6748 31602 6804 31612
rect 6972 32340 7028 32350
rect 6748 30996 6804 31006
rect 6748 25956 6804 30940
rect 6748 25890 6804 25900
rect 6860 26964 6916 26974
rect 6636 13570 6692 13580
rect 6748 19348 6804 19358
rect 6524 1586 6580 1596
rect 6748 1652 6804 19292
rect 6860 9044 6916 26908
rect 6972 26292 7028 32284
rect 6972 26226 7028 26236
rect 7084 27748 7140 45948
rect 7084 21924 7140 27692
rect 7420 24388 7476 49532
rect 7532 37380 7588 37390
rect 7532 36036 7588 37324
rect 7532 34468 7588 35980
rect 7532 34402 7588 34412
rect 7420 23604 7476 24332
rect 7420 23538 7476 23548
rect 7644 29316 7700 29326
rect 6860 8978 6916 8988
rect 6972 20916 7028 20926
rect 6748 1586 6804 1596
rect 6972 1652 7028 20860
rect 7084 17780 7140 21868
rect 7420 20132 7476 20142
rect 7084 17714 7140 17724
rect 7196 20020 7252 20030
rect 7196 17108 7252 19964
rect 7196 17042 7252 17052
rect 7084 9156 7140 9166
rect 7084 1764 7140 9100
rect 7084 1698 7140 1708
rect 6972 1586 7028 1596
rect 7420 1652 7476 20076
rect 7532 8372 7588 8382
rect 7532 5460 7588 8316
rect 7532 5394 7588 5404
rect 7420 1586 7476 1596
rect 7644 1652 7700 29260
rect 7644 1586 7700 1596
rect 7756 2772 7812 60620
rect 7868 53060 7924 89516
rect 7980 75908 8036 91420
rect 8092 82738 8148 102732
rect 8204 89348 8260 89358
rect 8204 84980 8260 89292
rect 8204 83972 8260 84924
rect 8204 83906 8260 83916
rect 8092 82682 8260 82738
rect 8092 82516 8148 82526
rect 8092 77252 8148 82460
rect 8204 80836 8260 82682
rect 8204 80770 8260 80780
rect 8092 77186 8148 77196
rect 7980 75842 8036 75852
rect 8204 68404 8260 68414
rect 8204 65492 8260 68348
rect 8204 65426 8260 65436
rect 7868 52994 7924 53004
rect 7980 63812 8036 63822
rect 7980 63140 8036 63756
rect 7756 1540 7812 2716
rect 7868 47236 7924 47246
rect 7868 1652 7924 47180
rect 7980 30324 8036 63084
rect 8316 55300 8372 106876
rect 8428 94388 8484 94398
rect 8428 87444 8484 94332
rect 8428 87378 8484 87388
rect 8428 82068 8484 82078
rect 8428 75236 8484 82012
rect 8428 75170 8484 75180
rect 8316 55234 8372 55244
rect 8316 52948 8372 52958
rect 8316 52164 8372 52892
rect 8204 50596 8260 50606
rect 8204 45108 8260 50540
rect 7980 30258 8036 30268
rect 8092 44548 8148 44558
rect 8092 44100 8148 44492
rect 7980 23604 8036 23614
rect 7980 22036 8036 23548
rect 7980 20468 8036 21980
rect 7980 20402 8036 20412
rect 8092 12964 8148 44044
rect 8204 33012 8260 45052
rect 8204 32946 8260 32956
rect 8204 31668 8260 31678
rect 8204 29092 8260 31612
rect 8204 16772 8260 29036
rect 8204 16706 8260 16716
rect 7980 7252 8036 7262
rect 7980 4116 8036 7196
rect 8092 6580 8148 12908
rect 8092 6514 8148 6524
rect 7980 4050 8036 4060
rect 7868 1586 7924 1596
rect 8316 1652 8372 52108
rect 8540 34692 8596 108668
rect 8764 107604 8820 113372
rect 9884 113428 9940 113438
rect 9324 113092 9380 113102
rect 8988 111412 9044 111422
rect 8764 107538 8820 107548
rect 8876 108612 8932 108622
rect 8764 106932 8820 106942
rect 8652 95732 8708 95742
rect 8652 94724 8708 95676
rect 8652 94658 8708 94668
rect 8764 89012 8820 106876
rect 8764 88946 8820 88956
rect 8876 70644 8932 108556
rect 8988 107578 9044 111356
rect 9324 107828 9380 113036
rect 9324 107762 9380 107772
rect 9548 109172 9604 109182
rect 9548 108612 9604 109116
rect 8988 107522 9268 107578
rect 9212 105700 9268 107522
rect 9212 105634 9268 105644
rect 9548 106932 9604 108556
rect 9884 107940 9940 113372
rect 10668 113092 10724 113102
rect 10668 112532 10724 113036
rect 10668 112466 10724 112476
rect 11676 112980 11732 112990
rect 11228 112420 11284 112430
rect 10556 111748 10612 111758
rect 10332 110180 10388 110190
rect 9884 107874 9940 107884
rect 9996 109396 10052 109406
rect 9324 104468 9380 104478
rect 9324 103124 9380 104412
rect 8988 94724 9044 94734
rect 8988 83636 9044 94668
rect 8988 83570 9044 83580
rect 9100 81508 9156 81518
rect 9100 79940 9156 81452
rect 9100 79874 9156 79884
rect 8876 70578 8932 70588
rect 9100 79380 9156 79390
rect 9100 66052 9156 79324
rect 9100 65986 9156 65996
rect 9212 77028 9268 77038
rect 9212 52948 9268 76972
rect 9324 68516 9380 103068
rect 9324 68450 9380 68460
rect 9212 52882 9268 52892
rect 9436 67508 9492 67518
rect 8988 45780 9044 45790
rect 8540 34626 8596 34636
rect 8876 40516 8932 40526
rect 8764 31332 8820 31342
rect 8540 25284 8596 25294
rect 8428 8596 8484 8606
rect 8428 4900 8484 8540
rect 8428 4834 8484 4844
rect 8316 1586 8372 1596
rect 8540 1652 8596 25228
rect 8652 8036 8708 8046
rect 8652 5124 8708 7980
rect 8652 5058 8708 5068
rect 8540 1586 8596 1596
rect 8764 1652 8820 31276
rect 8876 4340 8932 40460
rect 8988 18452 9044 45724
rect 9324 45332 9380 45342
rect 9212 33908 9268 33918
rect 9100 28196 9156 28206
rect 9100 27188 9156 28140
rect 9100 27122 9156 27132
rect 9212 26758 9268 33852
rect 9100 26702 9268 26758
rect 9100 19348 9156 26702
rect 9100 19282 9156 19292
rect 8988 18386 9044 18396
rect 8876 4274 8932 4284
rect 9212 6804 9268 6814
rect 9212 3556 9268 6748
rect 9212 3490 9268 3500
rect 8764 1586 8820 1596
rect 9324 1652 9380 45276
rect 9436 20132 9492 67452
rect 9548 55412 9604 106876
rect 9548 55346 9604 55356
rect 9660 104468 9716 104478
rect 9548 54404 9604 54414
rect 9548 29316 9604 54348
rect 9660 43652 9716 104412
rect 9884 96852 9940 96862
rect 9884 90132 9940 96796
rect 9884 88340 9940 90076
rect 9884 88274 9940 88284
rect 9884 84644 9940 84654
rect 9884 81172 9940 84588
rect 9884 62692 9940 81116
rect 9884 62626 9940 62636
rect 9884 45668 9940 45678
rect 9884 45444 9940 45612
rect 9884 45378 9940 45388
rect 9660 43586 9716 43596
rect 9884 44324 9940 44334
rect 9548 29250 9604 29260
rect 9548 26740 9604 26750
rect 9548 25396 9604 26684
rect 9548 25330 9604 25340
rect 9436 20066 9492 20076
rect 9548 19908 9604 19918
rect 9436 8596 9492 8606
rect 9436 7476 9492 8540
rect 9436 7410 9492 7420
rect 9548 6692 9604 19852
rect 9772 18676 9828 18686
rect 9548 6626 9604 6636
rect 9660 10724 9716 10734
rect 9660 4004 9716 10668
rect 9660 3938 9716 3948
rect 9772 3780 9828 18620
rect 9772 3714 9828 3724
rect 9324 1586 9380 1596
rect 7756 1474 7812 1484
rect 9212 1540 9268 1550
rect 5964 1362 6020 1372
rect 9212 980 9268 1484
rect 9212 914 9268 924
rect 9884 980 9940 44268
rect 9996 41860 10052 109340
rect 10220 109172 10276 109182
rect 10108 99764 10164 99774
rect 10108 56980 10164 99708
rect 10220 67508 10276 109116
rect 10332 98868 10388 110124
rect 10444 109060 10500 109070
rect 10444 108276 10500 109004
rect 10444 108210 10500 108220
rect 10332 98802 10388 98812
rect 10444 103572 10500 103582
rect 10444 102900 10500 103516
rect 10444 95396 10500 102844
rect 10444 95330 10500 95340
rect 10556 87780 10612 111692
rect 11228 111636 11284 112364
rect 11116 110964 11172 110974
rect 10556 87714 10612 87724
rect 10668 107828 10724 107838
rect 10332 80052 10388 80062
rect 10332 79604 10388 79996
rect 10332 77924 10388 79548
rect 10556 79940 10612 79950
rect 10556 79380 10612 79884
rect 10556 79314 10612 79324
rect 10332 77858 10388 77868
rect 10668 77028 10724 107772
rect 10668 76962 10724 76972
rect 10780 106932 10836 106942
rect 10220 67442 10276 67452
rect 10108 56914 10164 56924
rect 10668 50036 10724 50046
rect 9996 41794 10052 41804
rect 10108 46564 10164 46574
rect 10108 45668 10164 46508
rect 9996 25956 10052 25966
rect 9996 25732 10052 25900
rect 9996 25666 10052 25676
rect 10108 1652 10164 45612
rect 10556 46004 10612 46014
rect 10220 45108 10276 45118
rect 10220 35476 10276 45052
rect 10556 38500 10612 45948
rect 10556 38434 10612 38444
rect 10668 36596 10724 49980
rect 10668 36530 10724 36540
rect 10220 31892 10276 35420
rect 10668 34356 10724 34366
rect 10220 31826 10276 31836
rect 10332 33012 10388 33022
rect 10220 3332 10276 3342
rect 10220 2436 10276 3276
rect 10220 1876 10276 2380
rect 10220 1810 10276 1820
rect 10108 1586 10164 1596
rect 10332 1652 10388 32956
rect 10556 29764 10612 29774
rect 10556 23338 10612 29708
rect 10668 24612 10724 34300
rect 10668 24546 10724 24556
rect 10556 23282 10724 23338
rect 10668 14420 10724 23282
rect 10780 20244 10836 106876
rect 11116 97636 11172 110908
rect 11228 105924 11284 111580
rect 11452 111636 11508 111646
rect 11452 111188 11508 111580
rect 11452 111122 11508 111132
rect 11676 110740 11732 112924
rect 11900 112420 11956 113820
rect 15036 113540 15092 113550
rect 13692 113428 13748 113438
rect 11900 112354 11956 112364
rect 12684 112756 12740 112766
rect 12684 112196 12740 112700
rect 12684 112130 12740 112140
rect 13468 111412 13524 111422
rect 11676 110674 11732 110684
rect 12796 110964 12852 110974
rect 11340 110628 11396 110638
rect 11340 107828 11396 110572
rect 11340 107762 11396 107772
rect 11564 108388 11620 108398
rect 11228 105858 11284 105868
rect 11340 107604 11396 107614
rect 11116 97570 11172 97580
rect 10892 94052 10948 94062
rect 10892 84644 10948 93996
rect 11004 92932 11060 92942
rect 11004 86772 11060 92876
rect 11004 86706 11060 86716
rect 11228 90356 11284 90366
rect 11228 88340 11284 90300
rect 11228 84980 11284 88284
rect 11228 84914 11284 84924
rect 10892 84578 10948 84588
rect 11004 84420 11060 84430
rect 10892 77812 10948 77822
rect 10892 71652 10948 77756
rect 10892 71586 10948 71596
rect 11004 50036 11060 84364
rect 11228 79380 11284 79390
rect 11228 72548 11284 79324
rect 11228 72482 11284 72492
rect 11004 49970 11060 49980
rect 11228 68516 11284 68526
rect 11004 49812 11060 49822
rect 11004 46004 11060 49756
rect 11004 45938 11060 45948
rect 10780 20178 10836 20188
rect 10892 43652 10948 43662
rect 10668 14354 10724 14364
rect 10332 1586 10388 1596
rect 10556 13524 10612 13534
rect 10556 1540 10612 13468
rect 10668 9492 10724 9502
rect 10668 5460 10724 9436
rect 10668 5394 10724 5404
rect 10556 1474 10612 1484
rect 10892 1540 10948 43596
rect 11004 41972 11060 41982
rect 11004 3556 11060 41916
rect 11116 40964 11172 40974
rect 11116 36820 11172 40908
rect 11116 36754 11172 36764
rect 11116 36596 11172 36606
rect 11116 29764 11172 36540
rect 11116 29698 11172 29708
rect 11116 29316 11172 29326
rect 11116 16660 11172 29260
rect 11116 16594 11172 16604
rect 11004 3490 11060 3500
rect 11116 14420 11172 14430
rect 10892 1474 10948 1484
rect 9884 914 9940 924
rect 11116 980 11172 14364
rect 11228 1652 11284 68460
rect 11340 44548 11396 107548
rect 11452 104468 11508 104478
rect 11452 77252 11508 104412
rect 11452 77186 11508 77196
rect 11340 44482 11396 44492
rect 11452 44436 11508 44446
rect 11340 31892 11396 31902
rect 11340 4340 11396 31836
rect 11340 4274 11396 4284
rect 11228 1586 11284 1596
rect 11452 1652 11508 44380
rect 11564 41412 11620 108332
rect 11676 104468 11732 104478
rect 11676 104020 11732 104412
rect 11676 103954 11732 103964
rect 11900 104132 11956 104142
rect 11788 95844 11844 95854
rect 11676 90244 11732 90254
rect 11676 83188 11732 90188
rect 11788 87444 11844 95788
rect 11900 94612 11956 104076
rect 11900 94546 11956 94556
rect 12572 98532 12628 98542
rect 11788 87378 11844 87388
rect 11676 83122 11732 83132
rect 11676 79044 11732 79054
rect 11676 73220 11732 78988
rect 11676 73154 11732 73164
rect 12124 77252 12180 77262
rect 11900 55300 11956 55310
rect 11788 46452 11844 46462
rect 11564 41346 11620 41356
rect 11676 45108 11732 45118
rect 11564 40404 11620 40414
rect 11564 39508 11620 40348
rect 11564 39442 11620 39452
rect 11564 39060 11620 39070
rect 11564 38836 11620 39004
rect 11564 38770 11620 38780
rect 11564 4676 11620 4686
rect 11564 2660 11620 4620
rect 11564 2594 11620 2604
rect 11452 1586 11508 1596
rect 11116 914 11172 924
rect 11340 1316 11396 1326
rect 11340 980 11396 1260
rect 11340 914 11396 924
rect 4436 756 4464 812
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4728 756 4756 812
rect 4436 0 4756 756
rect 11676 644 11732 45052
rect 11788 38276 11844 46396
rect 11788 38210 11844 38220
rect 11788 34132 11844 34142
rect 11788 24500 11844 34076
rect 11788 24434 11844 24444
rect 11788 10500 11844 10510
rect 11788 7364 11844 10444
rect 11788 7298 11844 7308
rect 11900 1652 11956 55244
rect 12012 46564 12068 46574
rect 12012 45444 12068 46508
rect 12012 45378 12068 45388
rect 12012 31556 12068 31566
rect 12012 25172 12068 31500
rect 12012 25106 12068 25116
rect 12012 21028 12068 21038
rect 12012 20244 12068 20972
rect 12012 20178 12068 20188
rect 11900 1586 11956 1596
rect 12124 1652 12180 77196
rect 12572 64036 12628 98476
rect 12684 76580 12740 76590
rect 12684 73444 12740 76524
rect 12684 73378 12740 73388
rect 12572 62916 12628 63980
rect 12572 62850 12628 62860
rect 12348 55412 12404 55422
rect 12236 50708 12292 50718
rect 12236 4340 12292 50652
rect 12236 4274 12292 4284
rect 12124 1586 12180 1596
rect 12348 1652 12404 55356
rect 12572 41860 12628 41870
rect 12460 15876 12516 15886
rect 12460 15428 12516 15820
rect 12460 15362 12516 15372
rect 12348 1586 12404 1596
rect 12572 1652 12628 41804
rect 12684 23492 12740 23502
rect 12684 14196 12740 23436
rect 12684 14130 12740 14140
rect 12572 1586 12628 1596
rect 12796 1652 12852 110908
rect 12908 110068 12964 110078
rect 12908 74452 12964 110012
rect 13468 108948 13524 111356
rect 13468 108882 13524 108892
rect 13580 109508 13636 109518
rect 13468 107828 13524 107838
rect 13244 105924 13300 105934
rect 12908 74386 12964 74396
rect 13020 98868 13076 98878
rect 12908 62916 12964 62926
rect 12908 18340 12964 62860
rect 12908 18274 12964 18284
rect 12796 1586 12852 1596
rect 13020 1652 13076 98812
rect 13132 81396 13188 81406
rect 13132 55412 13188 81340
rect 13132 55346 13188 55356
rect 13132 27300 13188 27310
rect 13132 21700 13188 27244
rect 13132 21634 13188 21644
rect 13132 18564 13188 18574
rect 13132 14532 13188 18508
rect 13132 14466 13188 14476
rect 13020 1586 13076 1596
rect 13244 1652 13300 105868
rect 13468 104132 13524 107772
rect 13580 105252 13636 109452
rect 13580 105186 13636 105196
rect 13468 104066 13524 104076
rect 13580 103572 13636 103582
rect 13468 101444 13524 101454
rect 13468 86660 13524 101388
rect 13580 94164 13636 103516
rect 13692 97972 13748 113372
rect 14140 113428 14196 113438
rect 13916 110516 13972 110526
rect 13916 107828 13972 110460
rect 14028 110068 14084 110078
rect 14028 107940 14084 110012
rect 14028 107874 14084 107884
rect 13916 107762 13972 107772
rect 14028 107604 14084 107614
rect 13692 97906 13748 97916
rect 13804 107548 14028 107578
rect 13804 107522 14084 107548
rect 13580 94098 13636 94108
rect 13468 86324 13524 86604
rect 13468 86258 13524 86268
rect 13356 85316 13412 85326
rect 13356 84980 13412 85260
rect 13356 84914 13412 84924
rect 13692 84196 13748 84206
rect 13468 31892 13524 31902
rect 13468 30436 13524 31836
rect 13356 16996 13412 17006
rect 13356 4340 13412 16940
rect 13356 4274 13412 4284
rect 13468 3108 13524 30380
rect 13580 23380 13636 23390
rect 13580 21588 13636 23324
rect 13580 21522 13636 21532
rect 13580 19572 13636 19582
rect 13580 9156 13636 19516
rect 13580 9090 13636 9100
rect 13692 3556 13748 84140
rect 13804 34916 13860 107522
rect 14140 100018 14196 113372
rect 14588 113428 14644 113438
rect 14364 112644 14420 112654
rect 14028 99962 14196 100018
rect 14252 110180 14308 110190
rect 13916 99540 13972 99550
rect 13916 94388 13972 99484
rect 14028 95732 14084 99962
rect 14140 96964 14196 96974
rect 14140 96740 14196 96908
rect 14140 96674 14196 96684
rect 14028 95666 14084 95676
rect 13916 94322 13972 94332
rect 14140 85764 14196 85774
rect 14140 85540 14196 85708
rect 14140 85474 14196 85484
rect 14252 42980 14308 110124
rect 14364 98532 14420 112588
rect 14476 111636 14532 111646
rect 14476 106820 14532 111580
rect 14588 110628 14644 113372
rect 14812 112644 14868 112654
rect 14588 110562 14644 110572
rect 14700 112308 14756 112318
rect 14476 106754 14532 106764
rect 14588 107828 14644 107838
rect 14588 106932 14644 107772
rect 14700 107492 14756 112252
rect 14812 107604 14868 112588
rect 14812 107538 14868 107548
rect 14924 110180 14980 110190
rect 14924 109620 14980 110124
rect 14700 107426 14756 107436
rect 14364 98466 14420 98476
rect 14364 98084 14420 98094
rect 14364 97748 14420 98028
rect 14364 97678 14420 97692
rect 14364 97622 14532 97678
rect 14364 97188 14420 97198
rect 14364 95956 14420 97132
rect 14364 95890 14420 95900
rect 14364 87332 14420 87342
rect 14364 84868 14420 87276
rect 14364 83412 14420 84812
rect 14364 83346 14420 83356
rect 14364 81508 14420 81518
rect 14364 74788 14420 81452
rect 14364 74722 14420 74732
rect 14476 56196 14532 97622
rect 14476 56130 14532 56140
rect 14476 55412 14532 55422
rect 14252 42914 14308 42924
rect 14364 43316 14420 43326
rect 14252 39732 14308 39742
rect 14252 38836 14308 39676
rect 14252 38770 14308 38780
rect 13804 34468 13860 34860
rect 13804 34402 13860 34412
rect 14140 35140 14196 35150
rect 14140 33908 14196 35084
rect 14140 33842 14196 33852
rect 14364 28198 14420 43260
rect 14476 32788 14532 55356
rect 14588 36658 14644 106876
rect 14700 104132 14756 104142
rect 14700 38724 14756 104076
rect 14812 98084 14868 98094
rect 14812 95172 14868 98028
rect 14812 95106 14868 95116
rect 14812 85876 14868 85886
rect 14812 81172 14868 85820
rect 14812 81106 14868 81116
rect 14924 54516 14980 109564
rect 15036 107604 15092 113484
rect 19516 113540 19572 113550
rect 15036 107538 15092 107548
rect 15148 112644 15204 112654
rect 15148 85092 15204 112588
rect 16044 112644 16100 112654
rect 15260 112084 15316 112094
rect 15260 108948 15316 112028
rect 15260 108882 15316 108892
rect 15820 110628 15876 110638
rect 15820 109508 15876 110572
rect 15148 85026 15204 85036
rect 15260 108500 15316 108510
rect 15148 81284 15204 81294
rect 15036 81060 15092 81070
rect 15036 80724 15092 81004
rect 15036 80658 15092 80668
rect 15148 78036 15204 81228
rect 15148 77970 15204 77980
rect 14924 54450 14980 54460
rect 15148 52724 15204 52734
rect 14700 38658 14756 38668
rect 14924 48020 14980 48030
rect 14924 39284 14980 47964
rect 14812 37044 14868 37054
rect 14588 36602 14756 36658
rect 14476 32722 14532 32732
rect 14588 36372 14644 36382
rect 14252 28142 14420 28198
rect 14252 23518 14308 28142
rect 14588 28018 14644 36316
rect 14700 35140 14756 36602
rect 14700 35074 14756 35084
rect 13804 23462 14308 23518
rect 14364 27962 14644 28018
rect 14700 32788 14756 32798
rect 13804 16996 13860 23462
rect 14028 23380 14084 23390
rect 13916 22820 13972 22830
rect 13916 21028 13972 22764
rect 13916 20962 13972 20972
rect 13804 16930 13860 16940
rect 14028 14532 14084 23324
rect 14364 23044 14420 27962
rect 14700 27838 14756 32732
rect 14476 27782 14756 27838
rect 14476 23338 14532 27782
rect 14812 24052 14868 36988
rect 14924 26218 14980 39228
rect 15036 36820 15092 36830
rect 15036 35476 15092 36764
rect 15036 28532 15092 35420
rect 15036 28466 15092 28476
rect 14924 26162 15092 26218
rect 14476 23282 14756 23338
rect 14364 22978 14420 22988
rect 14364 22922 14532 22978
rect 14476 22618 14532 22922
rect 14364 22562 14532 22618
rect 14364 21538 14420 22562
rect 14700 22438 14756 23282
rect 14252 21482 14420 21538
rect 14476 22382 14756 22438
rect 14252 19572 14308 21482
rect 14252 19506 14308 19516
rect 14364 21252 14420 21262
rect 14364 16660 14420 21196
rect 14364 16594 14420 16604
rect 13804 14420 13860 14430
rect 13804 13300 13860 14364
rect 14028 13748 14084 14476
rect 14028 13682 14084 13692
rect 13804 13234 13860 13244
rect 14028 9828 14084 9838
rect 14028 8260 14084 9772
rect 14028 8194 14084 8204
rect 13692 3490 13748 3500
rect 14140 7028 14196 7038
rect 13468 2100 13524 3052
rect 14140 2548 14196 6972
rect 14140 2482 14196 2492
rect 14252 6580 14308 6590
rect 14252 5124 14308 6524
rect 13468 2034 13524 2044
rect 13244 1586 13300 1596
rect 11676 578 11732 588
rect 9324 420 9380 430
rect 9324 84 9380 364
rect 9324 18 9380 28
rect 14252 84 14308 5068
rect 14476 3556 14532 22382
rect 14700 22148 14756 22158
rect 14700 21476 14756 22092
rect 14700 21410 14756 21420
rect 14812 18340 14868 23996
rect 15036 26068 15092 26162
rect 14812 18274 14868 18284
rect 14924 23492 14980 23502
rect 14924 16100 14980 23436
rect 15036 21812 15092 26012
rect 15036 21746 15092 21756
rect 14924 16034 14980 16044
rect 14476 1988 14532 3500
rect 14476 1922 14532 1932
rect 15148 1204 15204 52668
rect 15260 50932 15316 108444
rect 15708 96628 15764 96638
rect 15596 93044 15652 93054
rect 15596 92596 15652 92988
rect 15596 92530 15652 92540
rect 15260 50866 15316 50876
rect 15596 54404 15652 54414
rect 15372 37044 15428 37054
rect 15372 5348 15428 36988
rect 15484 9044 15540 9054
rect 15484 7476 15540 8988
rect 15484 6804 15540 7420
rect 15484 5908 15540 6748
rect 15484 5842 15540 5852
rect 15372 5282 15428 5292
rect 15596 2772 15652 54348
rect 15708 36372 15764 96572
rect 15820 49812 15876 109452
rect 16044 72436 16100 112588
rect 17052 112644 17108 112654
rect 16156 112308 16212 112318
rect 16156 112084 16212 112252
rect 16156 112018 16212 112028
rect 16828 111524 16884 111534
rect 16156 104580 16212 104590
rect 16156 98308 16212 104524
rect 16156 98242 16212 98252
rect 16604 102900 16660 102910
rect 16044 72370 16100 72380
rect 16268 65716 16324 65726
rect 16268 60900 16324 65660
rect 16268 60834 16324 60844
rect 15820 49746 15876 49756
rect 16604 47348 16660 102844
rect 16828 100436 16884 111468
rect 16828 100370 16884 100380
rect 16940 97636 16996 97646
rect 16828 85092 16884 85102
rect 16604 47282 16660 47292
rect 16716 82628 16772 82638
rect 16716 46564 16772 82572
rect 16716 46498 16772 46508
rect 16828 43988 16884 85036
rect 16828 43922 16884 43932
rect 15708 36306 15764 36316
rect 16828 35252 16884 35262
rect 16828 34244 16884 35196
rect 16268 34132 16324 34142
rect 15596 2706 15652 2716
rect 15708 30324 15764 30334
rect 15708 2212 15764 30268
rect 16268 25172 16324 34076
rect 16716 32116 16772 32126
rect 16380 26292 16436 26302
rect 16380 25284 16436 26236
rect 16380 25218 16436 25228
rect 16268 25106 16324 25116
rect 16716 24612 16772 32060
rect 16828 29540 16884 34188
rect 16940 31220 16996 97580
rect 17052 85652 17108 112588
rect 17388 112308 17444 112318
rect 17388 101220 17444 112252
rect 17948 111860 18004 111870
rect 17724 111524 17780 111534
rect 17724 111188 17780 111468
rect 17724 111122 17780 111132
rect 17836 110964 17892 110974
rect 17388 101154 17444 101164
rect 17724 104244 17780 104254
rect 17724 99876 17780 104188
rect 17836 100212 17892 110908
rect 17836 100146 17892 100156
rect 17948 105588 18004 111804
rect 18620 110964 18676 110974
rect 18620 109508 18676 110908
rect 18620 109442 18676 109452
rect 19404 109172 19460 109182
rect 19404 108612 19460 109116
rect 19404 108546 19460 108556
rect 17724 99810 17780 99820
rect 17836 97972 17892 97982
rect 17836 96740 17892 97916
rect 17836 96180 17892 96684
rect 17836 96114 17892 96124
rect 17052 85586 17108 85596
rect 17164 94276 17220 94286
rect 17164 49700 17220 94220
rect 17836 93716 17892 93726
rect 17836 92372 17892 93660
rect 17276 92148 17332 92158
rect 17276 85428 17332 92092
rect 17836 90020 17892 92316
rect 17836 89954 17892 89964
rect 17948 93492 18004 105532
rect 19068 105588 19124 105598
rect 19068 104244 19124 105532
rect 19068 104178 19124 104188
rect 18396 98868 18452 98878
rect 18172 98420 18228 98430
rect 18172 96068 18228 98364
rect 18172 96002 18228 96012
rect 17276 85362 17332 85372
rect 17388 82404 17444 82414
rect 17388 72772 17444 82348
rect 17948 79380 18004 93436
rect 17948 79314 18004 79324
rect 17612 78932 17668 78942
rect 17612 74788 17668 78876
rect 17612 74004 17668 74732
rect 17612 73938 17668 73948
rect 17388 72706 17444 72716
rect 17164 49634 17220 49644
rect 17388 43652 17444 43662
rect 17164 41860 17220 41870
rect 16940 31154 16996 31164
rect 17052 33348 17108 33358
rect 16828 28084 16884 29484
rect 16828 28018 16884 28028
rect 16716 24546 16772 24556
rect 16492 23044 16548 23054
rect 16492 21028 16548 22988
rect 16492 20962 16548 20972
rect 16940 18340 16996 18350
rect 15932 16324 15988 16334
rect 15932 4004 15988 16268
rect 16940 13636 16996 18284
rect 17052 14980 17108 33292
rect 17052 14914 17108 14924
rect 16940 13570 16996 13580
rect 15932 3938 15988 3948
rect 16604 7812 16660 7822
rect 16604 2996 16660 7756
rect 17164 3556 17220 41804
rect 17276 32564 17332 32574
rect 17276 28420 17332 32508
rect 17388 29988 17444 43596
rect 18284 41972 18340 41982
rect 18172 40404 18228 40414
rect 18060 40180 18116 40190
rect 18060 39508 18116 40124
rect 17948 37268 18004 37278
rect 17724 36148 17780 36158
rect 17388 29922 17444 29932
rect 17500 35924 17556 35934
rect 17276 28354 17332 28364
rect 17500 26180 17556 35868
rect 17612 34804 17668 34814
rect 17612 31618 17668 34748
rect 17724 33124 17780 36092
rect 17724 33058 17780 33068
rect 17948 32116 18004 37212
rect 17948 32050 18004 32060
rect 17612 31562 17780 31618
rect 17500 26114 17556 26124
rect 17724 29316 17780 31562
rect 17164 3490 17220 3500
rect 17724 3444 17780 29260
rect 17836 28868 17892 28878
rect 17836 16660 17892 28812
rect 18060 28868 18116 39452
rect 18060 28802 18116 28812
rect 18172 28196 18228 40348
rect 18172 26964 18228 28140
rect 18172 26898 18228 26908
rect 18060 23044 18116 23054
rect 18060 20916 18116 22988
rect 18060 20850 18116 20860
rect 17836 16594 17892 16604
rect 18284 4340 18340 41916
rect 18396 40516 18452 98812
rect 18844 87220 18900 87230
rect 18732 86772 18788 86782
rect 18732 47460 18788 86716
rect 18844 83300 18900 87164
rect 18844 83234 18900 83244
rect 18732 47394 18788 47404
rect 19292 55524 19348 55534
rect 19292 47572 19348 55468
rect 18396 40450 18452 40460
rect 18844 43540 18900 43550
rect 18620 37604 18676 37614
rect 18508 36260 18564 36270
rect 18508 31220 18564 36204
rect 18620 33460 18676 37548
rect 18620 32228 18676 33404
rect 18620 32162 18676 32172
rect 18844 34132 18900 43484
rect 19292 36260 19348 47516
rect 19292 36194 19348 36204
rect 19404 44212 19460 44222
rect 18508 31154 18564 31164
rect 18844 29764 18900 34076
rect 19292 33348 19348 33358
rect 19292 32676 19348 33292
rect 19292 32610 19348 32620
rect 18844 29428 18900 29708
rect 18844 29362 18900 29372
rect 18956 30660 19012 30670
rect 18844 28756 18900 28766
rect 18732 27748 18788 27758
rect 18284 4274 18340 4284
rect 18620 26852 18676 26862
rect 17724 3378 17780 3388
rect 16604 2930 16660 2940
rect 18620 2772 18676 26796
rect 18732 26516 18788 27692
rect 18732 26450 18788 26460
rect 18732 23492 18788 23502
rect 18732 4452 18788 23436
rect 18844 22932 18900 28700
rect 18956 23044 19012 30604
rect 19404 23604 19460 44156
rect 19404 23538 19460 23548
rect 18956 22978 19012 22988
rect 18844 22866 18900 22876
rect 19516 14420 19572 113484
rect 19852 40404 19908 40414
rect 19852 38276 19908 40348
rect 19852 38210 19908 38220
rect 19628 33908 19684 33918
rect 19628 26964 19684 33852
rect 19740 33796 19796 33806
rect 19740 32452 19796 33740
rect 19852 33572 19908 33582
rect 19852 32564 19908 33516
rect 19852 32498 19908 32508
rect 19740 32386 19796 32396
rect 19852 28644 19908 28654
rect 19852 27748 19908 28588
rect 19852 27682 19908 27692
rect 19628 26898 19684 26908
rect 19516 14354 19572 14364
rect 19964 12628 20020 113932
rect 23776 112924 24096 114912
rect 23776 112868 23804 112924
rect 23860 112868 23908 112924
rect 23964 112868 24012 112924
rect 24068 112868 24096 112924
rect 21644 111860 21700 111870
rect 21308 106932 21364 106942
rect 20188 106708 20244 106718
rect 20076 98980 20132 98990
rect 20076 97860 20132 98924
rect 20076 92372 20132 97804
rect 20076 92306 20132 92316
rect 20076 73220 20132 73230
rect 20076 25732 20132 73164
rect 20188 56980 20244 106652
rect 20188 56914 20244 56924
rect 20300 103796 20356 103806
rect 20300 55524 20356 103740
rect 20748 67620 20804 67630
rect 20748 66500 20804 67564
rect 20748 66434 20804 66444
rect 21196 62468 21252 62478
rect 21196 62132 21252 62412
rect 21196 62066 21252 62076
rect 20300 55458 20356 55468
rect 20412 54628 20468 54638
rect 20188 36932 20244 36942
rect 20188 32004 20244 36876
rect 20412 34468 20468 54572
rect 20412 34402 20468 34412
rect 20524 39396 20580 39406
rect 20188 26404 20244 31948
rect 20524 30884 20580 39340
rect 20524 30818 20580 30828
rect 20188 26338 20244 26348
rect 20076 25666 20132 25676
rect 19964 12562 20020 12572
rect 19516 11956 19572 11966
rect 19516 8372 19572 11900
rect 19516 8306 19572 8316
rect 21308 7700 21364 106876
rect 21532 61236 21588 61246
rect 21420 41412 21476 41422
rect 21420 21476 21476 41356
rect 21420 21410 21476 21420
rect 21308 7634 21364 7644
rect 18732 4386 18788 4396
rect 18620 2706 18676 2716
rect 15708 2146 15764 2156
rect 21532 1540 21588 61180
rect 21644 17780 21700 111804
rect 22204 111860 22260 111870
rect 21980 91700 22036 91710
rect 21980 85652 22036 91644
rect 21980 85586 22036 85596
rect 21756 62244 21812 62254
rect 21756 22148 21812 62188
rect 21756 22082 21812 22092
rect 21644 17714 21700 17724
rect 21644 11284 21700 11294
rect 21644 7812 21700 11228
rect 21644 5572 21700 7756
rect 21644 5506 21700 5516
rect 22092 10724 22148 10734
rect 22092 2212 22148 10668
rect 22204 8036 22260 111804
rect 23776 111356 24096 112868
rect 23776 111300 23804 111356
rect 23860 111300 23908 111356
rect 23964 111300 24012 111356
rect 24068 111300 24096 111356
rect 22316 110964 22372 110974
rect 22316 16772 22372 110908
rect 23212 110964 23268 110974
rect 23212 109918 23268 110908
rect 23212 109862 23380 109918
rect 22652 87556 22708 87566
rect 22428 80948 22484 80958
rect 22428 79604 22484 80892
rect 22428 79538 22484 79548
rect 22316 16706 22372 16716
rect 22652 16660 22708 87500
rect 23100 86772 23156 86782
rect 23100 85316 23156 86716
rect 23100 85250 23156 85260
rect 22652 16594 22708 16604
rect 22988 77700 23044 77710
rect 22988 10388 23044 77644
rect 23100 23492 23156 23502
rect 23100 22932 23156 23436
rect 23100 22866 23156 22876
rect 22988 10322 23044 10332
rect 22204 7970 22260 7980
rect 23324 5348 23380 109862
rect 23776 109788 24096 111300
rect 23776 109732 23804 109788
rect 23860 109732 23908 109788
rect 23964 109732 24012 109788
rect 24068 109732 24096 109788
rect 23324 5282 23380 5292
rect 23436 108500 23492 108510
rect 22092 2146 22148 2156
rect 23100 3108 23156 3118
rect 23100 2212 23156 3052
rect 23100 2146 23156 2156
rect 21532 1474 21588 1484
rect 23436 1316 23492 108444
rect 23776 108220 24096 109732
rect 23776 108164 23804 108220
rect 23860 108164 23908 108220
rect 23964 108164 24012 108220
rect 24068 108164 24096 108220
rect 23776 106652 24096 108164
rect 23776 106596 23804 106652
rect 23860 106596 23908 106652
rect 23964 106596 24012 106652
rect 24068 106596 24096 106652
rect 23776 105084 24096 106596
rect 23776 105028 23804 105084
rect 23860 105028 23908 105084
rect 23964 105028 24012 105084
rect 24068 105028 24096 105084
rect 23776 103516 24096 105028
rect 23776 103460 23804 103516
rect 23860 103460 23908 103516
rect 23964 103460 24012 103516
rect 24068 103460 24096 103516
rect 23776 101948 24096 103460
rect 23776 101892 23804 101948
rect 23860 101892 23908 101948
rect 23964 101892 24012 101948
rect 24068 101892 24096 101948
rect 23776 100380 24096 101892
rect 23776 100324 23804 100380
rect 23860 100324 23908 100380
rect 23964 100324 24012 100380
rect 24068 100324 24096 100380
rect 23776 98812 24096 100324
rect 23776 98756 23804 98812
rect 23860 98756 23908 98812
rect 23964 98756 24012 98812
rect 24068 98756 24096 98812
rect 23776 97244 24096 98756
rect 23776 97188 23804 97244
rect 23860 97188 23908 97244
rect 23964 97188 24012 97244
rect 24068 97188 24096 97244
rect 23776 95676 24096 97188
rect 23776 95620 23804 95676
rect 23860 95620 23908 95676
rect 23964 95620 24012 95676
rect 24068 95620 24096 95676
rect 23776 94108 24096 95620
rect 23776 94052 23804 94108
rect 23860 94052 23908 94108
rect 23964 94052 24012 94108
rect 24068 94052 24096 94108
rect 23776 92540 24096 94052
rect 23776 92484 23804 92540
rect 23860 92484 23908 92540
rect 23964 92484 24012 92540
rect 24068 92484 24096 92540
rect 23776 90972 24096 92484
rect 23776 90916 23804 90972
rect 23860 90916 23908 90972
rect 23964 90916 24012 90972
rect 24068 90916 24096 90972
rect 23776 89404 24096 90916
rect 23776 89348 23804 89404
rect 23860 89348 23908 89404
rect 23964 89348 24012 89404
rect 24068 89348 24096 89404
rect 23776 87836 24096 89348
rect 23776 87780 23804 87836
rect 23860 87780 23908 87836
rect 23964 87780 24012 87836
rect 24068 87780 24096 87836
rect 23776 86268 24096 87780
rect 23776 86212 23804 86268
rect 23860 86212 23908 86268
rect 23964 86212 24012 86268
rect 24068 86212 24096 86268
rect 23548 86100 23604 86110
rect 23548 85540 23604 86044
rect 23548 85474 23604 85484
rect 23776 84700 24096 86212
rect 23776 84644 23804 84700
rect 23860 84644 23908 84700
rect 23964 84644 24012 84700
rect 24068 84644 24096 84700
rect 23776 83132 24096 84644
rect 23776 83076 23804 83132
rect 23860 83076 23908 83132
rect 23964 83076 24012 83132
rect 24068 83076 24096 83132
rect 23776 81564 24096 83076
rect 23776 81508 23804 81564
rect 23860 81508 23908 81564
rect 23964 81508 24012 81564
rect 24068 81508 24096 81564
rect 23776 79996 24096 81508
rect 23776 79940 23804 79996
rect 23860 79940 23908 79996
rect 23964 79940 24012 79996
rect 24068 79940 24096 79996
rect 23776 78428 24096 79940
rect 23776 78372 23804 78428
rect 23860 78372 23908 78428
rect 23964 78372 24012 78428
rect 24068 78372 24096 78428
rect 23776 76860 24096 78372
rect 23776 76804 23804 76860
rect 23860 76804 23908 76860
rect 23964 76804 24012 76860
rect 24068 76804 24096 76860
rect 23776 75292 24096 76804
rect 23776 75236 23804 75292
rect 23860 75236 23908 75292
rect 23964 75236 24012 75292
rect 24068 75236 24096 75292
rect 23776 73724 24096 75236
rect 23776 73668 23804 73724
rect 23860 73668 23908 73724
rect 23964 73668 24012 73724
rect 24068 73668 24096 73724
rect 23776 72156 24096 73668
rect 23776 72100 23804 72156
rect 23860 72100 23908 72156
rect 23964 72100 24012 72156
rect 24068 72100 24096 72156
rect 23776 70588 24096 72100
rect 23776 70532 23804 70588
rect 23860 70532 23908 70588
rect 23964 70532 24012 70588
rect 24068 70532 24096 70588
rect 23776 69020 24096 70532
rect 23776 68964 23804 69020
rect 23860 68964 23908 69020
rect 23964 68964 24012 69020
rect 24068 68964 24096 69020
rect 23776 67452 24096 68964
rect 23776 67396 23804 67452
rect 23860 67396 23908 67452
rect 23964 67396 24012 67452
rect 24068 67396 24096 67452
rect 23776 65884 24096 67396
rect 23776 65828 23804 65884
rect 23860 65828 23908 65884
rect 23964 65828 24012 65884
rect 24068 65828 24096 65884
rect 23776 64316 24096 65828
rect 23776 64260 23804 64316
rect 23860 64260 23908 64316
rect 23964 64260 24012 64316
rect 24068 64260 24096 64316
rect 23776 62748 24096 64260
rect 23776 62692 23804 62748
rect 23860 62692 23908 62748
rect 23964 62692 24012 62748
rect 24068 62692 24096 62748
rect 23776 61180 24096 62692
rect 23776 61124 23804 61180
rect 23860 61124 23908 61180
rect 23964 61124 24012 61180
rect 24068 61124 24096 61180
rect 23776 59612 24096 61124
rect 23776 59556 23804 59612
rect 23860 59556 23908 59612
rect 23964 59556 24012 59612
rect 24068 59556 24096 59612
rect 23776 58044 24096 59556
rect 23776 57988 23804 58044
rect 23860 57988 23908 58044
rect 23964 57988 24012 58044
rect 24068 57988 24096 58044
rect 23776 56476 24096 57988
rect 23776 56420 23804 56476
rect 23860 56420 23908 56476
rect 23964 56420 24012 56476
rect 24068 56420 24096 56476
rect 23776 54908 24096 56420
rect 23776 54852 23804 54908
rect 23860 54852 23908 54908
rect 23964 54852 24012 54908
rect 24068 54852 24096 54908
rect 23776 53340 24096 54852
rect 23776 53284 23804 53340
rect 23860 53284 23908 53340
rect 23964 53284 24012 53340
rect 24068 53284 24096 53340
rect 23776 51772 24096 53284
rect 23776 51716 23804 51772
rect 23860 51716 23908 51772
rect 23964 51716 24012 51772
rect 24068 51716 24096 51772
rect 23776 50204 24096 51716
rect 23776 50148 23804 50204
rect 23860 50148 23908 50204
rect 23964 50148 24012 50204
rect 24068 50148 24096 50204
rect 23776 48636 24096 50148
rect 23776 48580 23804 48636
rect 23860 48580 23908 48636
rect 23964 48580 24012 48636
rect 24068 48580 24096 48636
rect 23776 47068 24096 48580
rect 23548 47012 23604 47022
rect 23548 3780 23604 46956
rect 23776 47012 23804 47068
rect 23860 47012 23908 47068
rect 23964 47012 24012 47068
rect 24068 47012 24096 47068
rect 23776 45500 24096 47012
rect 23776 45444 23804 45500
rect 23860 45444 23908 45500
rect 23964 45444 24012 45500
rect 24068 45444 24096 45500
rect 23776 43932 24096 45444
rect 23776 43876 23804 43932
rect 23860 43876 23908 43932
rect 23964 43876 24012 43932
rect 24068 43876 24096 43932
rect 23776 42364 24096 43876
rect 23776 42308 23804 42364
rect 23860 42308 23908 42364
rect 23964 42308 24012 42364
rect 24068 42308 24096 42364
rect 23776 40796 24096 42308
rect 23776 40740 23804 40796
rect 23860 40740 23908 40796
rect 23964 40740 24012 40796
rect 24068 40740 24096 40796
rect 23776 39228 24096 40740
rect 23776 39172 23804 39228
rect 23860 39172 23908 39228
rect 23964 39172 24012 39228
rect 24068 39172 24096 39228
rect 23776 37660 24096 39172
rect 23776 37604 23804 37660
rect 23860 37604 23908 37660
rect 23964 37604 24012 37660
rect 24068 37604 24096 37660
rect 23776 36092 24096 37604
rect 23776 36036 23804 36092
rect 23860 36036 23908 36092
rect 23964 36036 24012 36092
rect 24068 36036 24096 36092
rect 23776 34524 24096 36036
rect 23776 34468 23804 34524
rect 23860 34468 23908 34524
rect 23964 34468 24012 34524
rect 24068 34468 24096 34524
rect 23776 32956 24096 34468
rect 23776 32900 23804 32956
rect 23860 32900 23908 32956
rect 23964 32900 24012 32956
rect 24068 32900 24096 32956
rect 23776 31388 24096 32900
rect 23776 31332 23804 31388
rect 23860 31332 23908 31388
rect 23964 31332 24012 31388
rect 24068 31332 24096 31388
rect 23776 29820 24096 31332
rect 23776 29764 23804 29820
rect 23860 29764 23908 29820
rect 23964 29764 24012 29820
rect 24068 29764 24096 29820
rect 23776 28252 24096 29764
rect 23776 28196 23804 28252
rect 23860 28196 23908 28252
rect 23964 28196 24012 28252
rect 24068 28196 24096 28252
rect 23776 26684 24096 28196
rect 23776 26628 23804 26684
rect 23860 26628 23908 26684
rect 23964 26628 24012 26684
rect 24068 26628 24096 26684
rect 23776 25116 24096 26628
rect 23776 25060 23804 25116
rect 23860 25060 23908 25116
rect 23964 25060 24012 25116
rect 24068 25060 24096 25116
rect 23776 23548 24096 25060
rect 23776 23492 23804 23548
rect 23860 23492 23908 23548
rect 23964 23492 24012 23548
rect 24068 23492 24096 23548
rect 23660 22260 23716 22270
rect 23660 18676 23716 22204
rect 23660 18610 23716 18620
rect 23776 21980 24096 23492
rect 23776 21924 23804 21980
rect 23860 21924 23908 21980
rect 23964 21924 24012 21980
rect 24068 21924 24096 21980
rect 23776 20412 24096 21924
rect 23776 20356 23804 20412
rect 23860 20356 23908 20412
rect 23964 20356 24012 20412
rect 24068 20356 24096 20412
rect 23776 18844 24096 20356
rect 23776 18788 23804 18844
rect 23860 18788 23908 18844
rect 23964 18788 24012 18844
rect 24068 18788 24096 18844
rect 23776 17276 24096 18788
rect 23776 17220 23804 17276
rect 23860 17220 23908 17276
rect 23964 17220 24012 17276
rect 24068 17220 24096 17276
rect 23776 15708 24096 17220
rect 23776 15652 23804 15708
rect 23860 15652 23908 15708
rect 23964 15652 24012 15708
rect 24068 15652 24096 15708
rect 23776 14140 24096 15652
rect 23776 14084 23804 14140
rect 23860 14084 23908 14140
rect 23964 14084 24012 14140
rect 24068 14084 24096 14140
rect 23776 12572 24096 14084
rect 23776 12516 23804 12572
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 24068 12516 24096 12572
rect 23776 11004 24096 12516
rect 23776 10948 23804 11004
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 24068 10948 24096 11004
rect 23776 9436 24096 10948
rect 23776 9380 23804 9436
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 24068 9380 24096 9436
rect 23776 7868 24096 9380
rect 23776 7812 23804 7868
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 24068 7812 24096 7868
rect 23548 3714 23604 3724
rect 23660 6916 23716 6926
rect 23548 2324 23604 2334
rect 23548 2100 23604 2268
rect 23548 2034 23604 2044
rect 23660 1428 23716 6860
rect 23660 1362 23716 1372
rect 23776 6300 24096 7812
rect 23776 6244 23804 6300
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 24068 6244 24096 6300
rect 23776 4732 24096 6244
rect 24436 113708 24756 114912
rect 24436 113652 24464 113708
rect 24520 113652 24568 113708
rect 24624 113652 24672 113708
rect 24728 113652 24756 113708
rect 24436 112140 24756 113652
rect 24436 112084 24464 112140
rect 24520 112084 24568 112140
rect 24624 112084 24672 112140
rect 24728 112084 24756 112140
rect 27356 113652 27412 113662
rect 24436 110572 24756 112084
rect 24436 110516 24464 110572
rect 24520 110516 24568 110572
rect 24624 110516 24672 110572
rect 24728 110516 24756 110572
rect 24436 109004 24756 110516
rect 25340 112084 25396 112094
rect 25340 110628 25396 112028
rect 27020 110852 27076 110862
rect 24436 108948 24464 109004
rect 24520 108948 24568 109004
rect 24624 108948 24672 109004
rect 24728 108948 24756 109004
rect 24436 107436 24756 108948
rect 25228 110292 25284 110302
rect 25228 107940 25284 110236
rect 25340 109060 25396 110572
rect 25340 108994 25396 109004
rect 26908 110740 26964 110750
rect 26908 108836 26964 110684
rect 26908 108770 26964 108780
rect 25228 107874 25284 107884
rect 26236 108612 26292 108622
rect 24436 107380 24464 107436
rect 24520 107380 24568 107436
rect 24624 107380 24672 107436
rect 24728 107380 24756 107436
rect 24436 105868 24756 107380
rect 24436 105812 24464 105868
rect 24520 105812 24568 105868
rect 24624 105812 24672 105868
rect 24728 105812 24756 105868
rect 24436 104300 24756 105812
rect 24436 104244 24464 104300
rect 24520 104244 24568 104300
rect 24624 104244 24672 104300
rect 24728 104244 24756 104300
rect 24436 102732 24756 104244
rect 24436 102676 24464 102732
rect 24520 102676 24568 102732
rect 24624 102676 24672 102732
rect 24728 102676 24756 102732
rect 24436 101164 24756 102676
rect 24436 101108 24464 101164
rect 24520 101108 24568 101164
rect 24624 101108 24672 101164
rect 24728 101108 24756 101164
rect 24436 99596 24756 101108
rect 24436 99540 24464 99596
rect 24520 99540 24568 99596
rect 24624 99540 24672 99596
rect 24728 99540 24756 99596
rect 24436 98028 24756 99540
rect 24436 97972 24464 98028
rect 24520 97972 24568 98028
rect 24624 97972 24672 98028
rect 24728 97972 24756 98028
rect 24436 96460 24756 97972
rect 24436 96404 24464 96460
rect 24520 96404 24568 96460
rect 24624 96404 24672 96460
rect 24728 96404 24756 96460
rect 24436 94892 24756 96404
rect 24436 94836 24464 94892
rect 24520 94836 24568 94892
rect 24624 94836 24672 94892
rect 24728 94836 24756 94892
rect 24436 93324 24756 94836
rect 24436 93268 24464 93324
rect 24520 93268 24568 93324
rect 24624 93268 24672 93324
rect 24728 93268 24756 93324
rect 24436 91756 24756 93268
rect 24436 91700 24464 91756
rect 24520 91700 24568 91756
rect 24624 91700 24672 91756
rect 24728 91700 24756 91756
rect 24436 90188 24756 91700
rect 24436 90132 24464 90188
rect 24520 90132 24568 90188
rect 24624 90132 24672 90188
rect 24728 90132 24756 90188
rect 24436 88620 24756 90132
rect 24436 88564 24464 88620
rect 24520 88564 24568 88620
rect 24624 88564 24672 88620
rect 24728 88564 24756 88620
rect 24436 87052 24756 88564
rect 24436 86996 24464 87052
rect 24520 86996 24568 87052
rect 24624 86996 24672 87052
rect 24728 86996 24756 87052
rect 24436 85484 24756 86996
rect 24436 85428 24464 85484
rect 24520 85428 24568 85484
rect 24624 85428 24672 85484
rect 24728 85428 24756 85484
rect 24436 83916 24756 85428
rect 24436 83860 24464 83916
rect 24520 83860 24568 83916
rect 24624 83860 24672 83916
rect 24728 83860 24756 83916
rect 24436 82348 24756 83860
rect 24436 82292 24464 82348
rect 24520 82292 24568 82348
rect 24624 82292 24672 82348
rect 24728 82292 24756 82348
rect 24436 80780 24756 82292
rect 24436 80724 24464 80780
rect 24520 80724 24568 80780
rect 24624 80724 24672 80780
rect 24728 80724 24756 80780
rect 24436 79212 24756 80724
rect 24436 79156 24464 79212
rect 24520 79156 24568 79212
rect 24624 79156 24672 79212
rect 24728 79156 24756 79212
rect 24436 77644 24756 79156
rect 24436 77588 24464 77644
rect 24520 77588 24568 77644
rect 24624 77588 24672 77644
rect 24728 77588 24756 77644
rect 24436 76076 24756 77588
rect 24436 76020 24464 76076
rect 24520 76020 24568 76076
rect 24624 76020 24672 76076
rect 24728 76020 24756 76076
rect 24436 74508 24756 76020
rect 24436 74452 24464 74508
rect 24520 74452 24568 74508
rect 24624 74452 24672 74508
rect 24728 74452 24756 74508
rect 24436 72940 24756 74452
rect 24436 72884 24464 72940
rect 24520 72884 24568 72940
rect 24624 72884 24672 72940
rect 24728 72884 24756 72940
rect 24436 71372 24756 72884
rect 24436 71316 24464 71372
rect 24520 71316 24568 71372
rect 24624 71316 24672 71372
rect 24728 71316 24756 71372
rect 24436 69804 24756 71316
rect 24436 69748 24464 69804
rect 24520 69748 24568 69804
rect 24624 69748 24672 69804
rect 24728 69748 24756 69804
rect 24436 68236 24756 69748
rect 24436 68180 24464 68236
rect 24520 68180 24568 68236
rect 24624 68180 24672 68236
rect 24728 68180 24756 68236
rect 24436 66668 24756 68180
rect 24436 66612 24464 66668
rect 24520 66612 24568 66668
rect 24624 66612 24672 66668
rect 24728 66612 24756 66668
rect 24436 65100 24756 66612
rect 24436 65044 24464 65100
rect 24520 65044 24568 65100
rect 24624 65044 24672 65100
rect 24728 65044 24756 65100
rect 24436 63532 24756 65044
rect 24436 63476 24464 63532
rect 24520 63476 24568 63532
rect 24624 63476 24672 63532
rect 24728 63476 24756 63532
rect 24436 61964 24756 63476
rect 24436 61908 24464 61964
rect 24520 61908 24568 61964
rect 24624 61908 24672 61964
rect 24728 61908 24756 61964
rect 24436 60396 24756 61908
rect 24436 60340 24464 60396
rect 24520 60340 24568 60396
rect 24624 60340 24672 60396
rect 24728 60340 24756 60396
rect 24436 58828 24756 60340
rect 24436 58772 24464 58828
rect 24520 58772 24568 58828
rect 24624 58772 24672 58828
rect 24728 58772 24756 58828
rect 24436 57260 24756 58772
rect 24436 57204 24464 57260
rect 24520 57204 24568 57260
rect 24624 57204 24672 57260
rect 24728 57204 24756 57260
rect 24436 55692 24756 57204
rect 24436 55636 24464 55692
rect 24520 55636 24568 55692
rect 24624 55636 24672 55692
rect 24728 55636 24756 55692
rect 24436 54124 24756 55636
rect 24436 54068 24464 54124
rect 24520 54068 24568 54124
rect 24624 54068 24672 54124
rect 24728 54068 24756 54124
rect 24436 52556 24756 54068
rect 24436 52500 24464 52556
rect 24520 52500 24568 52556
rect 24624 52500 24672 52556
rect 24728 52500 24756 52556
rect 24436 50988 24756 52500
rect 24436 50932 24464 50988
rect 24520 50932 24568 50988
rect 24624 50932 24672 50988
rect 24728 50932 24756 50988
rect 24436 49420 24756 50932
rect 24436 49364 24464 49420
rect 24520 49364 24568 49420
rect 24624 49364 24672 49420
rect 24728 49364 24756 49420
rect 24436 47852 24756 49364
rect 24436 47796 24464 47852
rect 24520 47796 24568 47852
rect 24624 47796 24672 47852
rect 24728 47796 24756 47852
rect 24436 46284 24756 47796
rect 24436 46228 24464 46284
rect 24520 46228 24568 46284
rect 24624 46228 24672 46284
rect 24728 46228 24756 46284
rect 24436 44716 24756 46228
rect 24436 44660 24464 44716
rect 24520 44660 24568 44716
rect 24624 44660 24672 44716
rect 24728 44660 24756 44716
rect 24436 43148 24756 44660
rect 24436 43092 24464 43148
rect 24520 43092 24568 43148
rect 24624 43092 24672 43148
rect 24728 43092 24756 43148
rect 24436 41580 24756 43092
rect 24436 41524 24464 41580
rect 24520 41524 24568 41580
rect 24624 41524 24672 41580
rect 24728 41524 24756 41580
rect 24436 40012 24756 41524
rect 24436 39956 24464 40012
rect 24520 39956 24568 40012
rect 24624 39956 24672 40012
rect 24728 39956 24756 40012
rect 24436 38444 24756 39956
rect 24436 38388 24464 38444
rect 24520 38388 24568 38444
rect 24624 38388 24672 38444
rect 24728 38388 24756 38444
rect 24436 36876 24756 38388
rect 24436 36820 24464 36876
rect 24520 36820 24568 36876
rect 24624 36820 24672 36876
rect 24728 36820 24756 36876
rect 24436 35308 24756 36820
rect 24436 35252 24464 35308
rect 24520 35252 24568 35308
rect 24624 35252 24672 35308
rect 24728 35252 24756 35308
rect 24436 33740 24756 35252
rect 24436 33684 24464 33740
rect 24520 33684 24568 33740
rect 24624 33684 24672 33740
rect 24728 33684 24756 33740
rect 24436 32172 24756 33684
rect 24436 32116 24464 32172
rect 24520 32116 24568 32172
rect 24624 32116 24672 32172
rect 24728 32116 24756 32172
rect 24436 30604 24756 32116
rect 24436 30548 24464 30604
rect 24520 30548 24568 30604
rect 24624 30548 24672 30604
rect 24728 30548 24756 30604
rect 24436 29036 24756 30548
rect 24436 28980 24464 29036
rect 24520 28980 24568 29036
rect 24624 28980 24672 29036
rect 24728 28980 24756 29036
rect 24436 27468 24756 28980
rect 24436 27412 24464 27468
rect 24520 27412 24568 27468
rect 24624 27412 24672 27468
rect 24728 27412 24756 27468
rect 24436 25900 24756 27412
rect 24436 25844 24464 25900
rect 24520 25844 24568 25900
rect 24624 25844 24672 25900
rect 24728 25844 24756 25900
rect 24436 24332 24756 25844
rect 24436 24276 24464 24332
rect 24520 24276 24568 24332
rect 24624 24276 24672 24332
rect 24728 24276 24756 24332
rect 24436 22764 24756 24276
rect 24436 22708 24464 22764
rect 24520 22708 24568 22764
rect 24624 22708 24672 22764
rect 24728 22708 24756 22764
rect 24436 21196 24756 22708
rect 24436 21140 24464 21196
rect 24520 21140 24568 21196
rect 24624 21140 24672 21196
rect 24728 21140 24756 21196
rect 24436 19628 24756 21140
rect 26124 106260 26180 106270
rect 24436 19572 24464 19628
rect 24520 19572 24568 19628
rect 24624 19572 24672 19628
rect 24728 19572 24756 19628
rect 24436 18060 24756 19572
rect 24436 18004 24464 18060
rect 24520 18004 24568 18060
rect 24624 18004 24672 18060
rect 24728 18004 24756 18060
rect 24436 16492 24756 18004
rect 24436 16436 24464 16492
rect 24520 16436 24568 16492
rect 24624 16436 24672 16492
rect 24728 16436 24756 16492
rect 24436 14924 24756 16436
rect 24436 14868 24464 14924
rect 24520 14868 24568 14924
rect 24624 14868 24672 14924
rect 24728 14868 24756 14924
rect 24436 13356 24756 14868
rect 26012 20244 26068 20254
rect 26012 14644 26068 20188
rect 26012 14578 26068 14588
rect 24436 13300 24464 13356
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24728 13300 24756 13356
rect 24436 11788 24756 13300
rect 24436 11732 24464 11788
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24728 11732 24756 11788
rect 24436 10220 24756 11732
rect 24436 10164 24464 10220
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24728 10164 24756 10220
rect 24436 8652 24756 10164
rect 24436 8596 24464 8652
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24728 8596 24756 8652
rect 24436 7084 24756 8596
rect 25116 10052 25172 10062
rect 25004 7700 25060 7710
rect 24436 7028 24464 7084
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 24728 7028 24756 7084
rect 24436 5516 24756 7028
rect 24436 5460 24464 5516
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24728 5460 24756 5516
rect 23776 4676 23804 4732
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 24068 4676 24096 4732
rect 23776 3164 24096 4676
rect 23776 3108 23804 3164
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 24068 3108 24096 3164
rect 23776 1596 24096 3108
rect 23776 1540 23804 1596
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 24068 1540 24096 1596
rect 23436 1250 23492 1260
rect 15148 1138 15204 1148
rect 14252 18 14308 28
rect 19964 308 20020 318
rect 19964 84 20020 252
rect 19964 18 20020 28
rect 23776 0 24096 1540
rect 24220 5124 24276 5134
rect 24220 644 24276 5068
rect 24220 578 24276 588
rect 24436 3948 24756 5460
rect 24436 3892 24464 3948
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24728 3892 24756 3948
rect 24436 2380 24756 3892
rect 24436 2324 24464 2380
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24728 2324 24756 2380
rect 24436 812 24756 2324
rect 24436 756 24464 812
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24728 756 24756 812
rect 24436 0 24756 756
rect 24892 7364 24948 7374
rect 24892 644 24948 7308
rect 25004 1652 25060 7644
rect 25116 5348 25172 9996
rect 25452 8036 25508 8046
rect 25116 5282 25172 5292
rect 25228 5460 25284 5470
rect 25228 2324 25284 5404
rect 25452 2772 25508 7980
rect 25788 7028 25844 7038
rect 25564 6580 25620 6590
rect 25564 5908 25620 6524
rect 25564 5842 25620 5852
rect 25452 2706 25508 2716
rect 25228 2258 25284 2268
rect 25004 1586 25060 1596
rect 24892 578 24948 588
rect 25116 1316 25172 1326
rect 25116 532 25172 1260
rect 25788 868 25844 6972
rect 25900 2996 25956 3006
rect 25900 1876 25956 2940
rect 26124 2772 26180 106204
rect 26124 2706 26180 2716
rect 25900 1810 25956 1820
rect 26236 1428 26292 108556
rect 26796 107604 26852 107614
rect 26572 80052 26628 80062
rect 26572 76468 26628 79996
rect 26572 76402 26628 76412
rect 26572 15988 26628 15998
rect 26572 14644 26628 15932
rect 26572 14578 26628 14588
rect 26348 5236 26404 5246
rect 26348 2212 26404 5180
rect 26684 3892 26740 3902
rect 26684 2324 26740 3836
rect 26796 3556 26852 107548
rect 26796 3490 26852 3500
rect 26684 2258 26740 2268
rect 26348 2146 26404 2156
rect 27020 1540 27076 110796
rect 27132 110404 27188 110414
rect 27132 109060 27188 110348
rect 27356 110404 27412 113596
rect 27356 110338 27412 110348
rect 27132 108994 27188 109004
rect 28028 109172 28084 109182
rect 27692 12404 27748 12414
rect 27692 4788 27748 12348
rect 27692 4722 27748 4732
rect 27020 1474 27076 1484
rect 26236 1362 26292 1372
rect 28028 1204 28084 109116
rect 28588 7588 28644 7598
rect 28588 2996 28644 7532
rect 28588 2930 28644 2940
rect 28028 1138 28084 1148
rect 25788 802 25844 812
rect 25116 466 25172 476
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0210_
timestamp 1486834041
transform 1 0 16576 0 -1 33712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0211_
timestamp 1486834041
transform 1 0 15904 0 -1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0212_
timestamp 1486834041
transform -1 0 19936 0 -1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0213_
timestamp 1486834041
transform 1 0 16576 0 -1 35280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0214_
timestamp 1486834041
transform -1 0 22176 0 1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0215_
timestamp 1486834041
transform -1 0 29904 0 1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0216_
timestamp 1486834041
transform 1 0 11984 0 1 102704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0217_
timestamp 1486834041
transform -1 0 8512 0 -1 99568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0218_
timestamp 1486834041
transform 1 0 22960 0 1 66640
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0219_
timestamp 1486834041
transform -1 0 24192 0 -1 87024
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0220_
timestamp 1486834041
transform -1 0 17920 0 -1 61936
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0221_
timestamp 1486834041
transform -1 0 11536 0 1 72912
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0222_
timestamp 1486834041
transform -1 0 12432 0 1 77616
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0223_
timestamp 1486834041
transform 1 0 14896 0 1 80752
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0224_
timestamp 1486834041
transform 1 0 22848 0 -1 85456
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0225_
timestamp 1486834041
transform 1 0 13776 0 1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0226_
timestamp 1486834041
transform -1 0 20160 0 1 98000
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0227_
timestamp 1486834041
transform -1 0 15456 0 -1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0228_
timestamp 1486834041
transform 1 0 9744 0 1 49392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0229_
timestamp 1486834041
transform -1 0 8400 0 -1 47824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0230_
timestamp 1486834041
transform 1 0 22848 0 1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0231_
timestamp 1486834041
transform -1 0 20944 0 1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0232_
timestamp 1486834041
transform -1 0 17920 0 1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0233_
timestamp 1486834041
transform -1 0 16688 0 1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0234_
timestamp 1486834041
transform 1 0 21504 0 -1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0235_
timestamp 1486834041
transform -1 0 19376 0 -1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0236_
timestamp 1486834041
transform 1 0 3136 0 -1 88592
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0237_
timestamp 1486834041
transform -1 0 11088 0 1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0238_
timestamp 1486834041
transform -1 0 8512 0 -1 29008
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0239_
timestamp 1486834041
transform 1 0 10752 0 -1 63504
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0240_
timestamp 1486834041
transform 1 0 16688 0 1 29008
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0241_
timestamp 1486834041
transform 1 0 15792 0 -1 30576
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0242_
timestamp 1486834041
transform -1 0 19488 0 -1 27440
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0243_
timestamp 1486834041
transform -1 0 17472 0 1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0244_
timestamp 1486834041
transform 1 0 16912 0 -1 30576
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0245_
timestamp 1486834041
transform -1 0 21168 0 -1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _0246_
timestamp 1486834041
transform 1 0 18480 0 -1 32144
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0247_
timestamp 1486834041
transform -1 0 19152 0 1 30576
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _0248_
timestamp 1486834041
transform 1 0 20496 0 1 29008
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0249_
timestamp 1486834041
transform 1 0 18368 0 -1 27440
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0250_
timestamp 1486834041
transform 1 0 21168 0 -1 30576
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0251_
timestamp 1486834041
transform -1 0 20384 0 -1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0252_
timestamp 1486834041
transform 1 0 19152 0 1 30576
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0253_
timestamp 1486834041
transform 1 0 21840 0 1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _0254_
timestamp 1486834041
transform -1 0 21728 0 1 27440
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0255_
timestamp 1486834041
transform 1 0 12656 0 1 102704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0256_
timestamp 1486834041
transform -1 0 12880 0 -1 104272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0257_
timestamp 1486834041
transform -1 0 16016 0 -1 104272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0258_
timestamp 1486834041
transform -1 0 12432 0 1 104272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0259_
timestamp 1486834041
transform 1 0 9408 0 -1 101136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0260_
timestamp 1486834041
transform 1 0 10192 0 -1 46256
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0261_
timestamp 1486834041
transform 1 0 11760 0 1 47824
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0262_
timestamp 1486834041
transform 1 0 11200 0 1 47824
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0263_
timestamp 1486834041
transform 1 0 12768 0 -1 47824
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0264_
timestamp 1486834041
transform 1 0 12880 0 1 47824
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0265_
timestamp 1486834041
transform 1 0 12656 0 1 50960
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0266_
timestamp 1486834041
transform 1 0 12768 0 -1 102704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0267_
timestamp 1486834041
transform 1 0 8512 0 1 101136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0268_
timestamp 1486834041
transform 1 0 4928 0 1 91728
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0269_
timestamp 1486834041
transform 1 0 4032 0 1 98000
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0270_
timestamp 1486834041
transform -1 0 8400 0 -1 98000
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0271_
timestamp 1486834041
transform 1 0 7168 0 -1 96432
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0272_
timestamp 1486834041
transform -1 0 7168 0 -1 101136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0273_
timestamp 1486834041
transform 1 0 5936 0 1 44688
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0274_
timestamp 1486834041
transform 1 0 9520 0 1 44688
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0275_
timestamp 1486834041
transform 1 0 8736 0 -1 44688
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0276_
timestamp 1486834041
transform 1 0 5376 0 1 44688
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0277_
timestamp 1486834041
transform 1 0 8736 0 -1 46256
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0278_
timestamp 1486834041
transform 1 0 9072 0 -1 47824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0279_
timestamp 1486834041
transform 1 0 5936 0 1 104272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0280_
timestamp 1486834041
transform -1 0 7280 0 -1 102704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0281_
timestamp 1486834041
transform 1 0 23296 0 -1 69776
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0282_
timestamp 1486834041
transform 1 0 18816 0 1 68208
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0283_
timestamp 1486834041
transform 1 0 19376 0 1 68208
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0284_
timestamp 1486834041
transform 1 0 24080 0 1 68208
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0285_
timestamp 1486834041
transform 1 0 20496 0 1 61936
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0286_
timestamp 1486834041
transform 1 0 20272 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0287_
timestamp 1486834041
transform 1 0 23072 0 -1 24304
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0288_
timestamp 1486834041
transform -1 0 24416 0 1 22736
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0289_
timestamp 1486834041
transform 1 0 23184 0 -1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0290_
timestamp 1486834041
transform -1 0 23856 0 1 22736
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0291_
timestamp 1486834041
transform 1 0 20496 0 1 43120
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0292_
timestamp 1486834041
transform 1 0 20496 0 1 60368
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0293_
timestamp 1486834041
transform 1 0 20272 0 -1 80752
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0294_
timestamp 1486834041
transform 1 0 2912 0 -1 90160
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0295_
timestamp 1486834041
transform -1 0 4592 0 1 99568
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0296_
timestamp 1486834041
transform -1 0 10304 0 1 52528
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0297_
timestamp 1486834041
transform 1 0 9744 0 -1 44688
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0298_
timestamp 1486834041
transform 1 0 8848 0 1 107408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0299_
timestamp 1486834041
transform -1 0 4592 0 1 101136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0300_
timestamp 1486834041
transform -1 0 4592 0 1 105840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0301_
timestamp 1486834041
transform 1 0 12768 0 -1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0302_
timestamp 1486834041
transform 1 0 9856 0 -1 41552
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0303_
timestamp 1486834041
transform 1 0 14560 0 1 107408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0304_
timestamp 1486834041
transform -1 0 5264 0 -1 107408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0305_
timestamp 1486834041
transform 1 0 18704 0 -1 87024
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0306_
timestamp 1486834041
transform 1 0 16576 0 -1 47824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0307_
timestamp 1486834041
transform 1 0 13552 0 1 38416
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0308_
timestamp 1486834041
transform -1 0 20160 0 -1 104272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0309_
timestamp 1486834041
transform 1 0 7840 0 1 85456
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0310_
timestamp 1486834041
transform 1 0 11872 0 -1 82320
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0311_
timestamp 1486834041
transform -1 0 14784 0 -1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0312_
timestamp 1486834041
transform 1 0 15008 0 1 32144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0313_
timestamp 1486834041
transform 1 0 12768 0 -1 85456
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0314_
timestamp 1486834041
transform 1 0 8736 0 -1 83888
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0315_
timestamp 1486834041
transform 1 0 8288 0 1 79184
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0316_
timestamp 1486834041
transform 1 0 8512 0 1 19600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0317_
timestamp 1486834041
transform 1 0 8624 0 1 33712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0318_
timestamp 1486834041
transform 1 0 10752 0 -1 108976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0319_
timestamp 1486834041
transform 1 0 5712 0 1 88592
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0320_
timestamp 1486834041
transform -1 0 10416 0 1 72912
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0321_
timestamp 1486834041
transform 1 0 14000 0 1 54096
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0322_
timestamp 1486834041
transform -1 0 16352 0 -1 43120
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0323_
timestamp 1486834041
transform 1 0 12768 0 -1 110544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0324_
timestamp 1486834041
transform 1 0 5936 0 1 90160
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0325_
timestamp 1486834041
transform 1 0 14112 0 1 61936
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0326_
timestamp 1486834041
transform 1 0 15232 0 1 49392
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0327_
timestamp 1486834041
transform 1 0 16016 0 1 39984
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0328_
timestamp 1486834041
transform 1 0 15344 0 1 108976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0329_
timestamp 1486834041
transform -1 0 12432 0 1 87024
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0330_
timestamp 1486834041
transform 1 0 18144 0 1 96432
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0331_
timestamp 1486834041
transform -1 0 17360 0 -1 96432
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0332_
timestamp 1486834041
transform 1 0 18816 0 -1 98000
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0333_
timestamp 1486834041
transform 1 0 18592 0 1 98000
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0334_
timestamp 1486834041
transform 1 0 14560 0 1 96432
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0335_
timestamp 1486834041
transform 1 0 14448 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0336_
timestamp 1486834041
transform 1 0 14224 0 1 22736
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0337_
timestamp 1486834041
transform -1 0 14112 0 -1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0338_
timestamp 1486834041
transform 1 0 13552 0 1 22736
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0339_
timestamp 1486834041
transform -1 0 15232 0 -1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0340_
timestamp 1486834041
transform 1 0 12992 0 1 22736
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0341_
timestamp 1486834041
transform 1 0 15120 0 1 22736
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0342_
timestamp 1486834041
transform 1 0 15456 0 -1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0343_
timestamp 1486834041
transform -1 0 18256 0 -1 25872
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0344_
timestamp 1486834041
transform 1 0 16464 0 1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _0345_
timestamp 1486834041
transform 1 0 16576 0 -1 25872
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0346_
timestamp 1486834041
transform 1 0 14448 0 1 57232
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0347_
timestamp 1486834041
transform 1 0 11424 0 -1 61936
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0348_
timestamp 1486834041
transform 1 0 5936 0 1 71344
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0349_
timestamp 1486834041
transform 1 0 16800 0 -1 60368
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0350_
timestamp 1486834041
transform 1 0 5488 0 1 60368
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0351_
timestamp 1486834041
transform 1 0 1008 0 1 83888
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0352_
timestamp 1486834041
transform 1 0 1008 0 1 82320
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0353_
timestamp 1486834041
transform 1 0 9184 0 -1 66640
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0354_
timestamp 1486834041
transform 1 0 8848 0 1 65072
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0355_
timestamp 1486834041
transform 1 0 1792 0 -1 63504
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0356_
timestamp 1486834041
transform 1 0 1344 0 -1 80752
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0357_
timestamp 1486834041
transform 1 0 4928 0 -1 66640
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0358_
timestamp 1486834041
transform 1 0 5488 0 1 61936
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0359_
timestamp 1486834041
transform 1 0 1792 0 -1 69776
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0360_
timestamp 1486834041
transform 1 0 1904 0 -1 65072
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0361_
timestamp 1486834041
transform 1 0 8848 0 1 69776
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0362_
timestamp 1486834041
transform 1 0 8848 0 -1 65072
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0363_
timestamp 1486834041
transform 1 0 1008 0 1 61936
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0364_
timestamp 1486834041
transform 1 0 1344 0 -1 71344
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0365_
timestamp 1486834041
transform 1 0 4928 0 -1 61936
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0366_
timestamp 1486834041
transform 1 0 18032 0 -1 61936
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0367_
timestamp 1486834041
transform 1 0 1680 0 -1 85456
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0368_
timestamp 1486834041
transform 1 0 4928 0 -1 83888
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0369_
timestamp 1486834041
transform 1 0 16352 0 1 76048
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0370_
timestamp 1486834041
transform 1 0 14000 0 1 66640
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0371_
timestamp 1486834041
transform 1 0 18032 0 -1 66640
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0372_
timestamp 1486834041
transform 1 0 16688 0 -1 68208
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0373_
timestamp 1486834041
transform 1 0 5936 0 1 110544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0374_
timestamp 1486834041
transform 1 0 4816 0 -1 68208
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0375_
timestamp 1486834041
transform 1 0 12656 0 1 104272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0376_
timestamp 1486834041
transform 1 0 3584 0 -1 82320
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0377_
timestamp 1486834041
transform 1 0 15456 0 1 79184
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0378_
timestamp 1486834041
transform 1 0 11984 0 -1 68208
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0379_
timestamp 1486834041
transform 1 0 20272 0 -1 68208
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0380_
timestamp 1486834041
transform 1 0 20496 0 1 68208
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0381_
timestamp 1486834041
transform 1 0 4592 0 -1 108976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0382_
timestamp 1486834041
transform 1 0 1904 0 -1 72912
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0383_
timestamp 1486834041
transform 1 0 13104 0 1 101136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0384_
timestamp 1486834041
transform 1 0 4928 0 -1 71344
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0385_
timestamp 1486834041
transform 1 0 16576 0 -1 83888
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0386_
timestamp 1486834041
transform 1 0 14448 0 1 71344
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0387_
timestamp 1486834041
transform 1 0 18928 0 -1 63504
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0388_
timestamp 1486834041
transform 1 0 20384 0 -1 72912
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0389_
timestamp 1486834041
transform 1 0 5936 0 1 108976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0390_
timestamp 1486834041
transform 1 0 2016 0 -1 76048
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0391_
timestamp 1486834041
transform 1 0 11312 0 -1 87024
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0392_
timestamp 1486834041
transform 1 0 6496 0 1 76048
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0393_
timestamp 1486834041
transform 1 0 16576 0 -1 79184
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0394_
timestamp 1486834041
transform 1 0 12656 0 1 72912
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0395_
timestamp 1486834041
transform 1 0 16576 0 1 74480
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0396_
timestamp 1486834041
transform 1 0 7280 0 1 83888
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0397_
timestamp 1486834041
transform 1 0 6160 0 1 102704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0398_
timestamp 1486834041
transform 1 0 15120 0 1 68208
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0399_
timestamp 1486834041
transform 1 0 17472 0 -1 74480
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0400_
timestamp 1486834041
transform 1 0 2800 0 -1 74480
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0401_
timestamp 1486834041
transform 1 0 4928 0 -1 80752
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0402_
timestamp 1486834041
transform 1 0 12656 0 1 74480
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0403_
timestamp 1486834041
transform 1 0 20608 0 -1 76048
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0404_
timestamp 1486834041
transform 1 0 2240 0 -1 77616
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0405_
timestamp 1486834041
transform 1 0 9744 0 -1 77616
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0406_
timestamp 1486834041
transform 1 0 12768 0 1 76048
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0407_
timestamp 1486834041
transform 1 0 15568 0 -1 63504
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0408_
timestamp 1486834041
transform -1 0 17472 0 -1 61936
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0409_
timestamp 1486834041
transform -1 0 15456 0 -1 63504
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0410_
timestamp 1486834041
transform 1 0 15232 0 -1 61936
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0411_
timestamp 1486834041
transform 1 0 10416 0 1 72912
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0412_
timestamp 1486834041
transform -1 0 9744 0 -1 72912
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0413_
timestamp 1486834041
transform -1 0 8512 0 -1 74480
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0414_
timestamp 1486834041
transform 1 0 9744 0 -1 72912
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0415_
timestamp 1486834041
transform 1 0 10416 0 1 80752
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0416_
timestamp 1486834041
transform -1 0 12992 0 -1 79184
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0417_
timestamp 1486834041
transform -1 0 12432 0 1 79184
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0418_
timestamp 1486834041
transform -1 0 12096 0 -1 79184
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0419_
timestamp 1486834041
transform 1 0 13888 0 1 79184
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0420_
timestamp 1486834041
transform -1 0 14112 0 -1 83888
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0421_
timestamp 1486834041
transform -1 0 16016 0 -1 82320
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0422_
timestamp 1486834041
transform -1 0 15456 0 -1 80752
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0423_
timestamp 1486834041
transform -1 0 23744 0 -1 87024
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0424_
timestamp 1486834041
transform -1 0 23184 0 -1 87024
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _0425_
timestamp 1486834041
transform 1 0 22736 0 1 85456
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0426_
timestamp 1486834041
transform 1 0 12768 0 -1 90160
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0427_
timestamp 1486834041
transform 1 0 12768 0 -1 91728
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0428_
timestamp 1486834041
transform -1 0 14112 0 -1 93296
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0429_
timestamp 1486834041
transform 1 0 8848 0 1 99568
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0430_
timestamp 1486834041
transform 1 0 9744 0 -1 99568
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0431_
timestamp 1486834041
transform 1 0 8848 0 -1 102704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0432_
timestamp 1486834041
transform -1 0 4592 0 -1 108976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0433_
timestamp 1486834041
transform -1 0 4592 0 1 107408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0434_
timestamp 1486834041
transform -1 0 5936 0 -1 110544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0435_
timestamp 1486834041
transform 1 0 19264 0 -1 85456
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0436_
timestamp 1486834041
transform 1 0 20496 0 1 83888
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0437_
timestamp 1486834041
transform -1 0 20272 0 1 85456
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0438_
timestamp 1486834041
transform 1 0 14896 0 1 83888
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0439_
timestamp 1486834041
transform 1 0 15008 0 1 85456
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0440_
timestamp 1486834041
transform 1 0 18480 0 1 83888
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0441_
timestamp 1486834041
transform 1 0 10864 0 -1 94864
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0442_
timestamp 1486834041
transform 1 0 10304 0 -1 96432
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0443_
timestamp 1486834041
transform -1 0 14336 0 1 96432
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0444_
timestamp 1486834041
transform 1 0 3920 0 -1 98000
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0445_
timestamp 1486834041
transform 1 0 3584 0 -1 96432
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0446_
timestamp 1486834041
transform -1 0 6272 0 -1 93296
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0447_
timestamp 1486834041
transform 1 0 20160 0 -1 79184
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0448_
timestamp 1486834041
transform 1 0 20496 0 1 79184
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0449_
timestamp 1486834041
transform 1 0 20384 0 -1 77616
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0450_
timestamp 1486834041
transform 1 0 15568 0 1 90160
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0451_
timestamp 1486834041
transform 1 0 15456 0 1 91728
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0452_
timestamp 1486834041
transform -1 0 18816 0 1 88592
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0453_
timestamp 1486834041
transform 1 0 8736 0 -1 93296
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0454_
timestamp 1486834041
transform 1 0 8064 0 1 91728
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0455_
timestamp 1486834041
transform -1 0 10528 0 -1 94864
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0456_
timestamp 1486834041
transform 1 0 1680 0 -1 94864
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0457_
timestamp 1486834041
transform 1 0 896 0 -1 93296
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0458_
timestamp 1486834041
transform -1 0 2912 0 -1 90160
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0459_
timestamp 1486834041
transform 1 0 20496 0 1 91728
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0460_
timestamp 1486834041
transform 1 0 19600 0 -1 94864
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0461_
timestamp 1486834041
transform -1 0 26096 0 -1 93296
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0462_
timestamp 1486834041
transform 1 0 16576 0 -1 91728
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0463_
timestamp 1486834041
transform 1 0 15456 0 1 93296
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0464_
timestamp 1486834041
transform -1 0 20832 0 -1 90160
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0465_
timestamp 1486834041
transform 1 0 8400 0 1 93296
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0466_
timestamp 1486834041
transform 1 0 7952 0 1 94864
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0467_
timestamp 1486834041
transform -1 0 16128 0 -1 94864
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0468_
timestamp 1486834041
transform -1 0 4592 0 1 93296
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0469_
timestamp 1486834041
transform 1 0 896 0 1 94864
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0470_
timestamp 1486834041
transform -1 0 8176 0 -1 90160
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0471_
timestamp 1486834041
transform 1 0 20496 0 1 94864
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0472_
timestamp 1486834041
transform 1 0 19600 0 -1 93296
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0473_
timestamp 1486834041
transform -1 0 22960 0 1 90160
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0474_
timestamp 1486834041
transform 1 0 15008 0 1 98000
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0475_
timestamp 1486834041
transform 1 0 12656 0 1 21168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0476_
timestamp 1486834041
transform 1 0 11648 0 -1 50960
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0477_
timestamp 1486834041
transform 1 0 9184 0 -1 43120
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0478_
timestamp 1486834041
transform 1 0 19600 0 -1 22736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0479_
timestamp 1486834041
transform -1 0 8512 0 -1 27440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0480_
timestamp 1486834041
transform 1 0 13888 0 1 43120
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0481_
timestamp 1486834041
transform 1 0 10752 0 -1 39984
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0482_
timestamp 1486834041
transform 1 0 14112 0 1 36848
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0483_
timestamp 1486834041
transform 1 0 14000 0 1 27440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0484_
timestamp 1486834041
transform 1 0 11536 0 -1 21168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0485_
timestamp 1486834041
transform 1 0 11424 0 -1 19600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0486_
timestamp 1486834041
transform 1 0 16688 0 1 21168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0487_
timestamp 1486834041
transform 1 0 11088 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0488_
timestamp 1486834041
transform 1 0 8848 0 1 18032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0489_
timestamp 1486834041
transform 1 0 4928 0 -1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0490_
timestamp 1486834041
transform 1 0 19264 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0491_
timestamp 1486834041
transform -1 0 6608 0 -1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0492_
timestamp 1486834041
transform -1 0 5376 0 -1 25872
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0493_
timestamp 1486834041
transform 1 0 1008 0 1 27440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0494_
timestamp 1486834041
transform 1 0 6608 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0495_
timestamp 1486834041
transform -1 0 10304 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0496_
timestamp 1486834041
transform 1 0 1008 0 1 19600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0497_
timestamp 1486834041
transform -1 0 4592 0 1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0498_
timestamp 1486834041
transform 1 0 2912 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0499_
timestamp 1486834041
transform 1 0 2912 0 -1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0500_
timestamp 1486834041
transform 1 0 1792 0 -1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0501_
timestamp 1486834041
transform 1 0 1792 0 -1 19600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0502_
timestamp 1486834041
transform 1 0 6272 0 1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0503_
timestamp 1486834041
transform -1 0 10304 0 1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0504_
timestamp 1486834041
transform -1 0 4928 0 -1 21168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0505_
timestamp 1486834041
transform -1 0 4928 0 -1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0506_
timestamp 1486834041
transform -1 0 6608 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0507_
timestamp 1486834041
transform 1 0 17584 0 -1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0508_
timestamp 1486834041
transform 1 0 1344 0 -1 27440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0509_
timestamp 1486834041
transform 1 0 2576 0 -1 30576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0510_
timestamp 1486834041
transform 1 0 11424 0 -1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0511_
timestamp 1486834041
transform 1 0 20048 0 -1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0512_
timestamp 1486834041
transform 1 0 20496 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0513_
timestamp 1486834041
transform 1 0 4928 0 -1 55664
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0514_
timestamp 1486834041
transform 1 0 1008 0 1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0515_
timestamp 1486834041
transform 1 0 8848 0 1 55664
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0516_
timestamp 1486834041
transform -1 0 4928 0 -1 14896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0517_
timestamp 1486834041
transform 1 0 13440 0 1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0518_
timestamp 1486834041
transform 1 0 10864 0 -1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0519_
timestamp 1486834041
transform 1 0 20608 0 -1 14896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0520_
timestamp 1486834041
transform 1 0 18032 0 -1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0521_
timestamp 1486834041
transform 1 0 5600 0 1 54096
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0522_
timestamp 1486834041
transform 1 0 1792 0 -1 32144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0523_
timestamp 1486834041
transform 1 0 9968 0 -1 57232
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0524_
timestamp 1486834041
transform 1 0 4928 0 1 19600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0525_
timestamp 1486834041
transform 1 0 14672 0 1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0526_
timestamp 1486834041
transform -1 0 12096 0 1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0527_
timestamp 1486834041
transform 1 0 20608 0 1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0528_
timestamp 1486834041
transform 1 0 17584 0 -1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0529_
timestamp 1486834041
transform 1 0 4816 0 1 50960
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0530_
timestamp 1486834041
transform -1 0 4928 0 -1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0531_
timestamp 1486834041
transform 1 0 9408 0 -1 54096
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0532_
timestamp 1486834041
transform 1 0 4928 0 -1 14896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0533_
timestamp 1486834041
transform 1 0 12768 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0534_
timestamp 1486834041
transform 1 0 8176 0 1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0535_
timestamp 1486834041
transform -1 0 20272 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0536_
timestamp 1486834041
transform 1 0 6608 0 1 46256
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0537_
timestamp 1486834041
transform 1 0 3920 0 -1 50960
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0538_
timestamp 1486834041
transform 1 0 12768 0 -1 14896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0539_
timestamp 1486834041
transform 1 0 18816 0 -1 18032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0540_
timestamp 1486834041
transform 1 0 1344 0 -1 36848
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0541_
timestamp 1486834041
transform 1 0 4928 0 -1 21168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0542_
timestamp 1486834041
transform 1 0 11760 0 -1 16464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0543_
timestamp 1486834041
transform 1 0 16576 0 -1 14896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0544_
timestamp 1486834041
transform 1 0 2464 0 -1 33712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0545_
timestamp 1486834041
transform 1 0 7056 0 1 22736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0546_
timestamp 1486834041
transform 1 0 8288 0 1 14896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0547_
timestamp 1486834041
transform 1 0 19264 0 -1 24304
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0548_
timestamp 1486834041
transform -1 0 20720 0 -1 24304
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0549_
timestamp 1486834041
transform -1 0 20272 0 -1 19600
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0550_
timestamp 1486834041
transform 1 0 21056 0 -1 21168
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0551_
timestamp 1486834041
transform 1 0 15568 0 -1 22736
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0552_
timestamp 1486834041
transform -1 0 18480 0 1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0553_
timestamp 1486834041
transform -1 0 17248 0 -1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0554_
timestamp 1486834041
transform -1 0 16352 0 -1 21168
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0555_
timestamp 1486834041
transform 1 0 15568 0 -1 19600
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0556_
timestamp 1486834041
transform 1 0 17136 0 1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0557_
timestamp 1486834041
transform 1 0 16576 0 -1 22736
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0558_
timestamp 1486834041
transform 1 0 16576 0 1 22736
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0559_
timestamp 1486834041
transform -1 0 22960 0 -1 25872
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0560_
timestamp 1486834041
transform -1 0 21168 0 1 24304
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0561_
timestamp 1486834041
transform -1 0 21504 0 -1 27440
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0562_
timestamp 1486834041
transform -1 0 22400 0 1 24304
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0563_
timestamp 1486834041
transform 1 0 11760 0 -1 25872
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0564_
timestamp 1486834041
transform 1 0 11648 0 -1 30576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0565_
timestamp 1486834041
transform 1 0 14896 0 1 30576
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0566_
timestamp 1486834041
transform 1 0 9968 0 -1 52528
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0567_
timestamp 1486834041
transform 1 0 8848 0 1 50960
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0568_
timestamp 1486834041
transform 1 0 10640 0 1 52528
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0569_
timestamp 1486834041
transform 1 0 4704 0 -1 41552
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0570_
timestamp 1486834041
transform 1 0 4816 0 1 41552
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0571_
timestamp 1486834041
transform 1 0 8400 0 1 41552
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0572_
timestamp 1486834041
transform 1 0 17696 0 -1 43120
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0573_
timestamp 1486834041
transform 1 0 17920 0 -1 41552
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0574_
timestamp 1486834041
transform 1 0 17584 0 -1 46256
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0575_
timestamp 1486834041
transform 1 0 12768 0 -1 29008
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0576_
timestamp 1486834041
transform -1 0 16352 0 -1 27440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0577_
timestamp 1486834041
transform -1 0 18256 0 -1 27440
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0578_
timestamp 1486834041
transform 1 0 10192 0 -1 36848
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0579_
timestamp 1486834041
transform -1 0 12432 0 1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0580_
timestamp 1486834041
transform -1 0 14336 0 1 32144
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0581_
timestamp 1486834041
transform 1 0 2576 0 -1 49392
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0582_
timestamp 1486834041
transform 1 0 2128 0 -1 47824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0583_
timestamp 1486834041
transform -1 0 2576 0 -1 49392
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0584_
timestamp 1486834041
transform 1 0 20496 0 1 41552
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0585_
timestamp 1486834041
transform 1 0 20496 0 1 39984
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0586_
timestamp 1486834041
transform -1 0 20272 0 1 41552
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0587_
timestamp 1486834041
transform -1 0 18928 0 -1 38416
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0588_
timestamp 1486834041
transform 1 0 18816 0 -1 36848
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _0589_
timestamp 1486834041
transform 1 0 17024 0 -1 35280
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0590_
timestamp 1486834041
transform -1 0 16240 0 1 35280
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _0591_
timestamp 1486834041
transform 1 0 17920 0 -1 33712
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0592_
timestamp 1486834041
transform 1 0 19152 0 -1 33712
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0593_
timestamp 1486834041
transform 1 0 19488 0 -1 38416
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0594_
timestamp 1486834041
transform 1 0 16688 0 1 33712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0595_
timestamp 1486834041
transform -1 0 17584 0 -1 32144
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0596_
timestamp 1486834041
transform 1 0 18592 0 1 32144
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0597_
timestamp 1486834041
transform 1 0 16240 0 1 35280
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0598_
timestamp 1486834041
transform -1 0 17920 0 -1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0599_
timestamp 1486834041
transform -1 0 18480 0 -1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0600_
timestamp 1486834041
transform 1 0 19600 0 1 35280
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0601_
timestamp 1486834041
transform -1 0 21392 0 1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0602_
timestamp 1486834041
transform 1 0 29456 0 -1 33712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0603_
timestamp 1486834041
transform 1 0 8624 0 1 25872
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0604_
timestamp 1486834041
transform 1 0 8176 0 1 27440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0605_
timestamp 1486834041
transform -1 0 8736 0 1 24304
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0606_
timestamp 1486834041
transform -1 0 8512 0 -1 36848
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0607_
timestamp 1486834041
transform 1 0 4928 0 -1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0608_
timestamp 1486834041
transform -1 0 10416 0 -1 35280
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0609_
timestamp 1486834041
transform 1 0 1792 0 -1 44688
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0610_
timestamp 1486834041
transform 1 0 1008 0 1 43120
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0611_
timestamp 1486834041
transform -1 0 6496 0 1 46256
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0612_
timestamp 1486834041
transform 1 0 20832 0 1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0613_
timestamp 1486834041
transform 1 0 20608 0 -1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0614_
timestamp 1486834041
transform -1 0 26096 0 -1 35280
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0615_
timestamp 1486834041
transform 1 0 8736 0 -1 27440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0616_
timestamp 1486834041
transform 1 0 8736 0 -1 29008
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0617_
timestamp 1486834041
transform -1 0 12320 0 1 22736
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0618_
timestamp 1486834041
transform 1 0 6272 0 1 36848
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0619_
timestamp 1486834041
transform 1 0 5264 0 1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0620_
timestamp 1486834041
transform -1 0 8512 0 -1 39984
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0621_
timestamp 1486834041
transform 1 0 1792 0 -1 43120
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0622_
timestamp 1486834041
transform 1 0 1008 0 1 41552
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0623_
timestamp 1486834041
transform -1 0 6496 0 1 39984
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0624_
timestamp 1486834041
transform 1 0 20832 0 1 33712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0625_
timestamp 1486834041
transform 1 0 20608 0 -1 33712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0626_
timestamp 1486834041
transform -1 0 26096 0 1 33712
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0627_
timestamp 1486834041
transform 1 0 20720 0 1 66640
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0628_
timestamp 1486834041
transform 1 0 20944 0 1 69776
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0629_
timestamp 1486834041
transform 1 0 5600 0 1 101136
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0630_
timestamp 1486834041
transform 1 0 5824 0 -1 99568
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0631_
timestamp 1486834041
transform -1 0 14112 0 -1 105840
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0632_
timestamp 1486834041
transform -1 0 15120 0 -1 104272
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0633_
timestamp 1486834041
transform 1 0 16576 0 -1 99568
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0634_
timestamp 1486834041
transform 1 0 16912 0 1 99568
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0635_
timestamp 1486834041
transform 1 0 14112 0 -1 112112
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0636_
timestamp 1486834041
transform 1 0 15456 0 1 110544
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0637_
timestamp 1486834041
transform 1 0 11648 0 -1 112112
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0638_
timestamp 1486834041
transform 1 0 13216 0 1 110544
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0639_
timestamp 1486834041
transform 1 0 8848 0 -1 113680
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0640_
timestamp 1486834041
transform 1 0 10528 0 -1 110544
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0641_
timestamp 1486834041
transform 1 0 10528 0 -1 85456
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0642_
timestamp 1486834041
transform 1 0 12880 0 -1 88592
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0643_
timestamp 1486834041
transform 1 0 16800 0 1 102704
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0644_
timestamp 1486834041
transform 1 0 16240 0 1 104272
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0645_
timestamp 1486834041
transform 1 0 14112 0 -1 105840
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0646_
timestamp 1486834041
transform 1 0 13104 0 1 108976
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0647_
timestamp 1486834041
transform 1 0 6048 0 -1 113680
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0648_
timestamp 1486834041
transform 1 0 5936 0 1 107408
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0649_
timestamp 1486834041
transform 1 0 9184 0 -1 60368
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0650_
timestamp 1486834041
transform 1 0 10192 0 1 60368
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0651_
timestamp 1486834041
transform 1 0 18704 0 -1 58800
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0652_
timestamp 1486834041
transform 1 0 17360 0 1 60368
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0653_
timestamp 1486834041
transform 1 0 5040 0 1 105840
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0654_
timestamp 1486834041
transform 1 0 5376 0 -1 112112
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0655_
timestamp 1486834041
transform 1 0 13328 0 1 102704
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0656_
timestamp 1486834041
transform 1 0 10528 0 -1 102704
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0657_
timestamp 1486834041
transform 1 0 16576 0 -1 77616
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0658_
timestamp 1486834041
transform 1 0 15120 0 1 77616
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0659_
timestamp 1486834041
transform 1 0 17920 0 1 65072
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0660_
timestamp 1486834041
transform -1 0 19824 0 1 66640
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0661_
timestamp 1486834041
transform 1 0 896 0 -1 112112
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0662_
timestamp 1486834041
transform 1 0 2352 0 1 112112
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0663_
timestamp 1486834041
transform 1 0 12656 0 1 105840
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0664_
timestamp 1486834041
transform 1 0 7280 0 1 105840
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0665_
timestamp 1486834041
transform 1 0 15344 0 1 80752
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0666_
timestamp 1486834041
transform 1 0 14000 0 -1 79184
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0667_
timestamp 1486834041
transform 1 0 18816 0 -1 69776
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0668_
timestamp 1486834041
transform 1 0 17360 0 1 69776
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0669_
timestamp 1486834041
transform -1 0 18368 0 -1 113680
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0670_
timestamp 1486834041
transform 1 0 2240 0 -1 113680
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0671_
timestamp 1486834041
transform 1 0 13552 0 -1 101136
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0672_
timestamp 1486834041
transform -1 0 14896 0 1 99568
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0673_
timestamp 1486834041
transform 1 0 16576 0 -1 85456
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0674_
timestamp 1486834041
transform 1 0 14112 0 -1 83888
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0675_
timestamp 1486834041
transform -1 0 22624 0 -1 60368
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0676_
timestamp 1486834041
transform 1 0 17696 0 1 61936
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0677_
timestamp 1486834041
transform 1 0 3136 0 -1 112112
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0678_
timestamp 1486834041
transform -1 0 8848 0 1 112112
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0679_
timestamp 1486834041
transform 1 0 10640 0 -1 88592
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0680_
timestamp 1486834041
transform 1 0 9072 0 -1 87024
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0681_
timestamp 1486834041
transform -1 0 19600 0 1 77616
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0682_
timestamp 1486834041
transform 1 0 14112 0 -1 77616
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0683_
timestamp 1486834041
transform 1 0 20944 0 -1 88592
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0684_
timestamp 1486834041
transform 1 0 21168 0 1 88592
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0685_
timestamp 1486834041
transform 1 0 12096 0 -1 80752
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0686_
timestamp 1486834041
transform 1 0 12656 0 1 80752
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0687_
timestamp 1486834041
transform 1 0 7504 0 1 77616
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0688_
timestamp 1486834041
transform 1 0 9184 0 -1 80752
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0689_
timestamp 1486834041
transform 1 0 8736 0 -1 74480
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0690_
timestamp 1486834041
transform -1 0 11760 0 1 71344
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0691_
timestamp 1486834041
transform 1 0 12880 0 1 60368
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0692_
timestamp 1486834041
transform 1 0 14000 0 -1 60368
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0693_
timestamp 1486834041
transform 1 0 20832 0 -1 91728
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0694_
timestamp 1486834041
transform 1 0 19152 0 -1 96432
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0695_
timestamp 1486834041
transform 1 0 17360 0 -1 94864
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0696_
timestamp 1486834041
transform 1 0 1008 0 -1 102704
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0697_
timestamp 1486834041
transform 1 0 896 0 1 110544
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0698_
timestamp 1486834041
transform 1 0 896 0 1 108976
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0699_
timestamp 1486834041
transform 1 0 6272 0 -1 93296
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0700_
timestamp 1486834041
transform 1 0 4928 0 1 98000
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0701_
timestamp 1486834041
transform -1 0 10976 0 -1 98000
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0702_
timestamp 1486834041
transform 1 0 16800 0 -1 93296
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0703_
timestamp 1486834041
transform 1 0 13216 0 1 93296
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0704_
timestamp 1486834041
transform 1 0 13328 0 1 90160
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0705_
timestamp 1486834041
transform 1 0 21392 0 -1 96432
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0706_
timestamp 1486834041
transform -1 0 22736 0 1 96432
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0707_
timestamp 1486834041
transform 1 0 18032 0 1 94864
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0708_
timestamp 1486834041
transform -1 0 3248 0 -1 101136
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0709_
timestamp 1486834041
transform 1 0 896 0 1 104272
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0710_
timestamp 1486834041
transform 1 0 896 0 1 102704
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0711_
timestamp 1486834041
transform -1 0 11984 0 1 90160
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0712_
timestamp 1486834041
transform 1 0 7392 0 1 96432
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0713_
timestamp 1486834041
transform 1 0 7168 0 1 98000
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0714_
timestamp 1486834041
transform -1 0 19152 0 -1 90160
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0715_
timestamp 1486834041
transform 1 0 14112 0 -1 93296
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0716_
timestamp 1486834041
transform 1 0 13216 0 1 91728
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0717_
timestamp 1486834041
transform 1 0 10192 0 1 76048
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0718_
timestamp 1486834041
transform 1 0 12656 0 1 77616
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0719_
timestamp 1486834041
transform 1 0 8736 0 -1 79184
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0720_
timestamp 1486834041
transform 1 0 9744 0 1 77616
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0721_
timestamp 1486834041
transform 1 0 896 0 -1 87024
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0722_
timestamp 1486834041
transform 1 0 1568 0 -1 83888
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0723_
timestamp 1486834041
transform -1 0 22736 0 1 76048
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0724_
timestamp 1486834041
transform 1 0 21056 0 -1 74480
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0725_
timestamp 1486834041
transform 1 0 12208 0 -1 76048
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0726_
timestamp 1486834041
transform 1 0 10192 0 1 74480
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0727_
timestamp 1486834041
transform 1 0 5488 0 1 82320
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0728_
timestamp 1486834041
transform -1 0 7504 0 -1 85456
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0729_
timestamp 1486834041
transform 1 0 3136 0 -1 79184
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0730_
timestamp 1486834041
transform 1 0 1344 0 1 80752
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0731_
timestamp 1486834041
transform 1 0 18032 0 1 71344
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0732_
timestamp 1486834041
transform 1 0 16464 0 1 72912
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0733_
timestamp 1486834041
transform 1 0 15008 0 1 69776
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0734_
timestamp 1486834041
transform 1 0 13776 0 -1 69776
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0735_
timestamp 1486834041
transform 1 0 5936 0 -1 110544
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0736_
timestamp 1486834041
transform -1 0 8176 0 -1 107408
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0737_
timestamp 1486834041
transform 1 0 5600 0 -1 87024
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0738_
timestamp 1486834041
transform 1 0 5936 0 1 87024
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0739_
timestamp 1486834041
transform 1 0 16688 0 -1 76048
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0740_
timestamp 1486834041
transform 1 0 14112 0 -1 74480
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0741_
timestamp 1486834041
transform 1 0 10864 0 -1 72912
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0742_
timestamp 1486834041
transform 1 0 11088 0 -1 74480
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0743_
timestamp 1486834041
transform 1 0 5264 0 1 77616
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0744_
timestamp 1486834041
transform 1 0 6160 0 -1 79184
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0745_
timestamp 1486834041
transform -1 0 7616 0 1 79184
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0746_
timestamp 1486834041
transform 1 0 1344 0 -1 82320
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0747_
timestamp 1486834041
transform 1 0 20720 0 1 71344
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0748_
timestamp 1486834041
transform 1 0 18144 0 -1 72912
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0749_
timestamp 1486834041
transform 1 0 14112 0 -1 71344
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0750_
timestamp 1486834041
transform 1 0 13104 0 -1 72912
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0751_
timestamp 1486834041
transform -1 0 7616 0 1 69776
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0752_
timestamp 1486834041
transform 1 0 5488 0 -1 72912
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0753_
timestamp 1486834041
transform 1 0 896 0 1 79184
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0754_
timestamp 1486834041
transform 1 0 1568 0 1 76048
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0755_
timestamp 1486834041
transform 1 0 20832 0 -1 71344
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0756_
timestamp 1486834041
transform -1 0 23296 0 -1 69776
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0757_
timestamp 1486834041
transform -1 0 14896 0 1 68208
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0758_
timestamp 1486834041
transform 1 0 10192 0 1 68208
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0759_
timestamp 1486834041
transform 1 0 1456 0 1 87024
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0760_
timestamp 1486834041
transform -1 0 7504 0 1 85456
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0761_
timestamp 1486834041
transform 1 0 5376 0 -1 69776
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0762_
timestamp 1486834041
transform 1 0 2576 0 -1 68208
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0763_
timestamp 1486834041
transform 1 0 16576 0 -1 69776
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0764_
timestamp 1486834041
transform 1 0 15456 0 1 65072
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0765_
timestamp 1486834041
transform 1 0 13888 0 -1 66640
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0766_
timestamp 1486834041
transform 1 0 12656 0 1 65072
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0767_
timestamp 1486834041
transform 1 0 2352 0 1 88592
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0768_
timestamp 1486834041
transform 1 0 2352 0 1 85456
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0769_
timestamp 1486834041
transform 1 0 896 0 -1 98000
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0770_
timestamp 1486834041
transform -1 0 10976 0 -1 82320
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0771_
timestamp 1486834041
transform 1 0 17920 0 1 63504
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0772_
timestamp 1486834041
transform 1 0 16688 0 -1 63504
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0773_
timestamp 1486834041
transform 1 0 5488 0 -1 63504
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0774_
timestamp 1486834041
transform 1 0 2688 0 -1 61936
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0775_
timestamp 1486834041
transform -1 0 3136 0 -1 79184
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0776_
timestamp 1486834041
transform 1 0 1456 0 1 74480
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0777_
timestamp 1486834041
transform -1 0 3136 0 -1 60368
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0778_
timestamp 1486834041
transform 1 0 1568 0 1 63504
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0779_
timestamp 1486834041
transform 1 0 6272 0 1 63504
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0780_
timestamp 1486834041
transform 1 0 6272 0 -1 65072
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0781_
timestamp 1486834041
transform -1 0 11760 0 -1 71344
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0782_
timestamp 1486834041
transform -1 0 10976 0 -1 69776
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0783_
timestamp 1486834041
transform 1 0 896 0 1 69776
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0784_
timestamp 1486834041
transform 1 0 1568 0 1 68208
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0785_
timestamp 1486834041
transform 1 0 896 0 1 77616
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0786_
timestamp 1486834041
transform 1 0 1456 0 1 72912
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0787_
timestamp 1486834041
transform 1 0 5488 0 1 65072
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0788_
timestamp 1486834041
transform 1 0 2352 0 1 60368
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0789_
timestamp 1486834041
transform 1 0 4816 0 1 68208
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0790_
timestamp 1486834041
transform 1 0 2352 0 1 66640
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0791_
timestamp 1486834041
transform -1 0 3136 0 1 90160
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0792_
timestamp 1486834041
transform 1 0 896 0 -1 88592
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0793_
timestamp 1486834041
transform 1 0 896 0 -1 66640
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0794_
timestamp 1486834041
transform 1 0 1568 0 1 65072
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0795_
timestamp 1486834041
transform 1 0 9184 0 -1 68208
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0796_
timestamp 1486834041
transform 1 0 6608 0 1 66640
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0797_
timestamp 1486834041
transform 1 0 9296 0 1 66640
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0798_
timestamp 1486834041
transform 1 0 7056 0 1 68208
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0799_
timestamp 1486834041
transform -1 0 3136 0 1 91728
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0800_
timestamp 1486834041
transform 1 0 896 0 -1 91728
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0801_
timestamp 1486834041
transform -1 0 5376 0 -1 91728
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0802_
timestamp 1486834041
transform 1 0 1008 0 -1 96432
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0803_
timestamp 1486834041
transform 1 0 5488 0 -1 60368
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0804_
timestamp 1486834041
transform 1 0 3248 0 -1 60368
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0805_
timestamp 1486834041
transform 1 0 15120 0 1 60368
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0806_
timestamp 1486834041
transform 1 0 16576 0 1 58800
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0807_
timestamp 1486834041
transform 1 0 2352 0 1 71344
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0808_
timestamp 1486834041
transform 1 0 5712 0 1 74480
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0809_
timestamp 1486834041
transform 1 0 8512 0 1 63504
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0810_
timestamp 1486834041
transform 1 0 9184 0 -1 61936
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0811_
timestamp 1486834041
transform 1 0 13328 0 -1 58800
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0812_
timestamp 1486834041
transform 1 0 14336 0 1 58800
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0813_
timestamp 1486834041
transform -1 0 22736 0 1 77616
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0814_
timestamp 1486834041
transform 1 0 18032 0 -1 80752
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0815_
timestamp 1486834041
transform 1 0 20496 0 1 80752
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0816_
timestamp 1486834041
transform 1 0 3584 0 -1 99568
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0817_
timestamp 1486834041
transform 1 0 1904 0 -1 110544
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0818_
timestamp 1486834041
transform 1 0 1792 0 -1 104272
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0819_
timestamp 1486834041
transform -1 0 14896 0 1 94864
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0820_
timestamp 1486834041
transform 1 0 9632 0 1 96432
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0821_
timestamp 1486834041
transform 1 0 10976 0 -1 98000
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0822_
timestamp 1486834041
transform 1 0 15792 0 1 82320
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0823_
timestamp 1486834041
transform 1 0 12656 0 1 85456
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0824_
timestamp 1486834041
transform 1 0 12768 0 1 87024
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0825_
timestamp 1486834041
transform 1 0 13888 0 1 63504
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0826_
timestamp 1486834041
transform 1 0 12768 0 -1 65072
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0827_
timestamp 1486834041
transform 1 0 6272 0 -1 76048
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0828_
timestamp 1486834041
transform 1 0 5824 0 -1 77616
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0829_
timestamp 1486834041
transform 1 0 8176 0 1 80752
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0830_
timestamp 1486834041
transform 1 0 5936 0 1 80752
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0831_
timestamp 1486834041
transform 1 0 10192 0 1 82320
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0832_
timestamp 1486834041
transform -1 0 14896 0 1 82320
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0833_
timestamp 1486834041
transform -1 0 22736 0 1 87024
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0834_
timestamp 1486834041
transform 1 0 17696 0 -1 88592
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0835_
timestamp 1486834041
transform -1 0 13552 0 -1 107408
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0836_
timestamp 1486834041
transform -1 0 17136 0 1 105840
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0837_
timestamp 1486834041
transform -1 0 18816 0 -1 112112
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0838_
timestamp 1486834041
transform -1 0 19936 0 1 110544
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0839_
timestamp 1486834041
transform -1 0 7504 0 1 94864
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0840_
timestamp 1486834041
transform 1 0 1456 0 1 98000
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0841_
timestamp 1486834041
transform 1 0 20608 0 1 63504
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0842_
timestamp 1486834041
transform 1 0 19376 0 -1 65072
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0843_
timestamp 1486834041
transform 1 0 1792 0 -1 105840
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0844_
timestamp 1486834041
transform -1 0 18816 0 -1 108976
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0845_
timestamp 1486834041
transform 1 0 9744 0 1 102704
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0846_
timestamp 1486834041
transform 1 0 6272 0 -1 104272
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0847_
timestamp 1486834041
transform 1 0 12768 0 1 98000
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0848_
timestamp 1486834041
transform 1 0 14112 0 -1 98000
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0849_
timestamp 1486834041
transform -1 0 22736 0 1 85456
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0850_
timestamp 1486834041
transform 1 0 18032 0 1 87024
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0851_
timestamp 1486834041
transform 1 0 20160 0 -1 83888
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0852_
timestamp 1486834041
transform -1 0 17136 0 1 112112
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0853_
timestamp 1486834041
transform -1 0 14560 0 -1 113680
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0854_
timestamp 1486834041
transform -1 0 14896 0 1 112112
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0855_
timestamp 1486834041
transform -1 0 12320 0 -1 104272
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0856_
timestamp 1486834041
transform 1 0 6272 0 -1 105840
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0857_
timestamp 1486834041
transform 1 0 9408 0 1 98000
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0858_
timestamp 1486834041
transform 1 0 6272 0 -1 91728
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0859_
timestamp 1486834041
transform 1 0 10192 0 -1 91728
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0860_
timestamp 1486834041
transform 1 0 12656 0 1 88592
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0861_
timestamp 1486834041
transform 1 0 9296 0 1 88592
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0862_
timestamp 1486834041
transform 1 0 9296 0 -1 90160
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0863_
timestamp 1486834041
transform 1 0 5152 0 1 96432
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0864_
timestamp 1486834041
transform 1 0 4816 0 1 99568
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0865_
timestamp 1486834041
transform 1 0 5376 0 1 93296
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0866_
timestamp 1486834041
transform -1 0 7504 0 -1 94864
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0867_
timestamp 1486834041
transform 1 0 7952 0 1 82320
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0868_
timestamp 1486834041
transform 1 0 5040 0 1 83888
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0869_
timestamp 1486834041
transform 1 0 3360 0 -1 87024
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0870_
timestamp 1486834041
transform 1 0 5824 0 1 91728
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0871_
timestamp 1486834041
transform -1 0 11088 0 1 112112
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0872_
timestamp 1486834041
transform -1 0 18816 0 -1 107408
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0873_
timestamp 1486834041
transform -1 0 21056 0 -1 112112
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0874_
timestamp 1486834041
transform -1 0 22176 0 -1 113680
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0875_
timestamp 1486834041
transform 1 0 2352 0 1 96432
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0876_
timestamp 1486834041
transform 1 0 1232 0 -1 99568
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0877_
timestamp 1486834041
transform -1 0 23632 0 -1 82320
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0878_
timestamp 1486834041
transform 1 0 19152 0 -1 82320
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0879_
timestamp 1486834041
transform -1 0 18816 0 -1 110544
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0880_
timestamp 1486834041
transform -1 0 19376 0 1 112112
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0881_
timestamp 1486834041
transform 1 0 4032 0 -1 104272
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0882_
timestamp 1486834041
transform 1 0 4032 0 -1 105840
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0883_
timestamp 1486834041
transform 1 0 14000 0 -1 99568
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0884_
timestamp 1486834041
transform -1 0 18816 0 -1 98000
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0885_
timestamp 1486834041
transform 1 0 20608 0 1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0886_
timestamp 1486834041
transform 1 0 20832 0 -1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0887_
timestamp 1486834041
transform 1 0 6272 0 -1 46256
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0888_
timestamp 1486834041
transform 1 0 6272 0 -1 44688
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0889_
timestamp 1486834041
transform 1 0 11872 0 -1 49392
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0890_
timestamp 1486834041
transform -1 0 14896 0 1 46256
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0891_
timestamp 1486834041
transform 1 0 12880 0 1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0892_
timestamp 1486834041
transform 1 0 12656 0 1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0893_
timestamp 1486834041
transform -1 0 18816 0 -1 50960
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0894_
timestamp 1486834041
transform 1 0 14000 0 1 47824
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0895_
timestamp 1486834041
transform 1 0 14112 0 1 52528
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0896_
timestamp 1486834041
transform 1 0 13328 0 -1 55664
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0897_
timestamp 1486834041
transform 1 0 6272 0 -1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0898_
timestamp 1486834041
transform 1 0 6272 0 -1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0899_
timestamp 1486834041
transform 1 0 9856 0 1 784
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0900_
timestamp 1486834041
transform 1 0 12320 0 1 784
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0901_
timestamp 1486834041
transform 1 0 14000 0 -1 47824
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0902_
timestamp 1486834041
transform 1 0 16240 0 1 47824
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0903_
timestamp 1486834041
transform 1 0 10528 0 -1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0904_
timestamp 1486834041
transform -1 0 15792 0 -1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0905_
timestamp 1486834041
transform 1 0 6272 0 -1 49392
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0906_
timestamp 1486834041
transform 1 0 2576 0 -1 52528
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0907_
timestamp 1486834041
transform -1 0 22736 0 1 2352
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0908_
timestamp 1486834041
transform -1 0 22176 0 1 784
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0909_
timestamp 1486834041
transform 1 0 21056 0 -1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0910_
timestamp 1486834041
transform 1 0 18032 0 1 7056
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0911_
timestamp 1486834041
transform 1 0 4032 0 -1 46256
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0912_
timestamp 1486834041
transform 1 0 4928 0 1 43120
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0913_
timestamp 1486834041
transform 1 0 10192 0 1 44688
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0914_
timestamp 1486834041
transform -1 0 12432 0 1 46256
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0915_
timestamp 1486834041
transform -1 0 18816 0 -1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0916_
timestamp 1486834041
transform 1 0 13104 0 -1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0917_
timestamp 1486834041
transform 1 0 20496 0 1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0918_
timestamp 1486834041
transform 1 0 18816 0 -1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0919_
timestamp 1486834041
transform 1 0 2688 0 -1 55664
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0920_
timestamp 1486834041
transform 1 0 1792 0 1 54096
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0921_
timestamp 1486834041
transform 1 0 9296 0 -1 58800
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0922_
timestamp 1486834041
transform 1 0 7952 0 1 58800
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0923_
timestamp 1486834041
transform 1 0 13328 0 1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0924_
timestamp 1486834041
transform 1 0 10192 0 1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0925_
timestamp 1486834041
transform 1 0 20832 0 1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0926_
timestamp 1486834041
transform -1 0 22736 0 1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0927_
timestamp 1486834041
transform 1 0 5488 0 1 55664
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0928_
timestamp 1486834041
transform 1 0 4032 0 -1 57232
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0929_
timestamp 1486834041
transform 1 0 9968 0 1 57232
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0930_
timestamp 1486834041
transform 1 0 7728 0 1 57232
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0931_
timestamp 1486834041
transform 1 0 13664 0 1 3920
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0932_
timestamp 1486834041
transform 1 0 13328 0 1 2352
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0933_
timestamp 1486834041
transform -1 0 23520 0 -1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0934_
timestamp 1486834041
transform -1 0 23408 0 -1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0935_
timestamp 1486834041
transform 1 0 2352 0 1 52528
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0936_
timestamp 1486834041
transform 1 0 2688 0 -1 54096
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0937_
timestamp 1486834041
transform 1 0 9072 0 -1 55664
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0938_
timestamp 1486834041
transform 1 0 6272 0 -1 57232
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0939_
timestamp 1486834041
transform 1 0 10528 0 -1 7056
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0940_
timestamp 1486834041
transform 1 0 11984 0 -1 2352
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0941_
timestamp 1486834041
transform 1 0 21280 0 -1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0942_
timestamp 1486834041
transform 1 0 20496 0 -1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0943_
timestamp 1486834041
transform 1 0 20608 0 1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0944_
timestamp 1486834041
transform 1 0 1344 0 1 39984
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0945_
timestamp 1486834041
transform 1 0 896 0 -1 39984
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0946_
timestamp 1486834041
transform 1 0 896 0 1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0947_
timestamp 1486834041
transform 1 0 5936 0 1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0948_
timestamp 1486834041
transform 1 0 5264 0 -1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0949_
timestamp 1486834041
transform 1 0 5264 0 1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0950_
timestamp 1486834041
transform 1 0 8736 0 -1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0951_
timestamp 1486834041
transform 1 0 5936 0 1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0952_
timestamp 1486834041
transform 1 0 7168 0 1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0953_
timestamp 1486834041
transform 1 0 19936 0 -1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0954_
timestamp 1486834041
transform -1 0 22736 0 1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0955_
timestamp 1486834041
transform 1 0 15232 0 1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0956_
timestamp 1486834041
transform 1 0 14896 0 1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0957_
timestamp 1486834041
transform 1 0 14112 0 -1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0958_
timestamp 1486834041
transform 1 0 16576 0 -1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0959_
timestamp 1486834041
transform 1 0 18032 0 1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0960_
timestamp 1486834041
transform 1 0 18816 0 -1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0961_
timestamp 1486834041
transform 1 0 21504 0 1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0962_
timestamp 1486834041
transform 1 0 20608 0 1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0963_
timestamp 1486834041
transform 1 0 20608 0 -1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0964_
timestamp 1486834041
transform 1 0 1120 0 -1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0965_
timestamp 1486834041
transform 1 0 896 0 -1 46256
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0966_
timestamp 1486834041
transform 1 0 896 0 1 44688
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0967_
timestamp 1486834041
transform 1 0 6048 0 1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0968_
timestamp 1486834041
transform 1 0 2352 0 1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0969_
timestamp 1486834041
transform -1 0 8288 0 -1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0970_
timestamp 1486834041
transform -1 0 10976 0 1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0971_
timestamp 1486834041
transform 1 0 6384 0 1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0972_
timestamp 1486834041
transform 1 0 6272 0 -1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0973_
timestamp 1486834041
transform 1 0 18368 0 -1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0974_
timestamp 1486834041
transform 1 0 17696 0 1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0975_
timestamp 1486834041
transform 1 0 17360 0 1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0976_
timestamp 1486834041
transform -1 0 18816 0 -1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0977_
timestamp 1486834041
transform 1 0 20496 0 -1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0978_
timestamp 1486834041
transform 1 0 18032 0 -1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0979_
timestamp 1486834041
transform 1 0 18032 0 1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0980_
timestamp 1486834041
transform -1 0 19488 0 -1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0981_
timestamp 1486834041
transform 1 0 5936 0 1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0982_
timestamp 1486834041
transform 1 0 8736 0 -1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0983_
timestamp 1486834041
transform 1 0 5824 0 -1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0984_
timestamp 1486834041
transform 1 0 6272 0 1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0985_
timestamp 1486834041
transform 1 0 896 0 1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0986_
timestamp 1486834041
transform -1 0 7056 0 1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0987_
timestamp 1486834041
transform 1 0 15568 0 1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0988_
timestamp 1486834041
transform 1 0 16240 0 1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0989_
timestamp 1486834041
transform 1 0 10528 0 -1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0990_
timestamp 1486834041
transform 1 0 9968 0 -1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0991_
timestamp 1486834041
transform 1 0 5152 0 -1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0992_
timestamp 1486834041
transform 1 0 3584 0 -1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0993_
timestamp 1486834041
transform -1 0 4368 0 1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0994_
timestamp 1486834041
transform -1 0 3136 0 1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0995_
timestamp 1486834041
transform 1 0 19040 0 -1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0996_
timestamp 1486834041
transform 1 0 17808 0 1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0997_
timestamp 1486834041
transform 1 0 13104 0 1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0998_
timestamp 1486834041
transform 1 0 12208 0 -1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _0999_
timestamp 1486834041
transform 1 0 2352 0 1 50960
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1000_
timestamp 1486834041
transform 1 0 1680 0 -1 50960
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1001_
timestamp 1486834041
transform 1 0 6384 0 1 47824
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1002_
timestamp 1486834041
transform 1 0 5712 0 -1 47824
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1003_
timestamp 1486834041
transform 1 0 16800 0 -1 5488
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1004_
timestamp 1486834041
transform 1 0 15904 0 1 3920
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1005_
timestamp 1486834041
transform 1 0 8176 0 1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1006_
timestamp 1486834041
transform 1 0 5936 0 1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1007_
timestamp 1486834041
transform 1 0 4032 0 -1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1008_
timestamp 1486834041
transform 1 0 5376 0 -1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1009_
timestamp 1486834041
transform -1 0 7616 0 -1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1010_
timestamp 1486834041
transform 1 0 1344 0 -1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1011_
timestamp 1486834041
transform 1 0 17808 0 1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1012_
timestamp 1486834041
transform 1 0 16352 0 1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1013_
timestamp 1486834041
transform 1 0 8736 0 -1 5488
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1014_
timestamp 1486834041
transform -1 0 14896 0 1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1015_
timestamp 1486834041
transform -1 0 7056 0 1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1016_
timestamp 1486834041
transform 1 0 5040 0 1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1017_
timestamp 1486834041
transform 1 0 896 0 1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1018_
timestamp 1486834041
transform -1 0 7056 0 1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1019_
timestamp 1486834041
transform 1 0 17808 0 -1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1020_
timestamp 1486834041
transform 1 0 16576 0 1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1021_
timestamp 1486834041
transform 1 0 10640 0 -1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1022_
timestamp 1486834041
transform 1 0 9184 0 -1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1023_
timestamp 1486834041
transform -1 0 11984 0 1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1024_
timestamp 1486834041
transform 1 0 1904 0 1 5488
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1025_
timestamp 1486834041
transform -1 0 3136 0 1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1026_
timestamp 1486834041
transform 1 0 1232 0 1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1027_
timestamp 1486834041
transform 1 0 20496 0 1 3920
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1028_
timestamp 1486834041
transform -1 0 22736 0 1 5488
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1029_
timestamp 1486834041
transform 1 0 10192 0 1 7056
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1030_
timestamp 1486834041
transform 1 0 6272 0 -1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1031_
timestamp 1486834041
transform 1 0 1008 0 1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1032_
timestamp 1486834041
transform 1 0 2352 0 1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1033_
timestamp 1486834041
transform -1 0 3136 0 1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1034_
timestamp 1486834041
transform 1 0 1792 0 -1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1035_
timestamp 1486834041
transform 1 0 17360 0 -1 2352
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1036_
timestamp 1486834041
transform 1 0 16240 0 1 2352
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1037_
timestamp 1486834041
transform -1 0 24976 0 1 5488
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1038_
timestamp 1486834041
transform 1 0 24976 0 1 5488
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1039_
timestamp 1486834041
transform -1 0 25984 0 1 784
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1040_
timestamp 1486834041
transform 1 0 1456 0 1 784
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1041_
timestamp 1486834041
transform -1 0 5376 0 -1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1042_
timestamp 1486834041
transform 1 0 1456 0 1 7056
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1043_
timestamp 1486834041
transform 1 0 3024 0 -1 2352
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1044_
timestamp 1486834041
transform -1 0 14896 0 1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1045_
timestamp 1486834041
transform 1 0 2352 0 1 3920
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1046_
timestamp 1486834041
transform 1 0 4928 0 1 2352
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1047_
timestamp 1486834041
transform 1 0 896 0 1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1048_
timestamp 1486834041
transform 1 0 1456 0 1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1049_
timestamp 1486834041
transform 1 0 896 0 1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1050_
timestamp 1486834041
transform 1 0 1344 0 -1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1051_
timestamp 1486834041
transform -1 0 14896 0 1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1052_
timestamp 1486834041
transform -1 0 24976 0 1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1053_
timestamp 1486834041
transform -1 0 19264 0 1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1054_
timestamp 1486834041
transform -1 0 22736 0 1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1055_
timestamp 1486834041
transform -1 0 26656 0 -1 2352
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1056_
timestamp 1486834041
transform 1 0 1456 0 1 2352
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1057_
timestamp 1486834041
transform -1 0 3136 0 -1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1058_
timestamp 1486834041
transform 1 0 896 0 -1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1059_
timestamp 1486834041
transform -1 0 23408 0 -1 3920
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1060_
timestamp 1486834041
transform -1 0 24976 0 1 3920
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1061_
timestamp 1486834041
transform 1 0 6048 0 1 784
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1062_
timestamp 1486834041
transform 1 0 5264 0 -1 2352
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1063_
timestamp 1486834041
transform -1 0 3136 0 -1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1064_
timestamp 1486834041
transform 1 0 1344 0 1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1065_
timestamp 1486834041
transform -1 0 6272 0 -1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1066_
timestamp 1486834041
transform -1 0 7728 0 1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1067_
timestamp 1486834041
transform -1 0 24080 0 -1 2352
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1068_
timestamp 1486834041
transform -1 0 24976 0 1 2352
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1069_
timestamp 1486834041
transform 1 0 17472 0 1 784
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1070_
timestamp 1486834041
transform 1 0 19600 0 -1 2352
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1071_
timestamp 1486834041
transform 1 0 2352 0 1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1072_
timestamp 1486834041
transform 1 0 5264 0 1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1073_
timestamp 1486834041
transform 1 0 7504 0 1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1074_
timestamp 1486834041
transform 1 0 8736 0 -1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1075_
timestamp 1486834041
transform 1 0 9744 0 -1 2352
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1076_
timestamp 1486834041
transform 1 0 8960 0 -1 3920
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1077_
timestamp 1486834041
transform -1 0 23744 0 -1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1078_
timestamp 1486834041
transform 1 0 19376 0 -1 46256
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1079_
timestamp 1486834041
transform -1 0 23520 0 -1 43120
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1080_
timestamp 1486834041
transform -1 0 4144 0 1 47824
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1081_
timestamp 1486834041
transform 1 0 1232 0 1 49392
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1082_
timestamp 1486834041
transform 1 0 1232 0 1 46256
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1083_
timestamp 1486834041
transform 1 0 10864 0 -1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1084_
timestamp 1486834041
transform 1 0 9856 0 1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1085_
timestamp 1486834041
transform -1 0 11872 0 1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1086_
timestamp 1486834041
transform 1 0 14224 0 1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1087_
timestamp 1486834041
transform 1 0 10192 0 1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1088_
timestamp 1486834041
transform 1 0 12656 0 1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1089_
timestamp 1486834041
transform -1 0 18816 0 -1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1090_
timestamp 1486834041
transform 1 0 17248 0 -1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1091_
timestamp 1486834041
transform 1 0 11088 0 -1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1092_
timestamp 1486834041
transform 1 0 9184 0 -1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1093_
timestamp 1486834041
transform 1 0 9296 0 -1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1094_
timestamp 1486834041
transform 1 0 10080 0 -1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1095_
timestamp 1486834041
transform 1 0 12656 0 1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1096_
timestamp 1486834041
transform 1 0 14000 0 1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1097_
timestamp 1486834041
transform 1 0 13104 0 1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1098_
timestamp 1486834041
transform 1 0 14112 0 -1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1099_
timestamp 1486834041
transform 1 0 7952 0 1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1100_
timestamp 1486834041
transform 1 0 10192 0 1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1101_
timestamp 1486834041
transform 1 0 14000 0 -1 44688
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1102_
timestamp 1486834041
transform 1 0 13104 0 1 44688
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1103_
timestamp 1486834041
transform 1 0 5488 0 -1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1104_
timestamp 1486834041
transform 1 0 4816 0 1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1105_
timestamp 1486834041
transform -1 0 22736 0 1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1106_
timestamp 1486834041
transform 1 0 18032 0 1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1107_
timestamp 1486834041
transform -1 0 12320 0 1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1108_
timestamp 1486834041
transform -1 0 10976 0 1 39984
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1109_
timestamp 1486834041
transform -1 0 15232 0 1 49392
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1110_
timestamp 1486834041
transform 1 0 10192 0 1 49392
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1111_
timestamp 1486834041
transform 1 0 11984 0 -1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1112_
timestamp 1486834041
transform 1 0 9744 0 -1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1113_
timestamp 1486834041
transform 1 0 17024 0 1 44688
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1114_
timestamp 1486834041
transform 1 0 16576 0 -1 44688
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1115_
timestamp 1486834041
transform 1 0 17472 0 1 43120
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1116_
timestamp 1486834041
transform 1 0 5376 0 -1 43120
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1117_
timestamp 1486834041
transform 1 0 2464 0 -1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1118_
timestamp 1486834041
transform 1 0 4592 0 -1 39984
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1119_
timestamp 1486834041
transform 1 0 10192 0 1 54096
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1120_
timestamp 1486834041
transform 1 0 6608 0 1 49392
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1121_
timestamp 1486834041
transform 1 0 9632 0 -1 49392
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1122_
timestamp 1486834041
transform 1 0 11200 0 -1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1123_
timestamp 1486834041
transform 1 0 10192 0 1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1124_
timestamp 1486834041
transform 1 0 9408 0 -1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1125_
timestamp 1486834041
transform 1 0 16128 0 1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1126_
timestamp 1486834041
transform 1 0 14112 0 -1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1127_
timestamp 1486834041
transform 1 0 12656 0 1 39984
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1128_
timestamp 1486834041
transform -1 0 15792 0 1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1129_
timestamp 1486834041
transform 1 0 7056 0 1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1130_
timestamp 1486834041
transform 1 0 8736 0 -1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1131_
timestamp 1486834041
transform 1 0 14448 0 1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1132_
timestamp 1486834041
transform 1 0 13888 0 -1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1133_
timestamp 1486834041
transform 1 0 11312 0 -1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1134_
timestamp 1486834041
transform 1 0 13552 0 -1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1135_
timestamp 1486834041
transform 1 0 6496 0 1 39984
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1136_
timestamp 1486834041
transform 1 0 9072 0 -1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1137_
timestamp 1486834041
transform 1 0 9632 0 1 43120
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1138_
timestamp 1486834041
transform 1 0 7392 0 1 43120
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1139_
timestamp 1486834041
transform 1 0 5376 0 -1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1140_
timestamp 1486834041
transform 1 0 4816 0 1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1141_
timestamp 1486834041
transform 1 0 19040 0 -1 44688
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1142_
timestamp 1486834041
transform -1 0 23520 0 -1 44688
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1143_
timestamp 1486834041
transform -1 0 11088 0 1 47824
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1144_
timestamp 1486834041
transform -1 0 11648 0 -1 50960
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1145_
timestamp 1486834041
transform -1 0 14896 0 1 55664
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1146_
timestamp 1486834041
transform -1 0 15792 0 -1 52528
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1147_
timestamp 1486834041
transform -1 0 17584 0 1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _1148_
timestamp 1486834041
transform 1 0 14112 0 -1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1149_
timestamp 1486834041
transform 1 0 23520 0 -1 36848
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1150_
timestamp 1486834041
transform 1 0 29344 0 1 77616
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1151_
timestamp 1486834041
transform 1 0 29344 0 1 79184
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1152_
timestamp 1486834041
transform 1 0 29344 0 -1 80752
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1153_
timestamp 1486834041
transform 1 0 29344 0 -1 82320
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1154_
timestamp 1486834041
transform 1 0 22400 0 1 82320
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1155_
timestamp 1486834041
transform 1 0 23184 0 -1 83888
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1156_
timestamp 1486834041
transform 1 0 23408 0 -1 85456
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1157_
timestamp 1486834041
transform 1 0 23968 0 1 85456
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1158_
timestamp 1486834041
transform 1 0 22736 0 1 87024
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1159_
timestamp 1486834041
transform 1 0 29344 0 -1 88592
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1160_
timestamp 1486834041
transform 1 0 12096 0 -1 90160
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1161_
timestamp 1486834041
transform 1 0 12656 0 1 90160
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1162_
timestamp 1486834041
transform 1 0 19040 0 1 91728
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1163_
timestamp 1486834041
transform 1 0 19040 0 1 93296
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1164_
timestamp 1486834041
transform 1 0 19376 0 1 96432
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1165_
timestamp 1486834041
transform 1 0 23184 0 -1 94864
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1166_
timestamp 1486834041
transform 1 0 29344 0 -1 96432
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1167_
timestamp 1486834041
transform 1 0 29344 0 -1 98000
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1168_
timestamp 1486834041
transform 1 0 18816 0 -1 99568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1169_
timestamp 1486834041
transform 1 0 17136 0 -1 101136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1170_
timestamp 1486834041
transform 1 0 29344 0 -1 101136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1171_
timestamp 1486834041
transform 1 0 17136 0 -1 102704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1172_
timestamp 1486834041
transform 1 0 19040 0 1 102704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1173_
timestamp 1486834041
transform 1 0 20384 0 -1 104272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1174_
timestamp 1486834041
transform 1 0 18928 0 -1 105840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1175_
timestamp 1486834041
transform 1 0 29344 0 1 105840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1176_
timestamp 1486834041
transform 1 0 15680 0 -1 108976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1177_
timestamp 1486834041
transform 1 0 29344 0 -1 108976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1178_
timestamp 1486834041
transform 1 0 29344 0 1 108976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1179_
timestamp 1486834041
transform 1 0 29344 0 1 110544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1180_
timestamp 1486834041
transform 1 0 23184 0 -1 112112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1181_
timestamp 1486834041
transform 1 0 24528 0 1 110544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1182_
timestamp 1486834041
transform 1 0 21504 0 -1 110544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1183_
timestamp 1486834041
transform 1 0 22176 0 -1 110544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1184_
timestamp 1486834041
transform 1 0 21504 0 -1 98000
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1185_
timestamp 1486834041
transform 1 0 21616 0 -1 105840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1186_
timestamp 1486834041
transform 1 0 23408 0 1 87024
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1187_
timestamp 1486834041
transform 1 0 22064 0 1 99568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1188_
timestamp 1486834041
transform 1 0 23184 0 1 110544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1189_
timestamp 1486834041
transform 1 0 23856 0 1 110544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1190_
timestamp 1486834041
transform 1 0 22736 0 1 108976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1191_
timestamp 1486834041
transform 1 0 23408 0 -1 110544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1192_
timestamp 1486834041
transform 1 0 24416 0 -1 112112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1193_
timestamp 1486834041
transform 1 0 26096 0 -1 112112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1194_
timestamp 1486834041
transform 1 0 24416 0 -1 110544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1195_
timestamp 1486834041
transform 1 0 25200 0 1 110544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1196_
timestamp 1486834041
transform 1 0 25088 0 -1 112112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1197_
timestamp 1486834041
transform 1 0 25088 0 -1 110544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1198_
timestamp 1486834041
transform 1 0 26320 0 1 110544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1199_
timestamp 1486834041
transform 1 0 26768 0 -1 112112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1200_
timestamp 1486834041
transform 1 0 26096 0 -1 110544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1201_
timestamp 1486834041
transform 1 0 26992 0 1 110544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1202_
timestamp 1486834041
transform 1 0 11760 0 1 110544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1203_
timestamp 1486834041
transform -1 0 10864 0 1 105840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1204_
timestamp 1486834041
transform 1 0 1120 0 -1 105840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1205_
timestamp 1486834041
transform -1 0 21504 0 -1 110544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1206_
timestamp 1486834041
transform -1 0 1680 0 -1 107408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1207_
timestamp 1486834041
transform 1 0 4816 0 1 102704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1208_
timestamp 1486834041
transform 1 0 3248 0 1 102704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1209_
timestamp 1486834041
transform -1 0 5936 0 1 108976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1210_
timestamp 1486834041
transform 1 0 1680 0 1 112112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1211_
timestamp 1486834041
transform -1 0 4592 0 1 104272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1212_
timestamp 1486834041
transform -1 0 5936 0 -1 107408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1213_
timestamp 1486834041
transform 1 0 5264 0 1 110544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1214_
timestamp 1486834041
transform -1 0 3920 0 1 108976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1215_
timestamp 1486834041
transform -1 0 6048 0 -1 113680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1216_
timestamp 1486834041
transform 1 0 4928 0 1 112112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1217_
timestamp 1486834041
transform 1 0 13216 0 1 107408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1218_
timestamp 1486834041
transform 1 0 10416 0 -1 112112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1219_
timestamp 1486834041
transform 1 0 3920 0 1 110544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1220_
timestamp 1486834041
transform 1 0 10752 0 1 110544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1221_
timestamp 1486834041
transform -1 0 19488 0 -1 110544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1222_
timestamp 1486834041
transform 1 0 9520 0 1 105840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1223_
timestamp 1486834041
transform 1 0 8176 0 1 107408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1224_
timestamp 1486834041
transform -1 0 11648 0 -1 105840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1225_
timestamp 1486834041
transform -1 0 10080 0 -1 108976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1226_
timestamp 1486834041
transform -1 0 10192 0 1 108976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1227_
timestamp 1486834041
transform -1 0 12096 0 -1 113680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1228_
timestamp 1486834041
transform -1 0 10528 0 -1 110544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1229_
timestamp 1486834041
transform -1 0 11760 0 1 112112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1230_
timestamp 1486834041
transform -1 0 10752 0 1 110544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1231_
timestamp 1486834041
transform 1 0 8736 0 -1 108976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1232_
timestamp 1486834041
transform 1 0 5600 0 1 112112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1233_
timestamp 1486834041
transform 1 0 15904 0 1 46256
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1234_
timestamp 1486834041
transform 1 0 13552 0 -1 107408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1235_
timestamp 1486834041
transform 1 0 8736 0 -1 110544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1236_
timestamp 1486834041
transform 1 0 10080 0 -1 108976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1237_
timestamp 1486834041
transform -1 0 21168 0 1 110544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1238_
timestamp 1486834041
transform 1 0 22400 0 -1 112112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1239_
timestamp 1486834041
transform -1 0 14448 0 1 57232
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1240_
timestamp 1486834041
transform -1 0 12096 0 -1 60368
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1241_
timestamp 1486834041
transform -1 0 2352 0 1 58800
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1242_
timestamp 1486834041
transform -1 0 17248 0 -1 58800
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1243_
timestamp 1486834041
transform -1 0 2352 0 1 60368
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1244_
timestamp 1486834041
transform -1 0 2352 0 -1 61936
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1245_
timestamp 1486834041
transform -1 0 1792 0 -1 63504
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1246_
timestamp 1486834041
transform -1 0 9744 0 1 61936
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1247_
timestamp 1486834041
transform -1 0 9408 0 -1 63504
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1248_
timestamp 1486834041
transform 1 0 1232 0 -1 65072
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1249_
timestamp 1486834041
transform -1 0 5488 0 1 63504
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1250_
timestamp 1486834041
transform -1 0 2352 0 -1 68208
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1251_
timestamp 1486834041
transform -1 0 5488 0 1 61936
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1252_
timestamp 1486834041
transform 1 0 3136 0 -1 66640
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1253_
timestamp 1486834041
transform -1 0 2352 0 1 66640
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1254_
timestamp 1486834041
transform -1 0 9968 0 1 68208
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1255_
timestamp 1486834041
transform -1 0 8512 0 -1 63504
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1256_
timestamp 1486834041
transform 1 0 3808 0 -1 66640
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1257_
timestamp 1486834041
transform -1 0 3808 0 1 69776
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1258_
timestamp 1486834041
transform 1 0 1008 0 1 66640
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1259_
timestamp 1486834041
transform -1 0 17248 0 -1 74480
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1260_
timestamp 1486834041
transform -1 0 8624 0 1 74480
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1261_
timestamp 1486834041
transform 1 0 1120 0 -1 104272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1262_
timestamp 1486834041
transform -1 0 15008 0 1 69776
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1263_
timestamp 1486834041
transform -1 0 17920 0 -1 72912
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1264_
timestamp 1486834041
transform 1 0 3136 0 1 77616
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1265_
timestamp 1486834041
transform 1 0 896 0 -1 83888
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1266_
timestamp 1486834041
transform -1 0 12208 0 -1 76048
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1267_
timestamp 1486834041
transform -1 0 20608 0 -1 76048
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1268_
timestamp 1486834041
transform 1 0 4816 0 1 82320
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1269_
timestamp 1486834041
transform -1 0 9744 0 -1 77616
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1270_
timestamp 1486834041
transform -1 0 14000 0 -1 77616
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1271_
timestamp 1486834041
transform -1 0 17920 0 1 63504
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1272_
timestamp 1486834041
transform -1 0 8288 0 1 69776
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1273_
timestamp 1486834041
transform 1 0 1680 0 -1 74480
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1274_
timestamp 1486834041
transform -1 0 14000 0 1 66640
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1275_
timestamp 1486834041
transform -1 0 16352 0 -1 68208
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1276_
timestamp 1486834041
transform 1 0 3808 0 1 69776
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1277_
timestamp 1486834041
transform -1 0 4368 0 1 72912
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1278_
timestamp 1486834041
transform -1 0 12432 0 -1 69776
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1279_
timestamp 1486834041
transform -1 0 20272 0 1 69776
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1280_
timestamp 1486834041
transform -1 0 5488 0 1 72912
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1281_
timestamp 1486834041
transform 1 0 3808 0 1 76048
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1282_
timestamp 1486834041
transform -1 0 14448 0 1 71344
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1283_
timestamp 1486834041
transform -1 0 21168 0 1 72912
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1284_
timestamp 1486834041
transform 1 0 3136 0 1 79184
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1285_
timestamp 1486834041
transform 1 0 4816 0 1 76048
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1286_
timestamp 1486834041
transform -1 0 12432 0 1 72912
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1287_
timestamp 1486834041
transform 1 0 29344 0 1 39984
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1288_
timestamp 1486834041
transform 1 0 29344 0 -1 41552
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1289_
timestamp 1486834041
transform 1 0 29344 0 1 41552
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1290_
timestamp 1486834041
transform 1 0 29344 0 1 43120
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1291_
timestamp 1486834041
transform 1 0 29344 0 -1 44688
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1292_
timestamp 1486834041
transform 1 0 29344 0 1 44688
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1293_
timestamp 1486834041
transform 1 0 22176 0 -1 46256
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1294_
timestamp 1486834041
transform 1 0 23072 0 1 46256
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1295_
timestamp 1486834041
transform 1 0 18480 0 1 47824
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1296_
timestamp 1486834041
transform 1 0 19264 0 -1 49392
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1297_
timestamp 1486834041
transform 1 0 16800 0 1 50960
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1298_
timestamp 1486834041
transform 1 0 16576 0 -1 52528
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1299_
timestamp 1486834041
transform 1 0 16352 0 1 52528
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1300_
timestamp 1486834041
transform 1 0 15120 0 -1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1301_
timestamp 1486834041
transform 1 0 21280 0 -1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1302_
timestamp 1486834041
transform 1 0 30016 0 -1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1303_
timestamp 1486834041
transform 1 0 20832 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1304_
timestamp 1486834041
transform 1 0 29344 0 1 57232
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1305_
timestamp 1486834041
transform 1 0 29344 0 -1 58800
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1306_
timestamp 1486834041
transform 1 0 29344 0 -1 60368
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1307_
timestamp 1486834041
transform 1 0 29344 0 1 60368
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1308_
timestamp 1486834041
transform 1 0 29344 0 -1 61936
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1309_
timestamp 1486834041
transform 1 0 29344 0 -1 63504
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1310_
timestamp 1486834041
transform 1 0 29344 0 1 63504
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1311_
timestamp 1486834041
transform 1 0 18592 0 -1 65072
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1312_
timestamp 1486834041
transform 1 0 20496 0 1 65072
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1313_
timestamp 1486834041
transform 1 0 29344 0 -1 68208
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1314_
timestamp 1486834041
transform 1 0 29344 0 1 68208
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1315_
timestamp 1486834041
transform 1 0 13104 0 1 57232
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1316_
timestamp 1486834041
transform 1 0 29344 0 -1 71344
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1317_
timestamp 1486834041
transform 1 0 22960 0 1 71344
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1318_
timestamp 1486834041
transform 1 0 22848 0 1 72912
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1319_
timestamp 1486834041
transform -1 0 13776 0 1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1320_
timestamp 1486834041
transform -1 0 12432 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1321_
timestamp 1486834041
transform 1 0 10416 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1322_
timestamp 1486834041
transform -1 0 19936 0 1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1323_
timestamp 1486834041
transform 1 0 11760 0 1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1324_
timestamp 1486834041
transform -1 0 13664 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1325_
timestamp 1486834041
transform -1 0 11760 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1326_
timestamp 1486834041
transform -1 0 15568 0 -1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1327_
timestamp 1486834041
transform -1 0 15568 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1328_
timestamp 1486834041
transform -1 0 14448 0 1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1329_
timestamp 1486834041
transform -1 0 13328 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1330_
timestamp 1486834041
transform -1 0 16352 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1331_
timestamp 1486834041
transform 1 0 15008 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1332_
timestamp 1486834041
transform 1 0 14560 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1333_
timestamp 1486834041
transform 1 0 15568 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1334_
timestamp 1486834041
transform 1 0 18144 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1335_
timestamp 1486834041
transform 1 0 14224 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1336_
timestamp 1486834041
transform 1 0 9856 0 -1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1337_
timestamp 1486834041
transform 1 0 15568 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1338_
timestamp 1486834041
transform 1 0 16576 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1339_
timestamp 1486834041
transform 1 0 20160 0 -1 110544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1340_
timestamp 1486834041
transform 1 0 21168 0 1 110544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1341_
timestamp 1486834041
transform 1 0 18928 0 1 108976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1342_
timestamp 1486834041
transform 1 0 21056 0 -1 112112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1343_
timestamp 1486834041
transform 1 0 19600 0 1 108976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1344_
timestamp 1486834041
transform 1 0 21840 0 1 110544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1345_
timestamp 1486834041
transform 1 0 21728 0 -1 112112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1346_
timestamp 1486834041
transform 1 0 22512 0 1 110544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1347_
timestamp 1486834041
transform 1 0 18032 0 1 82320
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1348_
timestamp 1486834041
transform 1 0 16688 0 -1 94864
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1349_
timestamp 1486834041
transform 1 0 18480 0 -1 96432
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1350_
timestamp 1486834041
transform 1 0 19712 0 -1 77616
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1351_
timestamp 1486834041
transform 1 0 18480 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1352_
timestamp 1486834041
transform 1 0 19488 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1353_
timestamp 1486834041
transform 1 0 23408 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1354_
timestamp 1486834041
transform 1 0 24416 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1355_
timestamp 1486834041
transform 1 0 7168 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1356_
timestamp 1486834041
transform 1 0 7840 0 -1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1357_
timestamp 1486834041
transform 1 0 4928 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1358_
timestamp 1486834041
transform -1 0 19488 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1359_
timestamp 1486834041
transform 1 0 11088 0 1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1360_
timestamp 1486834041
transform -1 0 13328 0 1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1361_
timestamp 1486834041
transform 1 0 8736 0 -1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1362_
timestamp 1486834041
transform 1 0 1680 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1363_
timestamp 1486834041
transform 1 0 12656 0 1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1364_
timestamp 1486834041
transform 1 0 1008 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1365_
timestamp 1486834041
transform 1 0 5600 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1366_
timestamp 1486834041
transform 1 0 7840 0 -1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1367_
timestamp 1486834041
transform 1 0 3696 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1368_
timestamp 1486834041
transform 1 0 3696 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1369_
timestamp 1486834041
transform 1 0 4816 0 1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1370_
timestamp 1486834041
transform -1 0 2912 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1371_
timestamp 1486834041
transform -1 0 7840 0 -1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1372_
timestamp 1486834041
transform 1 0 5488 0 1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1373_
timestamp 1486834041
transform 1 0 2240 0 -1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1374_
timestamp 1486834041
transform 1 0 5488 0 1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1375_
timestamp 1486834041
transform -1 0 16352 0 -1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1376_
timestamp 1486834041
transform 1 0 1456 0 -1 47824
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1377_
timestamp 1486834041
transform 1 0 1008 0 -1 50960
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1378_
timestamp 1486834041
transform -1 0 15568 0 1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1379_
timestamp 1486834041
transform -1 0 18816 0 -1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1380_
timestamp 1486834041
transform 1 0 1680 0 1 36848
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1381_
timestamp 1486834041
transform 1 0 1120 0 -1 19600
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1382_
timestamp 1486834041
transform -1 0 11760 0 -1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1383_
timestamp 1486834041
transform -1 0 17248 0 -1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1384_
timestamp 1486834041
transform -1 0 2352 0 -1 33712
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1385_
timestamp 1486834041
transform -1 0 8400 0 1 21168
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1386_
timestamp 1486834041
transform -1 0 8512 0 -1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1387_
timestamp 1486834041
transform -1 0 18928 0 1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1388_
timestamp 1486834041
transform -1 0 6160 0 1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1389_
timestamp 1486834041
transform -1 0 5488 0 1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1390_
timestamp 1486834041
transform -1 0 10864 0 -1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1391_
timestamp 1486834041
transform -1 0 20272 0 1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1392_
timestamp 1486834041
transform 1 0 1232 0 -1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1393_
timestamp 1486834041
transform -1 0 2352 0 -1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1394_
timestamp 1486834041
transform -1 0 10640 0 -1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1395_
timestamp 1486834041
transform -1 0 17584 0 -1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1396_
timestamp 1486834041
transform -1 0 3808 0 1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1397_
timestamp 1486834041
transform -1 0 4368 0 1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1398_
timestamp 1486834041
transform 1 0 1904 0 -1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1399_
timestamp 1486834041
transform -1 0 17920 0 -1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1400_
timestamp 1486834041
transform -1 0 4480 0 -1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1401_
timestamp 1486834041
transform -1 0 4592 0 1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1402_
timestamp 1486834041
transform -1 0 8288 0 1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_1
timestamp 1486834041
transform -1 0 10976 0 1 61936
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_2
timestamp 1486834041
transform -1 0 7728 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_3
timestamp 1486834041
transform 1 0 10752 0 1 63504
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_4
timestamp 1486834041
transform -1 0 11648 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_5
timestamp 1486834041
transform 1 0 12992 0 1 83888
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_6
timestamp 1486834041
transform -1 0 8736 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_7
timestamp 1486834041
transform 1 0 10752 0 1 108976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_8
timestamp 1486834041
transform 1 0 25200 0 1 108976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_9
timestamp 1486834041
transform -1 0 25424 0 1 112112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_10
timestamp 1486834041
transform -1 0 25312 0 -1 113680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_11
timestamp 1486834041
transform 1 0 25088 0 -1 108976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_12
timestamp 1486834041
transform 1 0 25088 0 1 107408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_13
timestamp 1486834041
transform 1 0 25088 0 -1 107408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_14
timestamp 1486834041
transform 1 0 25872 0 -1 110544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_15
timestamp 1486834041
transform -1 0 26096 0 -1 112112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_16
timestamp 1486834041
transform -1 0 23632 0 1 108976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_17
timestamp 1486834041
transform -1 0 6944 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_18
timestamp 1486834041
transform 1 0 14000 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_19
timestamp 1486834041
transform 1 0 15232 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_20
timestamp 1486834041
transform 1 0 6720 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_21
timestamp 1486834041
transform 1 0 8848 0 -1 107408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_22
timestamp 1486834041
transform 1 0 12768 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_23
timestamp 1486834041
transform 1 0 14560 0 -1 107408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_24
timestamp 1486834041
transform 1 0 16576 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_25
timestamp 1486834041
transform 1 0 16576 0 1 102704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_26
timestamp 1486834041
transform 1 0 8512 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_27
timestamp 1486834041
transform 1 0 10752 0 -1 107408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_28
timestamp 1486834041
transform 1 0 15232 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_29
timestamp 1486834041
transform 1 0 15344 0 -1 108976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_30
timestamp 1486834041
transform -1 0 11200 0 1 104272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_31
timestamp 1486834041
transform -1 0 11200 0 1 105840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_32
timestamp 1486834041
transform -1 0 9632 0 -1 107408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_33
timestamp 1486834041
transform -1 0 9632 0 -1 110544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_34
timestamp 1486834041
transform -1 0 9744 0 1 110544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_35
timestamp 1486834041
transform -1 0 9744 0 -1 112112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_36
timestamp 1486834041
transform -1 0 11648 0 -1 112112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_37
timestamp 1486834041
transform -1 0 11648 0 1 110544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_38
timestamp 1486834041
transform -1 0 10080 0 1 110544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_39
timestamp 1486834041
transform -1 0 10080 0 -1 112112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_40
timestamp 1486834041
transform -1 0 11312 0 -1 112112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_41
timestamp 1486834041
transform -1 0 11312 0 -1 113680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_42
timestamp 1486834041
transform -1 0 9744 0 -1 105840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_43
timestamp 1486834041
transform -1 0 9744 0 1 104272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_44
timestamp 1486834041
transform -1 0 8400 0 -1 107408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_45
timestamp 1486834041
transform -1 0 8400 0 -1 108976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_46
timestamp 1486834041
transform 1 0 26096 0 1 110544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_47
timestamp 1486834041
transform -1 0 26320 0 1 112112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_48
timestamp 1486834041
transform 1 0 11200 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_49
timestamp 1486834041
transform 1 0 12768 0 1 83888
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_50
timestamp 1486834041
transform 1 0 16576 0 -1 60368
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_51
timestamp 1486834041
transform 1 0 18928 0 1 58800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_52
timestamp 1486834041
transform 1 0 26768 0 -1 110544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_53
timestamp 1486834041
transform 1 0 26768 0 1 108976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_54
timestamp 1486834041
transform 1 0 26096 0 1 108976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_55
timestamp 1486834041
transform 1 0 26096 0 -1 108976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_56
timestamp 1486834041
transform 1 0 26992 0 -1 110544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_57
timestamp 1486834041
transform 1 0 26992 0 1 108976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_58
timestamp 1486834041
transform 1 0 23408 0 -1 108976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_59
timestamp 1486834041
transform 1 0 24416 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_60
timestamp 1486834041
transform 1 0 11312 0 1 83888
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_61
timestamp 1486834041
transform 1 0 7280 0 -1 88592
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_62
timestamp 1486834041
transform 1 0 25088 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_63
timestamp 1486834041
transform 1 0 26320 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_64
timestamp 1486834041
transform 1 0 26320 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_65
timestamp 1486834041
transform 1 0 30128 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_66
timestamp 1486834041
transform 1 0 18928 0 1 57232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_67
timestamp 1486834041
transform 1 0 18928 0 -1 57232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_68
timestamp 1486834041
transform 1 0 18928 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_69
timestamp 1486834041
transform 1 0 18928 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_70
timestamp 1486834041
transform 1 0 18928 0 -1 71344
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_Tile_X0Y1_UserCLK
timestamp 1486834041
transform 1 0 22512 0 1 74480
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_Tile_X0Y1_UserCLK
timestamp 1486834041
transform -1 0 30016 0 -1 55664
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_Tile_X0Y1_UserCLK
timestamp 1486834041
transform -1 0 28000 0 1 93296
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2
timestamp 1486834041
transform 1 0 896 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6
timestamp 1486834041
transform 1 0 1344 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33
timestamp 1486834041
transform 1 0 4368 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70
timestamp 1486834041
transform 1 0 8512 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74
timestamp 1486834041
transform 1 0 8960 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81
timestamp 1486834041
transform 1 0 9744 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_138
timestamp 1486834041
transform 1 0 16128 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_140
timestamp 1486834041
transform 1 0 16352 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_147
timestamp 1486834041
transform 1 0 17136 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_149
timestamp 1486834041
transform 1 0 17360 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_258
timestamp 1486834041
transform 1 0 29568 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_266
timestamp 1486834041
transform 1 0 30464 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_268
timestamp 1486834041
transform 1 0 30688 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_2
timestamp 1486834041
transform 1 0 896 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_63
timestamp 1486834041
transform 1 0 7728 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_72
timestamp 1486834041
transform 1 0 8736 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_74
timestamp 1486834041
transform 1 0 8960 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_139
timestamp 1486834041
transform 1 0 16240 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_142
timestamp 1486834041
transform 1 0 16576 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_209
timestamp 1486834041
transform 1 0 24080 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_250
timestamp 1486834041
transform 1 0 28672 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_266
timestamp 1486834041
transform 1 0 30464 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_268
timestamp 1486834041
transform 1 0 30688 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_2
timestamp 1486834041
transform 1 0 896 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_6
timestamp 1486834041
transform 1 0 1344 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_33
timestamp 1486834041
transform 1 0 4368 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_37
timestamp 1486834041
transform 1 0 4816 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_58
timestamp 1486834041
transform 1 0 7168 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_60
timestamp 1486834041
transform 1 0 7392 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_93
timestamp 1486834041
transform 1 0 11088 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_98
timestamp 1486834041
transform 1 0 11648 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_171
timestamp 1486834041
transform 1 0 19824 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_241
timestamp 1486834041
transform 1 0 27664 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_247
timestamp 1486834041
transform 1 0 28336 0 1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_263
timestamp 1486834041
transform 1 0 30128 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_267
timestamp 1486834041
transform 1 0 30576 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_20
timestamp 1486834041
transform 1 0 2912 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_53
timestamp 1486834041
transform 1 0 6608 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_57
timestamp 1486834041
transform 1 0 7056 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_72
timestamp 1486834041
transform 1 0 8736 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_126
timestamp 1486834041
transform 1 0 14784 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_148
timestamp 1486834041
transform 1 0 17248 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_150
timestamp 1486834041
transform 1 0 17472 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_209
timestamp 1486834041
transform 1 0 24080 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_236
timestamp 1486834041
transform 1 0 27104 0 -1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_268
timestamp 1486834041
transform 1 0 30688 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_14
timestamp 1486834041
transform 1 0 2240 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_37
timestamp 1486834041
transform 1 0 4816 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_50
timestamp 1486834041
transform 1 0 6272 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_86
timestamp 1486834041
transform 1 0 10304 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_107
timestamp 1486834041
transform 1 0 12656 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_109
timestamp 1486834041
transform 1 0 12880 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_174
timestamp 1486834041
transform 1 0 20160 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_223
timestamp 1486834041
transform 1 0 25648 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_227
timestamp 1486834041
transform 1 0 26096 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_231
timestamp 1486834041
transform 1 0 26544 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_239
timestamp 1486834041
transform 1 0 27440 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_243
timestamp 1486834041
transform 1 0 27888 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_247
timestamp 1486834041
transform 1 0 28336 0 1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_263
timestamp 1486834041
transform 1 0 30128 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_267
timestamp 1486834041
transform 1 0 30576 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_20
timestamp 1486834041
transform 1 0 2912 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_59
timestamp 1486834041
transform 1 0 7280 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_63
timestamp 1486834041
transform 1 0 7728 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_92
timestamp 1486834041
transform 1 0 10976 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_125
timestamp 1486834041
transform 1 0 14672 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_133
timestamp 1486834041
transform 1 0 15568 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_142
timestamp 1486834041
transform 1 0 16576 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_164
timestamp 1486834041
transform 1 0 19040 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_214
timestamp 1486834041
transform 1 0 24640 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_220
timestamp 1486834041
transform 1 0 25312 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_228
timestamp 1486834041
transform 1 0 26208 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_231
timestamp 1486834041
transform 1 0 26544 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_263
timestamp 1486834041
transform 1 0 30128 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_267
timestamp 1486834041
transform 1 0 30576 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_8
timestamp 1486834041
transform 1 0 1568 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_10
timestamp 1486834041
transform 1 0 1792 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_31
timestamp 1486834041
transform 1 0 4144 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_49
timestamp 1486834041
transform 1 0 6160 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_53
timestamp 1486834041
transform 1 0 6608 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_86
timestamp 1486834041
transform 1 0 10304 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_107
timestamp 1486834041
transform 1 0 12656 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_123
timestamp 1486834041
transform 1 0 14448 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_163
timestamp 1486834041
transform 1 0 18928 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_165
timestamp 1486834041
transform 1 0 19152 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_172
timestamp 1486834041
transform 1 0 19936 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_174
timestamp 1486834041
transform 1 0 20160 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_237
timestamp 1486834041
transform 1 0 27216 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_247
timestamp 1486834041
transform 1 0 28336 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_263
timestamp 1486834041
transform 1 0 30128 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_267
timestamp 1486834041
transform 1 0 30576 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_2
timestamp 1486834041
transform 1 0 896 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_4
timestamp 1486834041
transform 1 0 1120 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_17
timestamp 1486834041
transform 1 0 2576 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_19
timestamp 1486834041
transform 1 0 2800 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_78
timestamp 1486834041
transform 1 0 9408 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_142
timestamp 1486834041
transform 1 0 16576 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_207
timestamp 1486834041
transform 1 0 23856 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_209
timestamp 1486834041
transform 1 0 24080 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_212
timestamp 1486834041
transform 1 0 24416 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_244
timestamp 1486834041
transform 1 0 28000 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_260
timestamp 1486834041
transform 1 0 29792 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_268
timestamp 1486834041
transform 1 0 30688 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_2
timestamp 1486834041
transform 1 0 896 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_6
timestamp 1486834041
transform 1 0 1344 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_27
timestamp 1486834041
transform 1 0 3696 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_49
timestamp 1486834041
transform 1 0 6160 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_107
timestamp 1486834041
transform 1 0 12656 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_209
timestamp 1486834041
transform 1 0 24080 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_241
timestamp 1486834041
transform 1 0 27664 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_247
timestamp 1486834041
transform 1 0 28336 0 1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_263
timestamp 1486834041
transform 1 0 30128 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_267
timestamp 1486834041
transform 1 0 30576 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_8
timestamp 1486834041
transform 1 0 1568 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_15
timestamp 1486834041
transform 1 0 2352 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_19
timestamp 1486834041
transform 1 0 2800 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_72
timestamp 1486834041
transform 1 0 8736 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_202
timestamp 1486834041
transform 1 0 23296 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_212
timestamp 1486834041
transform 1 0 24416 0 -1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_244
timestamp 1486834041
transform 1 0 28000 0 -1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_260
timestamp 1486834041
transform 1 0 29792 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_268
timestamp 1486834041
transform 1 0 30688 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_14
timestamp 1486834041
transform 1 0 2240 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_49
timestamp 1486834041
transform 1 0 6160 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_82
timestamp 1486834041
transform 1 0 9856 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_84
timestamp 1486834041
transform 1 0 10080 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_113
timestamp 1486834041
transform 1 0 13328 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_166
timestamp 1486834041
transform 1 0 19264 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_168
timestamp 1486834041
transform 1 0 19488 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_217
timestamp 1486834041
transform 1 0 24976 0 1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_233
timestamp 1486834041
transform 1 0 26768 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_241
timestamp 1486834041
transform 1 0 27664 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_247
timestamp 1486834041
transform 1 0 28336 0 1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_263
timestamp 1486834041
transform 1 0 30128 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_267
timestamp 1486834041
transform 1 0 30576 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_22
timestamp 1486834041
transform 1 0 3136 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_84
timestamp 1486834041
transform 1 0 10080 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_135
timestamp 1486834041
transform 1 0 15792 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_139
timestamp 1486834041
transform 1 0 16240 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_148
timestamp 1486834041
transform 1 0 17248 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_152
timestamp 1486834041
transform 1 0 17696 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_205
timestamp 1486834041
transform 1 0 23632 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_209
timestamp 1486834041
transform 1 0 24080 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_212
timestamp 1486834041
transform 1 0 24416 0 -1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_244
timestamp 1486834041
transform 1 0 28000 0 -1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_260
timestamp 1486834041
transform 1 0 29792 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_268
timestamp 1486834041
transform 1 0 30688 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1486834041
transform 1 0 4480 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_37
timestamp 1486834041
transform 1 0 4816 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_67
timestamp 1486834041
transform 1 0 8176 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_69
timestamp 1486834041
transform 1 0 8400 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_102
timestamp 1486834041
transform 1 0 12096 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_104
timestamp 1486834041
transform 1 0 12320 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_139
timestamp 1486834041
transform 1 0 16240 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_141
timestamp 1486834041
transform 1 0 16464 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_162
timestamp 1486834041
transform 1 0 18816 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_170
timestamp 1486834041
transform 1 0 19712 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_174
timestamp 1486834041
transform 1 0 20160 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_197
timestamp 1486834041
transform 1 0 22736 0 1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_229
timestamp 1486834041
transform 1 0 26320 0 1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_247
timestamp 1486834041
transform 1 0 28336 0 1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_263
timestamp 1486834041
transform 1 0 30128 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_267
timestamp 1486834041
transform 1 0 30576 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_68
timestamp 1486834041
transform 1 0 8288 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_78
timestamp 1486834041
transform 1 0 9408 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_82
timestamp 1486834041
transform 1 0 9856 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_109
timestamp 1486834041
transform 1 0 12880 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_131
timestamp 1486834041
transform 1 0 15344 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_139
timestamp 1486834041
transform 1 0 16240 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_142
timestamp 1486834041
transform 1 0 16576 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_150
timestamp 1486834041
transform 1 0 17472 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_154
timestamp 1486834041
transform 1 0 17920 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_187
timestamp 1486834041
transform 1 0 21616 0 -1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_203
timestamp 1486834041
transform 1 0 23408 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_207
timestamp 1486834041
transform 1 0 23856 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_209
timestamp 1486834041
transform 1 0 24080 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_212
timestamp 1486834041
transform 1 0 24416 0 -1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_244
timestamp 1486834041
transform 1 0 28000 0 -1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_260
timestamp 1486834041
transform 1 0 29792 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_262
timestamp 1486834041
transform 1 0 30016 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_2
timestamp 1486834041
transform 1 0 896 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_6
timestamp 1486834041
transform 1 0 1344 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_33
timestamp 1486834041
transform 1 0 4368 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_43
timestamp 1486834041
transform 1 0 5488 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_127
timestamp 1486834041
transform 1 0 14896 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_135
timestamp 1486834041
transform 1 0 15792 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_139
timestamp 1486834041
transform 1 0 16240 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_160
timestamp 1486834041
transform 1 0 18592 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_168
timestamp 1486834041
transform 1 0 19488 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_172
timestamp 1486834041
transform 1 0 19936 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_174
timestamp 1486834041
transform 1 0 20160 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_197
timestamp 1486834041
transform 1 0 22736 0 1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_229
timestamp 1486834041
transform 1 0 26320 0 1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_247
timestamp 1486834041
transform 1 0 28336 0 1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_2
timestamp 1486834041
transform 1 0 896 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_78
timestamp 1486834041
transform 1 0 9408 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_82
timestamp 1486834041
transform 1 0 9856 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_123
timestamp 1486834041
transform 1 0 14448 0 -1 13328
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_139
timestamp 1486834041
transform 1 0 16240 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_142
timestamp 1486834041
transform 1 0 16576 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_144
timestamp 1486834041
transform 1 0 16800 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_203
timestamp 1486834041
transform 1 0 23408 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_207
timestamp 1486834041
transform 1 0 23856 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_209
timestamp 1486834041
transform 1 0 24080 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_212
timestamp 1486834041
transform 1 0 24416 0 -1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_244
timestamp 1486834041
transform 1 0 28000 0 -1 13328
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_260
timestamp 1486834041
transform 1 0 29792 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_262
timestamp 1486834041
transform 1 0 30016 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_2
timestamp 1486834041
transform 1 0 896 0 1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_43
timestamp 1486834041
transform 1 0 5488 0 1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_107
timestamp 1486834041
transform 1 0 12656 0 1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_131
timestamp 1486834041
transform 1 0 15344 0 1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_159
timestamp 1486834041
transform 1 0 18480 0 1 13328
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_177
timestamp 1486834041
transform 1 0 20496 0 1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_210
timestamp 1486834041
transform 1 0 24192 0 1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_242
timestamp 1486834041
transform 1 0 27776 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_244
timestamp 1486834041
transform 1 0 28000 0 1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_247
timestamp 1486834041
transform 1 0 28336 0 1 13328
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_265
timestamp 1486834041
transform 1 0 30352 0 1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_2
timestamp 1486834041
transform 1 0 896 0 -1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_84
timestamp 1486834041
transform 1 0 10080 0 -1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_174
timestamp 1486834041
transform 1 0 20160 0 -1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_17_212
timestamp 1486834041
transform 1 0 24416 0 -1 14896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_244
timestamp 1486834041
transform 1 0 28000 0 -1 14896
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_260
timestamp 1486834041
transform 1 0 29792 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_262
timestamp 1486834041
transform 1 0 30016 0 -1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_28
timestamp 1486834041
transform 1 0 3808 0 1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_57
timestamp 1486834041
transform 1 0 7056 0 1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_61
timestamp 1486834041
transform 1 0 7504 0 1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_100
timestamp 1486834041
transform 1 0 11872 0 1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_104
timestamp 1486834041
transform 1 0 12320 0 1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_173
timestamp 1486834041
transform 1 0 20048 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_177
timestamp 1486834041
transform 1 0 20496 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_179
timestamp 1486834041
transform 1 0 20720 0 1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_200
timestamp 1486834041
transform 1 0 23072 0 1 14896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_232
timestamp 1486834041
transform 1 0 26656 0 1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_240
timestamp 1486834041
transform 1 0 27552 0 1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_244
timestamp 1486834041
transform 1 0 28000 0 1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_247
timestamp 1486834041
transform 1 0 28336 0 1 14896
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_2
timestamp 1486834041
transform 1 0 896 0 -1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_26
timestamp 1486834041
transform 1 0 3584 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_60
timestamp 1486834041
transform 1 0 7392 0 -1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_92
timestamp 1486834041
transform 1 0 10976 0 -1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_131
timestamp 1486834041
transform 1 0 15344 0 -1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_139
timestamp 1486834041
transform 1 0 16240 0 -1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_154
timestamp 1486834041
transform 1 0 17920 0 -1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_162
timestamp 1486834041
transform 1 0 18816 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_204
timestamp 1486834041
transform 1 0 23520 0 -1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_208
timestamp 1486834041
transform 1 0 23968 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_19_212
timestamp 1486834041
transform 1 0 24416 0 -1 16464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_244
timestamp 1486834041
transform 1 0 28000 0 -1 16464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_260
timestamp 1486834041
transform 1 0 29792 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_262
timestamp 1486834041
transform 1 0 30016 0 -1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_34
timestamp 1486834041
transform 1 0 4480 0 1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_37
timestamp 1486834041
transform 1 0 4816 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_59
timestamp 1486834041
transform 1 0 7280 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_101
timestamp 1486834041
transform 1 0 11984 0 1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_127
timestamp 1486834041
transform 1 0 14896 0 1 16464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_143
timestamp 1486834041
transform 1 0 16688 0 1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_151
timestamp 1486834041
transform 1 0 17584 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_173
timestamp 1486834041
transform 1 0 20048 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_177
timestamp 1486834041
transform 1 0 20496 0 1 16464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_241
timestamp 1486834041
transform 1 0 27664 0 1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_247
timestamp 1486834041
transform 1 0 28336 0 1 16464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_22
timestamp 1486834041
transform 1 0 3136 0 -1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_66
timestamp 1486834041
transform 1 0 8064 0 -1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_92
timestamp 1486834041
transform 1 0 10976 0 -1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_113
timestamp 1486834041
transform 1 0 13328 0 -1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_148
timestamp 1486834041
transform 1 0 17248 0 -1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_194
timestamp 1486834041
transform 1 0 22400 0 -1 18032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_21_212
timestamp 1486834041
transform 1 0 24416 0 -1 18032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_244
timestamp 1486834041
transform 1 0 28000 0 -1 18032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_260
timestamp 1486834041
transform 1 0 29792 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_262
timestamp 1486834041
transform 1 0 30016 0 -1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_2
timestamp 1486834041
transform 1 0 896 0 1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_26
timestamp 1486834041
transform 1 0 3584 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_34
timestamp 1486834041
transform 1 0 4480 0 1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_49
timestamp 1486834041
transform 1 0 6160 0 1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_72
timestamp 1486834041
transform 1 0 8736 0 1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_159
timestamp 1486834041
transform 1 0 18480 0 1 18032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_177
timestamp 1486834041
transform 1 0 20496 0 1 18032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_241
timestamp 1486834041
transform 1 0 27664 0 1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_247
timestamp 1486834041
transform 1 0 28336 0 1 18032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_2
timestamp 1486834041
transform 1 0 896 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_48
timestamp 1486834041
transform 1 0 6048 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_72
timestamp 1486834041
transform 1 0 8736 0 -1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_132
timestamp 1486834041
transform 1 0 15456 0 -1 19600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_162
timestamp 1486834041
transform 1 0 18816 0 -1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_166
timestamp 1486834041
transform 1 0 19264 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_168
timestamp 1486834041
transform 1 0 19488 0 -1 19600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_23_175
timestamp 1486834041
transform 1 0 20272 0 -1 19600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_207
timestamp 1486834041
transform 1 0 23856 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_209
timestamp 1486834041
transform 1 0 24080 0 -1 19600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_23_212
timestamp 1486834041
transform 1 0 24416 0 -1 19600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_244
timestamp 1486834041
transform 1 0 28000 0 -1 19600
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_260
timestamp 1486834041
transform 1 0 29792 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_262
timestamp 1486834041
transform 1 0 30016 0 -1 19600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_2
timestamp 1486834041
transform 1 0 896 0 1 19600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_37
timestamp 1486834041
transform 1 0 4816 0 1 19600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_102
timestamp 1486834041
transform 1 0 12096 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_104
timestamp 1486834041
transform 1 0 12320 0 1 19600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_107
timestamp 1486834041
transform 1 0 12656 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_129
timestamp 1486834041
transform 1 0 15120 0 1 19600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_154
timestamp 1486834041
transform 1 0 17920 0 1 19600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_181
timestamp 1486834041
transform 1 0 20944 0 1 19600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_247
timestamp 1486834041
transform 1 0 28336 0 1 19600
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_263
timestamp 1486834041
transform 1 0 30128 0 1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_267
timestamp 1486834041
transform 1 0 30576 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_2
timestamp 1486834041
transform 1 0 896 0 -1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_72
timestamp 1486834041
transform 1 0 8736 0 -1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_76
timestamp 1486834041
transform 1 0 9184 0 -1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_193
timestamp 1486834041
transform 1 0 22288 0 -1 21168
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_209
timestamp 1486834041
transform 1 0 24080 0 -1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_25_212
timestamp 1486834041
transform 1 0 24416 0 -1 21168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_244
timestamp 1486834041
transform 1 0 28000 0 -1 21168
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_260
timestamp 1486834041
transform 1 0 29792 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_262
timestamp 1486834041
transform 1 0 30016 0 -1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_2
timestamp 1486834041
transform 1 0 896 0 1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_23
timestamp 1486834041
transform 1 0 3248 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_25
timestamp 1486834041
transform 1 0 3472 0 1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_32
timestamp 1486834041
transform 1 0 4256 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_34
timestamp 1486834041
transform 1 0 4480 0 1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_37
timestamp 1486834041
transform 1 0 4816 0 1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_41
timestamp 1486834041
transform 1 0 5264 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_69
timestamp 1486834041
transform 1 0 8400 0 1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_72
timestamp 1486834041
transform 1 0 8736 0 1 21168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_104
timestamp 1486834041
transform 1 0 12320 0 1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_177
timestamp 1486834041
transform 1 0 20496 0 1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_202
timestamp 1486834041
transform 1 0 23296 0 1 21168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_234
timestamp 1486834041
transform 1 0 26880 0 1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_242
timestamp 1486834041
transform 1 0 27776 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_244
timestamp 1486834041
transform 1 0 28000 0 1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_247
timestamp 1486834041
transform 1 0 28336 0 1 21168
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_2
timestamp 1486834041
transform 1 0 896 0 -1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_72
timestamp 1486834041
transform 1 0 8736 0 -1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_80
timestamp 1486834041
transform 1 0 9632 0 -1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_121
timestamp 1486834041
transform 1 0 14224 0 -1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_130
timestamp 1486834041
transform 1 0 15232 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_132
timestamp 1486834041
transform 1 0 15456 0 -1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_168
timestamp 1486834041
transform 1 0 19488 0 -1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_209
timestamp 1486834041
transform 1 0 24080 0 -1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_27_212
timestamp 1486834041
transform 1 0 24416 0 -1 22736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_244
timestamp 1486834041
transform 1 0 28000 0 -1 22736
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_260
timestamp 1486834041
transform 1 0 29792 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_262
timestamp 1486834041
transform 1 0 30016 0 -1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_14
timestamp 1486834041
transform 1 0 2240 0 1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_104
timestamp 1486834041
transform 1 0 12320 0 1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_107
timestamp 1486834041
transform 1 0 12656 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_109
timestamp 1486834041
transform 1 0 12880 0 1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_128
timestamp 1486834041
transform 1 0 15008 0 1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_139
timestamp 1486834041
transform 1 0 16240 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_141
timestamp 1486834041
transform 1 0 16464 0 1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_153
timestamp 1486834041
transform 1 0 17808 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_212
timestamp 1486834041
transform 1 0 24416 0 1 22736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_244
timestamp 1486834041
transform 1 0 28000 0 1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_247
timestamp 1486834041
transform 1 0 28336 0 1 22736
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_8
timestamp 1486834041
transform 1 0 1568 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_42
timestamp 1486834041
transform 1 0 5376 0 -1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_63
timestamp 1486834041
transform 1 0 7728 0 -1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_67
timestamp 1486834041
transform 1 0 8176 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_69
timestamp 1486834041
transform 1 0 8400 0 -1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_72
timestamp 1486834041
transform 1 0 8736 0 -1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_80
timestamp 1486834041
transform 1 0 9632 0 -1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_104
timestamp 1486834041
transform 1 0 12320 0 -1 24304
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_142
timestamp 1486834041
transform 1 0 16576 0 -1 24304
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_158
timestamp 1486834041
transform 1 0 18368 0 -1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_179
timestamp 1486834041
transform 1 0 20720 0 -1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_206
timestamp 1486834041
transform 1 0 23744 0 -1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_29_212
timestamp 1486834041
transform 1 0 24416 0 -1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_244
timestamp 1486834041
transform 1 0 28000 0 -1 24304
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_260
timestamp 1486834041
transform 1 0 29792 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_262
timestamp 1486834041
transform 1 0 30016 0 -1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_22
timestamp 1486834041
transform 1 0 3136 0 1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_30
timestamp 1486834041
transform 1 0 4032 0 1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_34
timestamp 1486834041
transform 1 0 4480 0 1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_92
timestamp 1486834041
transform 1 0 10976 0 1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_100
timestamp 1486834041
transform 1 0 11872 0 1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_104
timestamp 1486834041
transform 1 0 12320 0 1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_127
timestamp 1486834041
transform 1 0 14896 0 1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_151
timestamp 1486834041
transform 1 0 17584 0 1 24304
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_167
timestamp 1486834041
transform 1 0 19376 0 1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_194
timestamp 1486834041
transform 1 0 22400 0 1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_226
timestamp 1486834041
transform 1 0 25984 0 1 24304
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_242
timestamp 1486834041
transform 1 0 27776 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_244
timestamp 1486834041
transform 1 0 28000 0 1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_247
timestamp 1486834041
transform 1 0 28336 0 1 24304
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_2
timestamp 1486834041
transform 1 0 896 0 -1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_62
timestamp 1486834041
transform 1 0 7616 0 -1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_92
timestamp 1486834041
transform 1 0 10976 0 -1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_96
timestamp 1486834041
transform 1 0 11424 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_98
timestamp 1486834041
transform 1 0 11648 0 -1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_131
timestamp 1486834041
transform 1 0 15344 0 -1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_157
timestamp 1486834041
transform 1 0 18256 0 -1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_165
timestamp 1486834041
transform 1 0 19152 0 -1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_169
timestamp 1486834041
transform 1 0 19600 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_171
timestamp 1486834041
transform 1 0 19824 0 -1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_199
timestamp 1486834041
transform 1 0 22960 0 -1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_207
timestamp 1486834041
transform 1 0 23856 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_209
timestamp 1486834041
transform 1 0 24080 0 -1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_31_212
timestamp 1486834041
transform 1 0 24416 0 -1 25872
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_244
timestamp 1486834041
transform 1 0 28000 0 -1 25872
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_260
timestamp 1486834041
transform 1 0 29792 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_262
timestamp 1486834041
transform 1 0 30016 0 -1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_22
timestamp 1486834041
transform 1 0 3136 0 1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_30
timestamp 1486834041
transform 1 0 4032 0 1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_34
timestamp 1486834041
transform 1 0 4480 0 1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_37
timestamp 1486834041
transform 1 0 4816 0 1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_45
timestamp 1486834041
transform 1 0 5712 0 1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_49
timestamp 1486834041
transform 1 0 6160 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_103
timestamp 1486834041
transform 1 0 12208 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_107
timestamp 1486834041
transform 1 0 12656 0 1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_115
timestamp 1486834041
transform 1 0 13552 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_149
timestamp 1486834041
transform 1 0 17360 0 1 25872
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_165
timestamp 1486834041
transform 1 0 19152 0 1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_173
timestamp 1486834041
transform 1 0 20048 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_197
timestamp 1486834041
transform 1 0 22736 0 1 25872
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_229
timestamp 1486834041
transform 1 0 26320 0 1 25872
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_247
timestamp 1486834041
transform 1 0 28336 0 1 25872
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_263
timestamp 1486834041
transform 1 0 30128 0 1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_267
timestamp 1486834041
transform 1 0 30576 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_2
timestamp 1486834041
transform 1 0 896 0 -1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_104
timestamp 1486834041
transform 1 0 12320 0 -1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_157
timestamp 1486834041
transform 1 0 18256 0 -1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_172
timestamp 1486834041
transform 1 0 19936 0 -1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_190
timestamp 1486834041
transform 1 0 21952 0 -1 27440
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_206
timestamp 1486834041
transform 1 0 23744 0 -1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_33_212
timestamp 1486834041
transform 1 0 24416 0 -1 27440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_244
timestamp 1486834041
transform 1 0 28000 0 -1 27440
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_260
timestamp 1486834041
transform 1 0 29792 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_262
timestamp 1486834041
transform 1 0 30016 0 -1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_2
timestamp 1486834041
transform 1 0 896 0 1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_37
timestamp 1486834041
transform 1 0 4816 0 1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_45
timestamp 1486834041
transform 1 0 5712 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_99
timestamp 1486834041
transform 1 0 11760 0 1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_103
timestamp 1486834041
transform 1 0 12208 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_107
timestamp 1486834041
transform 1 0 12656 0 1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_115
timestamp 1486834041
transform 1 0 13552 0 1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_151
timestamp 1486834041
transform 1 0 17584 0 1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_192
timestamp 1486834041
transform 1 0 22176 0 1 27440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_224
timestamp 1486834041
transform 1 0 25760 0 1 27440
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_240
timestamp 1486834041
transform 1 0 27552 0 1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_244
timestamp 1486834041
transform 1 0 28000 0 1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_247
timestamp 1486834041
transform 1 0 28336 0 1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_255
timestamp 1486834041
transform 1 0 29232 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_261
timestamp 1486834041
transform 1 0 29904 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_2
timestamp 1486834041
transform 1 0 896 0 -1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_26
timestamp 1486834041
transform 1 0 3584 0 -1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_34
timestamp 1486834041
transform 1 0 4480 0 -1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_104
timestamp 1486834041
transform 1 0 12320 0 -1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_142
timestamp 1486834041
transform 1 0 16576 0 -1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_146
timestamp 1486834041
transform 1 0 17024 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_176
timestamp 1486834041
transform 1 0 20384 0 -1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_197
timestamp 1486834041
transform 1 0 22736 0 -1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_205
timestamp 1486834041
transform 1 0 23632 0 -1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_209
timestamp 1486834041
transform 1 0 24080 0 -1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_35_212
timestamp 1486834041
transform 1 0 24416 0 -1 29008
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_244
timestamp 1486834041
transform 1 0 28000 0 -1 29008
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_260
timestamp 1486834041
transform 1 0 29792 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_262
timestamp 1486834041
transform 1 0 30016 0 -1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_22
timestamp 1486834041
transform 1 0 3136 0 1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_30
timestamp 1486834041
transform 1 0 4032 0 1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_34
timestamp 1486834041
transform 1 0 4480 0 1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_57
timestamp 1486834041
transform 1 0 7056 0 1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_78
timestamp 1486834041
transform 1 0 9408 0 1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_82
timestamp 1486834041
transform 1 0 9856 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_84
timestamp 1486834041
transform 1 0 10080 0 1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_107
timestamp 1486834041
transform 1 0 12656 0 1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_115
timestamp 1486834041
transform 1 0 13552 0 1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_139
timestamp 1486834041
transform 1 0 16240 0 1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_197
timestamp 1486834041
transform 1 0 22736 0 1 29008
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_229
timestamp 1486834041
transform 1 0 26320 0 1 29008
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_247
timestamp 1486834041
transform 1 0 28336 0 1 29008
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_2
timestamp 1486834041
transform 1 0 896 0 -1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_10
timestamp 1486834041
transform 1 0 1792 0 -1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_14
timestamp 1486834041
transform 1 0 2240 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_16
timestamp 1486834041
transform 1 0 2464 0 -1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_49
timestamp 1486834041
transform 1 0 6160 0 -1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_72
timestamp 1486834041
transform 1 0 8736 0 -1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_76
timestamp 1486834041
transform 1 0 9184 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_130
timestamp 1486834041
transform 1 0 15232 0 -1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_134
timestamp 1486834041
transform 1 0 15680 0 -1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_142
timestamp 1486834041
transform 1 0 16576 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_144
timestamp 1486834041
transform 1 0 16800 0 -1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_188
timestamp 1486834041
transform 1 0 21728 0 -1 30576
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_204
timestamp 1486834041
transform 1 0 23520 0 -1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_208
timestamp 1486834041
transform 1 0 23968 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_212
timestamp 1486834041
transform 1 0 24416 0 -1 30576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_244
timestamp 1486834041
transform 1 0 28000 0 -1 30576
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_260
timestamp 1486834041
transform 1 0 29792 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_262
timestamp 1486834041
transform 1 0 30016 0 -1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_2
timestamp 1486834041
transform 1 0 896 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_4
timestamp 1486834041
transform 1 0 1120 0 1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_25
timestamp 1486834041
transform 1 0 3472 0 1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_33
timestamp 1486834041
transform 1 0 4368 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_77
timestamp 1486834041
transform 1 0 9296 0 1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_177
timestamp 1486834041
transform 1 0 20496 0 1 30576
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_241
timestamp 1486834041
transform 1 0 27664 0 1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_247
timestamp 1486834041
transform 1 0 28336 0 1 30576
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_2
timestamp 1486834041
transform 1 0 896 0 -1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_62
timestamp 1486834041
transform 1 0 7616 0 -1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_92
timestamp 1486834041
transform 1 0 10976 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_114
timestamp 1486834041
transform 1 0 13440 0 -1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_135
timestamp 1486834041
transform 1 0 15792 0 -1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_142
timestamp 1486834041
transform 1 0 16576 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_144
timestamp 1486834041
transform 1 0 16800 0 -1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_171
timestamp 1486834041
transform 1 0 19824 0 -1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_179
timestamp 1486834041
transform 1 0 20720 0 -1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_183
timestamp 1486834041
transform 1 0 21168 0 -1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_204
timestamp 1486834041
transform 1 0 23520 0 -1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_208
timestamp 1486834041
transform 1 0 23968 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_39_212
timestamp 1486834041
transform 1 0 24416 0 -1 32144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_244
timestamp 1486834041
transform 1 0 28000 0 -1 32144
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_260
timestamp 1486834041
transform 1 0 29792 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_262
timestamp 1486834041
transform 1 0 30016 0 -1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_22
timestamp 1486834041
transform 1 0 3136 0 1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_30
timestamp 1486834041
transform 1 0 4032 0 1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_34
timestamp 1486834041
transform 1 0 4480 0 1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_37
timestamp 1486834041
transform 1 0 4816 0 1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_45
timestamp 1486834041
transform 1 0 5712 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_47
timestamp 1486834041
transform 1 0 5936 0 1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_68
timestamp 1486834041
transform 1 0 8288 0 1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_76
timestamp 1486834041
transform 1 0 9184 0 1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_100
timestamp 1486834041
transform 1 0 11872 0 1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_104
timestamp 1486834041
transform 1 0 12320 0 1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_122
timestamp 1486834041
transform 1 0 14336 0 1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_126
timestamp 1486834041
transform 1 0 14784 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_170
timestamp 1486834041
transform 1 0 19712 0 1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_174
timestamp 1486834041
transform 1 0 20160 0 1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_185
timestamp 1486834041
transform 1 0 21392 0 1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_206
timestamp 1486834041
transform 1 0 23744 0 1 32144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_238
timestamp 1486834041
transform 1 0 27328 0 1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_242
timestamp 1486834041
transform 1 0 27776 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_244
timestamp 1486834041
transform 1 0 28000 0 1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_247
timestamp 1486834041
transform 1 0 28336 0 1 32144
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_263
timestamp 1486834041
transform 1 0 30128 0 1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_267
timestamp 1486834041
transform 1 0 30576 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_2
timestamp 1486834041
transform 1 0 896 0 -1 33712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_6
timestamp 1486834041
transform 1 0 1344 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_8
timestamp 1486834041
transform 1 0 1568 0 -1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_15
timestamp 1486834041
transform 1 0 2352 0 -1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_68
timestamp 1486834041
transform 1 0 8288 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_72
timestamp 1486834041
transform 1 0 8736 0 -1 33712
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_88
timestamp 1486834041
transform 1 0 10528 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_90
timestamp 1486834041
transform 1 0 10752 0 -1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_111
timestamp 1486834041
transform 1 0 13104 0 -1 33712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_115
timestamp 1486834041
transform 1 0 13552 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_117
timestamp 1486834041
transform 1 0 13776 0 -1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_138
timestamp 1486834041
transform 1 0 16128 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_176
timestamp 1486834041
transform 1 0 20384 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_41_212
timestamp 1486834041
transform 1 0 24416 0 -1 33712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_244
timestamp 1486834041
transform 1 0 28000 0 -1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_252
timestamp 1486834041
transform 1 0 28896 0 -1 33712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_256
timestamp 1486834041
transform 1 0 29344 0 -1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_261
timestamp 1486834041
transform 1 0 29904 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_2
timestamp 1486834041
transform 1 0 896 0 1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_10
timestamp 1486834041
transform 1 0 1792 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_12
timestamp 1486834041
transform 1 0 2016 0 1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_33
timestamp 1486834041
transform 1 0 4368 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_37
timestamp 1486834041
transform 1 0 4816 0 1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_45
timestamp 1486834041
transform 1 0 5712 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_67
timestamp 1486834041
transform 1 0 8176 0 1 33712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_103
timestamp 1486834041
transform 1 0 12208 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_107
timestamp 1486834041
transform 1 0 12656 0 1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_110
timestamp 1486834041
transform 1 0 12992 0 1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_118
timestamp 1486834041
transform 1 0 13888 0 1 33712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_122
timestamp 1486834041
transform 1 0 14336 0 1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_177
timestamp 1486834041
transform 1 0 20496 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_179
timestamp 1486834041
transform 1 0 20720 0 1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_227
timestamp 1486834041
transform 1 0 26096 0 1 33712
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_243
timestamp 1486834041
transform 1 0 27888 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_247
timestamp 1486834041
transform 1 0 28336 0 1 33712
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_2
timestamp 1486834041
transform 1 0 896 0 -1 35280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_87
timestamp 1486834041
transform 1 0 10416 0 -1 35280
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_43_227
timestamp 1486834041
transform 1 0 26096 0 -1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_259
timestamp 1486834041
transform 1 0 29680 0 -1 35280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_2
timestamp 1486834041
transform 1 0 896 0 1 35280
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_37
timestamp 1486834041
transform 1 0 4816 0 1 35280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_107
timestamp 1486834041
transform 1 0 12656 0 1 35280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_131
timestamp 1486834041
transform 1 0 15344 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_133
timestamp 1486834041
transform 1 0 15568 0 1 35280
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_177
timestamp 1486834041
transform 1 0 20496 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_179
timestamp 1486834041
transform 1 0 20720 0 1 35280
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_212
timestamp 1486834041
transform 1 0 24416 0 1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_244
timestamp 1486834041
transform 1 0 28000 0 1 35280
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_247
timestamp 1486834041
transform 1 0 28336 0 1 35280
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_2
timestamp 1486834041
transform 1 0 896 0 -1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_72
timestamp 1486834041
transform 1 0 8736 0 -1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_80
timestamp 1486834041
transform 1 0 9632 0 -1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_84
timestamp 1486834041
transform 1 0 10080 0 -1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_117
timestamp 1486834041
transform 1 0 13776 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_119
timestamp 1486834041
transform 1 0 14000 0 -1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_177
timestamp 1486834041
transform 1 0 20496 0 -1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_198
timestamp 1486834041
transform 1 0 22848 0 -1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_202
timestamp 1486834041
transform 1 0 23296 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_45_212
timestamp 1486834041
transform 1 0 24416 0 -1 36848
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_244
timestamp 1486834041
transform 1 0 28000 0 -1 36848
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_260
timestamp 1486834041
transform 1 0 29792 0 -1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_268
timestamp 1486834041
transform 1 0 30688 0 -1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_2
timestamp 1486834041
transform 1 0 896 0 1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_6
timestamp 1486834041
transform 1 0 1344 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_8
timestamp 1486834041
transform 1 0 1568 0 1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_37
timestamp 1486834041
transform 1 0 4816 0 1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_45
timestamp 1486834041
transform 1 0 5712 0 1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_49
timestamp 1486834041
transform 1 0 6160 0 1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_102
timestamp 1486834041
transform 1 0 12096 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_104
timestamp 1486834041
transform 1 0 12320 0 1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_107
timestamp 1486834041
transform 1 0 12656 0 1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_115
timestamp 1486834041
transform 1 0 13552 0 1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_119
timestamp 1486834041
transform 1 0 14000 0 1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_172
timestamp 1486834041
transform 1 0 19936 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_174
timestamp 1486834041
transform 1 0 20160 0 1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_177
timestamp 1486834041
transform 1 0 20496 0 1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_46_198
timestamp 1486834041
transform 1 0 22848 0 1 36848
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_230
timestamp 1486834041
transform 1 0 26432 0 1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_238
timestamp 1486834041
transform 1 0 27328 0 1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_242
timestamp 1486834041
transform 1 0 27776 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_244
timestamp 1486834041
transform 1 0 28000 0 1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_247
timestamp 1486834041
transform 1 0 28336 0 1 36848
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_263
timestamp 1486834041
transform 1 0 30128 0 1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_267
timestamp 1486834041
transform 1 0 30576 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_2
timestamp 1486834041
transform 1 0 896 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_24
timestamp 1486834041
transform 1 0 3360 0 -1 38416
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_40
timestamp 1486834041
transform 1 0 5152 0 -1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_61
timestamp 1486834041
transform 1 0 7504 0 -1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_69
timestamp 1486834041
transform 1 0 8400 0 -1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_72
timestamp 1486834041
transform 1 0 8736 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_74
timestamp 1486834041
transform 1 0 8960 0 -1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_135
timestamp 1486834041
transform 1 0 15792 0 -1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_139
timestamp 1486834041
transform 1 0 16240 0 -1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_142
timestamp 1486834041
transform 1 0 16576 0 -1 38416
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_167
timestamp 1486834041
transform 1 0 19376 0 -1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_175
timestamp 1486834041
transform 1 0 20272 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_197
timestamp 1486834041
transform 1 0 22736 0 -1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_205
timestamp 1486834041
transform 1 0 23632 0 -1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_209
timestamp 1486834041
transform 1 0 24080 0 -1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_212
timestamp 1486834041
transform 1 0 24416 0 -1 38416
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_244
timestamp 1486834041
transform 1 0 28000 0 -1 38416
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_260
timestamp 1486834041
transform 1 0 29792 0 -1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_268
timestamp 1486834041
transform 1 0 30688 0 -1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_22
timestamp 1486834041
transform 1 0 3136 0 1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_30
timestamp 1486834041
transform 1 0 4032 0 1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_34
timestamp 1486834041
transform 1 0 4480 0 1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_37
timestamp 1486834041
transform 1 0 4816 0 1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_61
timestamp 1486834041
transform 1 0 7504 0 1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_107
timestamp 1486834041
transform 1 0 12656 0 1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_147
timestamp 1486834041
transform 1 0 17136 0 1 38416
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_163
timestamp 1486834041
transform 1 0 18928 0 1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_171
timestamp 1486834041
transform 1 0 19824 0 1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_177
timestamp 1486834041
transform 1 0 20496 0 1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_48_198
timestamp 1486834041
transform 1 0 22848 0 1 38416
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_230
timestamp 1486834041
transform 1 0 26432 0 1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_238
timestamp 1486834041
transform 1 0 27328 0 1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_242
timestamp 1486834041
transform 1 0 27776 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_244
timestamp 1486834041
transform 1 0 28000 0 1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_247
timestamp 1486834041
transform 1 0 28336 0 1 38416
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_263
timestamp 1486834041
transform 1 0 30128 0 1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_267
timestamp 1486834041
transform 1 0 30576 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_22
timestamp 1486834041
transform 1 0 3136 0 -1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_30
timestamp 1486834041
transform 1 0 4032 0 -1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_34
timestamp 1486834041
transform 1 0 4480 0 -1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_72
timestamp 1486834041
transform 1 0 8736 0 -1 39984
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_88
timestamp 1486834041
transform 1 0 10528 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_122
timestamp 1486834041
transform 1 0 14336 0 -1 39984
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_138
timestamp 1486834041
transform 1 0 16128 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_142
timestamp 1486834041
transform 1 0 16576 0 -1 39984
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_206
timestamp 1486834041
transform 1 0 23744 0 -1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_49_212
timestamp 1486834041
transform 1 0 24416 0 -1 39984
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_244
timestamp 1486834041
transform 1 0 28000 0 -1 39984
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_260
timestamp 1486834041
transform 1 0 29792 0 -1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_268
timestamp 1486834041
transform 1 0 30688 0 -1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_2
timestamp 1486834041
transform 1 0 896 0 1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_26
timestamp 1486834041
transform 1 0 3584 0 1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_34
timestamp 1486834041
transform 1 0 4480 0 1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_92
timestamp 1486834041
transform 1 0 10976 0 1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_100
timestamp 1486834041
transform 1 0 11872 0 1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_104
timestamp 1486834041
transform 1 0 12320 0 1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_127
timestamp 1486834041
transform 1 0 14896 0 1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_135
timestamp 1486834041
transform 1 0 15792 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_169
timestamp 1486834041
transform 1 0 19600 0 1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_173
timestamp 1486834041
transform 1 0 20048 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_209
timestamp 1486834041
transform 1 0 24080 0 1 39984
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_241
timestamp 1486834041
transform 1 0 27664 0 1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_247
timestamp 1486834041
transform 1 0 28336 0 1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_255
timestamp 1486834041
transform 1 0 29232 0 1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_262
timestamp 1486834041
transform 1 0 30016 0 1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_2
timestamp 1486834041
transform 1 0 896 0 -1 41552
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_10
timestamp 1486834041
transform 1 0 1792 0 -1 41552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_14
timestamp 1486834041
transform 1 0 2240 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_68
timestamp 1486834041
transform 1 0 8288 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_72
timestamp 1486834041
transform 1 0 8736 0 -1 41552
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_80
timestamp 1486834041
transform 1 0 9632 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_114
timestamp 1486834041
transform 1 0 13440 0 -1 41552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_118
timestamp 1486834041
transform 1 0 13888 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_142
timestamp 1486834041
transform 1 0 16576 0 -1 41552
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_150
timestamp 1486834041
transform 1 0 17472 0 -1 41552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_206
timestamp 1486834041
transform 1 0 23744 0 -1 41552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_51_212
timestamp 1486834041
transform 1 0 24416 0 -1 41552
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_244
timestamp 1486834041
transform 1 0 28000 0 -1 41552
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_252
timestamp 1486834041
transform 1 0 28896 0 -1 41552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_262
timestamp 1486834041
transform 1 0 30016 0 -1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_2
timestamp 1486834041
transform 1 0 896 0 1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_104
timestamp 1486834041
transform 1 0 12320 0 1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_107
timestamp 1486834041
transform 1 0 12656 0 1 41552
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_135
timestamp 1486834041
transform 1 0 15792 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_137
timestamp 1486834041
transform 1 0 16016 0 1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_158
timestamp 1486834041
transform 1 0 18368 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_52_209
timestamp 1486834041
transform 1 0 24080 0 1 41552
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_241
timestamp 1486834041
transform 1 0 27664 0 1 41552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_247
timestamp 1486834041
transform 1 0 28336 0 1 41552
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_255
timestamp 1486834041
transform 1 0 29232 0 1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_262
timestamp 1486834041
transform 1 0 30016 0 1 41552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_266
timestamp 1486834041
transform 1 0 30464 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_268
timestamp 1486834041
transform 1 0 30688 0 1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_2
timestamp 1486834041
transform 1 0 896 0 -1 43120
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_62
timestamp 1486834041
transform 1 0 7616 0 -1 43120
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_72
timestamp 1486834041
transform 1 0 8736 0 -1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_142
timestamp 1486834041
transform 1 0 16576 0 -1 43120
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_150
timestamp 1486834041
transform 1 0 17472 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_204
timestamp 1486834041
transform 1 0 23520 0 -1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_208
timestamp 1486834041
transform 1 0 23968 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_53_212
timestamp 1486834041
transform 1 0 24416 0 -1 43120
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_244
timestamp 1486834041
transform 1 0 28000 0 -1 43120
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_260
timestamp 1486834041
transform 1 0 29792 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_262
timestamp 1486834041
transform 1 0 30016 0 -1 43120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_2
timestamp 1486834041
transform 1 0 896 0 1 43120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_37
timestamp 1486834041
transform 1 0 4816 0 1 43120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_58
timestamp 1486834041
transform 1 0 7168 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_100
timestamp 1486834041
transform 1 0 11872 0 1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_104
timestamp 1486834041
transform 1 0 12320 0 1 43120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_107
timestamp 1486834041
transform 1 0 12656 0 1 43120
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_115
timestamp 1486834041
transform 1 0 13552 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_117
timestamp 1486834041
transform 1 0 13776 0 1 43120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_170
timestamp 1486834041
transform 1 0 19712 0 1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_174
timestamp 1486834041
transform 1 0 20160 0 1 43120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_209
timestamp 1486834041
transform 1 0 24080 0 1 43120
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_241
timestamp 1486834041
transform 1 0 27664 0 1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_247
timestamp 1486834041
transform 1 0 28336 0 1 43120
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_255
timestamp 1486834041
transform 1 0 29232 0 1 43120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_262
timestamp 1486834041
transform 1 0 30016 0 1 43120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_2
timestamp 1486834041
transform 1 0 896 0 -1 44688
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_42
timestamp 1486834041
transform 1 0 5376 0 -1 44688
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_80
timestamp 1486834041
transform 1 0 9632 0 -1 44688
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_113
timestamp 1486834041
transform 1 0 13328 0 -1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_117
timestamp 1486834041
transform 1 0 13776 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_139
timestamp 1486834041
transform 1 0 16240 0 -1 44688
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_162
timestamp 1486834041
transform 1 0 18816 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_204
timestamp 1486834041
transform 1 0 23520 0 -1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_208
timestamp 1486834041
transform 1 0 23968 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_55_212
timestamp 1486834041
transform 1 0 24416 0 -1 44688
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_244
timestamp 1486834041
transform 1 0 28000 0 -1 44688
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_252
timestamp 1486834041
transform 1 0 28896 0 -1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_262
timestamp 1486834041
transform 1 0 30016 0 -1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_266
timestamp 1486834041
transform 1 0 30464 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_268
timestamp 1486834041
transform 1 0 30688 0 -1 44688
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_22
timestamp 1486834041
transform 1 0 3136 0 1 44688
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_30
timestamp 1486834041
transform 1 0 4032 0 1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_34
timestamp 1486834041
transform 1 0 4480 0 1 44688
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_37
timestamp 1486834041
transform 1 0 4816 0 1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_41
timestamp 1486834041
transform 1 0 5264 0 1 44688
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_107
timestamp 1486834041
transform 1 0 12656 0 1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_131
timestamp 1486834041
transform 1 0 15344 0 1 44688
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_139
timestamp 1486834041
transform 1 0 16240 0 1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_143
timestamp 1486834041
transform 1 0 16688 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_145
timestamp 1486834041
transform 1 0 16912 0 1 44688
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_166
timestamp 1486834041
transform 1 0 19264 0 1 44688
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_174
timestamp 1486834041
transform 1 0 20160 0 1 44688
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_177
timestamp 1486834041
transform 1 0 20496 0 1 44688
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_241
timestamp 1486834041
transform 1 0 27664 0 1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_247
timestamp 1486834041
transform 1 0 28336 0 1 44688
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_255
timestamp 1486834041
transform 1 0 29232 0 1 44688
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_262
timestamp 1486834041
transform 1 0 30016 0 1 44688
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_57_22
timestamp 1486834041
transform 1 0 3136 0 -1 46256
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_82
timestamp 1486834041
transform 1 0 9856 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_84
timestamp 1486834041
transform 1 0 10080 0 -1 46256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_57_117
timestamp 1486834041
transform 1 0 13776 0 -1 46256
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_133
timestamp 1486834041
transform 1 0 15568 0 -1 46256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_137
timestamp 1486834041
transform 1 0 16016 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_139
timestamp 1486834041
transform 1 0 16240 0 -1 46256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_57_142
timestamp 1486834041
transform 1 0 16576 0 -1 46256
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_150
timestamp 1486834041
transform 1 0 17472 0 -1 46256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_166
timestamp 1486834041
transform 1 0 19264 0 -1 46256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_187
timestamp 1486834041
transform 1 0 21616 0 -1 46256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_191
timestamp 1486834041
transform 1 0 22064 0 -1 46256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_57_198
timestamp 1486834041
transform 1 0 22848 0 -1 46256
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_206
timestamp 1486834041
transform 1 0 23744 0 -1 46256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_57_212
timestamp 1486834041
transform 1 0 24416 0 -1 46256
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_57_244
timestamp 1486834041
transform 1 0 28000 0 -1 46256
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_260
timestamp 1486834041
transform 1 0 29792 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_262
timestamp 1486834041
transform 1 0 30016 0 -1 46256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_2
timestamp 1486834041
transform 1 0 896 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_4
timestamp 1486834041
transform 1 0 1120 0 1 46256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_25
timestamp 1486834041
transform 1 0 3472 0 1 46256
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_33
timestamp 1486834041
transform 1 0 4368 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_52
timestamp 1486834041
transform 1 0 6496 0 1 46256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_127
timestamp 1486834041
transform 1 0 14896 0 1 46256
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_135
timestamp 1486834041
transform 1 0 15792 0 1 46256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_58_144
timestamp 1486834041
transform 1 0 16800 0 1 46256
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_160
timestamp 1486834041
transform 1 0 18592 0 1 46256
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_168
timestamp 1486834041
transform 1 0 19488 0 1 46256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_172
timestamp 1486834041
transform 1 0 19936 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_174
timestamp 1486834041
transform 1 0 20160 0 1 46256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_58_177
timestamp 1486834041
transform 1 0 20496 0 1 46256
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_193
timestamp 1486834041
transform 1 0 22288 0 1 46256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_197
timestamp 1486834041
transform 1 0 22736 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_199
timestamp 1486834041
transform 1 0 22960 0 1 46256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_58_206
timestamp 1486834041
transform 1 0 23744 0 1 46256
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_238
timestamp 1486834041
transform 1 0 27328 0 1 46256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_242
timestamp 1486834041
transform 1 0 27776 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_244
timestamp 1486834041
transform 1 0 28000 0 1 46256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_58_247
timestamp 1486834041
transform 1 0 28336 0 1 46256
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_263
timestamp 1486834041
transform 1 0 30128 0 1 46256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_267
timestamp 1486834041
transform 1 0 30576 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_2
timestamp 1486834041
transform 1 0 896 0 -1 47824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_6
timestamp 1486834041
transform 1 0 1344 0 -1 47824
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_69
timestamp 1486834041
transform 1 0 8400 0 -1 47824
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_72
timestamp 1486834041
transform 1 0 8736 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_74
timestamp 1486834041
transform 1 0 8960 0 -1 47824
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_107
timestamp 1486834041
transform 1 0 12656 0 -1 47824
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_116
timestamp 1486834041
transform 1 0 13664 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_118
timestamp 1486834041
transform 1 0 13888 0 -1 47824
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_139
timestamp 1486834041
transform 1 0 16240 0 -1 47824
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_59_174
timestamp 1486834041
transform 1 0 20160 0 -1 47824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_206
timestamp 1486834041
transform 1 0 23744 0 -1 47824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_59_212
timestamp 1486834041
transform 1 0 24416 0 -1 47824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_59_244
timestamp 1486834041
transform 1 0 28000 0 -1 47824
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_260
timestamp 1486834041
transform 1 0 29792 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_262
timestamp 1486834041
transform 1 0 30016 0 -1 47824
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_2
timestamp 1486834041
transform 1 0 896 0 1 47824
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_10
timestamp 1486834041
transform 1 0 1792 0 1 47824
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_31
timestamp 1486834041
transform 1 0 4144 0 1 47824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_37
timestamp 1486834041
transform 1 0 4816 0 1 47824
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_45
timestamp 1486834041
transform 1 0 5712 0 1 47824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_49
timestamp 1486834041
transform 1 0 6160 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_71
timestamp 1486834041
transform 1 0 8624 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_93
timestamp 1486834041
transform 1 0 11088 0 1 47824
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_107
timestamp 1486834041
transform 1 0 12656 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_165
timestamp 1486834041
transform 1 0 19152 0 1 47824
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_173
timestamp 1486834041
transform 1 0 20048 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_177
timestamp 1486834041
transform 1 0 20496 0 1 47824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_241
timestamp 1486834041
transform 1 0 27664 0 1 47824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_60_247
timestamp 1486834041
transform 1 0 28336 0 1 47824
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_49
timestamp 1486834041
transform 1 0 6160 0 -1 49392
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_72
timestamp 1486834041
transform 1 0 8736 0 -1 49392
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_120
timestamp 1486834041
transform 1 0 14112 0 -1 49392
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_128
timestamp 1486834041
transform 1 0 15008 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_132
timestamp 1486834041
transform 1 0 15456 0 -1 49392
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_61_142
timestamp 1486834041
transform 1 0 16576 0 -1 49392
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_158
timestamp 1486834041
transform 1 0 18368 0 -1 49392
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_61_172
timestamp 1486834041
transform 1 0 19936 0 -1 49392
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_204
timestamp 1486834041
transform 1 0 23520 0 -1 49392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_208
timestamp 1486834041
transform 1 0 23968 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_61_212
timestamp 1486834041
transform 1 0 24416 0 -1 49392
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_61_244
timestamp 1486834041
transform 1 0 28000 0 -1 49392
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_260
timestamp 1486834041
transform 1 0 29792 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_262
timestamp 1486834041
transform 1 0 30016 0 -1 49392
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_2
timestamp 1486834041
transform 1 0 896 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_4
timestamp 1486834041
transform 1 0 1120 0 1 49392
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_25
timestamp 1486834041
transform 1 0 3472 0 1 49392
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_33
timestamp 1486834041
transform 1 0 4368 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_62_37
timestamp 1486834041
transform 1 0 4816 0 1 49392
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_73
timestamp 1486834041
transform 1 0 8848 0 1 49392
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_107
timestamp 1486834041
transform 1 0 12656 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_109
timestamp 1486834041
transform 1 0 12880 0 1 49392
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_162
timestamp 1486834041
transform 1 0 18816 0 1 49392
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_170
timestamp 1486834041
transform 1 0 19712 0 1 49392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_174
timestamp 1486834041
transform 1 0 20160 0 1 49392
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_177
timestamp 1486834041
transform 1 0 20496 0 1 49392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_241
timestamp 1486834041
transform 1 0 27664 0 1 49392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_62_247
timestamp 1486834041
transform 1 0 28336 0 1 49392
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_263
timestamp 1486834041
transform 1 0 30128 0 1 49392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_267
timestamp 1486834041
transform 1 0 30576 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_2
timestamp 1486834041
transform 1 0 896 0 -1 50960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_61
timestamp 1486834041
transform 1 0 7504 0 -1 50960
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_69
timestamp 1486834041
transform 1 0 8400 0 -1 50960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_72
timestamp 1486834041
transform 1 0 8736 0 -1 50960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_76
timestamp 1486834041
transform 1 0 9184 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_132
timestamp 1486834041
transform 1 0 15456 0 -1 50960
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_63_162
timestamp 1486834041
transform 1 0 18816 0 -1 50960
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_63_194
timestamp 1486834041
transform 1 0 22400 0 -1 50960
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_63_212
timestamp 1486834041
transform 1 0 24416 0 -1 50960
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_63_244
timestamp 1486834041
transform 1 0 28000 0 -1 50960
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_260
timestamp 1486834041
transform 1 0 29792 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_262
timestamp 1486834041
transform 1 0 30016 0 -1 50960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_2
timestamp 1486834041
transform 1 0 896 0 1 50960
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_10
timestamp 1486834041
transform 1 0 1792 0 1 50960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_14
timestamp 1486834041
transform 1 0 2240 0 1 50960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_69
timestamp 1486834041
transform 1 0 8400 0 1 50960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_139
timestamp 1486834041
transform 1 0 16240 0 1 50960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_143
timestamp 1486834041
transform 1 0 16688 0 1 50960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_64_150
timestamp 1486834041
transform 1 0 17472 0 1 50960
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_166
timestamp 1486834041
transform 1 0 19264 0 1 50960
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_174
timestamp 1486834041
transform 1 0 20160 0 1 50960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_177
timestamp 1486834041
transform 1 0 20496 0 1 50960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_241
timestamp 1486834041
transform 1 0 27664 0 1 50960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_64_247
timestamp 1486834041
transform 1 0 28336 0 1 50960
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_2
timestamp 1486834041
transform 1 0 896 0 -1 52528
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_10
timestamp 1486834041
transform 1 0 1792 0 -1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_14
timestamp 1486834041
transform 1 0 2240 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_16
timestamp 1486834041
transform 1 0 2464 0 -1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_65_37
timestamp 1486834041
transform 1 0 4816 0 -1 52528
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_53
timestamp 1486834041
transform 1 0 6608 0 -1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_56
timestamp 1486834041
transform 1 0 6944 0 -1 52528
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_64
timestamp 1486834041
transform 1 0 7840 0 -1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_68
timestamp 1486834041
transform 1 0 8288 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_72
timestamp 1486834041
transform 1 0 8736 0 -1 52528
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_80
timestamp 1486834041
transform 1 0 9632 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_82
timestamp 1486834041
transform 1 0 9856 0 -1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_135
timestamp 1486834041
transform 1 0 15792 0 -1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_139
timestamp 1486834041
transform 1 0 16240 0 -1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_65_148
timestamp 1486834041
transform 1 0 17248 0 -1 52528
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_65_180
timestamp 1486834041
transform 1 0 20832 0 -1 52528
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_196
timestamp 1486834041
transform 1 0 22624 0 -1 52528
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_204
timestamp 1486834041
transform 1 0 23520 0 -1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_208
timestamp 1486834041
transform 1 0 23968 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_65_212
timestamp 1486834041
transform 1 0 24416 0 -1 52528
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_65_244
timestamp 1486834041
transform 1 0 28000 0 -1 52528
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_260
timestamp 1486834041
transform 1 0 29792 0 -1 52528
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_268
timestamp 1486834041
transform 1 0 30688 0 -1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_2
timestamp 1486834041
transform 1 0 896 0 1 52528
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_10
timestamp 1486834041
transform 1 0 1792 0 1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_14
timestamp 1486834041
transform 1 0 2240 0 1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_37
timestamp 1486834041
transform 1 0 4816 0 1 52528
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_53
timestamp 1486834041
transform 1 0 6608 0 1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_86
timestamp 1486834041
transform 1 0 10304 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_88
timestamp 1486834041
transform 1 0 10528 0 1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_104
timestamp 1486834041
transform 1 0 12320 0 1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_107
timestamp 1486834041
transform 1 0 12656 0 1 52528
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_115
timestamp 1486834041
transform 1 0 13552 0 1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_119
timestamp 1486834041
transform 1 0 14000 0 1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_146
timestamp 1486834041
transform 1 0 17024 0 1 52528
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_162
timestamp 1486834041
transform 1 0 18816 0 1 52528
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_170
timestamp 1486834041
transform 1 0 19712 0 1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_174
timestamp 1486834041
transform 1 0 20160 0 1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_177
timestamp 1486834041
transform 1 0 20496 0 1 52528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_241
timestamp 1486834041
transform 1 0 27664 0 1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_247
timestamp 1486834041
transform 1 0 28336 0 1 52528
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_2
timestamp 1486834041
transform 1 0 896 0 -1 54096
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_38
timestamp 1486834041
transform 1 0 4928 0 -1 54096
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_56
timestamp 1486834041
transform 1 0 6944 0 -1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_64
timestamp 1486834041
transform 1 0 7840 0 -1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_68
timestamp 1486834041
transform 1 0 8288 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_72
timestamp 1486834041
transform 1 0 8736 0 -1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_76
timestamp 1486834041
transform 1 0 9184 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_110
timestamp 1486834041
transform 1 0 12992 0 -1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_118
timestamp 1486834041
transform 1 0 13888 0 -1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_121
timestamp 1486834041
transform 1 0 14224 0 -1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_135
timestamp 1486834041
transform 1 0 15792 0 -1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_139
timestamp 1486834041
transform 1 0 16240 0 -1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_142
timestamp 1486834041
transform 1 0 16576 0 -1 54096
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_174
timestamp 1486834041
transform 1 0 20160 0 -1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_182
timestamp 1486834041
transform 1 0 21056 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_190
timestamp 1486834041
transform 1 0 21952 0 -1 54096
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_206
timestamp 1486834041
transform 1 0 23744 0 -1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_212
timestamp 1486834041
transform 1 0 24416 0 -1 54096
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_244
timestamp 1486834041
transform 1 0 28000 0 -1 54096
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_260
timestamp 1486834041
transform 1 0 29792 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_262
timestamp 1486834041
transform 1 0 30016 0 -1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_68_2
timestamp 1486834041
transform 1 0 896 0 1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_30
timestamp 1486834041
transform 1 0 4032 0 1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_34
timestamp 1486834041
transform 1 0 4480 0 1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_37
timestamp 1486834041
transform 1 0 4816 0 1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_41
timestamp 1486834041
transform 1 0 5264 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_43
timestamp 1486834041
transform 1 0 5488 0 1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_68_76
timestamp 1486834041
transform 1 0 9184 0 1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_84
timestamp 1486834041
transform 1 0 10080 0 1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_68_107
timestamp 1486834041
transform 1 0 12656 0 1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_115
timestamp 1486834041
transform 1 0 13552 0 1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_68_151
timestamp 1486834041
transform 1 0 17584 0 1 54096
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_68_167
timestamp 1486834041
transform 1 0 19376 0 1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_177
timestamp 1486834041
transform 1 0 20496 0 1 54096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_241
timestamp 1486834041
transform 1 0 27664 0 1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_68_247
timestamp 1486834041
transform 1 0 28336 0 1 54096
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_69_2
timestamp 1486834041
transform 1 0 896 0 -1 55664
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_72
timestamp 1486834041
transform 1 0 8736 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_74
timestamp 1486834041
transform 1 0 8960 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_69_95
timestamp 1486834041
transform 1 0 11312 0 -1 55664
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_111
timestamp 1486834041
transform 1 0 13104 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_133
timestamp 1486834041
transform 1 0 15568 0 -1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_137
timestamp 1486834041
transform 1 0 16016 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_139
timestamp 1486834041
transform 1 0 16240 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_69_142
timestamp 1486834041
transform 1 0 16576 0 -1 55664
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_158
timestamp 1486834041
transform 1 0 18368 0 -1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_162
timestamp 1486834041
transform 1 0 18816 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_69_165
timestamp 1486834041
transform 1 0 19152 0 -1 55664
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_69_197
timestamp 1486834041
transform 1 0 22736 0 -1 55664
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_205
timestamp 1486834041
transform 1 0 23632 0 -1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_209
timestamp 1486834041
transform 1 0 24080 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_268
timestamp 1486834041
transform 1 0 30688 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_70_2
timestamp 1486834041
transform 1 0 896 0 1 55664
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_34
timestamp 1486834041
transform 1 0 4480 0 1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_37
timestamp 1486834041
transform 1 0 4816 0 1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_41
timestamp 1486834041
transform 1 0 5264 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_70_63
timestamp 1486834041
transform 1 0 7728 0 1 55664
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_71
timestamp 1486834041
transform 1 0 8624 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_70_127
timestamp 1486834041
transform 1 0 14896 0 1 55664
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_159
timestamp 1486834041
transform 1 0 18480 0 1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_70_165
timestamp 1486834041
transform 1 0 19152 0 1 55664
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_173
timestamp 1486834041
transform 1 0 20048 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_177
timestamp 1486834041
transform 1 0 20496 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_179
timestamp 1486834041
transform 1 0 20720 0 1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_70_186
timestamp 1486834041
transform 1 0 21504 0 1 55664
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_70_218
timestamp 1486834041
transform 1 0 25088 0 1 55664
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_70_234
timestamp 1486834041
transform 1 0 26880 0 1 55664
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_242
timestamp 1486834041
transform 1 0 27776 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_244
timestamp 1486834041
transform 1 0 28000 0 1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_70_247
timestamp 1486834041
transform 1 0 28336 0 1 55664
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_71_2
timestamp 1486834041
transform 1 0 896 0 -1 57232
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_71_18
timestamp 1486834041
transform 1 0 2688 0 -1 57232
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_26
timestamp 1486834041
transform 1 0 3584 0 -1 57232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_71_72
timestamp 1486834041
transform 1 0 8736 0 -1 57232
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_80
timestamp 1486834041
transform 1 0 9632 0 -1 57232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_82
timestamp 1486834041
transform 1 0 9856 0 -1 57232
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_71_115
timestamp 1486834041
transform 1 0 13552 0 -1 57232
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_71_131
timestamp 1486834041
transform 1 0 15344 0 -1 57232
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_139
timestamp 1486834041
transform 1 0 16240 0 -1 57232
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_71_142
timestamp 1486834041
transform 1 0 16576 0 -1 57232
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_158
timestamp 1486834041
transform 1 0 18368 0 -1 57232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_162
timestamp 1486834041
transform 1 0 18816 0 -1 57232
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_71_165
timestamp 1486834041
transform 1 0 19152 0 -1 57232
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_71_197
timestamp 1486834041
transform 1 0 22736 0 -1 57232
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_205
timestamp 1486834041
transform 1 0 23632 0 -1 57232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_209
timestamp 1486834041
transform 1 0 24080 0 -1 57232
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_71_212
timestamp 1486834041
transform 1 0 24416 0 -1 57232
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_71_244
timestamp 1486834041
transform 1 0 28000 0 -1 57232
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_260
timestamp 1486834041
transform 1 0 29792 0 -1 57232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_262
timestamp 1486834041
transform 1 0 30016 0 -1 57232
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_72_8
timestamp 1486834041
transform 1 0 1568 0 1 57232
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_72_24
timestamp 1486834041
transform 1 0 3360 0 1 57232
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_32
timestamp 1486834041
transform 1 0 4256 0 1 57232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_34
timestamp 1486834041
transform 1 0 4480 0 1 57232
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_72_37
timestamp 1486834041
transform 1 0 4816 0 1 57232
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_72_53
timestamp 1486834041
transform 1 0 6608 0 1 57232
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_61
timestamp 1486834041
transform 1 0 7504 0 1 57232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_103
timestamp 1486834041
transform 1 0 12208 0 1 57232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_107
timestamp 1486834041
transform 1 0 12656 0 1 57232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_72_155
timestamp 1486834041
transform 1 0 18032 0 1 57232
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_72_165
timestamp 1486834041
transform 1 0 19152 0 1 57232
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_173
timestamp 1486834041
transform 1 0 20048 0 1 57232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_177
timestamp 1486834041
transform 1 0 20496 0 1 57232
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_241
timestamp 1486834041
transform 1 0 27664 0 1 57232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_72_247
timestamp 1486834041
transform 1 0 28336 0 1 57232
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_255
timestamp 1486834041
transform 1 0 29232 0 1 57232
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_262
timestamp 1486834041
transform 1 0 30016 0 1 57232
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_266
timestamp 1486834041
transform 1 0 30464 0 1 57232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_268
timestamp 1486834041
transform 1 0 30688 0 1 57232
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_73_14
timestamp 1486834041
transform 1 0 2240 0 -1 58800
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_73_46
timestamp 1486834041
transform 1 0 5824 0 -1 58800
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_73_62
timestamp 1486834041
transform 1 0 7616 0 -1 58800
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_72
timestamp 1486834041
transform 1 0 8736 0 -1 58800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_76
timestamp 1486834041
transform 1 0 9184 0 -1 58800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_73_97
timestamp 1486834041
transform 1 0 11536 0 -1 58800
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_133
timestamp 1486834041
transform 1 0 15568 0 -1 58800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_137
timestamp 1486834041
transform 1 0 16016 0 -1 58800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_139
timestamp 1486834041
transform 1 0 16240 0 -1 58800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_73_148
timestamp 1486834041
transform 1 0 17248 0 -1 58800
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_156
timestamp 1486834041
transform 1 0 18144 0 -1 58800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_160
timestamp 1486834041
transform 1 0 18592 0 -1 58800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_73_181
timestamp 1486834041
transform 1 0 20944 0 -1 58800
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_73_197
timestamp 1486834041
transform 1 0 22736 0 -1 58800
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_205
timestamp 1486834041
transform 1 0 23632 0 -1 58800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_209
timestamp 1486834041
transform 1 0 24080 0 -1 58800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_73_212
timestamp 1486834041
transform 1 0 24416 0 -1 58800
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_73_244
timestamp 1486834041
transform 1 0 28000 0 -1 58800
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_252
timestamp 1486834041
transform 1 0 28896 0 -1 58800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_262
timestamp 1486834041
transform 1 0 30016 0 -1 58800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_8
timestamp 1486834041
transform 1 0 1568 0 1 58800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_74_21
timestamp 1486834041
transform 1 0 3024 0 1 58800
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_29
timestamp 1486834041
transform 1 0 3920 0 1 58800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_33
timestamp 1486834041
transform 1 0 4368 0 1 58800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_74_37
timestamp 1486834041
transform 1 0 4816 0 1 58800
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_74_53
timestamp 1486834041
transform 1 0 6608 0 1 58800
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_61
timestamp 1486834041
transform 1 0 7504 0 1 58800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_74_85
timestamp 1486834041
transform 1 0 10192 0 1 58800
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_101
timestamp 1486834041
transform 1 0 11984 0 1 58800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_74_107
timestamp 1486834041
transform 1 0 12656 0 1 58800
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_115
timestamp 1486834041
transform 1 0 13552 0 1 58800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_119
timestamp 1486834041
transform 1 0 14000 0 1 58800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_121
timestamp 1486834041
transform 1 0 14224 0 1 58800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_162
timestamp 1486834041
transform 1 0 18816 0 1 58800
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_74_165
timestamp 1486834041
transform 1 0 19152 0 1 58800
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_173
timestamp 1486834041
transform 1 0 20048 0 1 58800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_177
timestamp 1486834041
transform 1 0 20496 0 1 58800
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_241
timestamp 1486834041
transform 1 0 27664 0 1 58800
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_74_247
timestamp 1486834041
transform 1 0 28336 0 1 58800
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_22
timestamp 1486834041
transform 1 0 3136 0 -1 60368
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_63
timestamp 1486834041
transform 1 0 7728 0 -1 60368
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_67
timestamp 1486834041
transform 1 0 8176 0 -1 60368
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_69
timestamp 1486834041
transform 1 0 8400 0 -1 60368
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_72
timestamp 1486834041
transform 1 0 8736 0 -1 60368
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_75_102
timestamp 1486834041
transform 1 0 12096 0 -1 60368
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_118
timestamp 1486834041
transform 1 0 13888 0 -1 60368
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_139
timestamp 1486834041
transform 1 0 16240 0 -1 60368
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_75_196
timestamp 1486834041
transform 1 0 22624 0 -1 60368
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_204
timestamp 1486834041
transform 1 0 23520 0 -1 60368
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_208
timestamp 1486834041
transform 1 0 23968 0 -1 60368
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_75_212
timestamp 1486834041
transform 1 0 24416 0 -1 60368
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_75_244
timestamp 1486834041
transform 1 0 28000 0 -1 60368
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_252
timestamp 1486834041
transform 1 0 28896 0 -1 60368
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_262
timestamp 1486834041
transform 1 0 30016 0 -1 60368
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_266
timestamp 1486834041
transform 1 0 30464 0 -1 60368
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_268
timestamp 1486834041
transform 1 0 30688 0 -1 60368
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_8
timestamp 1486834041
transform 1 0 1568 0 1 60368
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_37
timestamp 1486834041
transform 1 0 4816 0 1 60368
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_41
timestamp 1486834041
transform 1 0 5264 0 1 60368
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_76_75
timestamp 1486834041
transform 1 0 9072 0 1 60368
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_83
timestamp 1486834041
transform 1 0 9968 0 1 60368
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_107
timestamp 1486834041
transform 1 0 12656 0 1 60368
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_169
timestamp 1486834041
transform 1 0 19600 0 1 60368
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_173
timestamp 1486834041
transform 1 0 20048 0 1 60368
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_76_209
timestamp 1486834041
transform 1 0 24080 0 1 60368
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_241
timestamp 1486834041
transform 1 0 27664 0 1 60368
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_76_247
timestamp 1486834041
transform 1 0 28336 0 1 60368
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_255
timestamp 1486834041
transform 1 0 29232 0 1 60368
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_262
timestamp 1486834041
transform 1 0 30016 0 1 60368
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_8
timestamp 1486834041
transform 1 0 1568 0 -1 61936
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_15
timestamp 1486834041
transform 1 0 2352 0 -1 61936
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_17
timestamp 1486834041
transform 1 0 2576 0 -1 61936
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_72
timestamp 1486834041
transform 1 0 8736 0 -1 61936
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_128
timestamp 1486834041
transform 1 0 15008 0 -1 61936
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_154
timestamp 1486834041
transform 1 0 17920 0 -1 61936
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_77_187
timestamp 1486834041
transform 1 0 21616 0 -1 61936
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_203
timestamp 1486834041
transform 1 0 23408 0 -1 61936
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_207
timestamp 1486834041
transform 1 0 23856 0 -1 61936
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_209
timestamp 1486834041
transform 1 0 24080 0 -1 61936
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_77_212
timestamp 1486834041
transform 1 0 24416 0 -1 61936
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_77_244
timestamp 1486834041
transform 1 0 28000 0 -1 61936
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_252
timestamp 1486834041
transform 1 0 28896 0 -1 61936
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_262
timestamp 1486834041
transform 1 0 30016 0 -1 61936
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_2
timestamp 1486834041
transform 1 0 896 0 1 61936
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_78_81
timestamp 1486834041
transform 1 0 9744 0 1 61936
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_89
timestamp 1486834041
transform 1 0 10640 0 1 61936
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_78_92
timestamp 1486834041
transform 1 0 10976 0 1 61936
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_100
timestamp 1486834041
transform 1 0 11872 0 1 61936
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_104
timestamp 1486834041
transform 1 0 12320 0 1 61936
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_78_107
timestamp 1486834041
transform 1 0 12656 0 1 61936
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_115
timestamp 1486834041
transform 1 0 13552 0 1 61936
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_119
timestamp 1486834041
transform 1 0 14000 0 1 61936
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_172
timestamp 1486834041
transform 1 0 19936 0 1 61936
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_174
timestamp 1486834041
transform 1 0 20160 0 1 61936
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_78_209
timestamp 1486834041
transform 1 0 24080 0 1 61936
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_241
timestamp 1486834041
transform 1 0 27664 0 1 61936
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_78_247
timestamp 1486834041
transform 1 0 28336 0 1 61936
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_263
timestamp 1486834041
transform 1 0 30128 0 1 61936
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_267
timestamp 1486834041
transform 1 0 30576 0 1 61936
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_2
timestamp 1486834041
transform 1 0 896 0 -1 63504
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_42
timestamp 1486834041
transform 1 0 5376 0 -1 63504
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_63
timestamp 1486834041
transform 1 0 7728 0 -1 63504
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_79_78
timestamp 1486834041
transform 1 0 9408 0 -1 63504
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_86
timestamp 1486834041
transform 1 0 10304 0 -1 63504
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_122
timestamp 1486834041
transform 1 0 14336 0 -1 63504
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_126
timestamp 1486834041
transform 1 0 14784 0 -1 63504
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_132
timestamp 1486834041
transform 1 0 15456 0 -1 63504
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_139
timestamp 1486834041
transform 1 0 16240 0 -1 63504
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_142
timestamp 1486834041
transform 1 0 16576 0 -1 63504
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_79_195
timestamp 1486834041
transform 1 0 22512 0 -1 63504
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_203
timestamp 1486834041
transform 1 0 23408 0 -1 63504
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_207
timestamp 1486834041
transform 1 0 23856 0 -1 63504
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_209
timestamp 1486834041
transform 1 0 24080 0 -1 63504
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_79_212
timestamp 1486834041
transform 1 0 24416 0 -1 63504
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_79_244
timestamp 1486834041
transform 1 0 28000 0 -1 63504
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_252
timestamp 1486834041
transform 1 0 28896 0 -1 63504
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_262
timestamp 1486834041
transform 1 0 30016 0 -1 63504
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_34
timestamp 1486834041
transform 1 0 4480 0 1 63504
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_43
timestamp 1486834041
transform 1 0 5488 0 1 63504
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_47
timestamp 1486834041
transform 1 0 5936 0 1 63504
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_49
timestamp 1486834041
transform 1 0 6160 0 1 63504
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_80_92
timestamp 1486834041
transform 1 0 10976 0 1 63504
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_100
timestamp 1486834041
transform 1 0 11872 0 1 63504
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_104
timestamp 1486834041
transform 1 0 12320 0 1 63504
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_80_107
timestamp 1486834041
transform 1 0 12656 0 1 63504
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_115
timestamp 1486834041
transform 1 0 13552 0 1 63504
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_117
timestamp 1486834041
transform 1 0 13776 0 1 63504
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_80_138
timestamp 1486834041
transform 1 0 16128 0 1 63504
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_146
timestamp 1486834041
transform 1 0 17024 0 1 63504
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_174
timestamp 1486834041
transform 1 0 20160 0 1 63504
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_177
timestamp 1486834041
transform 1 0 20496 0 1 63504
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_80_198
timestamp 1486834041
transform 1 0 22848 0 1 63504
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_80_230
timestamp 1486834041
transform 1 0 26432 0 1 63504
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_238
timestamp 1486834041
transform 1 0 27328 0 1 63504
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_242
timestamp 1486834041
transform 1 0 27776 0 1 63504
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_244
timestamp 1486834041
transform 1 0 28000 0 1 63504
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_80_247
timestamp 1486834041
transform 1 0 28336 0 1 63504
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_255
timestamp 1486834041
transform 1 0 29232 0 1 63504
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_262
timestamp 1486834041
transform 1 0 30016 0 1 63504
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_2
timestamp 1486834041
transform 1 0 896 0 -1 65072
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_4
timestamp 1486834041
transform 1 0 1120 0 -1 65072
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_49
timestamp 1486834041
transform 1 0 6160 0 -1 65072
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_72
timestamp 1486834041
transform 1 0 8736 0 -1 65072
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_105
timestamp 1486834041
transform 1 0 12432 0 -1 65072
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_107
timestamp 1486834041
transform 1 0 12656 0 -1 65072
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_81_128
timestamp 1486834041
transform 1 0 15008 0 -1 65072
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_136
timestamp 1486834041
transform 1 0 15904 0 -1 65072
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_81_142
timestamp 1486834041
transform 1 0 16576 0 -1 65072
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_158
timestamp 1486834041
transform 1 0 18368 0 -1 65072
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_166
timestamp 1486834041
transform 1 0 19264 0 -1 65072
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_81_187
timestamp 1486834041
transform 1 0 21616 0 -1 65072
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_203
timestamp 1486834041
transform 1 0 23408 0 -1 65072
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_207
timestamp 1486834041
transform 1 0 23856 0 -1 65072
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_209
timestamp 1486834041
transform 1 0 24080 0 -1 65072
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_81_212
timestamp 1486834041
transform 1 0 24416 0 -1 65072
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_81_244
timestamp 1486834041
transform 1 0 28000 0 -1 65072
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_260
timestamp 1486834041
transform 1 0 29792 0 -1 65072
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_262
timestamp 1486834041
transform 1 0 30016 0 -1 65072
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_28
timestamp 1486834041
transform 1 0 3808 0 1 65072
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_82_63
timestamp 1486834041
transform 1 0 7728 0 1 65072
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_71
timestamp 1486834041
transform 1 0 8624 0 1 65072
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_127
timestamp 1486834041
transform 1 0 14896 0 1 65072
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_131
timestamp 1486834041
transform 1 0 15344 0 1 65072
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_152
timestamp 1486834041
transform 1 0 17696 0 1 65072
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_174
timestamp 1486834041
transform 1 0 20160 0 1 65072
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_82_183
timestamp 1486834041
transform 1 0 21168 0 1 65072
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_82_215
timestamp 1486834041
transform 1 0 24752 0 1 65072
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_82_231
timestamp 1486834041
transform 1 0 26544 0 1 65072
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_239
timestamp 1486834041
transform 1 0 27440 0 1 65072
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_243
timestamp 1486834041
transform 1 0 27888 0 1 65072
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_82_247
timestamp 1486834041
transform 1 0 28336 0 1 65072
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_263
timestamp 1486834041
transform 1 0 30128 0 1 65072
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_267
timestamp 1486834041
transform 1 0 30576 0 1 65072
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_34
timestamp 1486834041
transform 1 0 4480 0 -1 66640
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_72
timestamp 1486834041
transform 1 0 8736 0 -1 66640
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_83_108
timestamp 1486834041
transform 1 0 12768 0 -1 66640
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_116
timestamp 1486834041
transform 1 0 13664 0 -1 66640
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_138
timestamp 1486834041
transform 1 0 16128 0 -1 66640
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_83_142
timestamp 1486834041
transform 1 0 16576 0 -1 66640
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_150
timestamp 1486834041
transform 1 0 17472 0 -1 66640
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_154
timestamp 1486834041
transform 1 0 17920 0 -1 66640
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_83_187
timestamp 1486834041
transform 1 0 21616 0 -1 66640
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_203
timestamp 1486834041
transform 1 0 23408 0 -1 66640
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_207
timestamp 1486834041
transform 1 0 23856 0 -1 66640
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_209
timestamp 1486834041
transform 1 0 24080 0 -1 66640
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_83_212
timestamp 1486834041
transform 1 0 24416 0 -1 66640
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_83_244
timestamp 1486834041
transform 1 0 28000 0 -1 66640
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_260
timestamp 1486834041
transform 1 0 29792 0 -1 66640
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_262
timestamp 1486834041
transform 1 0 30016 0 -1 66640
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_2
timestamp 1486834041
transform 1 0 896 0 1 66640
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_84_37
timestamp 1486834041
transform 1 0 4816 0 1 66640
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_73
timestamp 1486834041
transform 1 0 8848 0 1 66640
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_84_97
timestamp 1486834041
transform 1 0 11536 0 1 66640
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_107
timestamp 1486834041
transform 1 0 12656 0 1 66640
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_111
timestamp 1486834041
transform 1 0 13104 0 1 66640
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_171
timestamp 1486834041
transform 1 0 19824 0 1 66640
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_177
timestamp 1486834041
transform 1 0 20496 0 1 66640
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_84_203
timestamp 1486834041
transform 1 0 23408 0 1 66640
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_84_235
timestamp 1486834041
transform 1 0 26992 0 1 66640
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_243
timestamp 1486834041
transform 1 0 27888 0 1 66640
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_84_247
timestamp 1486834041
transform 1 0 28336 0 1 66640
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_8
timestamp 1486834041
transform 1 0 1568 0 -1 68208
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_15
timestamp 1486834041
transform 1 0 2352 0 -1 68208
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_69
timestamp 1486834041
transform 1 0 8400 0 -1 68208
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_72
timestamp 1486834041
transform 1 0 8736 0 -1 68208
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_96
timestamp 1486834041
transform 1 0 11424 0 -1 68208
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_100
timestamp 1486834041
transform 1 0 11872 0 -1 68208
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_133
timestamp 1486834041
transform 1 0 15568 0 -1 68208
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_142
timestamp 1486834041
transform 1 0 16576 0 -1 68208
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_207
timestamp 1486834041
transform 1 0 23856 0 -1 68208
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_209
timestamp 1486834041
transform 1 0 24080 0 -1 68208
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_85_212
timestamp 1486834041
transform 1 0 24416 0 -1 68208
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_85_244
timestamp 1486834041
transform 1 0 28000 0 -1 68208
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_252
timestamp 1486834041
transform 1 0 28896 0 -1 68208
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_262
timestamp 1486834041
transform 1 0 30016 0 -1 68208
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_266
timestamp 1486834041
transform 1 0 30464 0 -1 68208
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_268
timestamp 1486834041
transform 1 0 30688 0 -1 68208
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_34
timestamp 1486834041
transform 1 0 4480 0 1 68208
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_83
timestamp 1486834041
transform 1 0 9968 0 1 68208
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_127
timestamp 1486834041
transform 1 0 14896 0 1 68208
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_161
timestamp 1486834041
transform 1 0 18704 0 1 68208
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_86_219
timestamp 1486834041
transform 1 0 25200 0 1 68208
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_86_235
timestamp 1486834041
transform 1 0 26992 0 1 68208
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_243
timestamp 1486834041
transform 1 0 27888 0 1 68208
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_86_247
timestamp 1486834041
transform 1 0 28336 0 1 68208
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_255
timestamp 1486834041
transform 1 0 29232 0 1 68208
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_262
timestamp 1486834041
transform 1 0 30016 0 1 68208
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_8
timestamp 1486834041
transform 1 0 1568 0 -1 69776
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_62
timestamp 1486834041
transform 1 0 7616 0 -1 69776
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_92
timestamp 1486834041
transform 1 0 10976 0 -1 69776
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_96
timestamp 1486834041
transform 1 0 11424 0 -1 69776
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_98
timestamp 1486834041
transform 1 0 11648 0 -1 69776
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_87_105
timestamp 1486834041
transform 1 0 12432 0 -1 69776
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_113
timestamp 1486834041
transform 1 0 13328 0 -1 69776
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_137
timestamp 1486834041
transform 1 0 16016 0 -1 69776
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_139
timestamp 1486834041
transform 1 0 16240 0 -1 69776
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_208
timestamp 1486834041
transform 1 0 23968 0 -1 69776
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_87_212
timestamp 1486834041
transform 1 0 24416 0 -1 69776
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_87_244
timestamp 1486834041
transform 1 0 28000 0 -1 69776
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_260
timestamp 1486834041
transform 1 0 29792 0 -1 69776
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_262
timestamp 1486834041
transform 1 0 30016 0 -1 69776
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_34
timestamp 1486834041
transform 1 0 4480 0 1 69776
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_37
timestamp 1486834041
transform 1 0 4816 0 1 69776
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_41
timestamp 1486834041
transform 1 0 5264 0 1 69776
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_68
timestamp 1486834041
transform 1 0 8288 0 1 69776
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_72
timestamp 1486834041
transform 1 0 8736 0 1 69776
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_88_107
timestamp 1486834041
transform 1 0 12656 0 1 69776
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_115
timestamp 1486834041
transform 1 0 13552 0 1 69776
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_119
timestamp 1486834041
transform 1 0 14000 0 1 69776
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_121
timestamp 1486834041
transform 1 0 14224 0 1 69776
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_148
timestamp 1486834041
transform 1 0 17248 0 1 69776
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_177
timestamp 1486834041
transform 1 0 20496 0 1 69776
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_88_201
timestamp 1486834041
transform 1 0 23184 0 1 69776
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_88_233
timestamp 1486834041
transform 1 0 26768 0 1 69776
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_241
timestamp 1486834041
transform 1 0 27664 0 1 69776
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_88_247
timestamp 1486834041
transform 1 0 28336 0 1 69776
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_263
timestamp 1486834041
transform 1 0 30128 0 1 69776
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_267
timestamp 1486834041
transform 1 0 30576 0 1 69776
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_2
timestamp 1486834041
transform 1 0 896 0 -1 71344
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_78
timestamp 1486834041
transform 1 0 9408 0 -1 71344
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_89_99
timestamp 1486834041
transform 1 0 11760 0 -1 71344
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_115
timestamp 1486834041
transform 1 0 13552 0 -1 71344
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_119
timestamp 1486834041
transform 1 0 14000 0 -1 71344
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_89_142
timestamp 1486834041
transform 1 0 16576 0 -1 71344
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_158
timestamp 1486834041
transform 1 0 18368 0 -1 71344
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_162
timestamp 1486834041
transform 1 0 18816 0 -1 71344
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_89_165
timestamp 1486834041
transform 1 0 19152 0 -1 71344
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_173
timestamp 1486834041
transform 1 0 20048 0 -1 71344
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_177
timestamp 1486834041
transform 1 0 20496 0 -1 71344
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_179
timestamp 1486834041
transform 1 0 20720 0 -1 71344
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_89_200
timestamp 1486834041
transform 1 0 23072 0 -1 71344
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_208
timestamp 1486834041
transform 1 0 23968 0 -1 71344
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_89_212
timestamp 1486834041
transform 1 0 24416 0 -1 71344
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_89_244
timestamp 1486834041
transform 1 0 28000 0 -1 71344
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_252
timestamp 1486834041
transform 1 0 28896 0 -1 71344
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_262
timestamp 1486834041
transform 1 0 30016 0 -1 71344
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_14
timestamp 1486834041
transform 1 0 2240 0 1 71344
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_43
timestamp 1486834041
transform 1 0 5488 0 1 71344
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_99
timestamp 1486834041
transform 1 0 11760 0 1 71344
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_103
timestamp 1486834041
transform 1 0 12208 0 1 71344
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_90_107
timestamp 1486834041
transform 1 0 12656 0 1 71344
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_115
timestamp 1486834041
transform 1 0 13552 0 1 71344
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_177
timestamp 1486834041
transform 1 0 20496 0 1 71344
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_90_205
timestamp 1486834041
transform 1 0 23632 0 1 71344
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_90_237
timestamp 1486834041
transform 1 0 27216 0 1 71344
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_90_247
timestamp 1486834041
transform 1 0 28336 0 1 71344
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_8
timestamp 1486834041
transform 1 0 1568 0 -1 72912
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_10
timestamp 1486834041
transform 1 0 1792 0 -1 72912
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_69
timestamp 1486834041
transform 1 0 8400 0 -1 72912
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_72
timestamp 1486834041
transform 1 0 8736 0 -1 72912
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_91_131
timestamp 1486834041
transform 1 0 15344 0 -1 72912
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_139
timestamp 1486834041
transform 1 0 16240 0 -1 72912
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_142
timestamp 1486834041
transform 1 0 16576 0 -1 72912
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_146
timestamp 1486834041
transform 1 0 17024 0 -1 72912
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_154
timestamp 1486834041
transform 1 0 17920 0 -1 72912
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_208
timestamp 1486834041
transform 1 0 23968 0 -1 72912
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_91_212
timestamp 1486834041
transform 1 0 24416 0 -1 72912
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_91_244
timestamp 1486834041
transform 1 0 28000 0 -1 72912
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_260
timestamp 1486834041
transform 1 0 29792 0 -1 72912
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_262
timestamp 1486834041
transform 1 0 30016 0 -1 72912
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_2
timestamp 1486834041
transform 1 0 896 0 1 72912
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_6
timestamp 1486834041
transform 1 0 1344 0 1 72912
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_33
timestamp 1486834041
transform 1 0 4368 0 1 72912
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_97
timestamp 1486834041
transform 1 0 11536 0 1 72912
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_139
timestamp 1486834041
transform 1 0 16240 0 1 72912
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_92_161
timestamp 1486834041
transform 1 0 18704 0 1 72912
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_169
timestamp 1486834041
transform 1 0 19600 0 1 72912
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_173
timestamp 1486834041
transform 1 0 20048 0 1 72912
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_92_183
timestamp 1486834041
transform 1 0 21168 0 1 72912
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_191
timestamp 1486834041
transform 1 0 22064 0 1 72912
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_195
timestamp 1486834041
transform 1 0 22512 0 1 72912
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_197
timestamp 1486834041
transform 1 0 22736 0 1 72912
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_92_204
timestamp 1486834041
transform 1 0 23520 0 1 72912
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_92_236
timestamp 1486834041
transform 1 0 27104 0 1 72912
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_244
timestamp 1486834041
transform 1 0 28000 0 1 72912
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_92_247
timestamp 1486834041
transform 1 0 28336 0 1 72912
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_263
timestamp 1486834041
transform 1 0 30128 0 1 72912
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_267
timestamp 1486834041
transform 1 0 30576 0 1 72912
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_8
timestamp 1486834041
transform 1 0 1568 0 -1 74480
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_15
timestamp 1486834041
transform 1 0 2352 0 -1 74480
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_63
timestamp 1486834041
transform 1 0 7728 0 -1 74480
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_92
timestamp 1486834041
transform 1 0 10976 0 -1 74480
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_113
timestamp 1486834041
transform 1 0 13328 0 -1 74480
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_117
timestamp 1486834041
transform 1 0 13776 0 -1 74480
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_119
timestamp 1486834041
transform 1 0 14000 0 -1 74480
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_148
timestamp 1486834041
transform 1 0 17248 0 -1 74480
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_93_202
timestamp 1486834041
transform 1 0 23296 0 -1 74480
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_212
timestamp 1486834041
transform 1 0 24416 0 -1 74480
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_93_244
timestamp 1486834041
transform 1 0 28000 0 -1 74480
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_260
timestamp 1486834041
transform 1 0 29792 0 -1 74480
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_262
timestamp 1486834041
transform 1 0 30016 0 -1 74480
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_2
timestamp 1486834041
transform 1 0 896 0 1 74480
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_6
timestamp 1486834041
transform 1 0 1344 0 1 74480
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_94_27
timestamp 1486834041
transform 1 0 3696 0 1 74480
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_94_37
timestamp 1486834041
transform 1 0 4816 0 1 74480
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_94_71
timestamp 1486834041
transform 1 0 8624 0 1 74480
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_79
timestamp 1486834041
transform 1 0 9520 0 1 74480
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_94_83
timestamp 1486834041
transform 1 0 9968 0 1 74480
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_94_139
timestamp 1486834041
transform 1 0 16240 0 1 74480
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_141
timestamp 1486834041
transform 1 0 16464 0 1 74480
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_174
timestamp 1486834041
transform 1 0 20160 0 1 74480
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_94_177
timestamp 1486834041
transform 1 0 20496 0 1 74480
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_94_193
timestamp 1486834041
transform 1 0 22288 0 1 74480
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_94_247
timestamp 1486834041
transform 1 0 28336 0 1 74480
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_8
timestamp 1486834041
transform 1 0 1568 0 -1 76048
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_44
timestamp 1486834041
transform 1 0 5600 0 -1 76048
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_95_48
timestamp 1486834041
transform 1 0 6048 0 -1 76048
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_95_72
timestamp 1486834041
transform 1 0 8736 0 -1 76048
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_95_88
timestamp 1486834041
transform 1 0 10528 0 -1 76048
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_96
timestamp 1486834041
transform 1 0 11424 0 -1 76048
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_95_123
timestamp 1486834041
transform 1 0 14448 0 -1 76048
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_139
timestamp 1486834041
transform 1 0 16240 0 -1 76048
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_142
timestamp 1486834041
transform 1 0 16576 0 -1 76048
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_95_163
timestamp 1486834041
transform 1 0 18928 0 -1 76048
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_171
timestamp 1486834041
transform 1 0 19824 0 -1 76048
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_95_212
timestamp 1486834041
transform 1 0 24416 0 -1 76048
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_95_244
timestamp 1486834041
transform 1 0 28000 0 -1 76048
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_95_260
timestamp 1486834041
transform 1 0 29792 0 -1 76048
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_268
timestamp 1486834041
transform 1 0 30688 0 -1 76048
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_34
timestamp 1486834041
transform 1 0 4480 0 1 76048
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_96_49
timestamp 1486834041
transform 1 0 6160 0 1 76048
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_51
timestamp 1486834041
transform 1 0 6384 0 1 76048
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_84
timestamp 1486834041
transform 1 0 10080 0 1 76048
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_107
timestamp 1486834041
transform 1 0 12656 0 1 76048
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_96_172
timestamp 1486834041
transform 1 0 19936 0 1 76048
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_174
timestamp 1486834041
transform 1 0 20160 0 1 76048
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_96_197
timestamp 1486834041
transform 1 0 22736 0 1 76048
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_96_229
timestamp 1486834041
transform 1 0 26320 0 1 76048
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_96_247
timestamp 1486834041
transform 1 0 28336 0 1 76048
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_263
timestamp 1486834041
transform 1 0 30128 0 1 76048
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_96_267
timestamp 1486834041
transform 1 0 30576 0 1 76048
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_66
timestamp 1486834041
transform 1 0 8064 0 -1 77616
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_97_72
timestamp 1486834041
transform 1 0 8736 0 -1 77616
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_74
timestamp 1486834041
transform 1 0 8960 0 -1 77616
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_119
timestamp 1486834041
transform 1 0 14000 0 -1 77616
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_97_162
timestamp 1486834041
transform 1 0 18816 0 -1 77616
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_97_191
timestamp 1486834041
transform 1 0 22064 0 -1 77616
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_97_207
timestamp 1486834041
transform 1 0 23856 0 -1 77616
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_209
timestamp 1486834041
transform 1 0 24080 0 -1 77616
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_97_212
timestamp 1486834041
transform 1 0 24416 0 -1 77616
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_97_244
timestamp 1486834041
transform 1 0 28000 0 -1 77616
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_97_260
timestamp 1486834041
transform 1 0 29792 0 -1 77616
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_268
timestamp 1486834041
transform 1 0 30688 0 -1 77616
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_34
timestamp 1486834041
transform 1 0 4480 0 1 77616
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_37
timestamp 1486834041
transform 1 0 4816 0 1 77616
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_98_127
timestamp 1486834041
transform 1 0 14896 0 1 77616
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_169
timestamp 1486834041
transform 1 0 19600 0 1 77616
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_98_173
timestamp 1486834041
transform 1 0 20048 0 1 77616
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_98_197
timestamp 1486834041
transform 1 0 22736 0 1 77616
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_98_229
timestamp 1486834041
transform 1 0 26320 0 1 77616
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_98_247
timestamp 1486834041
transform 1 0 28336 0 1 77616
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_255
timestamp 1486834041
transform 1 0 29232 0 1 77616
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_262
timestamp 1486834041
transform 1 0 30016 0 1 77616
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_98_266
timestamp 1486834041
transform 1 0 30464 0 1 77616
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_268
timestamp 1486834041
transform 1 0 30688 0 1 77616
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_48
timestamp 1486834041
transform 1 0 6048 0 -1 79184
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_69
timestamp 1486834041
transform 1 0 8400 0 -1 79184
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_99_110
timestamp 1486834041
transform 1 0 12992 0 -1 79184
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_118
timestamp 1486834041
transform 1 0 13888 0 -1 79184
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_139
timestamp 1486834041
transform 1 0 16240 0 -1 79184
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_206
timestamp 1486834041
transform 1 0 23744 0 -1 79184
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_99_212
timestamp 1486834041
transform 1 0 24416 0 -1 79184
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_99_244
timestamp 1486834041
transform 1 0 28000 0 -1 79184
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_99_260
timestamp 1486834041
transform 1 0 29792 0 -1 79184
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_262
timestamp 1486834041
transform 1 0 30016 0 -1 79184
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_28
timestamp 1486834041
transform 1 0 3808 0 1 79184
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_37
timestamp 1486834041
transform 1 0 4816 0 1 79184
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_41
timestamp 1486834041
transform 1 0 5264 0 1 79184
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_100_107
timestamp 1486834041
transform 1 0 12656 0 1 79184
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_100_115
timestamp 1486834041
transform 1 0 13552 0 1 79184
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_117
timestamp 1486834041
transform 1 0 13776 0 1 79184
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_100_124
timestamp 1486834041
transform 1 0 14560 0 1 79184
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_100_164
timestamp 1486834041
transform 1 0 19040 0 1 79184
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_100_172
timestamp 1486834041
transform 1 0 19936 0 1 79184
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_174
timestamp 1486834041
transform 1 0 20160 0 1 79184
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_100_209
timestamp 1486834041
transform 1 0 24080 0 1 79184
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_241
timestamp 1486834041
transform 1 0 27664 0 1 79184
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_100_247
timestamp 1486834041
transform 1 0 28336 0 1 79184
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_255
timestamp 1486834041
transform 1 0 29232 0 1 79184
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_262
timestamp 1486834041
transform 1 0 30016 0 1 79184
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_2
timestamp 1486834041
transform 1 0 896 0 -1 80752
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_72
timestamp 1486834041
transform 1 0 8736 0 -1 80752
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_96
timestamp 1486834041
transform 1 0 11424 0 -1 80752
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_101_100
timestamp 1486834041
transform 1 0 11872 0 -1 80752
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_101_132
timestamp 1486834041
transform 1 0 15456 0 -1 80752
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_101_142
timestamp 1486834041
transform 1 0 16576 0 -1 80752
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_150
timestamp 1486834041
transform 1 0 17472 0 -1 80752
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_154
timestamp 1486834041
transform 1 0 17920 0 -1 80752
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_101_207
timestamp 1486834041
transform 1 0 23856 0 -1 80752
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_209
timestamp 1486834041
transform 1 0 24080 0 -1 80752
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_101_212
timestamp 1486834041
transform 1 0 24416 0 -1 80752
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_101_244
timestamp 1486834041
transform 1 0 28000 0 -1 80752
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_252
timestamp 1486834041
transform 1 0 28896 0 -1 80752
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_262
timestamp 1486834041
transform 1 0 30016 0 -1 80752
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_101_266
timestamp 1486834041
transform 1 0 30464 0 -1 80752
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_268
timestamp 1486834041
transform 1 0 30688 0 -1 80752
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_2
timestamp 1486834041
transform 1 0 896 0 1 80752
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_102_26
timestamp 1486834041
transform 1 0 3584 0 1 80752
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_34
timestamp 1486834041
transform 1 0 4480 0 1 80752
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_43
timestamp 1486834041
transform 1 0 5488 0 1 80752
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_102_93
timestamp 1486834041
transform 1 0 11088 0 1 80752
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_101
timestamp 1486834041
transform 1 0 11984 0 1 80752
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_102_151
timestamp 1486834041
transform 1 0 17584 0 1 80752
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_102_167
timestamp 1486834041
transform 1 0 19376 0 1 80752
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_102_197
timestamp 1486834041
transform 1 0 22736 0 1 80752
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_102_229
timestamp 1486834041
transform 1 0 26320 0 1 80752
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_102_247
timestamp 1486834041
transform 1 0 28336 0 1 80752
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_2
timestamp 1486834041
transform 1 0 896 0 -1 82320
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_103_92
timestamp 1486834041
transform 1 0 10976 0 -1 82320
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_103_137
timestamp 1486834041
transform 1 0 16016 0 -1 82320
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_139
timestamp 1486834041
transform 1 0 16240 0 -1 82320
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_103_142
timestamp 1486834041
transform 1 0 16576 0 -1 82320
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_158
timestamp 1486834041
transform 1 0 18368 0 -1 82320
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_103_162
timestamp 1486834041
transform 1 0 18816 0 -1 82320
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_164
timestamp 1486834041
transform 1 0 19040 0 -1 82320
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_205
timestamp 1486834041
transform 1 0 23632 0 -1 82320
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_209
timestamp 1486834041
transform 1 0 24080 0 -1 82320
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_103_212
timestamp 1486834041
transform 1 0 24416 0 -1 82320
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_103_244
timestamp 1486834041
transform 1 0 28000 0 -1 82320
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_252
timestamp 1486834041
transform 1 0 28896 0 -1 82320
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_262
timestamp 1486834041
transform 1 0 30016 0 -1 82320
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_2
timestamp 1486834041
transform 1 0 896 0 1 82320
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_104_63
timestamp 1486834041
transform 1 0 7728 0 1 82320
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_104_127
timestamp 1486834041
transform 1 0 14896 0 1 82320
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_104_161
timestamp 1486834041
transform 1 0 18704 0 1 82320
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_169
timestamp 1486834041
transform 1 0 19600 0 1 82320
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_104_173
timestamp 1486834041
transform 1 0 20048 0 1 82320
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_104_177
timestamp 1486834041
transform 1 0 20496 0 1 82320
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_193
timestamp 1486834041
transform 1 0 22288 0 1 82320
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_104_200
timestamp 1486834041
transform 1 0 23072 0 1 82320
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_104_232
timestamp 1486834041
transform 1 0 26656 0 1 82320
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_240
timestamp 1486834041
transform 1 0 27552 0 1 82320
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_244
timestamp 1486834041
transform 1 0 28000 0 1 82320
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_104_247
timestamp 1486834041
transform 1 0 28336 0 1 82320
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_263
timestamp 1486834041
transform 1 0 30128 0 1 82320
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_104_267
timestamp 1486834041
transform 1 0 30576 0 1 82320
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_34
timestamp 1486834041
transform 1 0 4480 0 -1 83888
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_105_104
timestamp 1486834041
transform 1 0 12320 0 -1 83888
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_194
timestamp 1486834041
transform 1 0 22400 0 -1 83888
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_105_198
timestamp 1486834041
transform 1 0 22848 0 -1 83888
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_200
timestamp 1486834041
transform 1 0 23072 0 -1 83888
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_105_207
timestamp 1486834041
transform 1 0 23856 0 -1 83888
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_209
timestamp 1486834041
transform 1 0 24080 0 -1 83888
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_105_212
timestamp 1486834041
transform 1 0 24416 0 -1 83888
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_105_244
timestamp 1486834041
transform 1 0 28000 0 -1 83888
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_105_260
timestamp 1486834041
transform 1 0 29792 0 -1 83888
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_262
timestamp 1486834041
transform 1 0 30016 0 -1 83888
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_2
timestamp 1486834041
transform 1 0 896 0 1 83888
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_106_37
timestamp 1486834041
transform 1 0 4816 0 1 83888
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_91
timestamp 1486834041
transform 1 0 10864 0 1 83888
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_106_97
timestamp 1486834041
transform 1 0 11536 0 1 83888
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_107
timestamp 1486834041
transform 1 0 12656 0 1 83888
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_106_112
timestamp 1486834041
transform 1 0 13216 0 1 83888
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_120
timestamp 1486834041
transform 1 0 14112 0 1 83888
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_106_124
timestamp 1486834041
transform 1 0 14560 0 1 83888
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_126
timestamp 1486834041
transform 1 0 14784 0 1 83888
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_174
timestamp 1486834041
transform 1 0 20160 0 1 83888
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_106_209
timestamp 1486834041
transform 1 0 24080 0 1 83888
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_241
timestamp 1486834041
transform 1 0 27664 0 1 83888
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_106_247
timestamp 1486834041
transform 1 0 28336 0 1 83888
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_8
timestamp 1486834041
transform 1 0 1568 0 -1 85456
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_107_61
timestamp 1486834041
transform 1 0 7504 0 -1 85456
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_69
timestamp 1486834041
transform 1 0 8400 0 -1 85456
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_107_72
timestamp 1486834041
transform 1 0 8736 0 -1 85456
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_162
timestamp 1486834041
transform 1 0 18816 0 -1 85456
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_202
timestamp 1486834041
transform 1 0 23296 0 -1 85456
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_209
timestamp 1486834041
transform 1 0 24080 0 -1 85456
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_107_212
timestamp 1486834041
transform 1 0 24416 0 -1 85456
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_107_244
timestamp 1486834041
transform 1 0 28000 0 -1 85456
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_107_260
timestamp 1486834041
transform 1 0 29792 0 -1 85456
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_262
timestamp 1486834041
transform 1 0 30016 0 -1 85456
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_8
timestamp 1486834041
transform 1 0 1568 0 1 85456
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_37
timestamp 1486834041
transform 1 0 4816 0 1 85456
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_108_61
timestamp 1486834041
transform 1 0 7504 0 1 85456
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_63
timestamp 1486834041
transform 1 0 7728 0 1 85456
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_108_96
timestamp 1486834041
transform 1 0 11424 0 1 85456
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_104
timestamp 1486834041
transform 1 0 12320 0 1 85456
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_127
timestamp 1486834041
transform 1 0 14896 0 1 85456
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_108_214
timestamp 1486834041
transform 1 0 24640 0 1 85456
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_108_230
timestamp 1486834041
transform 1 0 26432 0 1 85456
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_238
timestamp 1486834041
transform 1 0 27328 0 1 85456
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_108_242
timestamp 1486834041
transform 1 0 27776 0 1 85456
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_244
timestamp 1486834041
transform 1 0 28000 0 1 85456
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_108_247
timestamp 1486834041
transform 1 0 28336 0 1 85456
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_263
timestamp 1486834041
transform 1 0 30128 0 1 85456
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_108_267
timestamp 1486834041
transform 1 0 30576 0 1 85456
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_109_22
timestamp 1486834041
transform 1 0 3136 0 -1 87024
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_64
timestamp 1486834041
transform 1 0 7840 0 -1 87024
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_109_68
timestamp 1486834041
transform 1 0 8288 0 -1 87024
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_109_72
timestamp 1486834041
transform 1 0 8736 0 -1 87024
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_74
timestamp 1486834041
transform 1 0 8960 0 -1 87024
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_109_127
timestamp 1486834041
transform 1 0 14896 0 -1 87024
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_135
timestamp 1486834041
transform 1 0 15792 0 -1 87024
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_139
timestamp 1486834041
transform 1 0 16240 0 -1 87024
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_109_142
timestamp 1486834041
transform 1 0 16576 0 -1 87024
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_109_158
timestamp 1486834041
transform 1 0 18368 0 -1 87024
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_160
timestamp 1486834041
transform 1 0 18592 0 -1 87024
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_109_212
timestamp 1486834041
transform 1 0 24416 0 -1 87024
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_109_244
timestamp 1486834041
transform 1 0 28000 0 -1 87024
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_109_260
timestamp 1486834041
transform 1 0 29792 0 -1 87024
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_262
timestamp 1486834041
transform 1 0 30016 0 -1 87024
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_2
timestamp 1486834041
transform 1 0 896 0 1 87024
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_6
timestamp 1486834041
transform 1 0 1344 0 1 87024
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_110_27
timestamp 1486834041
transform 1 0 3696 0 1 87024
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_110_37
timestamp 1486834041
transform 1 0 4816 0 1 87024
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_110_45
timestamp 1486834041
transform 1 0 5712 0 1 87024
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_67
timestamp 1486834041
transform 1 0 8176 0 1 87024
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_110_71
timestamp 1486834041
transform 1 0 8624 0 1 87024
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_107
timestamp 1486834041
transform 1 0 12656 0 1 87024
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_110_128
timestamp 1486834041
transform 1 0 15008 0 1 87024
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_110_144
timestamp 1486834041
transform 1 0 16800 0 1 87024
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_110_152
timestamp 1486834041
transform 1 0 17696 0 1 87024
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_154
timestamp 1486834041
transform 1 0 17920 0 1 87024
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_110_209
timestamp 1486834041
transform 1 0 24080 0 1 87024
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_241
timestamp 1486834041
transform 1 0 27664 0 1 87024
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_110_247
timestamp 1486834041
transform 1 0 28336 0 1 87024
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_54
timestamp 1486834041
transform 1 0 6720 0 -1 88592
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_58
timestamp 1486834041
transform 1 0 7168 0 -1 88592
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_111_61
timestamp 1486834041
transform 1 0 7504 0 -1 88592
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_69
timestamp 1486834041
transform 1 0 8400 0 -1 88592
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_111_72
timestamp 1486834041
transform 1 0 8736 0 -1 88592
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_88
timestamp 1486834041
transform 1 0 10528 0 -1 88592
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_111_129
timestamp 1486834041
transform 1 0 15120 0 -1 88592
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_111_137
timestamp 1486834041
transform 1 0 16016 0 -1 88592
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_139
timestamp 1486834041
transform 1 0 16240 0 -1 88592
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_111_142
timestamp 1486834041
transform 1 0 16576 0 -1 88592
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_111_150
timestamp 1486834041
transform 1 0 17472 0 -1 88592
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_111_172
timestamp 1486834041
transform 1 0 19936 0 -1 88592
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_180
timestamp 1486834041
transform 1 0 20832 0 -1 88592
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_111_201
timestamp 1486834041
transform 1 0 23184 0 -1 88592
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_209
timestamp 1486834041
transform 1 0 24080 0 -1 88592
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_111_212
timestamp 1486834041
transform 1 0 24416 0 -1 88592
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_111_244
timestamp 1486834041
transform 1 0 28000 0 -1 88592
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_252
timestamp 1486834041
transform 1 0 28896 0 -1 88592
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_262
timestamp 1486834041
transform 1 0 30016 0 -1 88592
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_111_266
timestamp 1486834041
transform 1 0 30464 0 -1 88592
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_268
timestamp 1486834041
transform 1 0 30688 0 -1 88592
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_112_2
timestamp 1486834041
transform 1 0 896 0 1 88592
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_10
timestamp 1486834041
transform 1 0 1792 0 1 88592
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_14
timestamp 1486834041
transform 1 0 2240 0 1 88592
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_112_37
timestamp 1486834041
transform 1 0 4816 0 1 88592
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_112_97
timestamp 1486834041
transform 1 0 11536 0 1 88592
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_112_127
timestamp 1486834041
transform 1 0 14896 0 1 88592
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_143
timestamp 1486834041
transform 1 0 16688 0 1 88592
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_112_162
timestamp 1486834041
transform 1 0 18816 0 1 88592
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_170
timestamp 1486834041
transform 1 0 19712 0 1 88592
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_174
timestamp 1486834041
transform 1 0 20160 0 1 88592
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_177
timestamp 1486834041
transform 1 0 20496 0 1 88592
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_112_181
timestamp 1486834041
transform 1 0 20944 0 1 88592
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_112_203
timestamp 1486834041
transform 1 0 23408 0 1 88592
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_112_235
timestamp 1486834041
transform 1 0 26992 0 1 88592
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_112_243
timestamp 1486834041
transform 1 0 27888 0 1 88592
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_112_247
timestamp 1486834041
transform 1 0 28336 0 1 88592
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_113_2
timestamp 1486834041
transform 1 0 896 0 -1 90160
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_4
timestamp 1486834041
transform 1 0 1120 0 -1 90160
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_113_67
timestamp 1486834041
transform 1 0 8176 0 -1 90160
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_69
timestamp 1486834041
transform 1 0 8400 0 -1 90160
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_72
timestamp 1486834041
transform 1 0 8736 0 -1 90160
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_76
timestamp 1486834041
transform 1 0 9184 0 -1 90160
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_97
timestamp 1486834041
transform 1 0 11536 0 -1 90160
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_101
timestamp 1486834041
transform 1 0 11984 0 -1 90160
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_113_142
timestamp 1486834041
transform 1 0 16576 0 -1 90160
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_144
timestamp 1486834041
transform 1 0 16800 0 -1 90160
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_113_180
timestamp 1486834041
transform 1 0 20832 0 -1 90160
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_113_196
timestamp 1486834041
transform 1 0 22624 0 -1 90160
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_204
timestamp 1486834041
transform 1 0 23520 0 -1 90160
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_113_208
timestamp 1486834041
transform 1 0 23968 0 -1 90160
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_113_212
timestamp 1486834041
transform 1 0 24416 0 -1 90160
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_113_244
timestamp 1486834041
transform 1 0 28000 0 -1 90160
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_113_260
timestamp 1486834041
transform 1 0 29792 0 -1 90160
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_262
timestamp 1486834041
transform 1 0 30016 0 -1 90160
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_114_22
timestamp 1486834041
transform 1 0 3136 0 1 90160
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_30
timestamp 1486834041
transform 1 0 4032 0 1 90160
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_34
timestamp 1486834041
transform 1 0 4480 0 1 90160
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_114_37
timestamp 1486834041
transform 1 0 4816 0 1 90160
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_114_45
timestamp 1486834041
transform 1 0 5712 0 1 90160
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_114_79
timestamp 1486834041
transform 1 0 9520 0 1 90160
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_101
timestamp 1486834041
transform 1 0 11984 0 1 90160
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_114_165
timestamp 1486834041
transform 1 0 19152 0 1 90160
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_114_173
timestamp 1486834041
transform 1 0 20048 0 1 90160
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_177
timestamp 1486834041
transform 1 0 20496 0 1 90160
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_114_181
timestamp 1486834041
transform 1 0 20944 0 1 90160
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_183
timestamp 1486834041
transform 1 0 21168 0 1 90160
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_114_199
timestamp 1486834041
transform 1 0 22960 0 1 90160
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_114_231
timestamp 1486834041
transform 1 0 26544 0 1 90160
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_239
timestamp 1486834041
transform 1 0 27440 0 1 90160
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_114_243
timestamp 1486834041
transform 1 0 27888 0 1 90160
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_114_247
timestamp 1486834041
transform 1 0 28336 0 1 90160
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_263
timestamp 1486834041
transform 1 0 30128 0 1 90160
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_114_267
timestamp 1486834041
transform 1 0 30576 0 1 90160
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_115_42
timestamp 1486834041
transform 1 0 5376 0 -1 91728
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_115_72
timestamp 1486834041
transform 1 0 8736 0 -1 91728
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_80
timestamp 1486834041
transform 1 0 9632 0 -1 91728
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_84
timestamp 1486834041
transform 1 0 10080 0 -1 91728
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_115_105
timestamp 1486834041
transform 1 0 12432 0 -1 91728
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_107
timestamp 1486834041
transform 1 0 12656 0 -1 91728
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_174
timestamp 1486834041
transform 1 0 20160 0 -1 91728
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_115_178
timestamp 1486834041
transform 1 0 20608 0 -1 91728
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_115_200
timestamp 1486834041
transform 1 0 23072 0 -1 91728
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_115_208
timestamp 1486834041
transform 1 0 23968 0 -1 91728
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_115_212
timestamp 1486834041
transform 1 0 24416 0 -1 91728
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_115_244
timestamp 1486834041
transform 1 0 28000 0 -1 91728
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_115_260
timestamp 1486834041
transform 1 0 29792 0 -1 91728
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_262
timestamp 1486834041
transform 1 0 30016 0 -1 91728
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_116_22
timestamp 1486834041
transform 1 0 3136 0 1 91728
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_30
timestamp 1486834041
transform 1 0 4032 0 1 91728
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_34
timestamp 1486834041
transform 1 0 4480 0 1 91728
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_37
timestamp 1486834041
transform 1 0 4816 0 1 91728
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_116_44
timestamp 1486834041
transform 1 0 5600 0 1 91728
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_98
timestamp 1486834041
transform 1 0 11648 0 1 91728
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_116_102
timestamp 1486834041
transform 1 0 12096 0 1 91728
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_104
timestamp 1486834041
transform 1 0 12320 0 1 91728
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_107
timestamp 1486834041
transform 1 0 12656 0 1 91728
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_111
timestamp 1486834041
transform 1 0 13104 0 1 91728
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_170
timestamp 1486834041
transform 1 0 19712 0 1 91728
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_174
timestamp 1486834041
transform 1 0 20160 0 1 91728
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_116_209
timestamp 1486834041
transform 1 0 24080 0 1 91728
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_241
timestamp 1486834041
transform 1 0 27664 0 1 91728
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_116_247
timestamp 1486834041
transform 1 0 28336 0 1 91728
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_34
timestamp 1486834041
transform 1 0 4480 0 -1 93296
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_104
timestamp 1486834041
transform 1 0 12320 0 -1 93296
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_117_142
timestamp 1486834041
transform 1 0 16576 0 -1 93296
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_164
timestamp 1486834041
transform 1 0 19040 0 -1 93296
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_168
timestamp 1486834041
transform 1 0 19488 0 -1 93296
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_117_201
timestamp 1486834041
transform 1 0 23184 0 -1 93296
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_209
timestamp 1486834041
transform 1 0 24080 0 -1 93296
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_117_227
timestamp 1486834041
transform 1 0 26096 0 -1 93296
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_259
timestamp 1486834041
transform 1 0 29680 0 -1 93296
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_2
timestamp 1486834041
transform 1 0 896 0 1 93296
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_37
timestamp 1486834041
transform 1 0 4816 0 1 93296
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_41
timestamp 1486834041
transform 1 0 5264 0 1 93296
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_62
timestamp 1486834041
transform 1 0 7616 0 1 93296
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_118_66
timestamp 1486834041
transform 1 0 8064 0 1 93296
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_68
timestamp 1486834041
transform 1 0 8288 0 1 93296
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_101
timestamp 1486834041
transform 1 0 11984 0 1 93296
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_107
timestamp 1486834041
transform 1 0 12656 0 1 93296
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_111
timestamp 1486834041
transform 1 0 13104 0 1 93296
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_170
timestamp 1486834041
transform 1 0 19712 0 1 93296
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_174
timestamp 1486834041
transform 1 0 20160 0 1 93296
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_118_177
timestamp 1486834041
transform 1 0 20496 0 1 93296
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_193
timestamp 1486834041
transform 1 0 22288 0 1 93296
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_244
timestamp 1486834041
transform 1 0 28000 0 1 93296
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_118_247
timestamp 1486834041
transform 1 0 28336 0 1 93296
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_263
timestamp 1486834041
transform 1 0 30128 0 1 93296
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_118_267
timestamp 1486834041
transform 1 0 30576 0 1 93296
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_119_2
timestamp 1486834041
transform 1 0 896 0 -1 94864
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_119_6
timestamp 1486834041
transform 1 0 1344 0 -1 94864
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_8
timestamp 1486834041
transform 1 0 1568 0 -1 94864
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_119_61
timestamp 1486834041
transform 1 0 7504 0 -1 94864
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_69
timestamp 1486834041
transform 1 0 8400 0 -1 94864
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_72
timestamp 1486834041
transform 1 0 8736 0 -1 94864
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_119_88
timestamp 1486834041
transform 1 0 10528 0 -1 94864
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_90
timestamp 1486834041
transform 1 0 10752 0 -1 94864
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_119_138
timestamp 1486834041
transform 1 0 16128 0 -1 94864
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_142
timestamp 1486834041
transform 1 0 16576 0 -1 94864
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_119_207
timestamp 1486834041
transform 1 0 23856 0 -1 94864
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_209
timestamp 1486834041
transform 1 0 24080 0 -1 94864
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_119_212
timestamp 1486834041
transform 1 0 24416 0 -1 94864
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_119_244
timestamp 1486834041
transform 1 0 28000 0 -1 94864
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_119_260
timestamp 1486834041
transform 1 0 29792 0 -1 94864
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_119_262
timestamp 1486834041
transform 1 0 30016 0 -1 94864
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_120_34
timestamp 1486834041
transform 1 0 4480 0 1 94864
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_37
timestamp 1486834041
transform 1 0 4816 0 1 94864
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_61
timestamp 1486834041
transform 1 0 7504 0 1 94864
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_120_97
timestamp 1486834041
transform 1 0 11536 0 1 94864
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_120_127
timestamp 1486834041
transform 1 0 14896 0 1 94864
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_120_143
timestamp 1486834041
transform 1 0 16688 0 1 94864
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_151
timestamp 1486834041
transform 1 0 17584 0 1 94864
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_120_209
timestamp 1486834041
transform 1 0 24080 0 1 94864
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_120_241
timestamp 1486834041
transform 1 0 27664 0 1 94864
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_120_247
timestamp 1486834041
transform 1 0 28336 0 1 94864
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_2
timestamp 1486834041
transform 1 0 896 0 -1 96432
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_121_23
timestamp 1486834041
transform 1 0 3248 0 -1 96432
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_25
timestamp 1486834041
transform 1 0 3472 0 -1 96432
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_121_68
timestamp 1486834041
transform 1 0 8288 0 -1 96432
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_121_72
timestamp 1486834041
transform 1 0 8736 0 -1 96432
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_80
timestamp 1486834041
transform 1 0 9632 0 -1 96432
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_121_84
timestamp 1486834041
transform 1 0 10080 0 -1 96432
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_121_118
timestamp 1486834041
transform 1 0 13888 0 -1 96432
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_134
timestamp 1486834041
transform 1 0 15680 0 -1 96432
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_121_138
timestamp 1486834041
transform 1 0 16128 0 -1 96432
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_121_142
timestamp 1486834041
transform 1 0 16576 0 -1 96432
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_121_149
timestamp 1486834041
transform 1 0 17360 0 -1 96432
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_121_157
timestamp 1486834041
transform 1 0 18256 0 -1 96432
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_205
timestamp 1486834041
transform 1 0 23632 0 -1 96432
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_209
timestamp 1486834041
transform 1 0 24080 0 -1 96432
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_121_212
timestamp 1486834041
transform 1 0 24416 0 -1 96432
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_121_244
timestamp 1486834041
transform 1 0 28000 0 -1 96432
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_252
timestamp 1486834041
transform 1 0 28896 0 -1 96432
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_121_262
timestamp 1486834041
transform 1 0 30016 0 -1 96432
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_121_266
timestamp 1486834041
transform 1 0 30464 0 -1 96432
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_121_268
timestamp 1486834041
transform 1 0 30688 0 -1 96432
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_122_2
timestamp 1486834041
transform 1 0 896 0 1 96432
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_10
timestamp 1486834041
transform 1 0 1792 0 1 96432
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_14
timestamp 1486834041
transform 1 0 2240 0 1 96432
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_122_37
timestamp 1486834041
transform 1 0 4816 0 1 96432
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_39
timestamp 1486834041
transform 1 0 5040 0 1 96432
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_100
timestamp 1486834041
transform 1 0 11872 0 1 96432
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_104
timestamp 1486834041
transform 1 0 12320 0 1 96432
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_122_122
timestamp 1486834041
transform 1 0 14336 0 1 96432
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_122_162
timestamp 1486834041
transform 1 0 18816 0 1 96432
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_122_166
timestamp 1486834041
transform 1 0 19264 0 1 96432
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_122_173
timestamp 1486834041
transform 1 0 20048 0 1 96432
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_122_197
timestamp 1486834041
transform 1 0 22736 0 1 96432
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_122_229
timestamp 1486834041
transform 1 0 26320 0 1 96432
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_122_247
timestamp 1486834041
transform 1 0 28336 0 1 96432
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_22
timestamp 1486834041
transform 1 0 3136 0 -1 98000
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_123_26
timestamp 1486834041
transform 1 0 3584 0 -1 98000
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_28
timestamp 1486834041
transform 1 0 3808 0 -1 98000
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_69
timestamp 1486834041
transform 1 0 8400 0 -1 98000
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_123_112
timestamp 1486834041
transform 1 0 13216 0 -1 98000
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_123_170
timestamp 1486834041
transform 1 0 19712 0 -1 98000
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_123_192
timestamp 1486834041
transform 1 0 22176 0 -1 98000
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_123_208
timestamp 1486834041
transform 1 0 23968 0 -1 98000
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_123_212
timestamp 1486834041
transform 1 0 24416 0 -1 98000
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_123_244
timestamp 1486834041
transform 1 0 28000 0 -1 98000
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_123_252
timestamp 1486834041
transform 1 0 28896 0 -1 98000
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_123_262
timestamp 1486834041
transform 1 0 30016 0 -1 98000
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_2
timestamp 1486834041
transform 1 0 896 0 1 98000
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_6
timestamp 1486834041
transform 1 0 1344 0 1 98000
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_124_27
timestamp 1486834041
transform 1 0 3696 0 1 98000
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_29
timestamp 1486834041
transform 1 0 3920 0 1 98000
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_37
timestamp 1486834041
transform 1 0 4816 0 1 98000
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_98
timestamp 1486834041
transform 1 0 11648 0 1 98000
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_124_102
timestamp 1486834041
transform 1 0 12096 0 1 98000
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_104
timestamp 1486834041
transform 1 0 12320 0 1 98000
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_107
timestamp 1486834041
transform 1 0 12656 0 1 98000
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_124_174
timestamp 1486834041
transform 1 0 20160 0 1 98000
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_124_177
timestamp 1486834041
transform 1 0 20496 0 1 98000
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_241
timestamp 1486834041
transform 1 0 27664 0 1 98000
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_124_247
timestamp 1486834041
transform 1 0 28336 0 1 98000
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_124_263
timestamp 1486834041
transform 1 0 30128 0 1 98000
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_124_267
timestamp 1486834041
transform 1 0 30576 0 1 98000
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_125_2
timestamp 1486834041
transform 1 0 896 0 -1 99568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_4
timestamp 1486834041
transform 1 0 1120 0 -1 99568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_25
timestamp 1486834041
transform 1 0 3472 0 -1 99568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_125_72
timestamp 1486834041
transform 1 0 8736 0 -1 99568
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_80
timestamp 1486834041
transform 1 0 9632 0 -1 99568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_125_113
timestamp 1486834041
transform 1 0 13328 0 -1 99568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_125_117
timestamp 1486834041
transform 1 0 13776 0 -1 99568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_139
timestamp 1486834041
transform 1 0 16240 0 -1 99568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_125_168
timestamp 1486834041
transform 1 0 19488 0 -1 99568
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_125_200
timestamp 1486834041
transform 1 0 23072 0 -1 99568
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_125_208
timestamp 1486834041
transform 1 0 23968 0 -1 99568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_125_212
timestamp 1486834041
transform 1 0 24416 0 -1 99568
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_125_244
timestamp 1486834041
transform 1 0 28000 0 -1 99568
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_125_260
timestamp 1486834041
transform 1 0 29792 0 -1 99568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_125_262
timestamp 1486834041
transform 1 0 30016 0 -1 99568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_126_2
timestamp 1486834041
transform 1 0 896 0 1 99568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_126_57
timestamp 1486834041
transform 1 0 7056 0 1 99568
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_126_127
timestamp 1486834041
transform 1 0 14896 0 1 99568
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_126_143
timestamp 1486834041
transform 1 0 16688 0 1 99568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_126_165
timestamp 1486834041
transform 1 0 19152 0 1 99568
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_126_173
timestamp 1486834041
transform 1 0 20048 0 1 99568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_126_177
timestamp 1486834041
transform 1 0 20496 0 1 99568
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_126_185
timestamp 1486834041
transform 1 0 21392 0 1 99568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_126_189
timestamp 1486834041
transform 1 0 21840 0 1 99568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_126_197
timestamp 1486834041
transform 1 0 22736 0 1 99568
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_126_229
timestamp 1486834041
transform 1 0 26320 0 1 99568
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_126_247
timestamp 1486834041
transform 1 0 28336 0 1 99568
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_2
timestamp 1486834041
transform 1 0 896 0 -1 101136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_127_23
timestamp 1486834041
transform 1 0 3248 0 -1 101136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_25
timestamp 1486834041
transform 1 0 3472 0 -1 101136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_64
timestamp 1486834041
transform 1 0 7840 0 -1 101136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_127_68
timestamp 1486834041
transform 1 0 8288 0 -1 101136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_72
timestamp 1486834041
transform 1 0 8736 0 -1 101136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_127_76
timestamp 1486834041
transform 1 0 9184 0 -1 101136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_110
timestamp 1486834041
transform 1 0 12992 0 -1 101136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_114
timestamp 1486834041
transform 1 0 13440 0 -1 101136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_135
timestamp 1486834041
transform 1 0 15792 0 -1 101136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_139
timestamp 1486834041
transform 1 0 16240 0 -1 101136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_142
timestamp 1486834041
transform 1 0 16576 0 -1 101136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_146
timestamp 1486834041
transform 1 0 17024 0 -1 101136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_127_153
timestamp 1486834041
transform 1 0 17808 0 -1 101136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_127_185
timestamp 1486834041
transform 1 0 21392 0 -1 101136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_127_201
timestamp 1486834041
transform 1 0 23184 0 -1 101136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_209
timestamp 1486834041
transform 1 0 24080 0 -1 101136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_127_212
timestamp 1486834041
transform 1 0 24416 0 -1 101136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_127_244
timestamp 1486834041
transform 1 0 28000 0 -1 101136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_127_252
timestamp 1486834041
transform 1 0 28896 0 -1 101136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_127_262
timestamp 1486834041
transform 1 0 30016 0 -1 101136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_2
timestamp 1486834041
transform 1 0 896 0 1 101136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_37
timestamp 1486834041
transform 1 0 4816 0 1 101136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_64
timestamp 1486834041
transform 1 0 7840 0 1 101136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_128_68
timestamp 1486834041
transform 1 0 8288 0 1 101136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_128_102
timestamp 1486834041
transform 1 0 12096 0 1 101136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_128_104
timestamp 1486834041
transform 1 0 12320 0 1 101136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_107
timestamp 1486834041
transform 1 0 12656 0 1 101136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_128_143
timestamp 1486834041
transform 1 0 16688 0 1 101136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_128_177
timestamp 1486834041
transform 1 0 20496 0 1 101136
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_241
timestamp 1486834041
transform 1 0 27664 0 1 101136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_128_247
timestamp 1486834041
transform 1 0 28336 0 1 101136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_128_263
timestamp 1486834041
transform 1 0 30128 0 1 101136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_128_267
timestamp 1486834041
transform 1 0 30576 0 1 101136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_2
timestamp 1486834041
transform 1 0 896 0 -1 102704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_23
timestamp 1486834041
transform 1 0 3248 0 -1 102704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_59
timestamp 1486834041
transform 1 0 7280 0 -1 102704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_63
timestamp 1486834041
transform 1 0 7728 0 -1 102704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_72
timestamp 1486834041
transform 1 0 8736 0 -1 102704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_129_142
timestamp 1486834041
transform 1 0 16576 0 -1 102704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_146
timestamp 1486834041
transform 1 0 17024 0 -1 102704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_129_153
timestamp 1486834041
transform 1 0 17808 0 -1 102704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_129_185
timestamp 1486834041
transform 1 0 21392 0 -1 102704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_129_201
timestamp 1486834041
transform 1 0 23184 0 -1 102704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_209
timestamp 1486834041
transform 1 0 24080 0 -1 102704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_129_212
timestamp 1486834041
transform 1 0 24416 0 -1 102704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_129_244
timestamp 1486834041
transform 1 0 28000 0 -1 102704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_129_260
timestamp 1486834041
transform 1 0 29792 0 -1 102704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_129_262
timestamp 1486834041
transform 1 0 30016 0 -1 102704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_22
timestamp 1486834041
transform 1 0 3136 0 1 102704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_130_133
timestamp 1486834041
transform 1 0 15568 0 1 102704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_141
timestamp 1486834041
transform 1 0 16464 0 1 102704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_170
timestamp 1486834041
transform 1 0 19712 0 1 102704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_130_174
timestamp 1486834041
transform 1 0 20160 0 1 102704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_130_177
timestamp 1486834041
transform 1 0 20496 0 1 102704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_130_241
timestamp 1486834041
transform 1 0 27664 0 1 102704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_130_247
timestamp 1486834041
transform 1 0 28336 0 1 102704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_131_2
timestamp 1486834041
transform 1 0 896 0 -1 104272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_131_72
timestamp 1486834041
transform 1 0 8736 0 -1 104272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_80
timestamp 1486834041
transform 1 0 9632 0 -1 104272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_131_137
timestamp 1486834041
transform 1 0 16016 0 -1 104272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_139
timestamp 1486834041
transform 1 0 16240 0 -1 104272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_131_174
timestamp 1486834041
transform 1 0 20160 0 -1 104272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_131_182
timestamp 1486834041
transform 1 0 21056 0 -1 104272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_131_198
timestamp 1486834041
transform 1 0 22848 0 -1 104272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_131_206
timestamp 1486834041
transform 1 0 23744 0 -1 104272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_131_212
timestamp 1486834041
transform 1 0 24416 0 -1 104272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_131_244
timestamp 1486834041
transform 1 0 28000 0 -1 104272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_131_260
timestamp 1486834041
transform 1 0 29792 0 -1 104272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_131_268
timestamp 1486834041
transform 1 0 30688 0 -1 104272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_22
timestamp 1486834041
transform 1 0 3136 0 1 104272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_43
timestamp 1486834041
transform 1 0 5488 0 1 104272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_132_81
timestamp 1486834041
transform 1 0 9744 0 1 104272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_132_89
timestamp 1486834041
transform 1 0 10640 0 1 104272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_91
timestamp 1486834041
transform 1 0 10864 0 1 104272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_132_94
timestamp 1486834041
transform 1 0 11200 0 1 104272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_132_159
timestamp 1486834041
transform 1 0 18480 0 1 104272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_132_177
timestamp 1486834041
transform 1 0 20496 0 1 104272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_132_241
timestamp 1486834041
transform 1 0 27664 0 1 104272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_132_247
timestamp 1486834041
transform 1 0 28336 0 1 104272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_133_2
timestamp 1486834041
transform 1 0 896 0 -1 105840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_78
timestamp 1486834041
transform 1 0 9408 0 -1 105840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_133_81
timestamp 1486834041
transform 1 0 9744 0 -1 105840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_133_89
timestamp 1486834041
transform 1 0 10640 0 -1 105840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_91
timestamp 1486834041
transform 1 0 10864 0 -1 105840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_133_98
timestamp 1486834041
transform 1 0 11648 0 -1 105840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_133_142
timestamp 1486834041
transform 1 0 16576 0 -1 105840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_133_158
timestamp 1486834041
transform 1 0 18368 0 -1 105840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_162
timestamp 1486834041
transform 1 0 18816 0 -1 105840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_133_169
timestamp 1486834041
transform 1 0 19600 0 -1 105840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_133_185
timestamp 1486834041
transform 1 0 21392 0 -1 105840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_133_193
timestamp 1486834041
transform 1 0 22288 0 -1 105840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_209
timestamp 1486834041
transform 1 0 24080 0 -1 105840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_133_212
timestamp 1486834041
transform 1 0 24416 0 -1 105840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_133_244
timestamp 1486834041
transform 1 0 28000 0 -1 105840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_133_260
timestamp 1486834041
transform 1 0 29792 0 -1 105840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_133_262
timestamp 1486834041
transform 1 0 30016 0 -1 105840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_2
timestamp 1486834041
transform 1 0 896 0 1 105840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_134_37
timestamp 1486834041
transform 1 0 4816 0 1 105840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_91
timestamp 1486834041
transform 1 0 10864 0 1 105840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_134_94
timestamp 1486834041
transform 1 0 11200 0 1 105840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_134_102
timestamp 1486834041
transform 1 0 12096 0 1 105840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_104
timestamp 1486834041
transform 1 0 12320 0 1 105840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_134_147
timestamp 1486834041
transform 1 0 17136 0 1 105840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_134_163
timestamp 1486834041
transform 1 0 18928 0 1 105840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_171
timestamp 1486834041
transform 1 0 19824 0 1 105840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_134_177
timestamp 1486834041
transform 1 0 20496 0 1 105840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_241
timestamp 1486834041
transform 1 0 27664 0 1 105840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_134_247
timestamp 1486834041
transform 1 0 28336 0 1 105840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_255
timestamp 1486834041
transform 1 0 29232 0 1 105840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_134_262
timestamp 1486834041
transform 1 0 30016 0 1 105840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_134_266
timestamp 1486834041
transform 1 0 30464 0 1 105840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_134_268
timestamp 1486834041
transform 1 0 30688 0 1 105840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_2
timestamp 1486834041
transform 1 0 896 0 -1 107408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_69
timestamp 1486834041
transform 1 0 8400 0 -1 107408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_72
timestamp 1486834041
transform 1 0 8736 0 -1 107408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_135_75
timestamp 1486834041
transform 1 0 9072 0 -1 107408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_77
timestamp 1486834041
transform 1 0 9296 0 -1 107408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_86
timestamp 1486834041
transform 1 0 10304 0 -1 107408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_135_92
timestamp 1486834041
transform 1 0 10976 0 -1 107408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_94
timestamp 1486834041
transform 1 0 11200 0 -1 107408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_135_121
timestamp 1486834041
transform 1 0 14224 0 -1 107408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_123
timestamp 1486834041
transform 1 0 14448 0 -1 107408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_135_126
timestamp 1486834041
transform 1 0 14784 0 -1 107408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_134
timestamp 1486834041
transform 1 0 15680 0 -1 107408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_135_138
timestamp 1486834041
transform 1 0 16128 0 -1 107408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_135_162
timestamp 1486834041
transform 1 0 18816 0 -1 107408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_135_194
timestamp 1486834041
transform 1 0 22400 0 -1 107408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_135_212
timestamp 1486834041
transform 1 0 24416 0 -1 107408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_135_216
timestamp 1486834041
transform 1 0 24864 0 -1 107408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_135_220
timestamp 1486834041
transform 1 0 25312 0 -1 107408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_135_252
timestamp 1486834041
transform 1 0 28896 0 -1 107408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_135_260
timestamp 1486834041
transform 1 0 29792 0 -1 107408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_135_262
timestamp 1486834041
transform 1 0 30016 0 -1 107408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_2
timestamp 1486834041
transform 1 0 896 0 1 107408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_37
timestamp 1486834041
transform 1 0 4816 0 1 107408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_136_44
timestamp 1486834041
transform 1 0 5600 0 1 107408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_46
timestamp 1486834041
transform 1 0 5824 0 1 107408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_136_107
timestamp 1486834041
transform 1 0 12656 0 1 107408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_111
timestamp 1486834041
transform 1 0 13104 0 1 107408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_136_156
timestamp 1486834041
transform 1 0 18144 0 1 107408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_136_172
timestamp 1486834041
transform 1 0 19936 0 1 107408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_174
timestamp 1486834041
transform 1 0 20160 0 1 107408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_136_177
timestamp 1486834041
transform 1 0 20496 0 1 107408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_136_209
timestamp 1486834041
transform 1 0 24080 0 1 107408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_217
timestamp 1486834041
transform 1 0 24976 0 1 107408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_136_220
timestamp 1486834041
transform 1 0 25312 0 1 107408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_136_236
timestamp 1486834041
transform 1 0 27104 0 1 107408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_136_244
timestamp 1486834041
transform 1 0 28000 0 1 107408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_136_247
timestamp 1486834041
transform 1 0 28336 0 1 107408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_2
timestamp 1486834041
transform 1 0 896 0 -1 108976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_69
timestamp 1486834041
transform 1 0 8400 0 -1 108976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_137_122
timestamp 1486834041
transform 1 0 14336 0 -1 108976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_124
timestamp 1486834041
transform 1 0 14560 0 -1 108976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_133
timestamp 1486834041
transform 1 0 15568 0 -1 108976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_137_162
timestamp 1486834041
transform 1 0 18816 0 -1 108976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_137_194
timestamp 1486834041
transform 1 0 22400 0 -1 108976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_202
timestamp 1486834041
transform 1 0 23296 0 -1 108976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_205
timestamp 1486834041
transform 1 0 23632 0 -1 108976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_209
timestamp 1486834041
transform 1 0 24080 0 -1 108976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_212
timestamp 1486834041
transform 1 0 24416 0 -1 108976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_137_216
timestamp 1486834041
transform 1 0 24864 0 -1 108976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_137_220
timestamp 1486834041
transform 1 0 25312 0 -1 108976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_137_224
timestamp 1486834041
transform 1 0 25760 0 -1 108976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_226
timestamp 1486834041
transform 1 0 25984 0 -1 108976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_137_229
timestamp 1486834041
transform 1 0 26320 0 -1 108976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_137_245
timestamp 1486834041
transform 1 0 28112 0 -1 108976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_137_253
timestamp 1486834041
transform 1 0 29008 0 -1 108976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_255
timestamp 1486834041
transform 1 0 29232 0 -1 108976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_137_262
timestamp 1486834041
transform 1 0 30016 0 -1 108976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_22
timestamp 1486834041
transform 1 0 3136 0 1 108976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_37
timestamp 1486834041
transform 1 0 4816 0 1 108976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_85
timestamp 1486834041
transform 1 0 10192 0 1 108976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_89
timestamp 1486834041
transform 1 0 10640 0 1 108976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_104
timestamp 1486834041
transform 1 0 12320 0 1 108976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_107
timestamp 1486834041
transform 1 0 12656 0 1 108976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_138_177
timestamp 1486834041
transform 1 0 20496 0 1 108976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_193
timestamp 1486834041
transform 1 0 22288 0 1 108976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_138_205
timestamp 1486834041
transform 1 0 23632 0 1 108976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_213
timestamp 1486834041
transform 1 0 24528 0 1 108976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_138_217
timestamp 1486834041
transform 1 0 24976 0 1 108976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_221
timestamp 1486834041
transform 1 0 25424 0 1 108976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_138_225
timestamp 1486834041
transform 1 0 25872 0 1 108976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_229
timestamp 1486834041
transform 1 0 26320 0 1 108976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_138_237
timestamp 1486834041
transform 1 0 27216 0 1 108976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_138_247
timestamp 1486834041
transform 1 0 28336 0 1 108976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_255
timestamp 1486834041
transform 1 0 29232 0 1 108976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_138_262
timestamp 1486834041
transform 1 0 30016 0 1 108976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_138_266
timestamp 1486834041
transform 1 0 30464 0 1 108976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_138_268
timestamp 1486834041
transform 1 0 30688 0 1 108976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_139_2
timestamp 1486834041
transform 1 0 896 0 -1 110544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_4
timestamp 1486834041
transform 1 0 1120 0 -1 110544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_31
timestamp 1486834041
transform 1 0 4144 0 -1 110544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_139_67
timestamp 1486834041
transform 1 0 8176 0 -1 110544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_69
timestamp 1486834041
transform 1 0 8400 0 -1 110544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_139_80
timestamp 1486834041
transform 1 0 9632 0 -1 110544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_198
timestamp 1486834041
transform 1 0 22848 0 -1 110544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_202
timestamp 1486834041
transform 1 0 23296 0 -1 110544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_209
timestamp 1486834041
transform 1 0 24080 0 -1 110544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_139_224
timestamp 1486834041
transform 1 0 25760 0 -1 110544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_139_243
timestamp 1486834041
transform 1 0 27888 0 -1 110544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_139_259
timestamp 1486834041
transform 1 0 29680 0 -1 110544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_22
timestamp 1486834041
transform 1 0 3136 0 1 110544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_37
timestamp 1486834041
transform 1 0 4816 0 1 110544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_81
timestamp 1486834041
transform 1 0 9744 0 1 110544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_98
timestamp 1486834041
transform 1 0 11648 0 1 110544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_107
timestamp 1486834041
transform 1 0 12656 0 1 110544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_111
timestamp 1486834041
transform 1 0 13104 0 1 110544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_140_172
timestamp 1486834041
transform 1 0 19936 0 1 110544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_174
timestamp 1486834041
transform 1 0 20160 0 1 110544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_140_225
timestamp 1486834041
transform 1 0 25872 0 1 110544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_140_241
timestamp 1486834041
transform 1 0 27664 0 1 110544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_140_247
timestamp 1486834041
transform 1 0 28336 0 1 110544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_255
timestamp 1486834041
transform 1 0 29232 0 1 110544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_140_262
timestamp 1486834041
transform 1 0 30016 0 1 110544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_141_68
timestamp 1486834041
transform 1 0 8288 0 -1 112112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_78
timestamp 1486834041
transform 1 0 9408 0 -1 112112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_81
timestamp 1486834041
transform 1 0 9744 0 -1 112112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_141_84
timestamp 1486834041
transform 1 0 10080 0 -1 112112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_86
timestamp 1486834041
transform 1 0 10304 0 -1 112112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_95
timestamp 1486834041
transform 1 0 11312 0 -1 112112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_141_118
timestamp 1486834041
transform 1 0 13888 0 -1 112112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_200
timestamp 1486834041
transform 1 0 23072 0 -1 112112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_141_207
timestamp 1486834041
transform 1 0 23856 0 -1 112112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_209
timestamp 1486834041
transform 1 0 24080 0 -1 112112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_141_224
timestamp 1486834041
transform 1 0 25760 0 -1 112112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_2
timestamp 1486834041
transform 1 0 896 0 1 112112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_37
timestamp 1486834041
transform 1 0 4816 0 1 112112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_142_50
timestamp 1486834041
transform 1 0 6272 0 1 112112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_142_52
timestamp 1486834041
transform 1 0 6496 0 1 112112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_142_173
timestamp 1486834041
transform 1 0 20048 0 1 112112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_241
timestamp 1486834041
transform 1 0 27664 0 1 112112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_142_265
timestamp 1486834041
transform 1 0 30352 0 1 112112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_2
timestamp 1486834041
transform 1 0 896 0 -1 113680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_9
timestamp 1486834041
transform 1 0 1680 0 -1 113680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_13
timestamp 1486834041
transform 1 0 2128 0 -1 113680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_143_70
timestamp 1486834041
transform 1 0 8512 0 -1 113680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_72
timestamp 1486834041
transform 1 0 8736 0 -1 113680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_95
timestamp 1486834041
transform 1 0 11312 0 -1 113680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_143_258
timestamp 1486834041
transform 1 0 29568 0 -1 113680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_143_265
timestamp 1486834041
transform 1 0 30352 0 -1 113680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output1
timestamp 1486834041
transform 1 0 30128 0 -1 21168
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output2
timestamp 1486834041
transform 1 0 30128 0 1 21168
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output3
timestamp 1486834041
transform 1 0 30128 0 -1 22736
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output4
timestamp 1486834041
transform 1 0 30128 0 1 22736
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output5
timestamp 1486834041
transform 1 0 30128 0 -1 24304
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output6
timestamp 1486834041
transform 1 0 30128 0 1 24304
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output7
timestamp 1486834041
transform 1 0 30128 0 -1 25872
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output8
timestamp 1486834041
transform 1 0 30128 0 -1 27440
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output9
timestamp 1486834041
transform 1 0 30128 0 1 27440
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output10
timestamp 1486834041
transform 1 0 30128 0 -1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output11
timestamp 1486834041
transform 1 0 30128 0 1 35280
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output12
timestamp 1486834041
transform 1 0 30128 0 -1 29008
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output13
timestamp 1486834041
transform 1 0 30128 0 1 29008
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output14
timestamp 1486834041
transform 1 0 30128 0 -1 30576
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output15
timestamp 1486834041
transform 1 0 30128 0 1 30576
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output16
timestamp 1486834041
transform 1 0 30128 0 -1 32144
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output17
timestamp 1486834041
transform 1 0 30128 0 -1 33712
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output18
timestamp 1486834041
transform 1 0 30128 0 1 33712
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output19
timestamp 1486834041
transform 1 0 30128 0 -1 35280
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output20
timestamp 1486834041
transform 1 0 30128 0 1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output21
timestamp 1486834041
transform 1 0 30128 0 -1 79184
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output22
timestamp 1486834041
transform 1 0 30128 0 -1 90160
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output23
timestamp 1486834041
transform 1 0 30128 0 -1 91728
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output24
timestamp 1486834041
transform 1 0 30128 0 1 91728
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output25
timestamp 1486834041
transform 1 0 30128 0 -1 93296
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output26
timestamp 1486834041
transform 1 0 30128 0 -1 94864
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output27
timestamp 1486834041
transform 1 0 30128 0 1 94864
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output28
timestamp 1486834041
transform 1 0 30128 0 1 96432
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output29
timestamp 1486834041
transform 1 0 30128 0 -1 98000
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output30
timestamp 1486834041
transform 1 0 30128 0 -1 99568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output31
timestamp 1486834041
transform 1 0 30128 0 1 99568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output32
timestamp 1486834041
transform 1 0 30128 0 1 79184
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output33
timestamp 1486834041
transform 1 0 30128 0 -1 101136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output34
timestamp 1486834041
transform 1 0 30128 0 -1 102704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output35
timestamp 1486834041
transform 1 0 30128 0 1 102704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output36
timestamp 1486834041
transform 1 0 30128 0 1 104272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output37
timestamp 1486834041
transform 1 0 30128 0 -1 105840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output38
timestamp 1486834041
transform 1 0 30128 0 -1 107408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output39
timestamp 1486834041
transform 1 0 30128 0 1 107408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output40
timestamp 1486834041
transform 1 0 30128 0 -1 108976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output41
timestamp 1486834041
transform 1 0 30128 0 -1 110544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output42
timestamp 1486834041
transform 1 0 30128 0 1 110544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output43
timestamp 1486834041
transform 1 0 30128 0 1 80752
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output44
timestamp 1486834041
transform 1 0 30128 0 -1 112112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output45
timestamp 1486834041
transform 1 0 29456 0 -1 112112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output46
timestamp 1486834041
transform 1 0 30128 0 -1 82320
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output47
timestamp 1486834041
transform 1 0 30128 0 -1 83888
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output48
timestamp 1486834041
transform 1 0 30128 0 1 83888
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output49
timestamp 1486834041
transform 1 0 30128 0 -1 85456
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output50
timestamp 1486834041
transform 1 0 30128 0 -1 87024
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output51
timestamp 1486834041
transform 1 0 30128 0 1 87024
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output52
timestamp 1486834041
transform 1 0 30128 0 1 88592
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output53
timestamp 1486834041
transform -1 0 25200 0 1 112112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output54
timestamp 1486834041
transform -1 0 29008 0 1 112112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output55
timestamp 1486834041
transform -1 0 29568 0 -1 113680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output56
timestamp 1486834041
transform -1 0 28224 0 -1 113680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output57
timestamp 1486834041
transform -1 0 29680 0 1 112112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output58
timestamp 1486834041
transform -1 0 29456 0 -1 112112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output59
timestamp 1486834041
transform -1 0 28112 0 -1 112112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output60
timestamp 1486834041
transform -1 0 28784 0 -1 112112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output61
timestamp 1486834041
transform -1 0 30352 0 1 112112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output62
timestamp 1486834041
transform -1 0 27888 0 -1 110544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output63
timestamp 1486834041
transform -1 0 30352 0 -1 113680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output64
timestamp 1486834041
transform -1 0 23856 0 1 112112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output65
timestamp 1486834041
transform -1 0 24528 0 1 112112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output66
timestamp 1486834041
transform -1 0 25984 0 -1 113680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output67
timestamp 1486834041
transform -1 0 26096 0 1 112112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output68
timestamp 1486834041
transform -1 0 26656 0 -1 113680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output69
timestamp 1486834041
transform -1 0 26992 0 1 112112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output70
timestamp 1486834041
transform -1 0 27328 0 -1 113680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output71
timestamp 1486834041
transform -1 0 27664 0 1 112112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output72
timestamp 1486834041
transform -1 0 28896 0 -1 113680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output73
timestamp 1486834041
transform -1 0 20160 0 -1 110544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output74
timestamp 1486834041
transform 1 0 4928 0 1 101136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output75
timestamp 1486834041
transform -1 0 23184 0 1 112112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output76
timestamp 1486834041
transform -1 0 7840 0 -1 101136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output77
timestamp 1486834041
transform 1 0 1232 0 -1 110544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output78
timestamp 1486834041
transform 1 0 5488 0 1 102704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output79
timestamp 1486834041
transform 1 0 4816 0 1 104272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output80
timestamp 1486834041
transform 1 0 1008 0 1 112112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output81
timestamp 1486834041
transform 1 0 3920 0 1 102704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output82
timestamp 1486834041
transform 1 0 3920 0 1 108976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output83
timestamp 1486834041
transform 1 0 3248 0 1 104272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output84
timestamp 1486834041
transform -1 0 8512 0 -1 102704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output85
timestamp 1486834041
transform 1 0 1008 0 -1 113680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output86
timestamp 1486834041
transform 1 0 4928 0 1 107408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output87
timestamp 1486834041
transform -1 0 24416 0 -1 113680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output88
timestamp 1486834041
transform -1 0 15344 0 -1 108976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output89
timestamp 1486834041
transform -1 0 20048 0 1 112112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output90
timestamp 1486834041
transform -1 0 22512 0 1 112112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output91
timestamp 1486834041
transform -1 0 14560 0 1 107408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output92
timestamp 1486834041
transform -1 0 19040 0 -1 113680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output93
timestamp 1486834041
transform -1 0 23520 0 -1 113680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output94
timestamp 1486834041
transform -1 0 15904 0 -1 113680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output95
timestamp 1486834041
transform -1 0 22848 0 -1 113680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output96
timestamp 1486834041
transform -1 0 19712 0 -1 113680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output97
timestamp 1486834041
transform -1 0 21840 0 1 112112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output98
timestamp 1486834041
transform -1 0 15232 0 -1 113680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output99
timestamp 1486834041
transform 1 0 11760 0 1 112112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output100
timestamp 1486834041
transform -1 0 12320 0 1 108976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output101
timestamp 1486834041
transform 1 0 4704 0 -1 113680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output102
timestamp 1486834041
transform 1 0 8736 0 -1 112112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output103
timestamp 1486834041
transform 1 0 8736 0 -1 105840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output104
timestamp 1486834041
transform 1 0 9632 0 -1 107408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output105
timestamp 1486834041
transform 1 0 3248 0 1 110544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output106
timestamp 1486834041
transform 1 0 10976 0 1 108976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output107
timestamp 1486834041
transform 1 0 7616 0 -1 112112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output108
timestamp 1486834041
transform -1 0 21168 0 1 112112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output109
timestamp 1486834041
transform -1 0 25088 0 -1 113680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output110
timestamp 1486834041
transform -1 0 2240 0 -1 58800
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output111
timestamp 1486834041
transform -1 0 1568 0 -1 58800
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output112
timestamp 1486834041
transform -1 0 1568 0 1 58800
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output113
timestamp 1486834041
transform -1 0 3024 0 1 58800
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output114
timestamp 1486834041
transform -1 0 1568 0 1 60368
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output115
timestamp 1486834041
transform -1 0 1568 0 -1 61936
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output116
timestamp 1486834041
transform -1 0 1568 0 1 63504
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output117
timestamp 1486834041
transform -1 0 1568 0 1 57232
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output118
timestamp 1486834041
transform -1 0 1568 0 1 65072
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output119
timestamp 1486834041
transform -1 0 4480 0 1 63504
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output120
timestamp 1486834041
transform -1 0 1568 0 -1 68208
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output121
timestamp 1486834041
transform -1 0 1568 0 1 68208
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output122
timestamp 1486834041
transform -1 0 1568 0 -1 69776
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output123
timestamp 1486834041
transform -1 0 6160 0 -1 65072
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output124
timestamp 1486834041
transform -1 0 1568 0 1 71344
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output125
timestamp 1486834041
transform -1 0 4592 0 1 65072
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output126
timestamp 1486834041
transform -1 0 5488 0 1 65072
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output127
timestamp 1486834041
transform -1 0 4480 0 1 68208
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output128
timestamp 1486834041
transform -1 0 1568 0 -1 72912
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output129
timestamp 1486834041
transform -1 0 2240 0 1 71344
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output130
timestamp 1486834041
transform -1 0 7728 0 -1 74480
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output131
timestamp 1486834041
transform -1 0 2352 0 1 85456
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output132
timestamp 1486834041
transform -1 0 7840 0 -1 82320
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output133
timestamp 1486834041
transform -1 0 6160 0 1 76048
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output134
timestamp 1486834041
transform -1 0 4480 0 -1 83888
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output135
timestamp 1486834041
transform -1 0 4480 0 1 80752
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output136
timestamp 1486834041
transform -1 0 1568 0 -1 85456
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output137
timestamp 1486834041
transform -1 0 4592 0 1 79184
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output138
timestamp 1486834041
transform -1 0 1568 0 1 85456
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output139
timestamp 1486834041
transform -1 0 5488 0 1 80752
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output140
timestamp 1486834041
transform -1 0 8288 0 1 79184
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output141
timestamp 1486834041
transform -1 0 8512 0 -1 82320
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output142
timestamp 1486834041
transform -1 0 1568 0 -1 74480
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output143
timestamp 1486834041
transform -1 0 6160 0 1 72912
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output144
timestamp 1486834041
transform -1 0 6832 0 1 72912
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output145
timestamp 1486834041
transform -1 0 4592 0 1 74480
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output146
timestamp 1486834041
transform -1 0 4480 0 1 77616
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output147
timestamp 1486834041
transform -1 0 5712 0 1 74480
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output148
timestamp 1486834041
transform -1 0 7056 0 -1 74480
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output149
timestamp 1486834041
transform -1 0 1568 0 -1 76048
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output150
timestamp 1486834041
transform -1 0 8512 0 -1 69776
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output151
timestamp 1486834041
transform -1 0 1568 0 1 76048
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output152
timestamp 1486834041
transform -1 0 5488 0 1 71344
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output153
timestamp 1486834041
transform -1 0 9408 0 -1 71344
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output154
timestamp 1486834041
transform -1 0 1568 0 -1 77616
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output155
timestamp 1486834041
transform -1 0 8400 0 -1 72912
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output156
timestamp 1486834041
transform -1 0 6048 0 -1 79184
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output157
timestamp 1486834041
transform -1 0 2240 0 -1 77616
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output158
timestamp 1486834041
transform 1 0 30128 0 1 39984
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output159
timestamp 1486834041
transform 1 0 30128 0 1 50960
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output160
timestamp 1486834041
transform 1 0 30128 0 1 52528
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output161
timestamp 1486834041
transform 1 0 30128 0 -1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output162
timestamp 1486834041
transform 1 0 30128 0 1 54096
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output163
timestamp 1486834041
transform 1 0 30128 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output164
timestamp 1486834041
transform 1 0 30128 0 -1 57232
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output165
timestamp 1486834041
transform 1 0 30128 0 -1 58800
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output166
timestamp 1486834041
transform 1 0 30128 0 1 58800
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output167
timestamp 1486834041
transform 1 0 30128 0 1 60368
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output168
timestamp 1486834041
transform 1 0 30128 0 -1 61936
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output169
timestamp 1486834041
transform 1 0 30128 0 -1 41552
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output170
timestamp 1486834041
transform 1 0 30128 0 -1 63504
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output171
timestamp 1486834041
transform 1 0 30128 0 1 63504
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output172
timestamp 1486834041
transform 1 0 30128 0 -1 65072
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output173
timestamp 1486834041
transform 1 0 30128 0 -1 66640
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output174
timestamp 1486834041
transform 1 0 30128 0 1 66640
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output175
timestamp 1486834041
transform 1 0 30128 0 1 68208
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output176
timestamp 1486834041
transform 1 0 30128 0 -1 69776
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output177
timestamp 1486834041
transform 1 0 30128 0 -1 71344
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output178
timestamp 1486834041
transform 1 0 30128 0 1 71344
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output179
timestamp 1486834041
transform 1 0 30128 0 -1 72912
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output180
timestamp 1486834041
transform 1 0 30128 0 -1 43120
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output181
timestamp 1486834041
transform 1 0 30128 0 -1 74480
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output182
timestamp 1486834041
transform 1 0 30128 0 1 74480
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output183
timestamp 1486834041
transform 1 0 30128 0 1 43120
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output184
timestamp 1486834041
transform 1 0 30128 0 1 44688
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output185
timestamp 1486834041
transform 1 0 30128 0 -1 46256
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output186
timestamp 1486834041
transform 1 0 30128 0 -1 47824
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output187
timestamp 1486834041
transform 1 0 30128 0 1 47824
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output188
timestamp 1486834041
transform 1 0 30128 0 -1 49392
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output189
timestamp 1486834041
transform 1 0 30128 0 -1 50960
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output190
timestamp 1486834041
transform 1 0 7840 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output191
timestamp 1486834041
transform 1 0 10416 0 1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output192
timestamp 1486834041
transform 1 0 11088 0 1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output193
timestamp 1486834041
transform 1 0 13104 0 1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output194
timestamp 1486834041
transform 1 0 13776 0 1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output195
timestamp 1486834041
transform 1 0 4704 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output196
timestamp 1486834041
transform 1 0 9072 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output197
timestamp 1486834041
transform 1 0 5376 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output198
timestamp 1486834041
transform 1 0 7840 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output199
timestamp 1486834041
transform 1 0 9072 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output200
timestamp 1486834041
transform 1 0 11760 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output201
timestamp 1486834041
transform 1 0 15680 0 -1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output202
timestamp 1486834041
transform 1 0 15232 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output203
timestamp 1486834041
transform -1 0 17136 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output204
timestamp 1486834041
transform -1 0 17360 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output205
timestamp 1486834041
transform -1 0 19824 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output206
timestamp 1486834041
transform -1 0 22848 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output207
timestamp 1486834041
transform -1 0 23520 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output208
timestamp 1486834041
transform -1 0 26656 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output209
timestamp 1486834041
transform -1 0 27328 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output210
timestamp 1486834041
transform -1 0 28224 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output211
timestamp 1486834041
transform -1 0 24192 0 -1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output212
timestamp 1486834041
transform -1 0 25760 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output213
timestamp 1486834041
transform -1 0 29568 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output214
timestamp 1486834041
transform -1 0 27664 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output215
timestamp 1486834041
transform -1 0 28672 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output216
timestamp 1486834041
transform -1 0 25648 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output217
timestamp 1486834041
transform -1 0 26320 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output218
timestamp 1486834041
transform -1 0 28896 0 1 784
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output219
timestamp 1486834041
transform -1 0 27328 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output220
timestamp 1486834041
transform -1 0 27104 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output221
timestamp 1486834041
transform -1 0 26432 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output222
timestamp 1486834041
transform -1 0 25648 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output223
timestamp 1486834041
transform -1 0 23520 0 -1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output224
timestamp 1486834041
transform -1 0 28000 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output225
timestamp 1486834041
transform -1 0 26992 0 1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output226
timestamp 1486834041
transform -1 0 16240 0 1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output227
timestamp 1486834041
transform -1 0 17248 0 -1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output228
timestamp 1486834041
transform -1 0 12432 0 1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output229
timestamp 1486834041
transform -1 0 15792 0 -1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output230
timestamp 1486834041
transform -1 0 15120 0 -1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output231
timestamp 1486834041
transform -1 0 10080 0 -1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output232
timestamp 1486834041
transform -1 0 12432 0 1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output233
timestamp 1486834041
transform -1 0 9408 0 -1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output234
timestamp 1486834041
transform -1 0 15680 0 -1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output235
timestamp 1486834041
transform -1 0 11088 0 1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output236
timestamp 1486834041
transform -1 0 9408 0 -1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output237
timestamp 1486834041
transform -1 0 10080 0 -1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output238
timestamp 1486834041
transform -1 0 9408 0 -1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output239
timestamp 1486834041
transform -1 0 9408 0 -1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output240
timestamp 1486834041
transform -1 0 7280 0 -1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output241
timestamp 1486834041
transform -1 0 3024 0 -1 2352
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output242
timestamp 1486834041
transform -1 0 7168 0 -1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output243
timestamp 1486834041
transform -1 0 8512 0 -1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output244
timestamp 1486834041
transform -1 0 7840 0 -1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output245
timestamp 1486834041
transform -1 0 7168 0 -1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output246
timestamp 1486834041
transform -1 0 6160 0 1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output247
timestamp 1486834041
transform -1 0 2240 0 1 22736
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output248
timestamp 1486834041
transform -1 0 1568 0 1 22736
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output249
timestamp 1486834041
transform -1 0 5152 0 -1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output250
timestamp 1486834041
transform -1 0 3808 0 1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output251
timestamp 1486834041
transform -1 0 4480 0 1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output252
timestamp 1486834041
transform -1 0 5488 0 1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output253
timestamp 1486834041
transform -1 0 6048 0 -1 19600
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output254
timestamp 1486834041
transform -1 0 4480 0 1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output255
timestamp 1486834041
transform -1 0 3808 0 1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output256
timestamp 1486834041
transform -1 0 4256 0 1 21168
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output257
timestamp 1486834041
transform -1 0 1568 0 -1 24304
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output258
timestamp 1486834041
transform -1 0 2240 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output259
timestamp 1486834041
transform -1 0 4480 0 1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output260
timestamp 1486834041
transform -1 0 5488 0 1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output261
timestamp 1486834041
transform -1 0 1568 0 -1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output262
timestamp 1486834041
transform -1 0 2240 0 1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output263
timestamp 1486834041
transform -1 0 1568 0 1 8624
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output264
timestamp 1486834041
transform -1 0 5488 0 1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output265
timestamp 1486834041
transform -1 0 5488 0 1 7056
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output266
timestamp 1486834041
transform -1 0 1568 0 -1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output267
timestamp 1486834041
transform -1 0 8176 0 1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output268
timestamp 1486834041
transform -1 0 2240 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output269
timestamp 1486834041
transform -1 0 8288 0 -1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output270
timestamp 1486834041
transform -1 0 1568 0 1 3920
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output271
timestamp 1486834041
transform -1 0 2240 0 -1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output272
timestamp 1486834041
transform -1 0 1568 0 -1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output273
timestamp 1486834041
transform -1 0 1568 0 1 5488
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output274
timestamp 1486834041
transform 1 0 30128 0 -1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output275
timestamp 1486834041
transform 1 0 30128 0 -1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output276
timestamp 1486834041
transform 1 0 30128 0 1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output277
timestamp 1486834041
transform 1 0 30128 0 -1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output278
timestamp 1486834041
transform 1 0 30128 0 1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output279
timestamp 1486834041
transform 1 0 30128 0 -1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output280
timestamp 1486834041
transform 1 0 30128 0 1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output281
timestamp 1486834041
transform 1 0 30128 0 -1 19600
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_144
timestamp 1486834041
transform 1 0 672 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1486834041
transform -1 0 31024 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_145
timestamp 1486834041
transform 1 0 672 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1486834041
transform -1 0 31024 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_146
timestamp 1486834041
transform 1 0 672 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1486834041
transform -1 0 31024 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_147
timestamp 1486834041
transform 1 0 672 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1486834041
transform -1 0 31024 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_148
timestamp 1486834041
transform 1 0 672 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1486834041
transform -1 0 31024 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_149
timestamp 1486834041
transform 1 0 672 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1486834041
transform -1 0 31024 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_150
timestamp 1486834041
transform 1 0 672 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1486834041
transform -1 0 31024 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_151
timestamp 1486834041
transform 1 0 672 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1486834041
transform -1 0 31024 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_152
timestamp 1486834041
transform 1 0 672 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1486834041
transform -1 0 31024 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_153
timestamp 1486834041
transform 1 0 672 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1486834041
transform -1 0 31024 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_154
timestamp 1486834041
transform 1 0 672 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1486834041
transform -1 0 31024 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_155
timestamp 1486834041
transform 1 0 672 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1486834041
transform -1 0 31024 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_156
timestamp 1486834041
transform 1 0 672 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1486834041
transform -1 0 31024 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_157
timestamp 1486834041
transform 1 0 672 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1486834041
transform -1 0 31024 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_158
timestamp 1486834041
transform 1 0 672 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1486834041
transform -1 0 31024 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_159
timestamp 1486834041
transform 1 0 672 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1486834041
transform -1 0 31024 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_160
timestamp 1486834041
transform 1 0 672 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1486834041
transform -1 0 31024 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_161
timestamp 1486834041
transform 1 0 672 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1486834041
transform -1 0 31024 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_162
timestamp 1486834041
transform 1 0 672 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1486834041
transform -1 0 31024 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_163
timestamp 1486834041
transform 1 0 672 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1486834041
transform -1 0 31024 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_164
timestamp 1486834041
transform 1 0 672 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1486834041
transform -1 0 31024 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_165
timestamp 1486834041
transform 1 0 672 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1486834041
transform -1 0 31024 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_166
timestamp 1486834041
transform 1 0 672 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1486834041
transform -1 0 31024 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_167
timestamp 1486834041
transform 1 0 672 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1486834041
transform -1 0 31024 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_168
timestamp 1486834041
transform 1 0 672 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1486834041
transform -1 0 31024 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_169
timestamp 1486834041
transform 1 0 672 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1486834041
transform -1 0 31024 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_170
timestamp 1486834041
transform 1 0 672 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1486834041
transform -1 0 31024 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_171
timestamp 1486834041
transform 1 0 672 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1486834041
transform -1 0 31024 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_172
timestamp 1486834041
transform 1 0 672 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1486834041
transform -1 0 31024 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_173
timestamp 1486834041
transform 1 0 672 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1486834041
transform -1 0 31024 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_174
timestamp 1486834041
transform 1 0 672 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1486834041
transform -1 0 31024 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_175
timestamp 1486834041
transform 1 0 672 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1486834041
transform -1 0 31024 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_176
timestamp 1486834041
transform 1 0 672 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1486834041
transform -1 0 31024 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_177
timestamp 1486834041
transform 1 0 672 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1486834041
transform -1 0 31024 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_178
timestamp 1486834041
transform 1 0 672 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1486834041
transform -1 0 31024 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_179
timestamp 1486834041
transform 1 0 672 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1486834041
transform -1 0 31024 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_180
timestamp 1486834041
transform 1 0 672 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1486834041
transform -1 0 31024 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_181
timestamp 1486834041
transform 1 0 672 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1486834041
transform -1 0 31024 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_182
timestamp 1486834041
transform 1 0 672 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1486834041
transform -1 0 31024 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_183
timestamp 1486834041
transform 1 0 672 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1486834041
transform -1 0 31024 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_184
timestamp 1486834041
transform 1 0 672 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1486834041
transform -1 0 31024 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_185
timestamp 1486834041
transform 1 0 672 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1486834041
transform -1 0 31024 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_186
timestamp 1486834041
transform 1 0 672 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1486834041
transform -1 0 31024 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_187
timestamp 1486834041
transform 1 0 672 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1486834041
transform -1 0 31024 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_188
timestamp 1486834041
transform 1 0 672 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1486834041
transform -1 0 31024 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_189
timestamp 1486834041
transform 1 0 672 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1486834041
transform -1 0 31024 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_190
timestamp 1486834041
transform 1 0 672 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1486834041
transform -1 0 31024 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_191
timestamp 1486834041
transform 1 0 672 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1486834041
transform -1 0 31024 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_192
timestamp 1486834041
transform 1 0 672 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1486834041
transform -1 0 31024 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_193
timestamp 1486834041
transform 1 0 672 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1486834041
transform -1 0 31024 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_194
timestamp 1486834041
transform 1 0 672 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1486834041
transform -1 0 31024 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_195
timestamp 1486834041
transform 1 0 672 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1486834041
transform -1 0 31024 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_196
timestamp 1486834041
transform 1 0 672 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1486834041
transform -1 0 31024 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_197
timestamp 1486834041
transform 1 0 672 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1486834041
transform -1 0 31024 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_198
timestamp 1486834041
transform 1 0 672 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1486834041
transform -1 0 31024 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_199
timestamp 1486834041
transform 1 0 672 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1486834041
transform -1 0 31024 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_200
timestamp 1486834041
transform 1 0 672 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1486834041
transform -1 0 31024 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_201
timestamp 1486834041
transform 1 0 672 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1486834041
transform -1 0 31024 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_202
timestamp 1486834041
transform 1 0 672 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1486834041
transform -1 0 31024 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_203
timestamp 1486834041
transform 1 0 672 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1486834041
transform -1 0 31024 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_204
timestamp 1486834041
transform 1 0 672 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1486834041
transform -1 0 31024 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_205
timestamp 1486834041
transform 1 0 672 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1486834041
transform -1 0 31024 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Left_206
timestamp 1486834041
transform 1 0 672 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Right_62
timestamp 1486834041
transform -1 0 31024 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Left_207
timestamp 1486834041
transform 1 0 672 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Right_63
timestamp 1486834041
transform -1 0 31024 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Left_208
timestamp 1486834041
transform 1 0 672 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Right_64
timestamp 1486834041
transform -1 0 31024 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Left_209
timestamp 1486834041
transform 1 0 672 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Right_65
timestamp 1486834041
transform -1 0 31024 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Left_210
timestamp 1486834041
transform 1 0 672 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Right_66
timestamp 1486834041
transform -1 0 31024 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Left_211
timestamp 1486834041
transform 1 0 672 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Right_67
timestamp 1486834041
transform -1 0 31024 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Left_212
timestamp 1486834041
transform 1 0 672 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Right_68
timestamp 1486834041
transform -1 0 31024 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Left_213
timestamp 1486834041
transform 1 0 672 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Right_69
timestamp 1486834041
transform -1 0 31024 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Left_214
timestamp 1486834041
transform 1 0 672 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Right_70
timestamp 1486834041
transform -1 0 31024 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_71_Left_215
timestamp 1486834041
transform 1 0 672 0 -1 57232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_71_Right_71
timestamp 1486834041
transform -1 0 31024 0 -1 57232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_72_Left_216
timestamp 1486834041
transform 1 0 672 0 1 57232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_72_Right_72
timestamp 1486834041
transform -1 0 31024 0 1 57232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_73_Left_217
timestamp 1486834041
transform 1 0 672 0 -1 58800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_73_Right_73
timestamp 1486834041
transform -1 0 31024 0 -1 58800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_74_Left_218
timestamp 1486834041
transform 1 0 672 0 1 58800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_74_Right_74
timestamp 1486834041
transform -1 0 31024 0 1 58800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_75_Left_219
timestamp 1486834041
transform 1 0 672 0 -1 60368
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_75_Right_75
timestamp 1486834041
transform -1 0 31024 0 -1 60368
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_76_Left_220
timestamp 1486834041
transform 1 0 672 0 1 60368
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_76_Right_76
timestamp 1486834041
transform -1 0 31024 0 1 60368
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_77_Left_221
timestamp 1486834041
transform 1 0 672 0 -1 61936
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_77_Right_77
timestamp 1486834041
transform -1 0 31024 0 -1 61936
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_78_Left_222
timestamp 1486834041
transform 1 0 672 0 1 61936
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_78_Right_78
timestamp 1486834041
transform -1 0 31024 0 1 61936
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_79_Left_223
timestamp 1486834041
transform 1 0 672 0 -1 63504
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_79_Right_79
timestamp 1486834041
transform -1 0 31024 0 -1 63504
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_80_Left_224
timestamp 1486834041
transform 1 0 672 0 1 63504
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_80_Right_80
timestamp 1486834041
transform -1 0 31024 0 1 63504
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_81_Left_225
timestamp 1486834041
transform 1 0 672 0 -1 65072
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_81_Right_81
timestamp 1486834041
transform -1 0 31024 0 -1 65072
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_82_Left_226
timestamp 1486834041
transform 1 0 672 0 1 65072
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_82_Right_82
timestamp 1486834041
transform -1 0 31024 0 1 65072
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_83_Left_227
timestamp 1486834041
transform 1 0 672 0 -1 66640
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_83_Right_83
timestamp 1486834041
transform -1 0 31024 0 -1 66640
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_84_Left_228
timestamp 1486834041
transform 1 0 672 0 1 66640
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_84_Right_84
timestamp 1486834041
transform -1 0 31024 0 1 66640
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_85_Left_229
timestamp 1486834041
transform 1 0 672 0 -1 68208
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_85_Right_85
timestamp 1486834041
transform -1 0 31024 0 -1 68208
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_86_Left_230
timestamp 1486834041
transform 1 0 672 0 1 68208
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_86_Right_86
timestamp 1486834041
transform -1 0 31024 0 1 68208
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_87_Left_231
timestamp 1486834041
transform 1 0 672 0 -1 69776
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_87_Right_87
timestamp 1486834041
transform -1 0 31024 0 -1 69776
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_88_Left_232
timestamp 1486834041
transform 1 0 672 0 1 69776
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_88_Right_88
timestamp 1486834041
transform -1 0 31024 0 1 69776
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_89_Left_233
timestamp 1486834041
transform 1 0 672 0 -1 71344
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_89_Right_89
timestamp 1486834041
transform -1 0 31024 0 -1 71344
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_90_Left_234
timestamp 1486834041
transform 1 0 672 0 1 71344
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_90_Right_90
timestamp 1486834041
transform -1 0 31024 0 1 71344
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_91_Left_235
timestamp 1486834041
transform 1 0 672 0 -1 72912
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_91_Right_91
timestamp 1486834041
transform -1 0 31024 0 -1 72912
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_92_Left_236
timestamp 1486834041
transform 1 0 672 0 1 72912
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_92_Right_92
timestamp 1486834041
transform -1 0 31024 0 1 72912
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_93_Left_237
timestamp 1486834041
transform 1 0 672 0 -1 74480
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_93_Right_93
timestamp 1486834041
transform -1 0 31024 0 -1 74480
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_94_Left_238
timestamp 1486834041
transform 1 0 672 0 1 74480
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_94_Right_94
timestamp 1486834041
transform -1 0 31024 0 1 74480
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_95_Left_239
timestamp 1486834041
transform 1 0 672 0 -1 76048
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_95_Right_95
timestamp 1486834041
transform -1 0 31024 0 -1 76048
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_96_Left_240
timestamp 1486834041
transform 1 0 672 0 1 76048
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_96_Right_96
timestamp 1486834041
transform -1 0 31024 0 1 76048
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_97_Left_241
timestamp 1486834041
transform 1 0 672 0 -1 77616
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_97_Right_97
timestamp 1486834041
transform -1 0 31024 0 -1 77616
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_98_Left_242
timestamp 1486834041
transform 1 0 672 0 1 77616
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_98_Right_98
timestamp 1486834041
transform -1 0 31024 0 1 77616
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_99_Left_243
timestamp 1486834041
transform 1 0 672 0 -1 79184
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_99_Right_99
timestamp 1486834041
transform -1 0 31024 0 -1 79184
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_100_Left_244
timestamp 1486834041
transform 1 0 672 0 1 79184
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_100_Right_100
timestamp 1486834041
transform -1 0 31024 0 1 79184
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_101_Left_245
timestamp 1486834041
transform 1 0 672 0 -1 80752
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_101_Right_101
timestamp 1486834041
transform -1 0 31024 0 -1 80752
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_102_Left_246
timestamp 1486834041
transform 1 0 672 0 1 80752
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_102_Right_102
timestamp 1486834041
transform -1 0 31024 0 1 80752
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_103_Left_247
timestamp 1486834041
transform 1 0 672 0 -1 82320
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_103_Right_103
timestamp 1486834041
transform -1 0 31024 0 -1 82320
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_104_Left_248
timestamp 1486834041
transform 1 0 672 0 1 82320
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_104_Right_104
timestamp 1486834041
transform -1 0 31024 0 1 82320
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_105_Left_249
timestamp 1486834041
transform 1 0 672 0 -1 83888
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_105_Right_105
timestamp 1486834041
transform -1 0 31024 0 -1 83888
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_106_Left_250
timestamp 1486834041
transform 1 0 672 0 1 83888
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_106_Right_106
timestamp 1486834041
transform -1 0 31024 0 1 83888
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_107_Left_251
timestamp 1486834041
transform 1 0 672 0 -1 85456
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_107_Right_107
timestamp 1486834041
transform -1 0 31024 0 -1 85456
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_108_Left_252
timestamp 1486834041
transform 1 0 672 0 1 85456
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_108_Right_108
timestamp 1486834041
transform -1 0 31024 0 1 85456
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_109_Left_253
timestamp 1486834041
transform 1 0 672 0 -1 87024
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_109_Right_109
timestamp 1486834041
transform -1 0 31024 0 -1 87024
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_110_Left_254
timestamp 1486834041
transform 1 0 672 0 1 87024
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_110_Right_110
timestamp 1486834041
transform -1 0 31024 0 1 87024
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_111_Left_255
timestamp 1486834041
transform 1 0 672 0 -1 88592
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_111_Right_111
timestamp 1486834041
transform -1 0 31024 0 -1 88592
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_112_Left_256
timestamp 1486834041
transform 1 0 672 0 1 88592
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_112_Right_112
timestamp 1486834041
transform -1 0 31024 0 1 88592
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_113_Left_257
timestamp 1486834041
transform 1 0 672 0 -1 90160
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_113_Right_113
timestamp 1486834041
transform -1 0 31024 0 -1 90160
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_114_Left_258
timestamp 1486834041
transform 1 0 672 0 1 90160
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_114_Right_114
timestamp 1486834041
transform -1 0 31024 0 1 90160
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_115_Left_259
timestamp 1486834041
transform 1 0 672 0 -1 91728
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_115_Right_115
timestamp 1486834041
transform -1 0 31024 0 -1 91728
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_116_Left_260
timestamp 1486834041
transform 1 0 672 0 1 91728
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_116_Right_116
timestamp 1486834041
transform -1 0 31024 0 1 91728
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_117_Left_261
timestamp 1486834041
transform 1 0 672 0 -1 93296
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_117_Right_117
timestamp 1486834041
transform -1 0 31024 0 -1 93296
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_118_Left_262
timestamp 1486834041
transform 1 0 672 0 1 93296
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_118_Right_118
timestamp 1486834041
transform -1 0 31024 0 1 93296
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_119_Left_263
timestamp 1486834041
transform 1 0 672 0 -1 94864
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_119_Right_119
timestamp 1486834041
transform -1 0 31024 0 -1 94864
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_120_Left_264
timestamp 1486834041
transform 1 0 672 0 1 94864
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_120_Right_120
timestamp 1486834041
transform -1 0 31024 0 1 94864
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_121_Left_265
timestamp 1486834041
transform 1 0 672 0 -1 96432
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_121_Right_121
timestamp 1486834041
transform -1 0 31024 0 -1 96432
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_122_Left_266
timestamp 1486834041
transform 1 0 672 0 1 96432
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_122_Right_122
timestamp 1486834041
transform -1 0 31024 0 1 96432
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_123_Left_267
timestamp 1486834041
transform 1 0 672 0 -1 98000
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_123_Right_123
timestamp 1486834041
transform -1 0 31024 0 -1 98000
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_124_Left_268
timestamp 1486834041
transform 1 0 672 0 1 98000
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_124_Right_124
timestamp 1486834041
transform -1 0 31024 0 1 98000
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_125_Left_269
timestamp 1486834041
transform 1 0 672 0 -1 99568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_125_Right_125
timestamp 1486834041
transform -1 0 31024 0 -1 99568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_126_Left_270
timestamp 1486834041
transform 1 0 672 0 1 99568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_126_Right_126
timestamp 1486834041
transform -1 0 31024 0 1 99568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_127_Left_271
timestamp 1486834041
transform 1 0 672 0 -1 101136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_127_Right_127
timestamp 1486834041
transform -1 0 31024 0 -1 101136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_128_Left_272
timestamp 1486834041
transform 1 0 672 0 1 101136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_128_Right_128
timestamp 1486834041
transform -1 0 31024 0 1 101136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_129_Left_273
timestamp 1486834041
transform 1 0 672 0 -1 102704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_129_Right_129
timestamp 1486834041
transform -1 0 31024 0 -1 102704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_130_Left_274
timestamp 1486834041
transform 1 0 672 0 1 102704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_130_Right_130
timestamp 1486834041
transform -1 0 31024 0 1 102704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_131_Left_275
timestamp 1486834041
transform 1 0 672 0 -1 104272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_131_Right_131
timestamp 1486834041
transform -1 0 31024 0 -1 104272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_132_Left_276
timestamp 1486834041
transform 1 0 672 0 1 104272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_132_Right_132
timestamp 1486834041
transform -1 0 31024 0 1 104272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_133_Left_277
timestamp 1486834041
transform 1 0 672 0 -1 105840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_133_Right_133
timestamp 1486834041
transform -1 0 31024 0 -1 105840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_134_Left_278
timestamp 1486834041
transform 1 0 672 0 1 105840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_134_Right_134
timestamp 1486834041
transform -1 0 31024 0 1 105840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_135_Left_279
timestamp 1486834041
transform 1 0 672 0 -1 107408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_135_Right_135
timestamp 1486834041
transform -1 0 31024 0 -1 107408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_136_Left_280
timestamp 1486834041
transform 1 0 672 0 1 107408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_136_Right_136
timestamp 1486834041
transform -1 0 31024 0 1 107408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_137_Left_281
timestamp 1486834041
transform 1 0 672 0 -1 108976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_137_Right_137
timestamp 1486834041
transform -1 0 31024 0 -1 108976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_138_Left_282
timestamp 1486834041
transform 1 0 672 0 1 108976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_138_Right_138
timestamp 1486834041
transform -1 0 31024 0 1 108976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_139_Left_283
timestamp 1486834041
transform 1 0 672 0 -1 110544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_139_Right_139
timestamp 1486834041
transform -1 0 31024 0 -1 110544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_140_Left_284
timestamp 1486834041
transform 1 0 672 0 1 110544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_140_Right_140
timestamp 1486834041
transform -1 0 31024 0 1 110544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_141_Left_285
timestamp 1486834041
transform 1 0 672 0 -1 112112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_141_Right_141
timestamp 1486834041
transform -1 0 31024 0 -1 112112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_142_Left_286
timestamp 1486834041
transform 1 0 672 0 1 112112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_142_Right_142
timestamp 1486834041
transform -1 0 31024 0 1 112112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_143_Left_287
timestamp 1486834041
transform 1 0 672 0 -1 113680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_143_Right_143
timestamp 1486834041
transform -1 0 31024 0 -1 113680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_288
timestamp 1486834041
transform 1 0 4480 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_289
timestamp 1486834041
transform 1 0 8288 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_290
timestamp 1486834041
transform 1 0 12096 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_291
timestamp 1486834041
transform 1 0 15904 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_292
timestamp 1486834041
transform 1 0 19712 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_293
timestamp 1486834041
transform 1 0 23520 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_294
timestamp 1486834041
transform 1 0 27328 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_295
timestamp 1486834041
transform 1 0 8512 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_296
timestamp 1486834041
transform 1 0 16352 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_297
timestamp 1486834041
transform 1 0 24192 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_298
timestamp 1486834041
transform 1 0 4592 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_299
timestamp 1486834041
transform 1 0 12432 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_300
timestamp 1486834041
transform 1 0 20272 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_301
timestamp 1486834041
transform 1 0 28112 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_302
timestamp 1486834041
transform 1 0 8512 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_303
timestamp 1486834041
transform 1 0 16352 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_304
timestamp 1486834041
transform 1 0 24192 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_305
timestamp 1486834041
transform 1 0 4592 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_306
timestamp 1486834041
transform 1 0 12432 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_307
timestamp 1486834041
transform 1 0 20272 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_308
timestamp 1486834041
transform 1 0 28112 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_309
timestamp 1486834041
transform 1 0 8512 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_310
timestamp 1486834041
transform 1 0 16352 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_311
timestamp 1486834041
transform 1 0 24192 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_312
timestamp 1486834041
transform 1 0 4592 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_313
timestamp 1486834041
transform 1 0 12432 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_314
timestamp 1486834041
transform 1 0 20272 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_315
timestamp 1486834041
transform 1 0 28112 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_316
timestamp 1486834041
transform 1 0 8512 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_317
timestamp 1486834041
transform 1 0 16352 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_318
timestamp 1486834041
transform 1 0 24192 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_319
timestamp 1486834041
transform 1 0 4592 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_320
timestamp 1486834041
transform 1 0 12432 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_321
timestamp 1486834041
transform 1 0 20272 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_322
timestamp 1486834041
transform 1 0 28112 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_323
timestamp 1486834041
transform 1 0 8512 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_324
timestamp 1486834041
transform 1 0 16352 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_325
timestamp 1486834041
transform 1 0 24192 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_326
timestamp 1486834041
transform 1 0 4592 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_327
timestamp 1486834041
transform 1 0 12432 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_328
timestamp 1486834041
transform 1 0 20272 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_329
timestamp 1486834041
transform 1 0 28112 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_330
timestamp 1486834041
transform 1 0 8512 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_331
timestamp 1486834041
transform 1 0 16352 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_332
timestamp 1486834041
transform 1 0 24192 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_333
timestamp 1486834041
transform 1 0 4592 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_334
timestamp 1486834041
transform 1 0 12432 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_335
timestamp 1486834041
transform 1 0 20272 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_336
timestamp 1486834041
transform 1 0 28112 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_337
timestamp 1486834041
transform 1 0 8512 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_338
timestamp 1486834041
transform 1 0 16352 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_339
timestamp 1486834041
transform 1 0 24192 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_340
timestamp 1486834041
transform 1 0 4592 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_341
timestamp 1486834041
transform 1 0 12432 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_342
timestamp 1486834041
transform 1 0 20272 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_343
timestamp 1486834041
transform 1 0 28112 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_344
timestamp 1486834041
transform 1 0 8512 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_345
timestamp 1486834041
transform 1 0 16352 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_346
timestamp 1486834041
transform 1 0 24192 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_347
timestamp 1486834041
transform 1 0 4592 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_348
timestamp 1486834041
transform 1 0 12432 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_349
timestamp 1486834041
transform 1 0 20272 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_350
timestamp 1486834041
transform 1 0 28112 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_351
timestamp 1486834041
transform 1 0 8512 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_352
timestamp 1486834041
transform 1 0 16352 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_353
timestamp 1486834041
transform 1 0 24192 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_354
timestamp 1486834041
transform 1 0 4592 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_355
timestamp 1486834041
transform 1 0 12432 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_356
timestamp 1486834041
transform 1 0 20272 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_357
timestamp 1486834041
transform 1 0 28112 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_358
timestamp 1486834041
transform 1 0 8512 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_359
timestamp 1486834041
transform 1 0 16352 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_360
timestamp 1486834041
transform 1 0 24192 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_361
timestamp 1486834041
transform 1 0 4592 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_362
timestamp 1486834041
transform 1 0 12432 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_363
timestamp 1486834041
transform 1 0 20272 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_364
timestamp 1486834041
transform 1 0 28112 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_365
timestamp 1486834041
transform 1 0 8512 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_366
timestamp 1486834041
transform 1 0 16352 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_367
timestamp 1486834041
transform 1 0 24192 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_368
timestamp 1486834041
transform 1 0 4592 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_369
timestamp 1486834041
transform 1 0 12432 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_370
timestamp 1486834041
transform 1 0 20272 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_371
timestamp 1486834041
transform 1 0 28112 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_372
timestamp 1486834041
transform 1 0 8512 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_373
timestamp 1486834041
transform 1 0 16352 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_374
timestamp 1486834041
transform 1 0 24192 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_375
timestamp 1486834041
transform 1 0 4592 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_376
timestamp 1486834041
transform 1 0 12432 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_377
timestamp 1486834041
transform 1 0 20272 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_378
timestamp 1486834041
transform 1 0 28112 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_379
timestamp 1486834041
transform 1 0 8512 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_380
timestamp 1486834041
transform 1 0 16352 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_381
timestamp 1486834041
transform 1 0 24192 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_382
timestamp 1486834041
transform 1 0 4592 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_383
timestamp 1486834041
transform 1 0 12432 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_384
timestamp 1486834041
transform 1 0 20272 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_385
timestamp 1486834041
transform 1 0 28112 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_386
timestamp 1486834041
transform 1 0 8512 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_387
timestamp 1486834041
transform 1 0 16352 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_388
timestamp 1486834041
transform 1 0 24192 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_389
timestamp 1486834041
transform 1 0 4592 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_390
timestamp 1486834041
transform 1 0 12432 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_391
timestamp 1486834041
transform 1 0 20272 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_392
timestamp 1486834041
transform 1 0 28112 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_393
timestamp 1486834041
transform 1 0 8512 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_394
timestamp 1486834041
transform 1 0 16352 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_395
timestamp 1486834041
transform 1 0 24192 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_396
timestamp 1486834041
transform 1 0 4592 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_397
timestamp 1486834041
transform 1 0 12432 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_398
timestamp 1486834041
transform 1 0 20272 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_399
timestamp 1486834041
transform 1 0 28112 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_400
timestamp 1486834041
transform 1 0 8512 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_401
timestamp 1486834041
transform 1 0 16352 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_402
timestamp 1486834041
transform 1 0 24192 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_403
timestamp 1486834041
transform 1 0 4592 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_404
timestamp 1486834041
transform 1 0 12432 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_405
timestamp 1486834041
transform 1 0 20272 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_406
timestamp 1486834041
transform 1 0 28112 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_407
timestamp 1486834041
transform 1 0 8512 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_408
timestamp 1486834041
transform 1 0 16352 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_409
timestamp 1486834041
transform 1 0 24192 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_410
timestamp 1486834041
transform 1 0 4592 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_411
timestamp 1486834041
transform 1 0 12432 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_412
timestamp 1486834041
transform 1 0 20272 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_413
timestamp 1486834041
transform 1 0 28112 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_414
timestamp 1486834041
transform 1 0 8512 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_415
timestamp 1486834041
transform 1 0 16352 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_416
timestamp 1486834041
transform 1 0 24192 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_417
timestamp 1486834041
transform 1 0 4592 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_418
timestamp 1486834041
transform 1 0 12432 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_419
timestamp 1486834041
transform 1 0 20272 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_420
timestamp 1486834041
transform 1 0 28112 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_421
timestamp 1486834041
transform 1 0 8512 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_422
timestamp 1486834041
transform 1 0 16352 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_423
timestamp 1486834041
transform 1 0 24192 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_424
timestamp 1486834041
transform 1 0 4592 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_425
timestamp 1486834041
transform 1 0 12432 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_426
timestamp 1486834041
transform 1 0 20272 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_427
timestamp 1486834041
transform 1 0 28112 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_428
timestamp 1486834041
transform 1 0 8512 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_429
timestamp 1486834041
transform 1 0 16352 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_430
timestamp 1486834041
transform 1 0 24192 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_431
timestamp 1486834041
transform 1 0 4592 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_432
timestamp 1486834041
transform 1 0 12432 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_433
timestamp 1486834041
transform 1 0 20272 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_434
timestamp 1486834041
transform 1 0 28112 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_435
timestamp 1486834041
transform 1 0 8512 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_436
timestamp 1486834041
transform 1 0 16352 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_437
timestamp 1486834041
transform 1 0 24192 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_438
timestamp 1486834041
transform 1 0 4592 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_439
timestamp 1486834041
transform 1 0 12432 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_440
timestamp 1486834041
transform 1 0 20272 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_441
timestamp 1486834041
transform 1 0 28112 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_442
timestamp 1486834041
transform 1 0 8512 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_443
timestamp 1486834041
transform 1 0 16352 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_444
timestamp 1486834041
transform 1 0 24192 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_445
timestamp 1486834041
transform 1 0 4592 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_446
timestamp 1486834041
transform 1 0 12432 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_447
timestamp 1486834041
transform 1 0 20272 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_448
timestamp 1486834041
transform 1 0 28112 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_449
timestamp 1486834041
transform 1 0 8512 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_450
timestamp 1486834041
transform 1 0 16352 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_451
timestamp 1486834041
transform 1 0 24192 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_452
timestamp 1486834041
transform 1 0 4592 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_453
timestamp 1486834041
transform 1 0 12432 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_454
timestamp 1486834041
transform 1 0 20272 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_455
timestamp 1486834041
transform 1 0 28112 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_456
timestamp 1486834041
transform 1 0 8512 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_457
timestamp 1486834041
transform 1 0 16352 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_458
timestamp 1486834041
transform 1 0 24192 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_459
timestamp 1486834041
transform 1 0 4592 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_460
timestamp 1486834041
transform 1 0 12432 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_461
timestamp 1486834041
transform 1 0 20272 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_462
timestamp 1486834041
transform 1 0 28112 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_463
timestamp 1486834041
transform 1 0 8512 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_464
timestamp 1486834041
transform 1 0 16352 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_465
timestamp 1486834041
transform 1 0 24192 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_466
timestamp 1486834041
transform 1 0 4592 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_467
timestamp 1486834041
transform 1 0 12432 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_468
timestamp 1486834041
transform 1 0 20272 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_469
timestamp 1486834041
transform 1 0 28112 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_470
timestamp 1486834041
transform 1 0 8512 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_471
timestamp 1486834041
transform 1 0 16352 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_472
timestamp 1486834041
transform 1 0 24192 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_473
timestamp 1486834041
transform 1 0 4592 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_474
timestamp 1486834041
transform 1 0 12432 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_475
timestamp 1486834041
transform 1 0 20272 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_476
timestamp 1486834041
transform 1 0 28112 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_477
timestamp 1486834041
transform 1 0 8512 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_478
timestamp 1486834041
transform 1 0 16352 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_479
timestamp 1486834041
transform 1 0 24192 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_480
timestamp 1486834041
transform 1 0 4592 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_481
timestamp 1486834041
transform 1 0 12432 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_482
timestamp 1486834041
transform 1 0 20272 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_483
timestamp 1486834041
transform 1 0 28112 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_484
timestamp 1486834041
transform 1 0 8512 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_485
timestamp 1486834041
transform 1 0 16352 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_486
timestamp 1486834041
transform 1 0 24192 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_487
timestamp 1486834041
transform 1 0 4592 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_488
timestamp 1486834041
transform 1 0 12432 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_489
timestamp 1486834041
transform 1 0 20272 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_490
timestamp 1486834041
transform 1 0 28112 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_491
timestamp 1486834041
transform 1 0 8512 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_492
timestamp 1486834041
transform 1 0 16352 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_493
timestamp 1486834041
transform 1 0 24192 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_494
timestamp 1486834041
transform 1 0 4592 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_495
timestamp 1486834041
transform 1 0 12432 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_496
timestamp 1486834041
transform 1 0 20272 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_497
timestamp 1486834041
transform 1 0 28112 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_498
timestamp 1486834041
transform 1 0 8512 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_499
timestamp 1486834041
transform 1 0 16352 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_500
timestamp 1486834041
transform 1 0 24192 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_501
timestamp 1486834041
transform 1 0 4592 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_502
timestamp 1486834041
transform 1 0 12432 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_503
timestamp 1486834041
transform 1 0 20272 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_504
timestamp 1486834041
transform 1 0 28112 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_505
timestamp 1486834041
transform 1 0 8512 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_506
timestamp 1486834041
transform 1 0 16352 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_507
timestamp 1486834041
transform 1 0 24192 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_508
timestamp 1486834041
transform 1 0 4592 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_509
timestamp 1486834041
transform 1 0 12432 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_510
timestamp 1486834041
transform 1 0 20272 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_511
timestamp 1486834041
transform 1 0 28112 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_512
timestamp 1486834041
transform 1 0 8512 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_513
timestamp 1486834041
transform 1 0 16352 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_514
timestamp 1486834041
transform 1 0 24192 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_515
timestamp 1486834041
transform 1 0 4592 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_516
timestamp 1486834041
transform 1 0 12432 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_517
timestamp 1486834041
transform 1 0 20272 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_518
timestamp 1486834041
transform 1 0 28112 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_519
timestamp 1486834041
transform 1 0 8512 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_520
timestamp 1486834041
transform 1 0 16352 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_521
timestamp 1486834041
transform 1 0 24192 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_522
timestamp 1486834041
transform 1 0 4592 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_523
timestamp 1486834041
transform 1 0 12432 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_524
timestamp 1486834041
transform 1 0 20272 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_525
timestamp 1486834041
transform 1 0 28112 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_526
timestamp 1486834041
transform 1 0 8512 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_527
timestamp 1486834041
transform 1 0 16352 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_528
timestamp 1486834041
transform 1 0 24192 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_529
timestamp 1486834041
transform 1 0 4592 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_530
timestamp 1486834041
transform 1 0 12432 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_531
timestamp 1486834041
transform 1 0 20272 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_532
timestamp 1486834041
transform 1 0 28112 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_533
timestamp 1486834041
transform 1 0 8512 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_534
timestamp 1486834041
transform 1 0 16352 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_535
timestamp 1486834041
transform 1 0 24192 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_536
timestamp 1486834041
transform 1 0 4592 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_537
timestamp 1486834041
transform 1 0 12432 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_538
timestamp 1486834041
transform 1 0 20272 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_539
timestamp 1486834041
transform 1 0 28112 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_540
timestamp 1486834041
transform 1 0 8512 0 -1 57232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_541
timestamp 1486834041
transform 1 0 16352 0 -1 57232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_542
timestamp 1486834041
transform 1 0 24192 0 -1 57232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_543
timestamp 1486834041
transform 1 0 4592 0 1 57232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_544
timestamp 1486834041
transform 1 0 12432 0 1 57232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_545
timestamp 1486834041
transform 1 0 20272 0 1 57232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_546
timestamp 1486834041
transform 1 0 28112 0 1 57232
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_547
timestamp 1486834041
transform 1 0 8512 0 -1 58800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_548
timestamp 1486834041
transform 1 0 16352 0 -1 58800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_549
timestamp 1486834041
transform 1 0 24192 0 -1 58800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_550
timestamp 1486834041
transform 1 0 4592 0 1 58800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_551
timestamp 1486834041
transform 1 0 12432 0 1 58800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_552
timestamp 1486834041
transform 1 0 20272 0 1 58800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_553
timestamp 1486834041
transform 1 0 28112 0 1 58800
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_554
timestamp 1486834041
transform 1 0 8512 0 -1 60368
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_555
timestamp 1486834041
transform 1 0 16352 0 -1 60368
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_556
timestamp 1486834041
transform 1 0 24192 0 -1 60368
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_557
timestamp 1486834041
transform 1 0 4592 0 1 60368
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_558
timestamp 1486834041
transform 1 0 12432 0 1 60368
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_559
timestamp 1486834041
transform 1 0 20272 0 1 60368
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_560
timestamp 1486834041
transform 1 0 28112 0 1 60368
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_561
timestamp 1486834041
transform 1 0 8512 0 -1 61936
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_562
timestamp 1486834041
transform 1 0 16352 0 -1 61936
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_563
timestamp 1486834041
transform 1 0 24192 0 -1 61936
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_564
timestamp 1486834041
transform 1 0 4592 0 1 61936
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_565
timestamp 1486834041
transform 1 0 12432 0 1 61936
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_566
timestamp 1486834041
transform 1 0 20272 0 1 61936
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_567
timestamp 1486834041
transform 1 0 28112 0 1 61936
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_568
timestamp 1486834041
transform 1 0 8512 0 -1 63504
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_569
timestamp 1486834041
transform 1 0 16352 0 -1 63504
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_570
timestamp 1486834041
transform 1 0 24192 0 -1 63504
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_571
timestamp 1486834041
transform 1 0 4592 0 1 63504
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_572
timestamp 1486834041
transform 1 0 12432 0 1 63504
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_573
timestamp 1486834041
transform 1 0 20272 0 1 63504
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_574
timestamp 1486834041
transform 1 0 28112 0 1 63504
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_575
timestamp 1486834041
transform 1 0 8512 0 -1 65072
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_576
timestamp 1486834041
transform 1 0 16352 0 -1 65072
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_577
timestamp 1486834041
transform 1 0 24192 0 -1 65072
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_578
timestamp 1486834041
transform 1 0 4592 0 1 65072
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_579
timestamp 1486834041
transform 1 0 12432 0 1 65072
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_580
timestamp 1486834041
transform 1 0 20272 0 1 65072
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_581
timestamp 1486834041
transform 1 0 28112 0 1 65072
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_582
timestamp 1486834041
transform 1 0 8512 0 -1 66640
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_583
timestamp 1486834041
transform 1 0 16352 0 -1 66640
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_584
timestamp 1486834041
transform 1 0 24192 0 -1 66640
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_585
timestamp 1486834041
transform 1 0 4592 0 1 66640
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_586
timestamp 1486834041
transform 1 0 12432 0 1 66640
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_587
timestamp 1486834041
transform 1 0 20272 0 1 66640
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_588
timestamp 1486834041
transform 1 0 28112 0 1 66640
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_589
timestamp 1486834041
transform 1 0 8512 0 -1 68208
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_590
timestamp 1486834041
transform 1 0 16352 0 -1 68208
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_591
timestamp 1486834041
transform 1 0 24192 0 -1 68208
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_592
timestamp 1486834041
transform 1 0 4592 0 1 68208
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_593
timestamp 1486834041
transform 1 0 12432 0 1 68208
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_594
timestamp 1486834041
transform 1 0 20272 0 1 68208
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_595
timestamp 1486834041
transform 1 0 28112 0 1 68208
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_596
timestamp 1486834041
transform 1 0 8512 0 -1 69776
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_597
timestamp 1486834041
transform 1 0 16352 0 -1 69776
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_598
timestamp 1486834041
transform 1 0 24192 0 -1 69776
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_599
timestamp 1486834041
transform 1 0 4592 0 1 69776
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_600
timestamp 1486834041
transform 1 0 12432 0 1 69776
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_601
timestamp 1486834041
transform 1 0 20272 0 1 69776
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_602
timestamp 1486834041
transform 1 0 28112 0 1 69776
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_603
timestamp 1486834041
transform 1 0 8512 0 -1 71344
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_604
timestamp 1486834041
transform 1 0 16352 0 -1 71344
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_605
timestamp 1486834041
transform 1 0 24192 0 -1 71344
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_606
timestamp 1486834041
transform 1 0 4592 0 1 71344
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_607
timestamp 1486834041
transform 1 0 12432 0 1 71344
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_608
timestamp 1486834041
transform 1 0 20272 0 1 71344
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_609
timestamp 1486834041
transform 1 0 28112 0 1 71344
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_610
timestamp 1486834041
transform 1 0 8512 0 -1 72912
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_611
timestamp 1486834041
transform 1 0 16352 0 -1 72912
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_612
timestamp 1486834041
transform 1 0 24192 0 -1 72912
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_613
timestamp 1486834041
transform 1 0 4592 0 1 72912
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_614
timestamp 1486834041
transform 1 0 12432 0 1 72912
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_615
timestamp 1486834041
transform 1 0 20272 0 1 72912
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_616
timestamp 1486834041
transform 1 0 28112 0 1 72912
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_617
timestamp 1486834041
transform 1 0 8512 0 -1 74480
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_618
timestamp 1486834041
transform 1 0 16352 0 -1 74480
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_619
timestamp 1486834041
transform 1 0 24192 0 -1 74480
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_94_620
timestamp 1486834041
transform 1 0 4592 0 1 74480
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_94_621
timestamp 1486834041
transform 1 0 12432 0 1 74480
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_94_622
timestamp 1486834041
transform 1 0 20272 0 1 74480
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_94_623
timestamp 1486834041
transform 1 0 28112 0 1 74480
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_95_624
timestamp 1486834041
transform 1 0 8512 0 -1 76048
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_95_625
timestamp 1486834041
transform 1 0 16352 0 -1 76048
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_95_626
timestamp 1486834041
transform 1 0 24192 0 -1 76048
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_96_627
timestamp 1486834041
transform 1 0 4592 0 1 76048
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_96_628
timestamp 1486834041
transform 1 0 12432 0 1 76048
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_96_629
timestamp 1486834041
transform 1 0 20272 0 1 76048
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_96_630
timestamp 1486834041
transform 1 0 28112 0 1 76048
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_97_631
timestamp 1486834041
transform 1 0 8512 0 -1 77616
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_97_632
timestamp 1486834041
transform 1 0 16352 0 -1 77616
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_97_633
timestamp 1486834041
transform 1 0 24192 0 -1 77616
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_98_634
timestamp 1486834041
transform 1 0 4592 0 1 77616
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_98_635
timestamp 1486834041
transform 1 0 12432 0 1 77616
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_98_636
timestamp 1486834041
transform 1 0 20272 0 1 77616
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_98_637
timestamp 1486834041
transform 1 0 28112 0 1 77616
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_99_638
timestamp 1486834041
transform 1 0 8512 0 -1 79184
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_99_639
timestamp 1486834041
transform 1 0 16352 0 -1 79184
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_99_640
timestamp 1486834041
transform 1 0 24192 0 -1 79184
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_100_641
timestamp 1486834041
transform 1 0 4592 0 1 79184
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_100_642
timestamp 1486834041
transform 1 0 12432 0 1 79184
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_100_643
timestamp 1486834041
transform 1 0 20272 0 1 79184
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_100_644
timestamp 1486834041
transform 1 0 28112 0 1 79184
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_101_645
timestamp 1486834041
transform 1 0 8512 0 -1 80752
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_101_646
timestamp 1486834041
transform 1 0 16352 0 -1 80752
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_101_647
timestamp 1486834041
transform 1 0 24192 0 -1 80752
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_102_648
timestamp 1486834041
transform 1 0 4592 0 1 80752
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_102_649
timestamp 1486834041
transform 1 0 12432 0 1 80752
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_102_650
timestamp 1486834041
transform 1 0 20272 0 1 80752
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_102_651
timestamp 1486834041
transform 1 0 28112 0 1 80752
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_103_652
timestamp 1486834041
transform 1 0 8512 0 -1 82320
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_103_653
timestamp 1486834041
transform 1 0 16352 0 -1 82320
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_103_654
timestamp 1486834041
transform 1 0 24192 0 -1 82320
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_104_655
timestamp 1486834041
transform 1 0 4592 0 1 82320
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_104_656
timestamp 1486834041
transform 1 0 12432 0 1 82320
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_104_657
timestamp 1486834041
transform 1 0 20272 0 1 82320
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_104_658
timestamp 1486834041
transform 1 0 28112 0 1 82320
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_105_659
timestamp 1486834041
transform 1 0 8512 0 -1 83888
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_105_660
timestamp 1486834041
transform 1 0 16352 0 -1 83888
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_105_661
timestamp 1486834041
transform 1 0 24192 0 -1 83888
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_106_662
timestamp 1486834041
transform 1 0 4592 0 1 83888
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_106_663
timestamp 1486834041
transform 1 0 12432 0 1 83888
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_106_664
timestamp 1486834041
transform 1 0 20272 0 1 83888
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_106_665
timestamp 1486834041
transform 1 0 28112 0 1 83888
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_107_666
timestamp 1486834041
transform 1 0 8512 0 -1 85456
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_107_667
timestamp 1486834041
transform 1 0 16352 0 -1 85456
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_107_668
timestamp 1486834041
transform 1 0 24192 0 -1 85456
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_108_669
timestamp 1486834041
transform 1 0 4592 0 1 85456
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_108_670
timestamp 1486834041
transform 1 0 12432 0 1 85456
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_108_671
timestamp 1486834041
transform 1 0 20272 0 1 85456
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_108_672
timestamp 1486834041
transform 1 0 28112 0 1 85456
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_109_673
timestamp 1486834041
transform 1 0 8512 0 -1 87024
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_109_674
timestamp 1486834041
transform 1 0 16352 0 -1 87024
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_109_675
timestamp 1486834041
transform 1 0 24192 0 -1 87024
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_110_676
timestamp 1486834041
transform 1 0 4592 0 1 87024
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_110_677
timestamp 1486834041
transform 1 0 12432 0 1 87024
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_110_678
timestamp 1486834041
transform 1 0 20272 0 1 87024
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_110_679
timestamp 1486834041
transform 1 0 28112 0 1 87024
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_111_680
timestamp 1486834041
transform 1 0 8512 0 -1 88592
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_111_681
timestamp 1486834041
transform 1 0 16352 0 -1 88592
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_111_682
timestamp 1486834041
transform 1 0 24192 0 -1 88592
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_112_683
timestamp 1486834041
transform 1 0 4592 0 1 88592
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_112_684
timestamp 1486834041
transform 1 0 12432 0 1 88592
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_112_685
timestamp 1486834041
transform 1 0 20272 0 1 88592
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_112_686
timestamp 1486834041
transform 1 0 28112 0 1 88592
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_113_687
timestamp 1486834041
transform 1 0 8512 0 -1 90160
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_113_688
timestamp 1486834041
transform 1 0 16352 0 -1 90160
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_113_689
timestamp 1486834041
transform 1 0 24192 0 -1 90160
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_114_690
timestamp 1486834041
transform 1 0 4592 0 1 90160
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_114_691
timestamp 1486834041
transform 1 0 12432 0 1 90160
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_114_692
timestamp 1486834041
transform 1 0 20272 0 1 90160
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_114_693
timestamp 1486834041
transform 1 0 28112 0 1 90160
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_115_694
timestamp 1486834041
transform 1 0 8512 0 -1 91728
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_115_695
timestamp 1486834041
transform 1 0 16352 0 -1 91728
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_115_696
timestamp 1486834041
transform 1 0 24192 0 -1 91728
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_116_697
timestamp 1486834041
transform 1 0 4592 0 1 91728
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_116_698
timestamp 1486834041
transform 1 0 12432 0 1 91728
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_116_699
timestamp 1486834041
transform 1 0 20272 0 1 91728
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_116_700
timestamp 1486834041
transform 1 0 28112 0 1 91728
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_117_701
timestamp 1486834041
transform 1 0 8512 0 -1 93296
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_117_702
timestamp 1486834041
transform 1 0 16352 0 -1 93296
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_117_703
timestamp 1486834041
transform 1 0 24192 0 -1 93296
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_118_704
timestamp 1486834041
transform 1 0 4592 0 1 93296
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_118_705
timestamp 1486834041
transform 1 0 12432 0 1 93296
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_118_706
timestamp 1486834041
transform 1 0 20272 0 1 93296
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_118_707
timestamp 1486834041
transform 1 0 28112 0 1 93296
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_119_708
timestamp 1486834041
transform 1 0 8512 0 -1 94864
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_119_709
timestamp 1486834041
transform 1 0 16352 0 -1 94864
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_119_710
timestamp 1486834041
transform 1 0 24192 0 -1 94864
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_120_711
timestamp 1486834041
transform 1 0 4592 0 1 94864
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_120_712
timestamp 1486834041
transform 1 0 12432 0 1 94864
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_120_713
timestamp 1486834041
transform 1 0 20272 0 1 94864
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_120_714
timestamp 1486834041
transform 1 0 28112 0 1 94864
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_121_715
timestamp 1486834041
transform 1 0 8512 0 -1 96432
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_121_716
timestamp 1486834041
transform 1 0 16352 0 -1 96432
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_121_717
timestamp 1486834041
transform 1 0 24192 0 -1 96432
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_122_718
timestamp 1486834041
transform 1 0 4592 0 1 96432
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_122_719
timestamp 1486834041
transform 1 0 12432 0 1 96432
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_122_720
timestamp 1486834041
transform 1 0 20272 0 1 96432
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_122_721
timestamp 1486834041
transform 1 0 28112 0 1 96432
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_123_722
timestamp 1486834041
transform 1 0 8512 0 -1 98000
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_123_723
timestamp 1486834041
transform 1 0 16352 0 -1 98000
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_123_724
timestamp 1486834041
transform 1 0 24192 0 -1 98000
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_124_725
timestamp 1486834041
transform 1 0 4592 0 1 98000
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_124_726
timestamp 1486834041
transform 1 0 12432 0 1 98000
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_124_727
timestamp 1486834041
transform 1 0 20272 0 1 98000
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_124_728
timestamp 1486834041
transform 1 0 28112 0 1 98000
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_125_729
timestamp 1486834041
transform 1 0 8512 0 -1 99568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_125_730
timestamp 1486834041
transform 1 0 16352 0 -1 99568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_125_731
timestamp 1486834041
transform 1 0 24192 0 -1 99568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_126_732
timestamp 1486834041
transform 1 0 4592 0 1 99568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_126_733
timestamp 1486834041
transform 1 0 12432 0 1 99568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_126_734
timestamp 1486834041
transform 1 0 20272 0 1 99568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_126_735
timestamp 1486834041
transform 1 0 28112 0 1 99568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_127_736
timestamp 1486834041
transform 1 0 8512 0 -1 101136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_127_737
timestamp 1486834041
transform 1 0 16352 0 -1 101136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_127_738
timestamp 1486834041
transform 1 0 24192 0 -1 101136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_128_739
timestamp 1486834041
transform 1 0 4592 0 1 101136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_128_740
timestamp 1486834041
transform 1 0 12432 0 1 101136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_128_741
timestamp 1486834041
transform 1 0 20272 0 1 101136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_128_742
timestamp 1486834041
transform 1 0 28112 0 1 101136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_129_743
timestamp 1486834041
transform 1 0 8512 0 -1 102704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_129_744
timestamp 1486834041
transform 1 0 16352 0 -1 102704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_129_745
timestamp 1486834041
transform 1 0 24192 0 -1 102704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_130_746
timestamp 1486834041
transform 1 0 4592 0 1 102704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_130_747
timestamp 1486834041
transform 1 0 12432 0 1 102704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_130_748
timestamp 1486834041
transform 1 0 20272 0 1 102704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_130_749
timestamp 1486834041
transform 1 0 28112 0 1 102704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_131_750
timestamp 1486834041
transform 1 0 8512 0 -1 104272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_131_751
timestamp 1486834041
transform 1 0 16352 0 -1 104272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_131_752
timestamp 1486834041
transform 1 0 24192 0 -1 104272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_132_753
timestamp 1486834041
transform 1 0 4592 0 1 104272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_132_754
timestamp 1486834041
transform 1 0 12432 0 1 104272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_132_755
timestamp 1486834041
transform 1 0 20272 0 1 104272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_132_756
timestamp 1486834041
transform 1 0 28112 0 1 104272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_133_757
timestamp 1486834041
transform 1 0 8512 0 -1 105840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_133_758
timestamp 1486834041
transform 1 0 16352 0 -1 105840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_133_759
timestamp 1486834041
transform 1 0 24192 0 -1 105840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_134_760
timestamp 1486834041
transform 1 0 4592 0 1 105840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_134_761
timestamp 1486834041
transform 1 0 12432 0 1 105840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_134_762
timestamp 1486834041
transform 1 0 20272 0 1 105840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_134_763
timestamp 1486834041
transform 1 0 28112 0 1 105840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_135_764
timestamp 1486834041
transform 1 0 8512 0 -1 107408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_135_765
timestamp 1486834041
transform 1 0 16352 0 -1 107408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_135_766
timestamp 1486834041
transform 1 0 24192 0 -1 107408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_136_767
timestamp 1486834041
transform 1 0 4592 0 1 107408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_136_768
timestamp 1486834041
transform 1 0 12432 0 1 107408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_136_769
timestamp 1486834041
transform 1 0 20272 0 1 107408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_136_770
timestamp 1486834041
transform 1 0 28112 0 1 107408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_137_771
timestamp 1486834041
transform 1 0 8512 0 -1 108976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_137_772
timestamp 1486834041
transform 1 0 16352 0 -1 108976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_137_773
timestamp 1486834041
transform 1 0 24192 0 -1 108976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_138_774
timestamp 1486834041
transform 1 0 4592 0 1 108976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_138_775
timestamp 1486834041
transform 1 0 12432 0 1 108976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_138_776
timestamp 1486834041
transform 1 0 20272 0 1 108976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_138_777
timestamp 1486834041
transform 1 0 28112 0 1 108976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_139_778
timestamp 1486834041
transform 1 0 8512 0 -1 110544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_139_779
timestamp 1486834041
transform 1 0 16352 0 -1 110544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_139_780
timestamp 1486834041
transform 1 0 24192 0 -1 110544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_140_781
timestamp 1486834041
transform 1 0 4592 0 1 110544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_140_782
timestamp 1486834041
transform 1 0 12432 0 1 110544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_140_783
timestamp 1486834041
transform 1 0 20272 0 1 110544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_140_784
timestamp 1486834041
transform 1 0 28112 0 1 110544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_141_785
timestamp 1486834041
transform 1 0 8512 0 -1 112112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_141_786
timestamp 1486834041
transform 1 0 16352 0 -1 112112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_141_787
timestamp 1486834041
transform 1 0 24192 0 -1 112112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_142_788
timestamp 1486834041
transform 1 0 4592 0 1 112112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_142_789
timestamp 1486834041
transform 1 0 12432 0 1 112112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_142_790
timestamp 1486834041
transform 1 0 20272 0 1 112112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_142_791
timestamp 1486834041
transform 1 0 28112 0 1 112112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_143_792
timestamp 1486834041
transform 1 0 4480 0 -1 113680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_143_793
timestamp 1486834041
transform 1 0 8288 0 -1 113680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_143_794
timestamp 1486834041
transform 1 0 12096 0 -1 113680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_143_795
timestamp 1486834041
transform 1 0 15904 0 -1 113680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_143_796
timestamp 1486834041
transform 1 0 19712 0 -1 113680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_143_797
timestamp 1486834041
transform 1 0 23520 0 -1 113680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_143_798
timestamp 1486834041
transform 1 0 27328 0 -1 113680
box -86 -86 310 870
<< labels >>
flabel metal3 s 31584 19936 31696 20048 0 FreeSans 448 0 0 0 A_SRAM0
port 0 nsew signal output
flabel metal3 s 31584 20832 31696 20944 0 FreeSans 448 0 0 0 A_SRAM1
port 1 nsew signal output
flabel metal3 s 31584 21728 31696 21840 0 FreeSans 448 0 0 0 A_SRAM2
port 2 nsew signal output
flabel metal3 s 31584 22624 31696 22736 0 FreeSans 448 0 0 0 A_SRAM3
port 3 nsew signal output
flabel metal3 s 31584 23520 31696 23632 0 FreeSans 448 0 0 0 A_SRAM4
port 4 nsew signal output
flabel metal3 s 31584 24416 31696 24528 0 FreeSans 448 0 0 0 A_SRAM5
port 5 nsew signal output
flabel metal3 s 31584 25312 31696 25424 0 FreeSans 448 0 0 0 A_SRAM6
port 6 nsew signal output
flabel metal3 s 31584 26208 31696 26320 0 FreeSans 448 0 0 0 A_SRAM7
port 7 nsew signal output
flabel metal3 s 31584 27104 31696 27216 0 FreeSans 448 0 0 0 A_SRAM8
port 8 nsew signal output
flabel metal3 s 31584 10976 31696 11088 0 FreeSans 448 0 0 0 CEN_SRAM
port 9 nsew signal output
flabel metal3 s 31584 35168 31696 35280 0 FreeSans 448 0 0 0 CLK_SRAM
port 10 nsew signal output
flabel metal3 s 31584 10080 31696 10192 0 FreeSans 448 0 0 0 CONFIGURED_top
port 11 nsew signal input
flabel metal3 s 31584 28000 31696 28112 0 FreeSans 448 0 0 0 D_SRAM0
port 12 nsew signal output
flabel metal3 s 31584 28896 31696 29008 0 FreeSans 448 0 0 0 D_SRAM1
port 13 nsew signal output
flabel metal3 s 31584 29792 31696 29904 0 FreeSans 448 0 0 0 D_SRAM2
port 14 nsew signal output
flabel metal3 s 31584 30688 31696 30800 0 FreeSans 448 0 0 0 D_SRAM3
port 15 nsew signal output
flabel metal3 s 31584 31584 31696 31696 0 FreeSans 448 0 0 0 D_SRAM4
port 16 nsew signal output
flabel metal3 s 31584 32480 31696 32592 0 FreeSans 448 0 0 0 D_SRAM5
port 17 nsew signal output
flabel metal3 s 31584 33376 31696 33488 0 FreeSans 448 0 0 0 D_SRAM6
port 18 nsew signal output
flabel metal3 s 31584 34272 31696 34384 0 FreeSans 448 0 0 0 D_SRAM7
port 19 nsew signal output
flabel metal3 s 31584 11872 31696 11984 0 FreeSans 448 0 0 0 GWEN_SRAM
port 20 nsew signal output
flabel metal3 s 31584 2912 31696 3024 0 FreeSans 448 0 0 0 Q_SRAM0
port 21 nsew signal input
flabel metal3 s 31584 3808 31696 3920 0 FreeSans 448 0 0 0 Q_SRAM1
port 22 nsew signal input
flabel metal3 s 31584 4704 31696 4816 0 FreeSans 448 0 0 0 Q_SRAM2
port 23 nsew signal input
flabel metal3 s 31584 5600 31696 5712 0 FreeSans 448 0 0 0 Q_SRAM3
port 24 nsew signal input
flabel metal3 s 31584 6496 31696 6608 0 FreeSans 448 0 0 0 Q_SRAM4
port 25 nsew signal input
flabel metal3 s 31584 7392 31696 7504 0 FreeSans 448 0 0 0 Q_SRAM5
port 26 nsew signal input
flabel metal3 s 31584 8288 31696 8400 0 FreeSans 448 0 0 0 Q_SRAM6
port 27 nsew signal input
flabel metal3 s 31584 9184 31696 9296 0 FreeSans 448 0 0 0 Q_SRAM7
port 28 nsew signal input
flabel metal3 s 0 79184 112 79296 0 FreeSans 448 0 0 0 Tile_X0Y0_E1END[0]
port 29 nsew signal input
flabel metal3 s 0 79632 112 79744 0 FreeSans 448 0 0 0 Tile_X0Y0_E1END[1]
port 30 nsew signal input
flabel metal3 s 0 80080 112 80192 0 FreeSans 448 0 0 0 Tile_X0Y0_E1END[2]
port 31 nsew signal input
flabel metal3 s 0 80528 112 80640 0 FreeSans 448 0 0 0 Tile_X0Y0_E1END[3]
port 32 nsew signal input
flabel metal3 s 0 84560 112 84672 0 FreeSans 448 0 0 0 Tile_X0Y0_E2END[0]
port 33 nsew signal input
flabel metal3 s 0 85008 112 85120 0 FreeSans 448 0 0 0 Tile_X0Y0_E2END[1]
port 34 nsew signal input
flabel metal3 s 0 85456 112 85568 0 FreeSans 448 0 0 0 Tile_X0Y0_E2END[2]
port 35 nsew signal input
flabel metal3 s 0 85904 112 86016 0 FreeSans 448 0 0 0 Tile_X0Y0_E2END[3]
port 36 nsew signal input
flabel metal3 s 0 86352 112 86464 0 FreeSans 448 0 0 0 Tile_X0Y0_E2END[4]
port 37 nsew signal input
flabel metal3 s 0 86800 112 86912 0 FreeSans 448 0 0 0 Tile_X0Y0_E2END[5]
port 38 nsew signal input
flabel metal3 s 0 87248 112 87360 0 FreeSans 448 0 0 0 Tile_X0Y0_E2END[6]
port 39 nsew signal input
flabel metal3 s 0 87696 112 87808 0 FreeSans 448 0 0 0 Tile_X0Y0_E2END[7]
port 40 nsew signal input
flabel metal3 s 0 80976 112 81088 0 FreeSans 448 0 0 0 Tile_X0Y0_E2MID[0]
port 41 nsew signal input
flabel metal3 s 0 81424 112 81536 0 FreeSans 448 0 0 0 Tile_X0Y0_E2MID[1]
port 42 nsew signal input
flabel metal3 s 0 81872 112 81984 0 FreeSans 448 0 0 0 Tile_X0Y0_E2MID[2]
port 43 nsew signal input
flabel metal3 s 0 82320 112 82432 0 FreeSans 448 0 0 0 Tile_X0Y0_E2MID[3]
port 44 nsew signal input
flabel metal3 s 0 82768 112 82880 0 FreeSans 448 0 0 0 Tile_X0Y0_E2MID[4]
port 45 nsew signal input
flabel metal3 s 0 83216 112 83328 0 FreeSans 448 0 0 0 Tile_X0Y0_E2MID[5]
port 46 nsew signal input
flabel metal3 s 0 83664 112 83776 0 FreeSans 448 0 0 0 Tile_X0Y0_E2MID[6]
port 47 nsew signal input
flabel metal3 s 0 84112 112 84224 0 FreeSans 448 0 0 0 Tile_X0Y0_E2MID[7]
port 48 nsew signal input
flabel metal3 s 0 95312 112 95424 0 FreeSans 448 0 0 0 Tile_X0Y0_E6END[0]
port 49 nsew signal input
flabel metal3 s 0 99792 112 99904 0 FreeSans 448 0 0 0 Tile_X0Y0_E6END[10]
port 50 nsew signal input
flabel metal3 s 0 100240 112 100352 0 FreeSans 448 0 0 0 Tile_X0Y0_E6END[11]
port 51 nsew signal input
flabel metal3 s 0 95760 112 95872 0 FreeSans 448 0 0 0 Tile_X0Y0_E6END[1]
port 52 nsew signal input
flabel metal3 s 0 96208 112 96320 0 FreeSans 448 0 0 0 Tile_X0Y0_E6END[2]
port 53 nsew signal input
flabel metal3 s 0 96656 112 96768 0 FreeSans 448 0 0 0 Tile_X0Y0_E6END[3]
port 54 nsew signal input
flabel metal3 s 0 97104 112 97216 0 FreeSans 448 0 0 0 Tile_X0Y0_E6END[4]
port 55 nsew signal input
flabel metal3 s 0 97552 112 97664 0 FreeSans 448 0 0 0 Tile_X0Y0_E6END[5]
port 56 nsew signal input
flabel metal3 s 0 98000 112 98112 0 FreeSans 448 0 0 0 Tile_X0Y0_E6END[6]
port 57 nsew signal input
flabel metal3 s 0 98448 112 98560 0 FreeSans 448 0 0 0 Tile_X0Y0_E6END[7]
port 58 nsew signal input
flabel metal3 s 0 98896 112 99008 0 FreeSans 448 0 0 0 Tile_X0Y0_E6END[8]
port 59 nsew signal input
flabel metal3 s 0 99344 112 99456 0 FreeSans 448 0 0 0 Tile_X0Y0_E6END[9]
port 60 nsew signal input
flabel metal3 s 0 88144 112 88256 0 FreeSans 448 0 0 0 Tile_X0Y0_EE4END[0]
port 61 nsew signal input
flabel metal3 s 0 92624 112 92736 0 FreeSans 448 0 0 0 Tile_X0Y0_EE4END[10]
port 62 nsew signal input
flabel metal3 s 0 93072 112 93184 0 FreeSans 448 0 0 0 Tile_X0Y0_EE4END[11]
port 63 nsew signal input
flabel metal3 s 0 93520 112 93632 0 FreeSans 448 0 0 0 Tile_X0Y0_EE4END[12]
port 64 nsew signal input
flabel metal3 s 0 93968 112 94080 0 FreeSans 448 0 0 0 Tile_X0Y0_EE4END[13]
port 65 nsew signal input
flabel metal3 s 0 94416 112 94528 0 FreeSans 448 0 0 0 Tile_X0Y0_EE4END[14]
port 66 nsew signal input
flabel metal3 s 0 94864 112 94976 0 FreeSans 448 0 0 0 Tile_X0Y0_EE4END[15]
port 67 nsew signal input
flabel metal3 s 0 88592 112 88704 0 FreeSans 448 0 0 0 Tile_X0Y0_EE4END[1]
port 68 nsew signal input
flabel metal3 s 0 89040 112 89152 0 FreeSans 448 0 0 0 Tile_X0Y0_EE4END[2]
port 69 nsew signal input
flabel metal3 s 0 89488 112 89600 0 FreeSans 448 0 0 0 Tile_X0Y0_EE4END[3]
port 70 nsew signal input
flabel metal3 s 0 89936 112 90048 0 FreeSans 448 0 0 0 Tile_X0Y0_EE4END[4]
port 71 nsew signal input
flabel metal3 s 0 90384 112 90496 0 FreeSans 448 0 0 0 Tile_X0Y0_EE4END[5]
port 72 nsew signal input
flabel metal3 s 0 90832 112 90944 0 FreeSans 448 0 0 0 Tile_X0Y0_EE4END[6]
port 73 nsew signal input
flabel metal3 s 0 91280 112 91392 0 FreeSans 448 0 0 0 Tile_X0Y0_EE4END[7]
port 74 nsew signal input
flabel metal3 s 0 91728 112 91840 0 FreeSans 448 0 0 0 Tile_X0Y0_EE4END[8]
port 75 nsew signal input
flabel metal3 s 0 92176 112 92288 0 FreeSans 448 0 0 0 Tile_X0Y0_EE4END[9]
port 76 nsew signal input
flabel metal3 s 0 100688 112 100800 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData[0]
port 77 nsew signal input
flabel metal3 s 0 105168 112 105280 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData[10]
port 78 nsew signal input
flabel metal3 s 0 105616 112 105728 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData[11]
port 79 nsew signal input
flabel metal3 s 0 106064 112 106176 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData[12]
port 80 nsew signal input
flabel metal3 s 0 106512 112 106624 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData[13]
port 81 nsew signal input
flabel metal3 s 0 106960 112 107072 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData[14]
port 82 nsew signal input
flabel metal3 s 0 107408 112 107520 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData[15]
port 83 nsew signal input
flabel metal3 s 0 107856 112 107968 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData[16]
port 84 nsew signal input
flabel metal3 s 0 108304 112 108416 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData[17]
port 85 nsew signal input
flabel metal3 s 0 108752 112 108864 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData[18]
port 86 nsew signal input
flabel metal3 s 0 109200 112 109312 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData[19]
port 87 nsew signal input
flabel metal3 s 0 101136 112 101248 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData[1]
port 88 nsew signal input
flabel metal3 s 0 109648 112 109760 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData[20]
port 89 nsew signal input
flabel metal3 s 0 110096 112 110208 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData[21]
port 90 nsew signal input
flabel metal3 s 0 110544 112 110656 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData[22]
port 91 nsew signal input
flabel metal3 s 0 110992 112 111104 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData[23]
port 92 nsew signal input
flabel metal3 s 0 111440 112 111552 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData[24]
port 93 nsew signal input
flabel metal3 s 0 111888 112 112000 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData[25]
port 94 nsew signal input
flabel metal3 s 0 112336 112 112448 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData[26]
port 95 nsew signal input
flabel metal3 s 0 112784 112 112896 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData[27]
port 96 nsew signal input
flabel metal3 s 0 113232 112 113344 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData[28]
port 97 nsew signal input
flabel metal3 s 0 113680 112 113792 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData[29]
port 98 nsew signal input
flabel metal3 s 0 101584 112 101696 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData[2]
port 99 nsew signal input
flabel metal3 s 0 114128 112 114240 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData[30]
port 100 nsew signal input
flabel metal3 s 0 114576 112 114688 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData[31]
port 101 nsew signal input
flabel metal3 s 0 102032 112 102144 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData[3]
port 102 nsew signal input
flabel metal3 s 0 102480 112 102592 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData[4]
port 103 nsew signal input
flabel metal3 s 0 102928 112 103040 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData[5]
port 104 nsew signal input
flabel metal3 s 0 103376 112 103488 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData[6]
port 105 nsew signal input
flabel metal3 s 0 103824 112 103936 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData[7]
port 106 nsew signal input
flabel metal3 s 0 104272 112 104384 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData[8]
port 107 nsew signal input
flabel metal3 s 0 104720 112 104832 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData[9]
port 108 nsew signal input
flabel metal3 s 31584 78176 31696 78288 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData_O[0]
port 109 nsew signal output
flabel metal3 s 31584 89376 31696 89488 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData_O[10]
port 110 nsew signal output
flabel metal3 s 31584 90496 31696 90608 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData_O[11]
port 111 nsew signal output
flabel metal3 s 31584 91616 31696 91728 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData_O[12]
port 112 nsew signal output
flabel metal3 s 31584 92736 31696 92848 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData_O[13]
port 113 nsew signal output
flabel metal3 s 31584 93856 31696 93968 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData_O[14]
port 114 nsew signal output
flabel metal3 s 31584 94976 31696 95088 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData_O[15]
port 115 nsew signal output
flabel metal3 s 31584 96096 31696 96208 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData_O[16]
port 116 nsew signal output
flabel metal3 s 31584 97216 31696 97328 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData_O[17]
port 117 nsew signal output
flabel metal3 s 31584 98336 31696 98448 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData_O[18]
port 118 nsew signal output
flabel metal3 s 31584 99456 31696 99568 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData_O[19]
port 119 nsew signal output
flabel metal3 s 31584 79296 31696 79408 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData_O[1]
port 120 nsew signal output
flabel metal3 s 31584 100576 31696 100688 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData_O[20]
port 121 nsew signal output
flabel metal3 s 31584 101696 31696 101808 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData_O[21]
port 122 nsew signal output
flabel metal3 s 31584 102816 31696 102928 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData_O[22]
port 123 nsew signal output
flabel metal3 s 31584 103936 31696 104048 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData_O[23]
port 124 nsew signal output
flabel metal3 s 31584 105056 31696 105168 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData_O[24]
port 125 nsew signal output
flabel metal3 s 31584 106176 31696 106288 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData_O[25]
port 126 nsew signal output
flabel metal3 s 31584 107296 31696 107408 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData_O[26]
port 127 nsew signal output
flabel metal3 s 31584 108416 31696 108528 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData_O[27]
port 128 nsew signal output
flabel metal3 s 31584 109536 31696 109648 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData_O[28]
port 129 nsew signal output
flabel metal3 s 31584 110656 31696 110768 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData_O[29]
port 130 nsew signal output
flabel metal3 s 31584 80416 31696 80528 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData_O[2]
port 131 nsew signal output
flabel metal3 s 31584 111776 31696 111888 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData_O[30]
port 132 nsew signal output
flabel metal3 s 31584 112896 31696 113008 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData_O[31]
port 133 nsew signal output
flabel metal3 s 31584 81536 31696 81648 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData_O[3]
port 134 nsew signal output
flabel metal3 s 31584 82656 31696 82768 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData_O[4]
port 135 nsew signal output
flabel metal3 s 31584 83776 31696 83888 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData_O[5]
port 136 nsew signal output
flabel metal3 s 31584 84896 31696 85008 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData_O[6]
port 137 nsew signal output
flabel metal3 s 31584 86016 31696 86128 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData_O[7]
port 138 nsew signal output
flabel metal3 s 31584 87136 31696 87248 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData_O[8]
port 139 nsew signal output
flabel metal3 s 31584 88256 31696 88368 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameData_O[9]
port 140 nsew signal output
flabel metal2 s 21728 114800 21840 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameStrobe_O[0]
port 141 nsew signal output
flabel metal2 s 23968 114800 24080 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameStrobe_O[10]
port 142 nsew signal output
flabel metal2 s 24192 114800 24304 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameStrobe_O[11]
port 143 nsew signal output
flabel metal2 s 24416 114800 24528 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameStrobe_O[12]
port 144 nsew signal output
flabel metal2 s 24640 114800 24752 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameStrobe_O[13]
port 145 nsew signal output
flabel metal2 s 24864 114800 24976 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameStrobe_O[14]
port 146 nsew signal output
flabel metal2 s 25088 114800 25200 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameStrobe_O[15]
port 147 nsew signal output
flabel metal2 s 25312 114800 25424 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameStrobe_O[16]
port 148 nsew signal output
flabel metal2 s 25536 114800 25648 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameStrobe_O[17]
port 149 nsew signal output
flabel metal2 s 25760 114800 25872 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameStrobe_O[18]
port 150 nsew signal output
flabel metal2 s 25984 114800 26096 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameStrobe_O[19]
port 151 nsew signal output
flabel metal2 s 21952 114800 22064 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameStrobe_O[1]
port 152 nsew signal output
flabel metal2 s 22176 114800 22288 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameStrobe_O[2]
port 153 nsew signal output
flabel metal2 s 22400 114800 22512 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameStrobe_O[3]
port 154 nsew signal output
flabel metal2 s 22624 114800 22736 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameStrobe_O[4]
port 155 nsew signal output
flabel metal2 s 22848 114800 22960 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameStrobe_O[5]
port 156 nsew signal output
flabel metal2 s 23072 114800 23184 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameStrobe_O[6]
port 157 nsew signal output
flabel metal2 s 23296 114800 23408 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameStrobe_O[7]
port 158 nsew signal output
flabel metal2 s 23520 114800 23632 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameStrobe_O[8]
port 159 nsew signal output
flabel metal2 s 23744 114800 23856 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_FrameStrobe_O[9]
port 160 nsew signal output
flabel metal2 s 5376 114800 5488 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_N1BEG[0]
port 161 nsew signal output
flabel metal2 s 5600 114800 5712 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_N1BEG[1]
port 162 nsew signal output
flabel metal2 s 5824 114800 5936 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_N1BEG[2]
port 163 nsew signal output
flabel metal2 s 6048 114800 6160 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_N1BEG[3]
port 164 nsew signal output
flabel metal2 s 6272 114800 6384 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_N2BEG[0]
port 165 nsew signal output
flabel metal2 s 6496 114800 6608 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_N2BEG[1]
port 166 nsew signal output
flabel metal2 s 6720 114800 6832 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_N2BEG[2]
port 167 nsew signal output
flabel metal2 s 6944 114800 7056 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_N2BEG[3]
port 168 nsew signal output
flabel metal2 s 7168 114800 7280 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_N2BEG[4]
port 169 nsew signal output
flabel metal2 s 7392 114800 7504 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_N2BEG[5]
port 170 nsew signal output
flabel metal2 s 7616 114800 7728 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_N2BEG[6]
port 171 nsew signal output
flabel metal2 s 7840 114800 7952 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_N2BEG[7]
port 172 nsew signal output
flabel metal2 s 8064 114800 8176 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_N2BEGb[0]
port 173 nsew signal output
flabel metal2 s 8288 114800 8400 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_N2BEGb[1]
port 174 nsew signal output
flabel metal2 s 8512 114800 8624 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_N2BEGb[2]
port 175 nsew signal output
flabel metal2 s 8736 114800 8848 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_N2BEGb[3]
port 176 nsew signal output
flabel metal2 s 8960 114800 9072 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_N2BEGb[4]
port 177 nsew signal output
flabel metal2 s 9184 114800 9296 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_N2BEGb[5]
port 178 nsew signal output
flabel metal2 s 9408 114800 9520 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_N2BEGb[6]
port 179 nsew signal output
flabel metal2 s 9632 114800 9744 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_N2BEGb[7]
port 180 nsew signal output
flabel metal2 s 9856 114800 9968 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_N4BEG[0]
port 181 nsew signal output
flabel metal2 s 12096 114800 12208 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_N4BEG[10]
port 182 nsew signal output
flabel metal2 s 12320 114800 12432 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_N4BEG[11]
port 183 nsew signal output
flabel metal2 s 12544 114800 12656 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_N4BEG[12]
port 184 nsew signal output
flabel metal2 s 12768 114800 12880 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_N4BEG[13]
port 185 nsew signal output
flabel metal2 s 12992 114800 13104 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_N4BEG[14]
port 186 nsew signal output
flabel metal2 s 13216 114800 13328 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_N4BEG[15]
port 187 nsew signal output
flabel metal2 s 10080 114800 10192 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_N4BEG[1]
port 188 nsew signal output
flabel metal2 s 10304 114800 10416 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_N4BEG[2]
port 189 nsew signal output
flabel metal2 s 10528 114800 10640 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_N4BEG[3]
port 190 nsew signal output
flabel metal2 s 10752 114800 10864 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_N4BEG[4]
port 191 nsew signal output
flabel metal2 s 10976 114800 11088 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_N4BEG[5]
port 192 nsew signal output
flabel metal2 s 11200 114800 11312 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_N4BEG[6]
port 193 nsew signal output
flabel metal2 s 11424 114800 11536 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_N4BEG[7]
port 194 nsew signal output
flabel metal2 s 11648 114800 11760 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_N4BEG[8]
port 195 nsew signal output
flabel metal2 s 11872 114800 11984 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_N4BEG[9]
port 196 nsew signal output
flabel metal2 s 13440 114800 13552 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_S1END[0]
port 197 nsew signal input
flabel metal2 s 13664 114800 13776 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_S1END[1]
port 198 nsew signal input
flabel metal2 s 13888 114800 14000 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_S1END[2]
port 199 nsew signal input
flabel metal2 s 14112 114800 14224 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_S1END[3]
port 200 nsew signal input
flabel metal2 s 16128 114800 16240 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_S2END[0]
port 201 nsew signal input
flabel metal2 s 16352 114800 16464 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_S2END[1]
port 202 nsew signal input
flabel metal2 s 16576 114800 16688 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_S2END[2]
port 203 nsew signal input
flabel metal2 s 16800 114800 16912 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_S2END[3]
port 204 nsew signal input
flabel metal2 s 17024 114800 17136 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_S2END[4]
port 205 nsew signal input
flabel metal2 s 17248 114800 17360 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_S2END[5]
port 206 nsew signal input
flabel metal2 s 17472 114800 17584 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_S2END[6]
port 207 nsew signal input
flabel metal2 s 17696 114800 17808 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_S2END[7]
port 208 nsew signal input
flabel metal2 s 14336 114800 14448 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_S2MID[0]
port 209 nsew signal input
flabel metal2 s 14560 114800 14672 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_S2MID[1]
port 210 nsew signal input
flabel metal2 s 14784 114800 14896 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_S2MID[2]
port 211 nsew signal input
flabel metal2 s 15008 114800 15120 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_S2MID[3]
port 212 nsew signal input
flabel metal2 s 15232 114800 15344 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_S2MID[4]
port 213 nsew signal input
flabel metal2 s 15456 114800 15568 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_S2MID[5]
port 214 nsew signal input
flabel metal2 s 15680 114800 15792 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_S2MID[6]
port 215 nsew signal input
flabel metal2 s 15904 114800 16016 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_S2MID[7]
port 216 nsew signal input
flabel metal2 s 17920 114800 18032 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_S4END[0]
port 217 nsew signal input
flabel metal2 s 20160 114800 20272 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_S4END[10]
port 218 nsew signal input
flabel metal2 s 20384 114800 20496 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_S4END[11]
port 219 nsew signal input
flabel metal2 s 20608 114800 20720 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_S4END[12]
port 220 nsew signal input
flabel metal2 s 20832 114800 20944 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_S4END[13]
port 221 nsew signal input
flabel metal2 s 21056 114800 21168 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_S4END[14]
port 222 nsew signal input
flabel metal2 s 21280 114800 21392 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_S4END[15]
port 223 nsew signal input
flabel metal2 s 18144 114800 18256 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_S4END[1]
port 224 nsew signal input
flabel metal2 s 18368 114800 18480 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_S4END[2]
port 225 nsew signal input
flabel metal2 s 18592 114800 18704 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_S4END[3]
port 226 nsew signal input
flabel metal2 s 18816 114800 18928 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_S4END[4]
port 227 nsew signal input
flabel metal2 s 19040 114800 19152 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_S4END[5]
port 228 nsew signal input
flabel metal2 s 19264 114800 19376 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_S4END[6]
port 229 nsew signal input
flabel metal2 s 19488 114800 19600 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_S4END[7]
port 230 nsew signal input
flabel metal2 s 19712 114800 19824 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_S4END[8]
port 231 nsew signal input
flabel metal2 s 19936 114800 20048 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_S4END[9]
port 232 nsew signal input
flabel metal2 s 21504 114800 21616 114912 0 FreeSans 448 0 0 0 Tile_X0Y0_UserCLKo
port 233 nsew signal output
flabel metal3 s 0 57680 112 57792 0 FreeSans 448 0 0 0 Tile_X0Y0_W1BEG[0]
port 234 nsew signal output
flabel metal3 s 0 58128 112 58240 0 FreeSans 448 0 0 0 Tile_X0Y0_W1BEG[1]
port 235 nsew signal output
flabel metal3 s 0 58576 112 58688 0 FreeSans 448 0 0 0 Tile_X0Y0_W1BEG[2]
port 236 nsew signal output
flabel metal3 s 0 59024 112 59136 0 FreeSans 448 0 0 0 Tile_X0Y0_W1BEG[3]
port 237 nsew signal output
flabel metal3 s 0 59472 112 59584 0 FreeSans 448 0 0 0 Tile_X0Y0_W2BEG[0]
port 238 nsew signal output
flabel metal3 s 0 59920 112 60032 0 FreeSans 448 0 0 0 Tile_X0Y0_W2BEG[1]
port 239 nsew signal output
flabel metal3 s 0 60368 112 60480 0 FreeSans 448 0 0 0 Tile_X0Y0_W2BEG[2]
port 240 nsew signal output
flabel metal3 s 0 60816 112 60928 0 FreeSans 448 0 0 0 Tile_X0Y0_W2BEG[3]
port 241 nsew signal output
flabel metal3 s 0 61264 112 61376 0 FreeSans 448 0 0 0 Tile_X0Y0_W2BEG[4]
port 242 nsew signal output
flabel metal3 s 0 61712 112 61824 0 FreeSans 448 0 0 0 Tile_X0Y0_W2BEG[5]
port 243 nsew signal output
flabel metal3 s 0 62160 112 62272 0 FreeSans 448 0 0 0 Tile_X0Y0_W2BEG[6]
port 244 nsew signal output
flabel metal3 s 0 62608 112 62720 0 FreeSans 448 0 0 0 Tile_X0Y0_W2BEG[7]
port 245 nsew signal output
flabel metal3 s 0 63056 112 63168 0 FreeSans 448 0 0 0 Tile_X0Y0_W2BEGb[0]
port 246 nsew signal output
flabel metal3 s 0 63504 112 63616 0 FreeSans 448 0 0 0 Tile_X0Y0_W2BEGb[1]
port 247 nsew signal output
flabel metal3 s 0 63952 112 64064 0 FreeSans 448 0 0 0 Tile_X0Y0_W2BEGb[2]
port 248 nsew signal output
flabel metal3 s 0 64400 112 64512 0 FreeSans 448 0 0 0 Tile_X0Y0_W2BEGb[3]
port 249 nsew signal output
flabel metal3 s 0 64848 112 64960 0 FreeSans 448 0 0 0 Tile_X0Y0_W2BEGb[4]
port 250 nsew signal output
flabel metal3 s 0 65296 112 65408 0 FreeSans 448 0 0 0 Tile_X0Y0_W2BEGb[5]
port 251 nsew signal output
flabel metal3 s 0 65744 112 65856 0 FreeSans 448 0 0 0 Tile_X0Y0_W2BEGb[6]
port 252 nsew signal output
flabel metal3 s 0 66192 112 66304 0 FreeSans 448 0 0 0 Tile_X0Y0_W2BEGb[7]
port 253 nsew signal output
flabel metal3 s 0 73808 112 73920 0 FreeSans 448 0 0 0 Tile_X0Y0_W6BEG[0]
port 254 nsew signal output
flabel metal3 s 0 78288 112 78400 0 FreeSans 448 0 0 0 Tile_X0Y0_W6BEG[10]
port 255 nsew signal output
flabel metal3 s 0 78736 112 78848 0 FreeSans 448 0 0 0 Tile_X0Y0_W6BEG[11]
port 256 nsew signal output
flabel metal3 s 0 74256 112 74368 0 FreeSans 448 0 0 0 Tile_X0Y0_W6BEG[1]
port 257 nsew signal output
flabel metal3 s 0 74704 112 74816 0 FreeSans 448 0 0 0 Tile_X0Y0_W6BEG[2]
port 258 nsew signal output
flabel metal3 s 0 75152 112 75264 0 FreeSans 448 0 0 0 Tile_X0Y0_W6BEG[3]
port 259 nsew signal output
flabel metal3 s 0 75600 112 75712 0 FreeSans 448 0 0 0 Tile_X0Y0_W6BEG[4]
port 260 nsew signal output
flabel metal3 s 0 76048 112 76160 0 FreeSans 448 0 0 0 Tile_X0Y0_W6BEG[5]
port 261 nsew signal output
flabel metal3 s 0 76496 112 76608 0 FreeSans 448 0 0 0 Tile_X0Y0_W6BEG[6]
port 262 nsew signal output
flabel metal3 s 0 76944 112 77056 0 FreeSans 448 0 0 0 Tile_X0Y0_W6BEG[7]
port 263 nsew signal output
flabel metal3 s 0 77392 112 77504 0 FreeSans 448 0 0 0 Tile_X0Y0_W6BEG[8]
port 264 nsew signal output
flabel metal3 s 0 77840 112 77952 0 FreeSans 448 0 0 0 Tile_X0Y0_W6BEG[9]
port 265 nsew signal output
flabel metal3 s 0 66640 112 66752 0 FreeSans 448 0 0 0 Tile_X0Y0_WW4BEG[0]
port 266 nsew signal output
flabel metal3 s 0 71120 112 71232 0 FreeSans 448 0 0 0 Tile_X0Y0_WW4BEG[10]
port 267 nsew signal output
flabel metal3 s 0 71568 112 71680 0 FreeSans 448 0 0 0 Tile_X0Y0_WW4BEG[11]
port 268 nsew signal output
flabel metal3 s 0 72016 112 72128 0 FreeSans 448 0 0 0 Tile_X0Y0_WW4BEG[12]
port 269 nsew signal output
flabel metal3 s 0 72464 112 72576 0 FreeSans 448 0 0 0 Tile_X0Y0_WW4BEG[13]
port 270 nsew signal output
flabel metal3 s 0 72912 112 73024 0 FreeSans 448 0 0 0 Tile_X0Y0_WW4BEG[14]
port 271 nsew signal output
flabel metal3 s 0 73360 112 73472 0 FreeSans 448 0 0 0 Tile_X0Y0_WW4BEG[15]
port 272 nsew signal output
flabel metal3 s 0 67088 112 67200 0 FreeSans 448 0 0 0 Tile_X0Y0_WW4BEG[1]
port 273 nsew signal output
flabel metal3 s 0 67536 112 67648 0 FreeSans 448 0 0 0 Tile_X0Y0_WW4BEG[2]
port 274 nsew signal output
flabel metal3 s 0 67984 112 68096 0 FreeSans 448 0 0 0 Tile_X0Y0_WW4BEG[3]
port 275 nsew signal output
flabel metal3 s 0 68432 112 68544 0 FreeSans 448 0 0 0 Tile_X0Y0_WW4BEG[4]
port 276 nsew signal output
flabel metal3 s 0 68880 112 68992 0 FreeSans 448 0 0 0 Tile_X0Y0_WW4BEG[5]
port 277 nsew signal output
flabel metal3 s 0 69328 112 69440 0 FreeSans 448 0 0 0 Tile_X0Y0_WW4BEG[6]
port 278 nsew signal output
flabel metal3 s 0 69776 112 69888 0 FreeSans 448 0 0 0 Tile_X0Y0_WW4BEG[7]
port 279 nsew signal output
flabel metal3 s 0 70224 112 70336 0 FreeSans 448 0 0 0 Tile_X0Y0_WW4BEG[8]
port 280 nsew signal output
flabel metal3 s 0 70672 112 70784 0 FreeSans 448 0 0 0 Tile_X0Y0_WW4BEG[9]
port 281 nsew signal output
flabel metal3 s 0 21728 112 21840 0 FreeSans 448 0 0 0 Tile_X0Y1_E1END[0]
port 282 nsew signal input
flabel metal3 s 0 22176 112 22288 0 FreeSans 448 0 0 0 Tile_X0Y1_E1END[1]
port 283 nsew signal input
flabel metal3 s 0 22624 112 22736 0 FreeSans 448 0 0 0 Tile_X0Y1_E1END[2]
port 284 nsew signal input
flabel metal3 s 0 23072 112 23184 0 FreeSans 448 0 0 0 Tile_X0Y1_E1END[3]
port 285 nsew signal input
flabel metal3 s 0 27104 112 27216 0 FreeSans 448 0 0 0 Tile_X0Y1_E2END[0]
port 286 nsew signal input
flabel metal3 s 0 27552 112 27664 0 FreeSans 448 0 0 0 Tile_X0Y1_E2END[1]
port 287 nsew signal input
flabel metal3 s 0 28000 112 28112 0 FreeSans 448 0 0 0 Tile_X0Y1_E2END[2]
port 288 nsew signal input
flabel metal3 s 0 28448 112 28560 0 FreeSans 448 0 0 0 Tile_X0Y1_E2END[3]
port 289 nsew signal input
flabel metal3 s 0 28896 112 29008 0 FreeSans 448 0 0 0 Tile_X0Y1_E2END[4]
port 290 nsew signal input
flabel metal3 s 0 29344 112 29456 0 FreeSans 448 0 0 0 Tile_X0Y1_E2END[5]
port 291 nsew signal input
flabel metal3 s 0 29792 112 29904 0 FreeSans 448 0 0 0 Tile_X0Y1_E2END[6]
port 292 nsew signal input
flabel metal3 s 0 30240 112 30352 0 FreeSans 448 0 0 0 Tile_X0Y1_E2END[7]
port 293 nsew signal input
flabel metal3 s 0 23520 112 23632 0 FreeSans 448 0 0 0 Tile_X0Y1_E2MID[0]
port 294 nsew signal input
flabel metal3 s 0 23968 112 24080 0 FreeSans 448 0 0 0 Tile_X0Y1_E2MID[1]
port 295 nsew signal input
flabel metal3 s 0 24416 112 24528 0 FreeSans 448 0 0 0 Tile_X0Y1_E2MID[2]
port 296 nsew signal input
flabel metal3 s 0 24864 112 24976 0 FreeSans 448 0 0 0 Tile_X0Y1_E2MID[3]
port 297 nsew signal input
flabel metal3 s 0 25312 112 25424 0 FreeSans 448 0 0 0 Tile_X0Y1_E2MID[4]
port 298 nsew signal input
flabel metal3 s 0 25760 112 25872 0 FreeSans 448 0 0 0 Tile_X0Y1_E2MID[5]
port 299 nsew signal input
flabel metal3 s 0 26208 112 26320 0 FreeSans 448 0 0 0 Tile_X0Y1_E2MID[6]
port 300 nsew signal input
flabel metal3 s 0 26656 112 26768 0 FreeSans 448 0 0 0 Tile_X0Y1_E2MID[7]
port 301 nsew signal input
flabel metal3 s 0 37856 112 37968 0 FreeSans 448 0 0 0 Tile_X0Y1_E6END[0]
port 302 nsew signal input
flabel metal3 s 0 42336 112 42448 0 FreeSans 448 0 0 0 Tile_X0Y1_E6END[10]
port 303 nsew signal input
flabel metal3 s 0 42784 112 42896 0 FreeSans 448 0 0 0 Tile_X0Y1_E6END[11]
port 304 nsew signal input
flabel metal3 s 0 38304 112 38416 0 FreeSans 448 0 0 0 Tile_X0Y1_E6END[1]
port 305 nsew signal input
flabel metal3 s 0 38752 112 38864 0 FreeSans 448 0 0 0 Tile_X0Y1_E6END[2]
port 306 nsew signal input
flabel metal3 s 0 39200 112 39312 0 FreeSans 448 0 0 0 Tile_X0Y1_E6END[3]
port 307 nsew signal input
flabel metal3 s 0 39648 112 39760 0 FreeSans 448 0 0 0 Tile_X0Y1_E6END[4]
port 308 nsew signal input
flabel metal3 s 0 40096 112 40208 0 FreeSans 448 0 0 0 Tile_X0Y1_E6END[5]
port 309 nsew signal input
flabel metal3 s 0 40544 112 40656 0 FreeSans 448 0 0 0 Tile_X0Y1_E6END[6]
port 310 nsew signal input
flabel metal3 s 0 40992 112 41104 0 FreeSans 448 0 0 0 Tile_X0Y1_E6END[7]
port 311 nsew signal input
flabel metal3 s 0 41440 112 41552 0 FreeSans 448 0 0 0 Tile_X0Y1_E6END[8]
port 312 nsew signal input
flabel metal3 s 0 41888 112 42000 0 FreeSans 448 0 0 0 Tile_X0Y1_E6END[9]
port 313 nsew signal input
flabel metal3 s 0 30688 112 30800 0 FreeSans 448 0 0 0 Tile_X0Y1_EE4END[0]
port 314 nsew signal input
flabel metal3 s 0 35168 112 35280 0 FreeSans 448 0 0 0 Tile_X0Y1_EE4END[10]
port 315 nsew signal input
flabel metal3 s 0 35616 112 35728 0 FreeSans 448 0 0 0 Tile_X0Y1_EE4END[11]
port 316 nsew signal input
flabel metal3 s 0 36064 112 36176 0 FreeSans 448 0 0 0 Tile_X0Y1_EE4END[12]
port 317 nsew signal input
flabel metal3 s 0 36512 112 36624 0 FreeSans 448 0 0 0 Tile_X0Y1_EE4END[13]
port 318 nsew signal input
flabel metal3 s 0 36960 112 37072 0 FreeSans 448 0 0 0 Tile_X0Y1_EE4END[14]
port 319 nsew signal input
flabel metal3 s 0 37408 112 37520 0 FreeSans 448 0 0 0 Tile_X0Y1_EE4END[15]
port 320 nsew signal input
flabel metal3 s 0 31136 112 31248 0 FreeSans 448 0 0 0 Tile_X0Y1_EE4END[1]
port 321 nsew signal input
flabel metal3 s 0 31584 112 31696 0 FreeSans 448 0 0 0 Tile_X0Y1_EE4END[2]
port 322 nsew signal input
flabel metal3 s 0 32032 112 32144 0 FreeSans 448 0 0 0 Tile_X0Y1_EE4END[3]
port 323 nsew signal input
flabel metal3 s 0 32480 112 32592 0 FreeSans 448 0 0 0 Tile_X0Y1_EE4END[4]
port 324 nsew signal input
flabel metal3 s 0 32928 112 33040 0 FreeSans 448 0 0 0 Tile_X0Y1_EE4END[5]
port 325 nsew signal input
flabel metal3 s 0 33376 112 33488 0 FreeSans 448 0 0 0 Tile_X0Y1_EE4END[6]
port 326 nsew signal input
flabel metal3 s 0 33824 112 33936 0 FreeSans 448 0 0 0 Tile_X0Y1_EE4END[7]
port 327 nsew signal input
flabel metal3 s 0 34272 112 34384 0 FreeSans 448 0 0 0 Tile_X0Y1_EE4END[8]
port 328 nsew signal input
flabel metal3 s 0 34720 112 34832 0 FreeSans 448 0 0 0 Tile_X0Y1_EE4END[9]
port 329 nsew signal input
flabel metal3 s 0 43232 112 43344 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData[0]
port 330 nsew signal input
flabel metal3 s 0 47712 112 47824 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData[10]
port 331 nsew signal input
flabel metal3 s 0 48160 112 48272 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData[11]
port 332 nsew signal input
flabel metal3 s 0 48608 112 48720 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData[12]
port 333 nsew signal input
flabel metal3 s 0 49056 112 49168 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData[13]
port 334 nsew signal input
flabel metal3 s 0 49504 112 49616 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData[14]
port 335 nsew signal input
flabel metal3 s 0 49952 112 50064 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData[15]
port 336 nsew signal input
flabel metal3 s 0 50400 112 50512 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData[16]
port 337 nsew signal input
flabel metal3 s 0 50848 112 50960 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData[17]
port 338 nsew signal input
flabel metal3 s 0 51296 112 51408 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData[18]
port 339 nsew signal input
flabel metal3 s 0 51744 112 51856 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData[19]
port 340 nsew signal input
flabel metal3 s 0 43680 112 43792 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData[1]
port 341 nsew signal input
flabel metal3 s 0 52192 112 52304 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData[20]
port 342 nsew signal input
flabel metal3 s 0 52640 112 52752 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData[21]
port 343 nsew signal input
flabel metal3 s 0 53088 112 53200 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData[22]
port 344 nsew signal input
flabel metal3 s 0 53536 112 53648 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData[23]
port 345 nsew signal input
flabel metal3 s 0 53984 112 54096 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData[24]
port 346 nsew signal input
flabel metal3 s 0 54432 112 54544 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData[25]
port 347 nsew signal input
flabel metal3 s 0 54880 112 54992 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData[26]
port 348 nsew signal input
flabel metal3 s 0 55328 112 55440 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData[27]
port 349 nsew signal input
flabel metal3 s 0 55776 112 55888 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData[28]
port 350 nsew signal input
flabel metal3 s 0 56224 112 56336 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData[29]
port 351 nsew signal input
flabel metal3 s 0 44128 112 44240 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData[2]
port 352 nsew signal input
flabel metal3 s 0 56672 112 56784 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData[30]
port 353 nsew signal input
flabel metal3 s 0 57120 112 57232 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData[31]
port 354 nsew signal input
flabel metal3 s 0 44576 112 44688 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData[3]
port 355 nsew signal input
flabel metal3 s 0 45024 112 45136 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData[4]
port 356 nsew signal input
flabel metal3 s 0 45472 112 45584 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData[5]
port 357 nsew signal input
flabel metal3 s 0 45920 112 46032 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData[6]
port 358 nsew signal input
flabel metal3 s 0 46368 112 46480 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData[7]
port 359 nsew signal input
flabel metal3 s 0 46816 112 46928 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData[8]
port 360 nsew signal input
flabel metal3 s 0 47264 112 47376 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData[9]
port 361 nsew signal input
flabel metal3 s 31584 39872 31696 39984 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData_O[0]
port 362 nsew signal output
flabel metal3 s 31584 51072 31696 51184 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData_O[10]
port 363 nsew signal output
flabel metal3 s 31584 52192 31696 52304 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData_O[11]
port 364 nsew signal output
flabel metal3 s 31584 53312 31696 53424 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData_O[12]
port 365 nsew signal output
flabel metal3 s 31584 54432 31696 54544 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData_O[13]
port 366 nsew signal output
flabel metal3 s 31584 55552 31696 55664 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData_O[14]
port 367 nsew signal output
flabel metal3 s 31584 56672 31696 56784 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData_O[15]
port 368 nsew signal output
flabel metal3 s 31584 57792 31696 57904 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData_O[16]
port 369 nsew signal output
flabel metal3 s 31584 58912 31696 59024 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData_O[17]
port 370 nsew signal output
flabel metal3 s 31584 60032 31696 60144 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData_O[18]
port 371 nsew signal output
flabel metal3 s 31584 61152 31696 61264 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData_O[19]
port 372 nsew signal output
flabel metal3 s 31584 40992 31696 41104 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData_O[1]
port 373 nsew signal output
flabel metal3 s 31584 62272 31696 62384 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData_O[20]
port 374 nsew signal output
flabel metal3 s 31584 63392 31696 63504 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData_O[21]
port 375 nsew signal output
flabel metal3 s 31584 64512 31696 64624 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData_O[22]
port 376 nsew signal output
flabel metal3 s 31584 65632 31696 65744 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData_O[23]
port 377 nsew signal output
flabel metal3 s 31584 66752 31696 66864 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData_O[24]
port 378 nsew signal output
flabel metal3 s 31584 67872 31696 67984 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData_O[25]
port 379 nsew signal output
flabel metal3 s 31584 68992 31696 69104 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData_O[26]
port 380 nsew signal output
flabel metal3 s 31584 70112 31696 70224 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData_O[27]
port 381 nsew signal output
flabel metal3 s 31584 71232 31696 71344 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData_O[28]
port 382 nsew signal output
flabel metal3 s 31584 72352 31696 72464 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData_O[29]
port 383 nsew signal output
flabel metal3 s 31584 42112 31696 42224 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData_O[2]
port 384 nsew signal output
flabel metal3 s 31584 73472 31696 73584 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData_O[30]
port 385 nsew signal output
flabel metal3 s 31584 74592 31696 74704 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData_O[31]
port 386 nsew signal output
flabel metal3 s 31584 43232 31696 43344 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData_O[3]
port 387 nsew signal output
flabel metal3 s 31584 44352 31696 44464 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData_O[4]
port 388 nsew signal output
flabel metal3 s 31584 45472 31696 45584 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData_O[5]
port 389 nsew signal output
flabel metal3 s 31584 46592 31696 46704 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData_O[6]
port 390 nsew signal output
flabel metal3 s 31584 47712 31696 47824 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData_O[7]
port 391 nsew signal output
flabel metal3 s 31584 48832 31696 48944 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData_O[8]
port 392 nsew signal output
flabel metal3 s 31584 49952 31696 50064 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameData_O[9]
port 393 nsew signal output
flabel metal2 s 21728 0 21840 112 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameStrobe[0]
port 394 nsew signal input
flabel metal2 s 23968 0 24080 112 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameStrobe[10]
port 395 nsew signal input
flabel metal2 s 24192 0 24304 112 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameStrobe[11]
port 396 nsew signal input
flabel metal2 s 24416 0 24528 112 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameStrobe[12]
port 397 nsew signal input
flabel metal2 s 24640 0 24752 112 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameStrobe[13]
port 398 nsew signal input
flabel metal2 s 24864 0 24976 112 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameStrobe[14]
port 399 nsew signal input
flabel metal2 s 25088 0 25200 112 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameStrobe[15]
port 400 nsew signal input
flabel metal2 s 25312 0 25424 112 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameStrobe[16]
port 401 nsew signal input
flabel metal2 s 25536 0 25648 112 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameStrobe[17]
port 402 nsew signal input
flabel metal2 s 25760 0 25872 112 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameStrobe[18]
port 403 nsew signal input
flabel metal2 s 25984 0 26096 112 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameStrobe[19]
port 404 nsew signal input
flabel metal2 s 21952 0 22064 112 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameStrobe[1]
port 405 nsew signal input
flabel metal2 s 22176 0 22288 112 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameStrobe[2]
port 406 nsew signal input
flabel metal2 s 22400 0 22512 112 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameStrobe[3]
port 407 nsew signal input
flabel metal2 s 22624 0 22736 112 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameStrobe[4]
port 408 nsew signal input
flabel metal2 s 22848 0 22960 112 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameStrobe[5]
port 409 nsew signal input
flabel metal2 s 23072 0 23184 112 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameStrobe[6]
port 410 nsew signal input
flabel metal2 s 23296 0 23408 112 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameStrobe[7]
port 411 nsew signal input
flabel metal2 s 23520 0 23632 112 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameStrobe[8]
port 412 nsew signal input
flabel metal2 s 23744 0 23856 112 0 FreeSans 448 0 0 0 Tile_X0Y1_FrameStrobe[9]
port 413 nsew signal input
flabel metal2 s 5376 0 5488 112 0 FreeSans 448 0 0 0 Tile_X0Y1_N1END[0]
port 414 nsew signal input
flabel metal2 s 5600 0 5712 112 0 FreeSans 448 0 0 0 Tile_X0Y1_N1END[1]
port 415 nsew signal input
flabel metal2 s 5824 0 5936 112 0 FreeSans 448 0 0 0 Tile_X0Y1_N1END[2]
port 416 nsew signal input
flabel metal2 s 6048 0 6160 112 0 FreeSans 448 0 0 0 Tile_X0Y1_N1END[3]
port 417 nsew signal input
flabel metal2 s 8064 0 8176 112 0 FreeSans 448 0 0 0 Tile_X0Y1_N2END[0]
port 418 nsew signal input
flabel metal2 s 8288 0 8400 112 0 FreeSans 448 0 0 0 Tile_X0Y1_N2END[1]
port 419 nsew signal input
flabel metal2 s 8512 0 8624 112 0 FreeSans 448 0 0 0 Tile_X0Y1_N2END[2]
port 420 nsew signal input
flabel metal2 s 8736 0 8848 112 0 FreeSans 448 0 0 0 Tile_X0Y1_N2END[3]
port 421 nsew signal input
flabel metal2 s 8960 0 9072 112 0 FreeSans 448 0 0 0 Tile_X0Y1_N2END[4]
port 422 nsew signal input
flabel metal2 s 9184 0 9296 112 0 FreeSans 448 0 0 0 Tile_X0Y1_N2END[5]
port 423 nsew signal input
flabel metal2 s 9408 0 9520 112 0 FreeSans 448 0 0 0 Tile_X0Y1_N2END[6]
port 424 nsew signal input
flabel metal2 s 9632 0 9744 112 0 FreeSans 448 0 0 0 Tile_X0Y1_N2END[7]
port 425 nsew signal input
flabel metal2 s 6272 0 6384 112 0 FreeSans 448 0 0 0 Tile_X0Y1_N2MID[0]
port 426 nsew signal input
flabel metal2 s 6496 0 6608 112 0 FreeSans 448 0 0 0 Tile_X0Y1_N2MID[1]
port 427 nsew signal input
flabel metal2 s 6720 0 6832 112 0 FreeSans 448 0 0 0 Tile_X0Y1_N2MID[2]
port 428 nsew signal input
flabel metal2 s 6944 0 7056 112 0 FreeSans 448 0 0 0 Tile_X0Y1_N2MID[3]
port 429 nsew signal input
flabel metal2 s 7168 0 7280 112 0 FreeSans 448 0 0 0 Tile_X0Y1_N2MID[4]
port 430 nsew signal input
flabel metal2 s 7392 0 7504 112 0 FreeSans 448 0 0 0 Tile_X0Y1_N2MID[5]
port 431 nsew signal input
flabel metal2 s 7616 0 7728 112 0 FreeSans 448 0 0 0 Tile_X0Y1_N2MID[6]
port 432 nsew signal input
flabel metal2 s 7840 0 7952 112 0 FreeSans 448 0 0 0 Tile_X0Y1_N2MID[7]
port 433 nsew signal input
flabel metal2 s 9856 0 9968 112 0 FreeSans 448 0 0 0 Tile_X0Y1_N4END[0]
port 434 nsew signal input
flabel metal2 s 12096 0 12208 112 0 FreeSans 448 0 0 0 Tile_X0Y1_N4END[10]
port 435 nsew signal input
flabel metal2 s 12320 0 12432 112 0 FreeSans 448 0 0 0 Tile_X0Y1_N4END[11]
port 436 nsew signal input
flabel metal2 s 12544 0 12656 112 0 FreeSans 448 0 0 0 Tile_X0Y1_N4END[12]
port 437 nsew signal input
flabel metal2 s 12768 0 12880 112 0 FreeSans 448 0 0 0 Tile_X0Y1_N4END[13]
port 438 nsew signal input
flabel metal2 s 12992 0 13104 112 0 FreeSans 448 0 0 0 Tile_X0Y1_N4END[14]
port 439 nsew signal input
flabel metal2 s 13216 0 13328 112 0 FreeSans 448 0 0 0 Tile_X0Y1_N4END[15]
port 440 nsew signal input
flabel metal2 s 10080 0 10192 112 0 FreeSans 448 0 0 0 Tile_X0Y1_N4END[1]
port 441 nsew signal input
flabel metal2 s 10304 0 10416 112 0 FreeSans 448 0 0 0 Tile_X0Y1_N4END[2]
port 442 nsew signal input
flabel metal2 s 10528 0 10640 112 0 FreeSans 448 0 0 0 Tile_X0Y1_N4END[3]
port 443 nsew signal input
flabel metal2 s 10752 0 10864 112 0 FreeSans 448 0 0 0 Tile_X0Y1_N4END[4]
port 444 nsew signal input
flabel metal2 s 10976 0 11088 112 0 FreeSans 448 0 0 0 Tile_X0Y1_N4END[5]
port 445 nsew signal input
flabel metal2 s 11200 0 11312 112 0 FreeSans 448 0 0 0 Tile_X0Y1_N4END[6]
port 446 nsew signal input
flabel metal2 s 11424 0 11536 112 0 FreeSans 448 0 0 0 Tile_X0Y1_N4END[7]
port 447 nsew signal input
flabel metal2 s 11648 0 11760 112 0 FreeSans 448 0 0 0 Tile_X0Y1_N4END[8]
port 448 nsew signal input
flabel metal2 s 11872 0 11984 112 0 FreeSans 448 0 0 0 Tile_X0Y1_N4END[9]
port 449 nsew signal input
flabel metal2 s 13440 0 13552 112 0 FreeSans 448 0 0 0 Tile_X0Y1_S1BEG[0]
port 450 nsew signal output
flabel metal2 s 13664 0 13776 112 0 FreeSans 448 0 0 0 Tile_X0Y1_S1BEG[1]
port 451 nsew signal output
flabel metal2 s 13888 0 14000 112 0 FreeSans 448 0 0 0 Tile_X0Y1_S1BEG[2]
port 452 nsew signal output
flabel metal2 s 14112 0 14224 112 0 FreeSans 448 0 0 0 Tile_X0Y1_S1BEG[3]
port 453 nsew signal output
flabel metal2 s 14336 0 14448 112 0 FreeSans 448 0 0 0 Tile_X0Y1_S2BEG[0]
port 454 nsew signal output
flabel metal2 s 14560 0 14672 112 0 FreeSans 448 0 0 0 Tile_X0Y1_S2BEG[1]
port 455 nsew signal output
flabel metal2 s 14784 0 14896 112 0 FreeSans 448 0 0 0 Tile_X0Y1_S2BEG[2]
port 456 nsew signal output
flabel metal2 s 15008 0 15120 112 0 FreeSans 448 0 0 0 Tile_X0Y1_S2BEG[3]
port 457 nsew signal output
flabel metal2 s 15232 0 15344 112 0 FreeSans 448 0 0 0 Tile_X0Y1_S2BEG[4]
port 458 nsew signal output
flabel metal2 s 15456 0 15568 112 0 FreeSans 448 0 0 0 Tile_X0Y1_S2BEG[5]
port 459 nsew signal output
flabel metal2 s 15680 0 15792 112 0 FreeSans 448 0 0 0 Tile_X0Y1_S2BEG[6]
port 460 nsew signal output
flabel metal2 s 15904 0 16016 112 0 FreeSans 448 0 0 0 Tile_X0Y1_S2BEG[7]
port 461 nsew signal output
flabel metal2 s 16128 0 16240 112 0 FreeSans 448 0 0 0 Tile_X0Y1_S2BEGb[0]
port 462 nsew signal output
flabel metal2 s 16352 0 16464 112 0 FreeSans 448 0 0 0 Tile_X0Y1_S2BEGb[1]
port 463 nsew signal output
flabel metal2 s 16576 0 16688 112 0 FreeSans 448 0 0 0 Tile_X0Y1_S2BEGb[2]
port 464 nsew signal output
flabel metal2 s 16800 0 16912 112 0 FreeSans 448 0 0 0 Tile_X0Y1_S2BEGb[3]
port 465 nsew signal output
flabel metal2 s 17024 0 17136 112 0 FreeSans 448 0 0 0 Tile_X0Y1_S2BEGb[4]
port 466 nsew signal output
flabel metal2 s 17248 0 17360 112 0 FreeSans 448 0 0 0 Tile_X0Y1_S2BEGb[5]
port 467 nsew signal output
flabel metal2 s 17472 0 17584 112 0 FreeSans 448 0 0 0 Tile_X0Y1_S2BEGb[6]
port 468 nsew signal output
flabel metal2 s 17696 0 17808 112 0 FreeSans 448 0 0 0 Tile_X0Y1_S2BEGb[7]
port 469 nsew signal output
flabel metal2 s 17920 0 18032 112 0 FreeSans 448 0 0 0 Tile_X0Y1_S4BEG[0]
port 470 nsew signal output
flabel metal2 s 20160 0 20272 112 0 FreeSans 448 0 0 0 Tile_X0Y1_S4BEG[10]
port 471 nsew signal output
flabel metal2 s 20384 0 20496 112 0 FreeSans 448 0 0 0 Tile_X0Y1_S4BEG[11]
port 472 nsew signal output
flabel metal2 s 20608 0 20720 112 0 FreeSans 448 0 0 0 Tile_X0Y1_S4BEG[12]
port 473 nsew signal output
flabel metal2 s 20832 0 20944 112 0 FreeSans 448 0 0 0 Tile_X0Y1_S4BEG[13]
port 474 nsew signal output
flabel metal2 s 21056 0 21168 112 0 FreeSans 448 0 0 0 Tile_X0Y1_S4BEG[14]
port 475 nsew signal output
flabel metal2 s 21280 0 21392 112 0 FreeSans 448 0 0 0 Tile_X0Y1_S4BEG[15]
port 476 nsew signal output
flabel metal2 s 18144 0 18256 112 0 FreeSans 448 0 0 0 Tile_X0Y1_S4BEG[1]
port 477 nsew signal output
flabel metal2 s 18368 0 18480 112 0 FreeSans 448 0 0 0 Tile_X0Y1_S4BEG[2]
port 478 nsew signal output
flabel metal2 s 18592 0 18704 112 0 FreeSans 448 0 0 0 Tile_X0Y1_S4BEG[3]
port 479 nsew signal output
flabel metal2 s 18816 0 18928 112 0 FreeSans 448 0 0 0 Tile_X0Y1_S4BEG[4]
port 480 nsew signal output
flabel metal2 s 19040 0 19152 112 0 FreeSans 448 0 0 0 Tile_X0Y1_S4BEG[5]
port 481 nsew signal output
flabel metal2 s 19264 0 19376 112 0 FreeSans 448 0 0 0 Tile_X0Y1_S4BEG[6]
port 482 nsew signal output
flabel metal2 s 19488 0 19600 112 0 FreeSans 448 0 0 0 Tile_X0Y1_S4BEG[7]
port 483 nsew signal output
flabel metal2 s 19712 0 19824 112 0 FreeSans 448 0 0 0 Tile_X0Y1_S4BEG[8]
port 484 nsew signal output
flabel metal2 s 19936 0 20048 112 0 FreeSans 448 0 0 0 Tile_X0Y1_S4BEG[9]
port 485 nsew signal output
flabel metal2 s 21504 0 21616 112 0 FreeSans 448 0 0 0 Tile_X0Y1_UserCLK
port 486 nsew signal input
flabel metal3 s 0 224 112 336 0 FreeSans 448 0 0 0 Tile_X0Y1_W1BEG[0]
port 487 nsew signal output
flabel metal3 s 0 672 112 784 0 FreeSans 448 0 0 0 Tile_X0Y1_W1BEG[1]
port 488 nsew signal output
flabel metal3 s 0 1120 112 1232 0 FreeSans 448 0 0 0 Tile_X0Y1_W1BEG[2]
port 489 nsew signal output
flabel metal3 s 0 1568 112 1680 0 FreeSans 448 0 0 0 Tile_X0Y1_W1BEG[3]
port 490 nsew signal output
flabel metal3 s 0 2016 112 2128 0 FreeSans 448 0 0 0 Tile_X0Y1_W2BEG[0]
port 491 nsew signal output
flabel metal3 s 0 2464 112 2576 0 FreeSans 448 0 0 0 Tile_X0Y1_W2BEG[1]
port 492 nsew signal output
flabel metal3 s 0 2912 112 3024 0 FreeSans 448 0 0 0 Tile_X0Y1_W2BEG[2]
port 493 nsew signal output
flabel metal3 s 0 3360 112 3472 0 FreeSans 448 0 0 0 Tile_X0Y1_W2BEG[3]
port 494 nsew signal output
flabel metal3 s 0 3808 112 3920 0 FreeSans 448 0 0 0 Tile_X0Y1_W2BEG[4]
port 495 nsew signal output
flabel metal3 s 0 4256 112 4368 0 FreeSans 448 0 0 0 Tile_X0Y1_W2BEG[5]
port 496 nsew signal output
flabel metal3 s 0 4704 112 4816 0 FreeSans 448 0 0 0 Tile_X0Y1_W2BEG[6]
port 497 nsew signal output
flabel metal3 s 0 5152 112 5264 0 FreeSans 448 0 0 0 Tile_X0Y1_W2BEG[7]
port 498 nsew signal output
flabel metal3 s 0 5600 112 5712 0 FreeSans 448 0 0 0 Tile_X0Y1_W2BEGb[0]
port 499 nsew signal output
flabel metal3 s 0 6048 112 6160 0 FreeSans 448 0 0 0 Tile_X0Y1_W2BEGb[1]
port 500 nsew signal output
flabel metal3 s 0 6496 112 6608 0 FreeSans 448 0 0 0 Tile_X0Y1_W2BEGb[2]
port 501 nsew signal output
flabel metal3 s 0 6944 112 7056 0 FreeSans 448 0 0 0 Tile_X0Y1_W2BEGb[3]
port 502 nsew signal output
flabel metal3 s 0 7392 112 7504 0 FreeSans 448 0 0 0 Tile_X0Y1_W2BEGb[4]
port 503 nsew signal output
flabel metal3 s 0 7840 112 7952 0 FreeSans 448 0 0 0 Tile_X0Y1_W2BEGb[5]
port 504 nsew signal output
flabel metal3 s 0 8288 112 8400 0 FreeSans 448 0 0 0 Tile_X0Y1_W2BEGb[6]
port 505 nsew signal output
flabel metal3 s 0 8736 112 8848 0 FreeSans 448 0 0 0 Tile_X0Y1_W2BEGb[7]
port 506 nsew signal output
flabel metal3 s 0 16352 112 16464 0 FreeSans 448 0 0 0 Tile_X0Y1_W6BEG[0]
port 507 nsew signal output
flabel metal3 s 0 20832 112 20944 0 FreeSans 448 0 0 0 Tile_X0Y1_W6BEG[10]
port 508 nsew signal output
flabel metal3 s 0 21280 112 21392 0 FreeSans 448 0 0 0 Tile_X0Y1_W6BEG[11]
port 509 nsew signal output
flabel metal3 s 0 16800 112 16912 0 FreeSans 448 0 0 0 Tile_X0Y1_W6BEG[1]
port 510 nsew signal output
flabel metal3 s 0 17248 112 17360 0 FreeSans 448 0 0 0 Tile_X0Y1_W6BEG[2]
port 511 nsew signal output
flabel metal3 s 0 17696 112 17808 0 FreeSans 448 0 0 0 Tile_X0Y1_W6BEG[3]
port 512 nsew signal output
flabel metal3 s 0 18144 112 18256 0 FreeSans 448 0 0 0 Tile_X0Y1_W6BEG[4]
port 513 nsew signal output
flabel metal3 s 0 18592 112 18704 0 FreeSans 448 0 0 0 Tile_X0Y1_W6BEG[5]
port 514 nsew signal output
flabel metal3 s 0 19040 112 19152 0 FreeSans 448 0 0 0 Tile_X0Y1_W6BEG[6]
port 515 nsew signal output
flabel metal3 s 0 19488 112 19600 0 FreeSans 448 0 0 0 Tile_X0Y1_W6BEG[7]
port 516 nsew signal output
flabel metal3 s 0 19936 112 20048 0 FreeSans 448 0 0 0 Tile_X0Y1_W6BEG[8]
port 517 nsew signal output
flabel metal3 s 0 20384 112 20496 0 FreeSans 448 0 0 0 Tile_X0Y1_W6BEG[9]
port 518 nsew signal output
flabel metal3 s 0 9184 112 9296 0 FreeSans 448 0 0 0 Tile_X0Y1_WW4BEG[0]
port 519 nsew signal output
flabel metal3 s 0 13664 112 13776 0 FreeSans 448 0 0 0 Tile_X0Y1_WW4BEG[10]
port 520 nsew signal output
flabel metal3 s 0 14112 112 14224 0 FreeSans 448 0 0 0 Tile_X0Y1_WW4BEG[11]
port 521 nsew signal output
flabel metal3 s 0 14560 112 14672 0 FreeSans 448 0 0 0 Tile_X0Y1_WW4BEG[12]
port 522 nsew signal output
flabel metal3 s 0 15008 112 15120 0 FreeSans 448 0 0 0 Tile_X0Y1_WW4BEG[13]
port 523 nsew signal output
flabel metal3 s 0 15456 112 15568 0 FreeSans 448 0 0 0 Tile_X0Y1_WW4BEG[14]
port 524 nsew signal output
flabel metal3 s 0 15904 112 16016 0 FreeSans 448 0 0 0 Tile_X0Y1_WW4BEG[15]
port 525 nsew signal output
flabel metal3 s 0 9632 112 9744 0 FreeSans 448 0 0 0 Tile_X0Y1_WW4BEG[1]
port 526 nsew signal output
flabel metal3 s 0 10080 112 10192 0 FreeSans 448 0 0 0 Tile_X0Y1_WW4BEG[2]
port 527 nsew signal output
flabel metal3 s 0 10528 112 10640 0 FreeSans 448 0 0 0 Tile_X0Y1_WW4BEG[3]
port 528 nsew signal output
flabel metal3 s 0 10976 112 11088 0 FreeSans 448 0 0 0 Tile_X0Y1_WW4BEG[4]
port 529 nsew signal output
flabel metal3 s 0 11424 112 11536 0 FreeSans 448 0 0 0 Tile_X0Y1_WW4BEG[5]
port 530 nsew signal output
flabel metal3 s 0 11872 112 11984 0 FreeSans 448 0 0 0 Tile_X0Y1_WW4BEG[6]
port 531 nsew signal output
flabel metal3 s 0 12320 112 12432 0 FreeSans 448 0 0 0 Tile_X0Y1_WW4BEG[7]
port 532 nsew signal output
flabel metal3 s 0 12768 112 12880 0 FreeSans 448 0 0 0 Tile_X0Y1_WW4BEG[8]
port 533 nsew signal output
flabel metal3 s 0 13216 112 13328 0 FreeSans 448 0 0 0 Tile_X0Y1_WW4BEG[9]
port 534 nsew signal output
flabel metal4 s 3776 0 4096 114912 0 FreeSans 1472 90 0 0 VDD
port 535 nsew power bidirectional
flabel metal4 s 3776 0 4096 56 0 FreeSans 368 0 0 0 VDD
port 535 nsew power bidirectional
flabel metal4 s 3776 114856 4096 114912 0 FreeSans 368 0 0 0 VDD
port 535 nsew power bidirectional
flabel metal4 s 23776 0 24096 114912 0 FreeSans 1472 90 0 0 VDD
port 535 nsew power bidirectional
flabel metal4 s 23776 0 24096 56 0 FreeSans 368 0 0 0 VDD
port 535 nsew power bidirectional
flabel metal4 s 23776 114856 24096 114912 0 FreeSans 368 0 0 0 VDD
port 535 nsew power bidirectional
flabel metal4 s 4436 0 4756 114912 0 FreeSans 1472 90 0 0 VSS
port 536 nsew ground bidirectional
flabel metal4 s 4436 0 4756 56 0 FreeSans 368 0 0 0 VSS
port 536 nsew ground bidirectional
flabel metal4 s 4436 114856 4756 114912 0 FreeSans 368 0 0 0 VSS
port 536 nsew ground bidirectional
flabel metal4 s 24436 0 24756 114912 0 FreeSans 1472 90 0 0 VSS
port 536 nsew ground bidirectional
flabel metal4 s 24436 0 24756 56 0 FreeSans 368 0 0 0 VSS
port 536 nsew ground bidirectional
flabel metal4 s 24436 114856 24756 114912 0 FreeSans 368 0 0 0 VSS
port 536 nsew ground bidirectional
flabel metal3 s 31584 12768 31696 12880 0 FreeSans 448 0 0 0 WEN_SRAM0
port 537 nsew signal output
flabel metal3 s 31584 13664 31696 13776 0 FreeSans 448 0 0 0 WEN_SRAM1
port 538 nsew signal output
flabel metal3 s 31584 14560 31696 14672 0 FreeSans 448 0 0 0 WEN_SRAM2
port 539 nsew signal output
flabel metal3 s 31584 15456 31696 15568 0 FreeSans 448 0 0 0 WEN_SRAM3
port 540 nsew signal output
flabel metal3 s 31584 16352 31696 16464 0 FreeSans 448 0 0 0 WEN_SRAM4
port 541 nsew signal output
flabel metal3 s 31584 17248 31696 17360 0 FreeSans 448 0 0 0 WEN_SRAM5
port 542 nsew signal output
flabel metal3 s 31584 18144 31696 18256 0 FreeSans 448 0 0 0 WEN_SRAM6
port 543 nsew signal output
flabel metal3 s 31584 19040 31696 19152 0 FreeSans 448 0 0 0 WEN_SRAM7
port 544 nsew signal output
rlabel metal1 15848 112896 15848 112896 0 VDD
rlabel metal1 15848 113680 15848 113680 0 VSS
rlabel metal3 31122 19992 31122 19992 0 A_SRAM0
rlabel metal3 31178 20888 31178 20888 0 A_SRAM1
rlabel metal3 31122 21784 31122 21784 0 A_SRAM2
rlabel metal3 31122 22680 31122 22680 0 A_SRAM3
rlabel metal3 31122 23576 31122 23576 0 A_SRAM4
rlabel metal3 31122 24472 31122 24472 0 A_SRAM5
rlabel metal3 31122 25368 31122 25368 0 A_SRAM6
rlabel metal3 31122 26264 31122 26264 0 A_SRAM7
rlabel metal3 31178 27160 31178 27160 0 A_SRAM8
rlabel metal3 31122 11032 31122 11032 0 CEN_SRAM
rlabel metal3 31122 35224 31122 35224 0 CLK_SRAM
rlabel metal3 30632 27720 30632 27720 0 CONFIGURED_top
rlabel metal3 31122 28056 31122 28056 0 D_SRAM0
rlabel metal3 31122 28952 31122 28952 0 D_SRAM1
rlabel metal3 31122 29848 31122 29848 0 D_SRAM2
rlabel metal3 31122 30744 31122 30744 0 D_SRAM3
rlabel metal3 31122 31640 31122 31640 0 D_SRAM4
rlabel metal3 31122 32536 31122 32536 0 D_SRAM5
rlabel metal3 31178 33432 31178 33432 0 D_SRAM6
rlabel metal3 31122 34328 31122 34328 0 D_SRAM7
rlabel metal3 31122 11928 31122 11928 0 GWEN_SRAM
rlabel metal4 28616 5264 28616 5264 0 Q_SRAM0
rlabel metal3 31640 4256 31640 4256 0 Q_SRAM1
rlabel metal3 29666 4760 29666 4760 0 Q_SRAM2
rlabel metal3 29512 5768 29512 5768 0 Q_SRAM3
rlabel metal3 29666 6552 29666 6552 0 Q_SRAM4
rlabel metal2 5432 77672 5432 77672 0 Q_SRAM5
rlabel metal3 31514 8344 31514 8344 0 Q_SRAM6
rlabel metal3 29946 9240 29946 9240 0 Q_SRAM7
rlabel metal2 15960 91280 15960 91280 0 Tile_X0Y0_E1END[0]
rlabel metal3 11032 93016 11032 93016 0 Tile_X0Y0_E1END[1]
rlabel metal2 1288 107632 1288 107632 0 Tile_X0Y0_E1END[2]
rlabel metal3 24416 62328 24416 62328 0 Tile_X0Y0_E1END[3]
rlabel metal2 15288 63336 15288 63336 0 Tile_X0Y0_E2END[0]
rlabel metal2 8232 74760 8232 74760 0 Tile_X0Y0_E2END[1]
rlabel metal3 1722 85512 1722 85512 0 Tile_X0Y0_E2END[2]
rlabel metal3 5096 86016 5096 86016 0 Tile_X0Y0_E2END[3]
rlabel metal2 20888 86520 20888 86520 0 Tile_X0Y0_E2END[4]
rlabel metal3 1078 86856 1078 86856 0 Tile_X0Y0_E2END[5]
rlabel metal3 126 87304 126 87304 0 Tile_X0Y0_E2END[6]
rlabel metal3 1722 87752 1722 87752 0 Tile_X0Y0_E2END[7]
rlabel metal2 16296 62496 16296 62496 0 Tile_X0Y0_E2MID[0]
rlabel metal2 8120 72800 8120 72800 0 Tile_X0Y0_E2MID[1]
rlabel metal3 9184 88984 9184 88984 0 Tile_X0Y0_E2MID[2]
rlabel metal3 910 82376 910 82376 0 Tile_X0Y0_E2MID[3]
rlabel metal2 21896 86408 21896 86408 0 Tile_X0Y0_E2MID[4]
rlabel metal3 238 83272 238 83272 0 Tile_X0Y0_E2MID[5]
rlabel metal3 182 83720 182 83720 0 Tile_X0Y0_E2MID[6]
rlabel metal2 6440 87696 6440 87696 0 Tile_X0Y0_E2MID[7]
rlabel metal2 18872 91728 18872 91728 0 Tile_X0Y0_E6END[0]
rlabel metal2 4760 100296 4760 100296 0 Tile_X0Y0_E6END[10]
rlabel metal2 22344 72744 22344 72744 0 Tile_X0Y0_E6END[11]
rlabel metal3 294 95816 294 95816 0 Tile_X0Y0_E6END[1]
rlabel metal2 1288 94976 1288 94976 0 Tile_X0Y0_E6END[2]
rlabel metal2 24024 69384 24024 69384 0 Tile_X0Y0_E6END[3]
rlabel metal2 15736 88200 15736 88200 0 Tile_X0Y0_E6END[4]
rlabel metal3 8400 97272 8400 97272 0 Tile_X0Y0_E6END[5]
rlabel metal2 1848 94640 1848 94640 0 Tile_X0Y0_E6END[6]
rlabel metal2 3080 89600 3080 89600 0 Tile_X0Y0_E6END[7]
rlabel metal4 3304 92568 3304 92568 0 Tile_X0Y0_E6END[8]
rlabel metal2 4368 99848 4368 99848 0 Tile_X0Y0_E6END[9]
rlabel metal2 18648 91840 18648 91840 0 Tile_X0Y0_EE4END[0]
rlabel metal2 1064 94080 1064 94080 0 Tile_X0Y0_EE4END[10]
rlabel metal2 19768 93072 19768 93072 0 Tile_X0Y0_EE4END[11]
rlabel metal2 16408 88984 16408 88984 0 Tile_X0Y0_EE4END[12]
rlabel metal3 1722 94024 1722 94024 0 Tile_X0Y0_EE4END[13]
rlabel metal2 1960 95480 1960 95480 0 Tile_X0Y0_EE4END[14]
rlabel metal2 20552 91728 20552 91728 0 Tile_X0Y0_EE4END[15]
rlabel metal3 1722 88648 1722 88648 0 Tile_X0Y0_EE4END[1]
rlabel metal2 4200 91000 4200 91000 0 Tile_X0Y0_EE4END[2]
rlabel metal3 910 89544 910 89544 0 Tile_X0Y0_EE4END[3]
rlabel metal4 17864 91840 17864 91840 0 Tile_X0Y0_EE4END[4]
rlabel metal2 10248 91280 10248 91280 0 Tile_X0Y0_EE4END[5]
rlabel metal2 3080 92008 3080 92008 0 Tile_X0Y0_EE4END[6]
rlabel metal2 21896 92568 21896 92568 0 Tile_X0Y0_EE4END[7]
rlabel metal2 15624 92904 15624 92904 0 Tile_X0Y0_EE4END[8]
rlabel metal3 1722 92232 1722 92232 0 Tile_X0Y0_EE4END[9]
rlabel metal3 2576 83608 2576 83608 0 Tile_X0Y0_FrameData[0]
rlabel metal2 2296 74816 2296 74816 0 Tile_X0Y0_FrameData[10]
rlabel metal2 3192 72772 3192 72772 0 Tile_X0Y0_FrameData[11]
rlabel metal3 2408 109256 2408 109256 0 Tile_X0Y0_FrameData[12]
rlabel metal2 15568 61320 15568 61320 0 Tile_X0Y0_FrameData[13]
rlabel metal2 18424 62776 18424 62776 0 Tile_X0Y0_FrameData[14]
rlabel metal2 21896 60032 21896 60032 0 Tile_X0Y0_FrameData[15]
rlabel metal2 29512 96432 29512 96432 0 Tile_X0Y0_FrameData[16]
rlabel metal2 29512 97216 29512 97216 0 Tile_X0Y0_FrameData[17]
rlabel metal3 1904 87192 1904 87192 0 Tile_X0Y0_FrameData[18]
rlabel metal3 518 109256 518 109256 0 Tile_X0Y0_FrameData[19]
rlabel metal2 29512 79128 29512 79128 0 Tile_X0Y0_FrameData[1]
rlabel metal3 966 109704 966 109704 0 Tile_X0Y0_FrameData[20]
rlabel metal2 15960 68544 15960 68544 0 Tile_X0Y0_FrameData[21]
rlabel metal3 3192 110432 3192 110432 0 Tile_X0Y0_FrameData[22]
rlabel metal3 18424 69496 18424 69496 0 Tile_X0Y0_FrameData[23]
rlabel metal2 1624 109424 1624 109424 0 Tile_X0Y0_FrameData[24]
rlabel metal2 1624 110880 1624 110880 0 Tile_X0Y0_FrameData[25]
rlabel metal2 1680 110152 1680 110152 0 Tile_X0Y0_FrameData[26]
rlabel metal2 29624 107296 29624 107296 0 Tile_X0Y0_FrameData[27]
rlabel metal2 3192 111888 3192 111888 0 Tile_X0Y0_FrameData[28]
rlabel metal3 1232 111832 1232 111832 0 Tile_X0Y0_FrameData[29]
rlabel metal2 29512 80024 29512 80024 0 Tile_X0Y0_FrameData[2]
rlabel metal3 126 114184 126 114184 0 Tile_X0Y0_FrameData[30]
rlabel metal2 18760 65184 18760 65184 0 Tile_X0Y0_FrameData[31]
rlabel metal2 1736 69776 1736 69776 0 Tile_X0Y0_FrameData[3]
rlabel metal3 910 102536 910 102536 0 Tile_X0Y0_FrameData[4]
rlabel metal2 22792 81256 22792 81256 0 Tile_X0Y0_FrameData[5]
rlabel metal3 18480 60648 18480 60648 0 Tile_X0Y0_FrameData[6]
rlabel metal3 20160 58520 20160 58520 0 Tile_X0Y0_FrameData[7]
rlabel metal3 2464 63784 2464 63784 0 Tile_X0Y0_FrameData[8]
rlabel metal2 2408 60032 2408 60032 0 Tile_X0Y0_FrameData[9]
rlabel metal3 31122 78232 31122 78232 0 Tile_X0Y0_FrameData_O[0]
rlabel metal3 31122 89432 31122 89432 0 Tile_X0Y0_FrameData_O[10]
rlabel metal3 31122 90552 31122 90552 0 Tile_X0Y0_FrameData_O[11]
rlabel metal3 31122 91672 31122 91672 0 Tile_X0Y0_FrameData_O[12]
rlabel metal3 31122 92792 31122 92792 0 Tile_X0Y0_FrameData_O[13]
rlabel metal3 31122 93912 31122 93912 0 Tile_X0Y0_FrameData_O[14]
rlabel metal3 31122 95032 31122 95032 0 Tile_X0Y0_FrameData_O[15]
rlabel metal3 31122 96152 31122 96152 0 Tile_X0Y0_FrameData_O[16]
rlabel metal3 31122 97272 31122 97272 0 Tile_X0Y0_FrameData_O[17]
rlabel metal3 31122 98392 31122 98392 0 Tile_X0Y0_FrameData_O[18]
rlabel metal3 31122 99512 31122 99512 0 Tile_X0Y0_FrameData_O[19]
rlabel metal3 31122 79352 31122 79352 0 Tile_X0Y0_FrameData_O[1]
rlabel metal3 31122 100632 31122 100632 0 Tile_X0Y0_FrameData_O[20]
rlabel metal3 31122 101752 31122 101752 0 Tile_X0Y0_FrameData_O[21]
rlabel metal3 31122 102872 31122 102872 0 Tile_X0Y0_FrameData_O[22]
rlabel metal3 31122 103992 31122 103992 0 Tile_X0Y0_FrameData_O[23]
rlabel metal3 31122 105112 31122 105112 0 Tile_X0Y0_FrameData_O[24]
rlabel metal3 31122 106232 31122 106232 0 Tile_X0Y0_FrameData_O[25]
rlabel metal3 31122 107352 31122 107352 0 Tile_X0Y0_FrameData_O[26]
rlabel metal3 31122 108472 31122 108472 0 Tile_X0Y0_FrameData_O[27]
rlabel metal3 31122 109592 31122 109592 0 Tile_X0Y0_FrameData_O[28]
rlabel metal3 31122 110712 31122 110712 0 Tile_X0Y0_FrameData_O[29]
rlabel metal3 31122 80472 31122 80472 0 Tile_X0Y0_FrameData_O[2]
rlabel metal3 31122 111832 31122 111832 0 Tile_X0Y0_FrameData_O[30]
rlabel metal2 29960 112448 29960 112448 0 Tile_X0Y0_FrameData_O[31]
rlabel metal3 31122 81592 31122 81592 0 Tile_X0Y0_FrameData_O[3]
rlabel metal3 31122 82712 31122 82712 0 Tile_X0Y0_FrameData_O[4]
rlabel metal3 31122 83832 31122 83832 0 Tile_X0Y0_FrameData_O[5]
rlabel metal3 31122 84952 31122 84952 0 Tile_X0Y0_FrameData_O[6]
rlabel metal3 31122 86072 31122 86072 0 Tile_X0Y0_FrameData_O[7]
rlabel metal3 31122 87192 31122 87192 0 Tile_X0Y0_FrameData_O[8]
rlabel metal3 31122 88312 31122 88312 0 Tile_X0Y0_FrameData_O[9]
rlabel metal2 24696 112896 24696 112896 0 Tile_X0Y0_FrameStrobe_O[0]
rlabel metal2 28504 113568 28504 113568 0 Tile_X0Y0_FrameStrobe_O[10]
rlabel metal2 29064 113848 29064 113848 0 Tile_X0Y0_FrameStrobe_O[11]
rlabel metal2 27720 113736 27720 113736 0 Tile_X0Y0_FrameStrobe_O[12]
rlabel metal2 29176 113512 29176 113512 0 Tile_X0Y0_FrameStrobe_O[13]
rlabel metal2 28952 112224 28952 112224 0 Tile_X0Y0_FrameStrobe_O[14]
rlabel metal2 27608 112504 27608 112504 0 Tile_X0Y0_FrameStrobe_O[15]
rlabel metal2 28280 112280 28280 112280 0 Tile_X0Y0_FrameStrobe_O[16]
rlabel metal2 29848 112560 29848 112560 0 Tile_X0Y0_FrameStrobe_O[17]
rlabel metal4 27384 112000 27384 112000 0 Tile_X0Y0_FrameStrobe_O[18]
rlabel metal2 26040 114170 26040 114170 0 Tile_X0Y0_FrameStrobe_O[19]
rlabel metal2 23352 112672 23352 112672 0 Tile_X0Y0_FrameStrobe_O[1]
rlabel metal2 24024 112560 24024 112560 0 Tile_X0Y0_FrameStrobe_O[2]
rlabel metal2 25480 113792 25480 113792 0 Tile_X0Y0_FrameStrobe_O[3]
rlabel metal2 25648 112392 25648 112392 0 Tile_X0Y0_FrameStrobe_O[4]
rlabel metal2 26152 114016 26152 114016 0 Tile_X0Y0_FrameStrobe_O[5]
rlabel metal2 26488 112672 26488 112672 0 Tile_X0Y0_FrameStrobe_O[6]
rlabel metal2 26824 113960 26824 113960 0 Tile_X0Y0_FrameStrobe_O[7]
rlabel metal2 27160 112784 27160 112784 0 Tile_X0Y0_FrameStrobe_O[8]
rlabel metal2 28392 113904 28392 113904 0 Tile_X0Y0_FrameStrobe_O[9]
rlabel metal2 16968 76384 16968 76384 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit0.Q
rlabel metal2 18200 76720 18200 76720 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit1.Q
rlabel metal3 9184 107688 9184 107688 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit10.Q
rlabel metal4 9352 110432 9352 110432 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit11.Q
rlabel metal2 15288 109228 15288 109228 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit12.Q
rlabel metal2 16128 105672 16128 105672 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit13.Q
rlabel metal2 19544 104160 19544 104160 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit14.Q
rlabel metal2 18536 103600 18536 103600 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit15.Q
rlabel metal2 14728 85064 14728 85064 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit16.Q
rlabel metal3 12880 85064 12880 85064 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit17.Q
rlabel metal2 12488 109256 12488 109256 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit18.Q
rlabel metal2 10920 113064 10920 113064 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit19.Q
rlabel metal2 12488 101976 12488 101976 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit2.Q
rlabel metal2 14616 110544 14616 110544 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit20.Q
rlabel metal2 13440 110152 13440 110152 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit21.Q
rlabel metal2 17192 110040 17192 110040 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit22.Q
rlabel metal2 16016 109368 16016 109368 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit23.Q
rlabel metal2 19432 97412 19432 97412 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit24.Q
rlabel metal2 18984 98672 18984 98672 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit25.Q
rlabel metal2 12152 103432 12152 103432 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit26.Q
rlabel metal2 12040 104216 12040 104216 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit27.Q
rlabel metal2 7896 99064 7896 99064 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit28.Q
rlabel metal2 7672 96376 7672 96376 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit29.Q
rlabel metal2 15288 102592 15288 102592 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit3.Q
rlabel metal2 23128 67928 23128 67928 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit30.Q
rlabel metal2 22680 67256 22680 67256 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit31.Q
rlabel metal3 6888 107576 6888 107576 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit4.Q
rlabel metal2 7560 105336 7560 105336 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit5.Q
rlabel metal3 20160 60760 20160 60760 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit6.Q
rlabel metal2 20664 58968 20664 58968 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit7.Q
rlabel metal2 12320 63112 12320 63112 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit8.Q
rlabel metal2 11200 60200 11200 60200 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame0_bit9.Q
rlabel metal3 9744 72408 9744 72408 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit0.Q
rlabel metal3 10136 73864 10136 73864 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit1.Q
rlabel metal3 11424 86632 11424 86632 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit10.Q
rlabel metal2 12936 87360 12936 87360 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit11.Q
rlabel metal2 6552 110096 6552 110096 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit12.Q
rlabel metal2 7672 110600 7672 110600 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit13.Q
rlabel metal2 19600 62552 19600 62552 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit14.Q
rlabel metal2 20720 60200 20720 60200 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit15.Q
rlabel metal3 16576 83496 16576 83496 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit16.Q
rlabel metal2 18424 84168 18424 84168 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit17.Q
rlabel metal2 12936 100856 12936 100856 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit18.Q
rlabel metal2 15512 101136 15512 101136 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit19.Q
rlabel metal3 11480 78904 11480 78904 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit2.Q
rlabel metal2 4144 109592 4144 109592 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit20.Q
rlabel metal2 6272 110264 6272 110264 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit21.Q
rlabel metal3 20104 67816 20104 67816 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit22.Q
rlabel metal2 21896 67984 21896 67984 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit23.Q
rlabel metal2 15960 79296 15960 79296 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit24.Q
rlabel metal2 17304 80248 17304 80248 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit25.Q
rlabel metal2 13160 105224 13160 105224 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit26.Q
rlabel metal2 14560 104664 14560 104664 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit27.Q
rlabel metal2 6440 111048 6440 111048 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit28.Q
rlabel metal2 2856 111216 2856 111216 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit29.Q
rlabel metal3 10864 78120 10864 78120 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit3.Q
rlabel metal3 18200 66248 18200 66248 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit30.Q
rlabel metal2 19880 65968 19880 65968 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit31.Q
rlabel metal3 14168 81144 14168 81144 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit4.Q
rlabel metal2 14000 80584 14000 80584 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit5.Q
rlabel metal2 22792 87696 22792 87696 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit6.Q
rlabel metal2 23016 87304 23016 87304 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit7.Q
rlabel metal2 16072 78008 16072 78008 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit8.Q
rlabel metal3 17920 78792 17920 78792 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame1_bit9.Q
rlabel metal2 3864 77616 3864 77616 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit0.Q
rlabel metal2 2856 86044 2856 86044 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit1.Q
rlabel metal2 9408 92904 9408 92904 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit10.Q
rlabel metal2 9744 94584 9744 94584 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit11.Q
rlabel metal2 1512 93632 1512 93632 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit12.Q
rlabel metal2 2520 93240 2520 93240 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit13.Q
rlabel metal3 1064 90664 1064 90664 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit14.Q
rlabel metal3 21168 94472 21168 94472 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit15.Q
rlabel metal2 21336 95536 21336 95536 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit16.Q
rlabel metal2 24920 93968 24920 93968 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit17.Q
rlabel metal3 16744 91336 16744 91336 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit18.Q
rlabel metal3 16128 93688 16128 93688 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit19.Q
rlabel metal2 11592 77504 11592 77504 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit2.Q
rlabel metal2 19432 91224 19432 91224 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit20.Q
rlabel metal2 8568 95032 8568 95032 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit21.Q
rlabel metal2 9016 94472 9016 94472 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit22.Q
rlabel metal2 8232 93800 8232 93800 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit23.Q
rlabel metal3 2184 95256 2184 95256 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit24.Q
rlabel metal2 2688 110712 2688 110712 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit25.Q
rlabel metal3 7448 89880 7448 89880 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit26.Q
rlabel metal3 20776 94248 20776 94248 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit27.Q
rlabel metal2 21168 95256 21168 95256 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit28.Q
rlabel metal2 22120 90776 22120 90776 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit29.Q
rlabel metal2 10360 77840 10360 77840 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit3.Q
rlabel metal3 16352 61544 16352 61544 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit30.Q
rlabel metal2 17192 61152 17192 61152 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit31.Q
rlabel metal2 14616 77112 14616 77112 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit4.Q
rlabel metal3 12712 76440 12712 76440 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit5.Q
rlabel metal2 15960 92064 15960 92064 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit6.Q
rlabel metal3 16576 92120 16576 92120 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit7.Q
rlabel metal2 17528 89264 17528 89264 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit8.Q
rlabel metal2 10472 93408 10472 93408 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame2_bit9.Q
rlabel metal2 3528 74424 3528 74424 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit0.Q
rlabel metal2 2464 75992 2464 75992 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit1.Q
rlabel metal2 8120 77504 8120 77504 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit10.Q
rlabel metal2 7168 76440 7168 76440 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit11.Q
rlabel metal2 13104 73864 13104 73864 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit12.Q
rlabel metal3 13552 72744 13552 72744 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit13.Q
rlabel metal2 16072 74592 16072 74592 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit14.Q
rlabel metal2 18424 75264 18424 75264 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit15.Q
rlabel metal2 7896 85736 7896 85736 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit16.Q
rlabel metal3 8232 84280 8232 84280 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit17.Q
rlabel metal3 6496 103096 6496 103096 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit18.Q
rlabel metal2 7896 109564 7896 109564 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit19.Q
rlabel metal2 6664 71624 6664 71624 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit2.Q
rlabel metal2 15736 68880 15736 68880 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit20.Q
rlabel metal2 16856 69272 16856 69272 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit21.Q
rlabel metal3 18256 73528 18256 73528 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit22.Q
rlabel metal3 19656 71960 19656 71960 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit23.Q
rlabel metal2 3304 75768 3304 75768 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit24.Q
rlabel metal2 4760 74088 4760 74088 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit25.Q
rlabel metal2 5544 82600 5544 82600 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit26.Q
rlabel metal3 6888 80472 6888 80472 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit27.Q
rlabel metal3 12656 74872 12656 74872 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit28.Q
rlabel metal2 14224 74872 14224 74872 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit29.Q
rlabel metal2 5600 70392 5600 70392 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit3.Q
rlabel metal3 22736 74312 22736 74312 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit30.Q
rlabel metal2 21112 75936 21112 75936 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit31.Q
rlabel metal2 15064 72016 15064 72016 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit4.Q
rlabel metal2 16072 71400 16072 71400 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit5.Q
rlabel metal3 20496 72520 20496 72520 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit6.Q
rlabel metal2 22568 71960 22568 71960 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit7.Q
rlabel metal2 3080 79800 3080 79800 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit8.Q
rlabel metal2 2632 76160 2632 76160 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame3_bit9.Q
rlabel metal2 3416 71288 3416 71288 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit0.Q
rlabel metal2 2800 72744 2800 72744 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit1.Q
rlabel metal2 3304 72408 3304 72408 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit10.Q
rlabel metal3 1512 72408 1512 72408 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit11.Q
rlabel metal3 5040 61544 5040 61544 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit12.Q
rlabel metal3 7000 62888 7000 62888 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit13.Q
rlabel metal2 18648 62216 18648 62216 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit14.Q
rlabel metal2 19824 63672 19824 63672 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit15.Q
rlabel metal2 9016 83608 9016 83608 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit16.Q
rlabel metal2 2744 97384 2744 97384 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit17.Q
rlabel metal2 6552 84616 6552 84616 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit18.Q
rlabel metal2 4144 86520 4144 86520 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit19.Q
rlabel metal2 3640 65296 3640 65296 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit2.Q
rlabel metal2 14616 66360 14616 66360 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit20.Q
rlabel metal2 15848 66752 15848 66752 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit21.Q
rlabel metal2 17360 65464 17360 65464 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit22.Q
rlabel metal2 18480 67816 18480 67816 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit23.Q
rlabel metal3 4928 67816 4928 67816 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit24.Q
rlabel metal2 6664 68488 6664 68488 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit25.Q
rlabel metal2 5376 85624 5376 85624 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit26.Q
rlabel metal2 3528 87080 3528 87080 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit27.Q
rlabel metal2 12488 68096 12488 68096 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit28.Q
rlabel metal2 13608 68152 13608 68152 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit29.Q
rlabel metal2 2352 64680 2352 64680 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit3.Q
rlabel metal2 21112 68768 21112 68768 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit30.Q
rlabel metal2 22344 69664 22344 69664 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit31.Q
rlabel metal2 9128 69608 9128 69608 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit4.Q
rlabel metal2 10472 70448 10472 70448 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit5.Q
rlabel metal3 8792 64680 8792 64680 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit6.Q
rlabel metal2 10472 64400 10472 64400 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit7.Q
rlabel metal2 2856 63112 2856 63112 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit8.Q
rlabel metal2 1232 60200 1232 60200 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame4_bit9.Q
rlabel metal2 5656 98392 5656 98392 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit0.Q
rlabel metal2 3752 109928 3752 109928 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit1.Q
rlabel metal2 7672 73192 7672 73192 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit10.Q
rlabel metal3 5376 71736 5376 71736 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit11.Q
rlabel metal2 18536 59696 18536 59696 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit12.Q
rlabel metal2 17304 60256 17304 60256 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit13.Q
rlabel metal3 5600 60200 5600 60200 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit14.Q
rlabel metal2 7392 60200 7392 60200 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit15.Q
rlabel metal2 3248 86856 3248 86856 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit16.Q
rlabel metal2 1512 84840 1512 84840 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit17.Q
rlabel metal2 3024 88424 3024 88424 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit18.Q
rlabel metal3 1512 86520 1512 86520 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit19.Q
rlabel metal2 5320 94640 5320 94640 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit2.Q
rlabel metal2 9632 66248 9632 66248 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit20.Q
rlabel metal2 11032 66528 11032 66528 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit21.Q
rlabel metal3 8960 65464 8960 65464 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit22.Q
rlabel metal2 10696 66360 10696 66360 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit23.Q
rlabel metal2 3416 64232 3416 64232 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit24.Q
rlabel metal2 2464 63112 2464 63112 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit25.Q
rlabel metal2 2912 87976 2912 87976 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit26.Q
rlabel metal3 896 90328 896 90328 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit27.Q
rlabel metal2 5432 66528 5432 66528 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit28.Q
rlabel metal2 6664 66752 6664 66752 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit29.Q
rlabel metal3 22400 79576 22400 79576 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit3.Q
rlabel metal3 5096 62328 5096 62328 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit30.Q
rlabel metal2 7336 63784 7336 63784 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit31.Q
rlabel metal3 20496 79576 20496 79576 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit4.Q
rlabel metal2 21224 77448 21224 77448 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit5.Q
rlabel metal2 16296 58296 16296 58296 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit6.Q
rlabel metal2 15064 57904 15064 57904 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit7.Q
rlabel metal3 12096 61544 12096 61544 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit8.Q
rlabel metal3 11200 62888 11200 62888 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame5_bit9.Q
rlabel metal2 19936 86408 19936 86408 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit0.Q
rlabel metal3 20104 85736 20104 85736 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit1.Q
rlabel metal2 3528 94696 3528 94696 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit10.Q
rlabel metal2 4872 90328 4872 90328 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit11.Q
rlabel metal3 17920 110936 17920 110936 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit12.Q
rlabel metal2 2968 100072 2968 100072 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit13.Q
rlabel metal2 4312 106344 4312 106344 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit14.Q
rlabel metal2 2968 106344 2968 106344 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit15.Q
rlabel metal2 19320 87304 19320 87304 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit16.Q
rlabel metal2 20552 86912 20552 86912 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit17.Q
rlabel metal3 13216 82040 13216 82040 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit18.Q
rlabel metal2 12376 82208 12376 82208 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit19.Q
rlabel metal2 16072 97104 16072 97104 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit2.Q
rlabel metal3 8344 79576 8344 79576 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit20.Q
rlabel metal2 10080 79576 10080 79576 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit21.Q
rlabel metal3 8792 73304 8792 73304 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit22.Q
rlabel metal3 8400 75656 8400 75656 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit23.Q
rlabel metal2 14616 63392 14616 63392 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit24.Q
rlabel metal2 15848 63000 15848 63000 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit25.Q
rlabel metal2 15512 86632 15512 86632 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit26.Q
rlabel metal3 16016 85736 16016 85736 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit27.Q
rlabel metal2 17808 82936 17808 82936 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit28.Q
rlabel metal2 12152 96656 12152 96656 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit29.Q
rlabel metal2 15064 97160 15064 97160 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit3.Q
rlabel metal2 10920 96432 10920 96432 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit30.Q
rlabel metal2 12992 95480 12992 95480 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit31.Q
rlabel metal3 9072 100744 9072 100744 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit4.Q
rlabel metal2 11256 102200 11256 102200 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit5.Q
rlabel metal2 16968 101976 16968 101976 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit6.Q
rlabel metal2 5320 101024 5320 101024 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit7.Q
rlabel metal2 21168 62328 21168 62328 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit8.Q
rlabel metal2 22344 63000 22344 63000 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame6_bit9.Q
rlabel metal2 9016 101976 9016 101976 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit0.Q
rlabel metal3 8120 101416 8120 101416 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit1.Q
rlabel metal3 10808 107016 10808 107016 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit10.Q
rlabel metal3 8848 112280 8848 112280 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit11.Q
rlabel metal2 8400 85848 8400 85848 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit12.Q
rlabel metal2 9464 85904 9464 85904 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit13.Q
rlabel metal3 8120 83496 8120 83496 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit14.Q
rlabel metal3 10136 83496 10136 83496 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit15.Q
rlabel metal2 6216 89152 6216 89152 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit16.Q
rlabel metal2 7336 91224 7336 91224 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit17.Q
rlabel metal2 6776 92344 6776 92344 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit18.Q
rlabel metal2 7560 92120 7560 92120 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit19.Q
rlabel metal4 17416 106736 17416 106736 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit2.Q
rlabel metal2 11816 88480 11816 88480 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit20.Q
rlabel metal2 10808 88088 10808 88088 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit21.Q
rlabel metal2 14392 89992 14392 89992 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit22.Q
rlabel via2 13272 91336 13272 91336 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit23.Q
rlabel metal3 10472 91560 10472 91560 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit24.Q
rlabel metal2 11480 99568 11480 99568 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit25.Q
rlabel metal3 8736 99960 8736 99960 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit26.Q
rlabel metal2 10248 102984 10248 102984 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit27.Q
rlabel metal2 2968 108192 2968 108192 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit28.Q
rlabel metal3 8400 114520 8400 114520 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit29.Q
rlabel metal2 17416 105280 17416 105280 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit3.Q
rlabel metal2 15176 112896 15176 112896 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit30.Q
rlabel metal3 21616 84280 21616 84280 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit31.Q
rlabel metal2 20944 80360 20944 80360 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit4.Q
rlabel metal2 21840 80472 21840 80472 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit5.Q
rlabel metal3 3304 99176 3304 99176 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit6.Q
rlabel metal2 4536 89936 4536 89936 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit7.Q
rlabel metal3 20776 111048 20776 111048 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit8.Q
rlabel metal2 19152 111496 19152 111496 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame7_bit9.Q
rlabel metal2 16856 98112 16856 98112 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame8_bit30.Q
rlabel metal2 15624 98672 15624 98672 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_ConfigMem.Inst_frame8_bit31.Q
rlabel metal2 18424 74144 18424 74144 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG0
rlabel metal2 3808 69384 3808 69384 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG1
rlabel metal2 2296 77896 2296 77896 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG2
rlabel metal2 17640 67648 17640 67648 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG3
rlabel metal2 15512 69384 15512 69384 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG4
rlabel metal2 2856 71680 2856 71680 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG5
rlabel metal3 2632 70952 2632 70952 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG6
rlabel metal2 21392 68600 21392 68600 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS2_BEG7
rlabel metal2 17752 90832 17752 90832 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG0
rlabel metal2 11032 98280 11032 98280 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG1
rlabel metal2 16072 67984 16072 67984 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG12
rlabel metal2 13048 92568 13048 92568 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG13
rlabel metal2 2296 108136 2296 108136 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG14
rlabel metal3 21168 61992 21168 61992 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG15
rlabel metal2 2184 92848 2184 92848 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG2
rlabel metal2 20552 69216 20552 69216 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG3
rlabel metal2 17528 90776 17528 90776 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG4
rlabel metal3 9240 92904 9240 92904 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG5
rlabel metal2 2744 94808 2744 94808 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG6
rlabel metal2 20664 69384 20664 69384 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.J_NS4_BEG7
rlabel metal2 12208 110936 12208 110936 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1BEG0
rlabel metal2 9688 101976 9688 101976 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1BEG1
rlabel metal2 1176 103880 1176 103880 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1BEG2
rlabel metal3 20888 80584 20888 80584 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1BEG3
rlabel metal2 17752 58968 17752 58968 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END0
rlabel metal2 16296 93408 16296 93408 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END1
rlabel metal2 10192 47656 10192 47656 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END2
rlabel metal2 20216 59752 20216 59752 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N1END3
rlabel metal3 1960 95816 1960 95816 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG0
rlabel metal2 3304 101920 3304 101920 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG1
rlabel metal2 3304 104440 3304 104440 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG2
rlabel metal3 7448 88760 7448 88760 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG3
rlabel metal4 1848 99064 1848 99064 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG4
rlabel metal3 5880 88872 5880 88872 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG5
rlabel metal2 7112 90608 7112 90608 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG6
rlabel metal2 11256 87360 11256 87360 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEG7
rlabel metal3 7840 63784 7840 63784 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb0
rlabel metal3 11144 44520 11144 44520 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb1
rlabel metal2 17752 108080 17752 108080 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb2
rlabel metal2 16856 103992 16856 103992 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb3
rlabel metal3 16184 43960 16184 43960 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb4
rlabel metal3 4480 110712 4480 110712 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb5
rlabel metal2 15960 110096 15960 110096 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb6
rlabel metal2 17192 40376 17192 40376 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N2BEGb7
rlabel metal2 13888 107016 13888 107016 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N4BEG0
rlabel metal2 8904 109676 8904 109676 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N4BEG1
rlabel metal3 10248 109984 10248 109984 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N4BEG2
rlabel metal2 20048 86072 20048 86072 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.N4BEG3
rlabel metal2 10920 3080 10920 3080 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG0
rlabel metal3 1960 58744 1960 58744 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG1
rlabel metal3 1680 58184 1680 58184 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG2
rlabel metal2 18760 44688 18760 44688 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG3
rlabel metal3 14448 1960 14448 1960 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG4
rlabel metal2 448 55440 448 55440 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG5
rlabel metal3 15680 2744 15680 2744 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG6
rlabel metal2 16240 55440 16240 55440 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S2BEG7
rlabel metal2 18312 82992 18312 82992 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S4BEG0
rlabel metal2 16856 95256 16856 95256 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S4BEG1
rlabel metal2 18536 94416 18536 94416 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S4BEG2
rlabel metal3 20328 77224 20328 77224 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.S4BEG3
rlabel metal3 14952 57400 14952 57400 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W1BEG0
rlabel metal2 12600 60928 12600 60928 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W1BEG1
rlabel metal2 2240 59192 2240 59192 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W1BEG2
rlabel metal2 17976 59360 17976 59360 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W1BEG3
rlabel metal3 4424 60648 4424 60648 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG0
rlabel metal3 2128 61768 2128 61768 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG1
rlabel metal2 1456 68600 1456 68600 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG2
rlabel metal2 9576 63112 9576 63112 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG3
rlabel metal2 10024 65128 10024 65128 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG4
rlabel metal3 2184 63336 2184 63336 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG5
rlabel metal4 3640 78711 3640 78711 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG6
rlabel metal2 2184 67704 2184 67704 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEG7
rlabel metal3 5992 62216 5992 62216 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb0
rlabel metal2 3304 67984 3304 67984 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb1
rlabel metal2 3080 65744 3080 65744 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb2
rlabel metal2 9800 69272 9800 69272 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb3
rlabel metal3 9184 64792 9184 64792 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb4
rlabel metal2 2184 64232 2184 64232 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb5
rlabel metal2 2520 70840 2520 70840 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb6
rlabel metal3 896 66808 896 66808 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W2BEGb7
rlabel metal3 17416 74648 17416 74648 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG0
rlabel metal2 8344 76216 8344 76216 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG1
rlabel metal2 10920 77280 10920 77280 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG10
rlabel metal2 13888 76328 13888 76328 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG11
rlabel metal2 7336 103432 7336 103432 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG2
rlabel metal2 14840 69216 14840 69216 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG3
rlabel metal3 18200 74088 18200 74088 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG4
rlabel metal2 3976 74368 3976 74368 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG5
rlabel metal2 1064 81872 1064 81872 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG6
rlabel metal3 12936 74760 12936 74760 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG7
rlabel metal3 21112 75768 21112 75768 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG8
rlabel metal2 3416 77280 3416 77280 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.W6BEG9
rlabel metal3 18480 63672 18480 63672 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG0
rlabel metal3 2912 85176 2912 85176 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG1
rlabel metal2 6160 71176 6160 71176 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG10
rlabel metal3 14952 71512 14952 71512 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG11
rlabel metal2 21560 72912 21560 72912 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG12
rlabel metal2 3192 76160 3192 76160 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG13
rlabel metal3 6384 76328 6384 76328 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG14
rlabel metal3 13048 73080 13048 73080 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG15
rlabel metal2 1960 74928 1960 74928 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG2
rlabel metal3 14504 66808 14504 66808 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG3
rlabel metal3 17024 67928 17024 67928 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG4
rlabel metal2 5992 68432 5992 68432 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG5
rlabel metal3 4592 75432 4592 75432 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG6
rlabel metal2 13160 68712 13160 68712 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG7
rlabel metal2 21672 69216 21672 69216 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG8
rlabel metal2 5320 72912 5320 72912 0 Tile_X0Y0_GF_SRAM_top.Inst_GF_SRAM_top_switch_matrix.WW4BEG9
rlabel metal3 7560 41944 7560 41944 0 Tile_X0Y0_GF_SRAM_top.N4BEG_outbuf_10.A
rlabel metal3 16968 46088 16968 46088 0 Tile_X0Y0_GF_SRAM_top.N4BEG_outbuf_11.A
rlabel metal3 16072 31192 16072 31192 0 Tile_X0Y0_GF_SRAM_top.N4BEG_outbuf_8.A
rlabel metal2 5432 68040 5432 68040 0 Tile_X0Y0_GF_SRAM_top.N4BEG_outbuf_9.A
rlabel metal2 19656 109648 19656 109648 0 Tile_X0Y0_N1BEG[0]
rlabel metal2 5656 113442 5656 113442 0 Tile_X0Y0_N1BEG[1]
rlabel metal2 22680 112224 22680 112224 0 Tile_X0Y0_N1BEG[2]
rlabel metal2 6104 114058 6104 114058 0 Tile_X0Y0_N1BEG[3]
rlabel metal2 1736 110432 1736 110432 0 Tile_X0Y0_N2BEG[0]
rlabel metal2 6552 113442 6552 113442 0 Tile_X0Y0_N2BEG[1]
rlabel metal2 6776 114282 6776 114282 0 Tile_X0Y0_N2BEG[2]
rlabel metal2 1512 112784 1512 112784 0 Tile_X0Y0_N2BEG[3]
rlabel metal2 7224 113722 7224 113722 0 Tile_X0Y0_N2BEG[4]
rlabel metal2 7448 113890 7448 113890 0 Tile_X0Y0_N2BEG[5]
rlabel metal2 7672 113666 7672 113666 0 Tile_X0Y0_N2BEG[6]
rlabel metal2 7896 113162 7896 113162 0 Tile_X0Y0_N2BEG[7]
rlabel metal2 8120 114170 8120 114170 0 Tile_X0Y0_N2BEGb[0]
rlabel metal2 5376 107688 5376 107688 0 Tile_X0Y0_N2BEGb[1]
rlabel metal3 19544 112448 19544 112448 0 Tile_X0Y0_N2BEGb[2]
rlabel metal2 8792 113218 8792 113218 0 Tile_X0Y0_N2BEGb[3]
rlabel metal2 19544 112616 19544 112616 0 Tile_X0Y0_N2BEGb[4]
rlabel metal2 22008 112560 22008 112560 0 Tile_X0Y0_N2BEGb[5]
rlabel metal2 9464 113442 9464 113442 0 Tile_X0Y0_N2BEGb[6]
rlabel metal2 18536 113736 18536 113736 0 Tile_X0Y0_N2BEGb[7]
rlabel metal2 23016 114072 23016 114072 0 Tile_X0Y0_N4BEG[0]
rlabel metal2 15400 113848 15400 113848 0 Tile_X0Y0_N4BEG[10]
rlabel metal2 22344 113680 22344 113680 0 Tile_X0Y0_N4BEG[11]
rlabel metal2 19208 113568 19208 113568 0 Tile_X0Y0_N4BEG[12]
rlabel metal2 21336 112616 21336 112616 0 Tile_X0Y0_N4BEG[13]
rlabel metal3 13888 113512 13888 113512 0 Tile_X0Y0_N4BEG[14]
rlabel metal2 12264 112728 12264 112728 0 Tile_X0Y0_N4BEG[15]
rlabel metal2 10136 113722 10136 113722 0 Tile_X0Y0_N4BEG[1]
rlabel metal2 5208 113568 5208 113568 0 Tile_X0Y0_N4BEG[2]
rlabel metal2 9240 112448 9240 112448 0 Tile_X0Y0_N4BEG[3]
rlabel metal2 10808 114114 10808 114114 0 Tile_X0Y0_N4BEG[4]
rlabel metal2 11032 114058 11032 114058 0 Tile_X0Y0_N4BEG[5]
rlabel metal2 3752 110936 3752 110936 0 Tile_X0Y0_N4BEG[6]
rlabel metal2 11480 112042 11480 112042 0 Tile_X0Y0_N4BEG[7]
rlabel metal2 8120 112336 8120 112336 0 Tile_X0Y0_N4BEG[8]
rlabel metal2 20608 112392 20608 112392 0 Tile_X0Y0_N4BEG[9]
rlabel metal3 16800 96152 16800 96152 0 Tile_X0Y0_S1END[0]
rlabel metal2 11536 86744 11536 86744 0 Tile_X0Y0_S1END[1]
rlabel metal2 6104 110152 6104 110152 0 Tile_X0Y0_S1END[2]
rlabel metal2 20664 61320 20664 61320 0 Tile_X0Y0_S1END[3]
rlabel metal2 16184 113722 16184 113722 0 Tile_X0Y0_S2END[0]
rlabel metal2 16408 114058 16408 114058 0 Tile_X0Y0_S2END[1]
rlabel metal2 16632 113722 16632 113722 0 Tile_X0Y0_S2END[2]
rlabel metal2 16856 113554 16856 113554 0 Tile_X0Y0_S2END[3]
rlabel metal2 17080 113722 17080 113722 0 Tile_X0Y0_S2END[4]
rlabel metal2 17304 114002 17304 114002 0 Tile_X0Y0_S2END[5]
rlabel metal2 17528 114114 17528 114114 0 Tile_X0Y0_S2END[6]
rlabel metal2 17752 112098 17752 112098 0 Tile_X0Y0_S2END[7]
rlabel metal2 10136 2856 10136 2856 0 Tile_X0Y0_S2MID[0]
rlabel metal2 14616 114114 14616 114114 0 Tile_X0Y0_S2MID[1]
rlabel metal2 16744 34608 16744 34608 0 Tile_X0Y0_S2MID[2]
rlabel metal3 19824 55496 19824 55496 0 Tile_X0Y0_S2MID[3]
rlabel metal3 11704 2520 11704 2520 0 Tile_X0Y0_S2MID[4]
rlabel metal2 15512 112266 15512 112266 0 Tile_X0Y0_S2MID[5]
rlabel metal2 15736 112490 15736 112490 0 Tile_X0Y0_S2MID[6]
rlabel metal3 16016 49784 16016 49784 0 Tile_X0Y0_S2MID[7]
rlabel metal2 17976 114114 17976 114114 0 Tile_X0Y0_S4END[0]
rlabel metal2 19096 109984 19096 109984 0 Tile_X0Y0_S4END[10]
rlabel metal2 20440 114058 20440 114058 0 Tile_X0Y0_S4END[11]
rlabel metal2 19880 110544 19880 110544 0 Tile_X0Y0_S4END[12]
rlabel metal2 22008 111048 22008 111048 0 Tile_X0Y0_S4END[13]
rlabel metal2 21112 113386 21112 113386 0 Tile_X0Y0_S4END[14]
rlabel metal2 22792 111496 22792 111496 0 Tile_X0Y0_S4END[15]
rlabel metal2 18200 111482 18200 111482 0 Tile_X0Y0_S4END[1]
rlabel metal2 18424 114002 18424 114002 0 Tile_X0Y0_S4END[2]
rlabel metal3 21000 67592 21000 67592 0 Tile_X0Y0_S4END[3]
rlabel metal2 18872 114394 18872 114394 0 Tile_X0Y0_S4END[4]
rlabel metal2 19096 114170 19096 114170 0 Tile_X0Y0_S4END[5]
rlabel metal2 18872 68432 18872 68432 0 Tile_X0Y0_S4END[6]
rlabel metal2 19544 114170 19544 114170 0 Tile_X0Y0_S4END[7]
rlabel metal2 19768 113666 19768 113666 0 Tile_X0Y0_S4END[8]
rlabel metal3 20720 110936 20720 110936 0 Tile_X0Y0_S4END[9]
rlabel metal3 23072 113512 23072 113512 0 Tile_X0Y0_UserCLKo
rlabel metal3 910 57736 910 57736 0 Tile_X0Y0_W1BEG[0]
rlabel metal3 574 58184 574 58184 0 Tile_X0Y0_W1BEG[1]
rlabel metal3 518 58632 518 58632 0 Tile_X0Y0_W1BEG[2]
rlabel metal3 1302 59080 1302 59080 0 Tile_X0Y0_W1BEG[3]
rlabel metal3 574 59528 574 59528 0 Tile_X0Y0_W2BEG[0]
rlabel metal3 518 59976 518 59976 0 Tile_X0Y0_W2BEG[1]
rlabel metal3 462 60424 462 60424 0 Tile_X0Y0_W2BEG[2]
rlabel metal2 1064 57680 1064 57680 0 Tile_X0Y0_W2BEG[3]
rlabel metal3 406 61320 406 61320 0 Tile_X0Y0_W2BEG[4]
rlabel metal3 966 61768 966 61768 0 Tile_X0Y0_W2BEG[5]
rlabel metal3 294 62216 294 62216 0 Tile_X0Y0_W2BEG[6]
rlabel metal3 238 62664 238 62664 0 Tile_X0Y0_W2BEG[7]
rlabel metal3 126 63112 126 63112 0 Tile_X0Y0_W2BEGb[0]
rlabel metal3 1722 63560 1722 63560 0 Tile_X0Y0_W2BEGb[1]
rlabel metal3 462 64008 462 64008 0 Tile_X0Y0_W2BEGb[2]
rlabel metal2 3976 64848 3976 64848 0 Tile_X0Y0_W2BEGb[3]
rlabel metal2 4984 65072 4984 65072 0 Tile_X0Y0_W2BEGb[4]
rlabel metal3 1806 65352 1806 65352 0 Tile_X0Y0_W2BEGb[5]
rlabel metal3 406 65800 406 65800 0 Tile_X0Y0_W2BEGb[6]
rlabel metal3 462 66248 462 66248 0 Tile_X0Y0_W2BEGb[7]
rlabel metal3 3598 73864 3598 73864 0 Tile_X0Y0_W6BEG[0]
rlabel metal3 966 78344 966 78344 0 Tile_X0Y0_W6BEG[10]
rlabel metal3 1722 78792 1722 78792 0 Tile_X0Y0_W6BEG[11]
rlabel metal2 5656 75264 5656 75264 0 Tile_X0Y0_W6BEG[1]
rlabel metal3 406 74760 406 74760 0 Tile_X0Y0_W6BEG[2]
rlabel metal3 462 75208 462 75208 0 Tile_X0Y0_W6BEG[3]
rlabel metal3 686 75656 686 75656 0 Tile_X0Y0_W6BEG[4]
rlabel metal3 518 76104 518 76104 0 Tile_X0Y0_W6BEG[5]
rlabel metal3 616 85736 616 85736 0 Tile_X0Y0_W6BEG[6]
rlabel metal3 350 77000 350 77000 0 Tile_X0Y0_W6BEG[7]
rlabel metal3 5544 77504 5544 77504 0 Tile_X0Y0_W6BEG[8]
rlabel metal3 910 77896 910 77896 0 Tile_X0Y0_W6BEG[9]
rlabel metal3 182 66696 182 66696 0 Tile_X0Y0_WW4BEG[0]
rlabel metal2 5656 72128 5656 72128 0 Tile_X0Y0_WW4BEG[10]
rlabel metal2 6328 71792 6328 71792 0 Tile_X0Y0_WW4BEG[11]
rlabel metal3 518 72072 518 72072 0 Tile_X0Y0_WW4BEG[12]
rlabel metal3 854 72520 854 72520 0 Tile_X0Y0_WW4BEG[13]
rlabel metal3 1358 72968 1358 72968 0 Tile_X0Y0_WW4BEG[14]
rlabel metal3 3318 73416 3318 73416 0 Tile_X0Y0_WW4BEG[15]
rlabel metal3 350 67144 350 67144 0 Tile_X0Y0_WW4BEG[1]
rlabel metal3 910 67592 910 67592 0 Tile_X0Y0_WW4BEG[2]
rlabel metal3 126 68040 126 68040 0 Tile_X0Y0_WW4BEG[3]
rlabel metal2 4872 70000 4872 70000 0 Tile_X0Y0_WW4BEG[4]
rlabel metal3 3640 69104 3640 69104 0 Tile_X0Y0_WW4BEG[5]
rlabel metal3 126 69384 126 69384 0 Tile_X0Y0_WW4BEG[6]
rlabel metal3 1722 69832 1722 69832 0 Tile_X0Y0_WW4BEG[7]
rlabel metal2 5432 70728 5432 70728 0 Tile_X0Y0_WW4BEG[8]
rlabel metal3 462 70728 462 70728 0 Tile_X0Y0_WW4BEG[9]
rlabel metal2 16856 26096 16856 26096 0 Tile_X0Y1_E1END[0]
rlabel metal2 15848 50904 15848 50904 0 Tile_X0Y1_E1END[1]
rlabel metal3 7840 23576 7840 23576 0 Tile_X0Y1_E1END[2]
rlabel metal2 23016 24024 23016 24024 0 Tile_X0Y1_E1END[3]
rlabel metal2 19096 24192 19096 24192 0 Tile_X0Y1_E2END[0]
rlabel metal2 16744 17752 16744 17752 0 Tile_X0Y1_E2END[1]
rlabel metal2 16968 23240 16968 23240 0 Tile_X0Y1_E2END[2]
rlabel metal3 1722 28504 1722 28504 0 Tile_X0Y1_E2END[3]
rlabel metal2 19992 36344 19992 36344 0 Tile_X0Y1_E2END[4]
rlabel metal2 18536 27832 18536 27832 0 Tile_X0Y1_E2END[5]
rlabel metal2 16072 43344 16072 43344 0 Tile_X0Y1_E2END[6]
rlabel metal3 1722 30296 1722 30296 0 Tile_X0Y1_E2END[7]
rlabel metal2 17192 22736 17192 22736 0 Tile_X0Y1_E2MID[0]
rlabel metal2 17976 18760 17976 18760 0 Tile_X0Y1_E2MID[1]
rlabel metal2 17472 18312 17472 18312 0 Tile_X0Y1_E2MID[2]
rlabel metal2 20608 24696 20608 24696 0 Tile_X0Y1_E2MID[3]
rlabel metal3 17024 37240 17024 37240 0 Tile_X0Y1_E2MID[4]
rlabel metal3 1722 25816 1722 25816 0 Tile_X0Y1_E2MID[5]
rlabel metal3 238 26264 238 26264 0 Tile_X0Y1_E2MID[6]
rlabel metal3 1722 26712 1722 26712 0 Tile_X0Y1_E2MID[7]
rlabel metal2 16184 38808 16184 38808 0 Tile_X0Y1_E6END[0]
rlabel metal3 1722 42392 1722 42392 0 Tile_X0Y1_E6END[10]
rlabel metal2 20216 41944 20216 41944 0 Tile_X0Y1_E6END[11]
rlabel metal2 13944 42616 13944 42616 0 Tile_X0Y1_E6END[1]
rlabel metal2 4928 42728 4928 42728 0 Tile_X0Y1_E6END[2]
rlabel metal2 23576 25396 23576 25396 0 Tile_X0Y1_E6END[3]
rlabel metal3 15512 38808 15512 38808 0 Tile_X0Y1_E6END[4]
rlabel metal2 12264 43624 12264 43624 0 Tile_X0Y1_E6END[5]
rlabel metal3 2296 47600 2296 47600 0 Tile_X0Y1_E6END[6]
rlabel metal3 910 41048 910 41048 0 Tile_X0Y1_E6END[7]
rlabel metal3 1358 41496 1358 41496 0 Tile_X0Y1_E6END[8]
rlabel metal3 966 41944 966 41944 0 Tile_X0Y1_E6END[9]
rlabel metal3 1722 30744 1722 30744 0 Tile_X0Y1_EE4END[0]
rlabel metal2 1120 41832 1120 41832 0 Tile_X0Y1_EE4END[10]
rlabel metal2 20776 35224 20776 35224 0 Tile_X0Y1_EE4END[11]
rlabel metal3 1722 36120 1722 36120 0 Tile_X0Y1_EE4END[12]
rlabel metal3 9296 35672 9296 35672 0 Tile_X0Y1_EE4END[13]
rlabel metal2 1904 41944 1904 41944 0 Tile_X0Y1_EE4END[14]
rlabel metal2 21448 34888 21448 34888 0 Tile_X0Y1_EE4END[15]
rlabel metal2 8512 41384 8512 41384 0 Tile_X0Y1_EE4END[1]
rlabel metal3 182 31640 182 31640 0 Tile_X0Y1_EE4END[2]
rlabel metal3 18368 37576 18368 37576 0 Tile_X0Y1_EE4END[3]
rlabel metal2 11144 30576 11144 30576 0 Tile_X0Y1_EE4END[4]
rlabel metal3 1722 32984 1722 32984 0 Tile_X0Y1_EE4END[5]
rlabel metal2 3192 41888 3192 41888 0 Tile_X0Y1_EE4END[6]
rlabel metal2 22792 33600 22792 33600 0 Tile_X0Y1_EE4END[7]
rlabel metal2 8904 28560 8904 28560 0 Tile_X0Y1_EE4END[8]
rlabel metal2 5376 35560 5376 35560 0 Tile_X0Y1_EE4END[9]
rlabel metal2 29512 39816 29512 39816 0 Tile_X0Y1_FrameData[0]
rlabel metal2 2296 47936 2296 47936 0 Tile_X0Y1_FrameData[10]
rlabel metal2 16856 52304 16856 52304 0 Tile_X0Y1_FrameData[11]
rlabel metal2 2520 52136 2520 52136 0 Tile_X0Y1_FrameData[12]
rlabel metal2 3080 52024 3080 52024 0 Tile_X0Y1_FrameData[13]
rlabel metal3 6664 3304 6664 3304 0 Tile_X0Y1_FrameData[14]
rlabel metal2 6888 1904 6888 1904 0 Tile_X0Y1_FrameData[15]
rlabel metal2 21000 53816 21000 53816 0 Tile_X0Y1_FrameData[16]
rlabel metal3 1638 50904 1638 50904 0 Tile_X0Y1_FrameData[17]
rlabel metal3 1526 51352 1526 51352 0 Tile_X0Y1_FrameData[18]
rlabel metal3 3080 51912 3080 51912 0 Tile_X0Y1_FrameData[19]
rlabel metal2 3864 1960 3864 1960 0 Tile_X0Y1_FrameData[1]
rlabel metal2 29288 58464 29288 58464 0 Tile_X0Y1_FrameData[20]
rlabel metal2 1512 53312 1512 53312 0 Tile_X0Y1_FrameData[21]
rlabel metal3 29176 63112 29176 63112 0 Tile_X0Y1_FrameData[22]
rlabel metal4 3304 52581 3304 52581 0 Tile_X0Y1_FrameData[23]
rlabel metal3 686 54040 686 54040 0 Tile_X0Y1_FrameData[24]
rlabel metal3 20244 53928 20244 53928 0 Tile_X0Y1_FrameData[25]
rlabel metal3 966 54936 966 54936 0 Tile_X0Y1_FrameData[26]
rlabel metal3 1022 55384 1022 55384 0 Tile_X0Y1_FrameData[27]
rlabel metal3 1302 55832 1302 55832 0 Tile_X0Y1_FrameData[28]
rlabel metal2 22792 44520 22792 44520 0 Tile_X0Y1_FrameData[29]
rlabel metal2 29456 41720 29456 41720 0 Tile_X0Y1_FrameData[2]
rlabel metal3 686 56728 686 56728 0 Tile_X0Y1_FrameData[30]
rlabel metal2 19488 59976 19488 59976 0 Tile_X0Y1_FrameData[31]
rlabel metal2 29344 43288 29344 43288 0 Tile_X0Y1_FrameData[3]
rlabel metal2 2296 1232 2296 1232 0 Tile_X0Y1_FrameData[4]
rlabel metal3 910 45528 910 45528 0 Tile_X0Y1_FrameData[5]
rlabel metal2 22176 42392 22176 42392 0 Tile_X0Y1_FrameData[6]
rlabel metal2 18144 1064 18144 1064 0 Tile_X0Y1_FrameData[7]
rlabel metal3 13160 2072 13160 2072 0 Tile_X0Y1_FrameData[8]
rlabel metal3 17864 2184 17864 2184 0 Tile_X0Y1_FrameData[9]
rlabel metal3 31122 39928 31122 39928 0 Tile_X0Y1_FrameData_O[0]
rlabel metal3 31122 51128 31122 51128 0 Tile_X0Y1_FrameData_O[10]
rlabel metal3 31122 52248 31122 52248 0 Tile_X0Y1_FrameData_O[11]
rlabel metal3 31122 53368 31122 53368 0 Tile_X0Y1_FrameData_O[12]
rlabel metal2 30632 54432 30632 54432 0 Tile_X0Y1_FrameData_O[13]
rlabel metal3 31122 55608 31122 55608 0 Tile_X0Y1_FrameData_O[14]
rlabel metal3 31122 56728 31122 56728 0 Tile_X0Y1_FrameData_O[15]
rlabel metal3 31122 57848 31122 57848 0 Tile_X0Y1_FrameData_O[16]
rlabel metal3 31122 58968 31122 58968 0 Tile_X0Y1_FrameData_O[17]
rlabel metal3 31122 60088 31122 60088 0 Tile_X0Y1_FrameData_O[18]
rlabel metal3 31122 61208 31122 61208 0 Tile_X0Y1_FrameData_O[19]
rlabel metal3 31122 41048 31122 41048 0 Tile_X0Y1_FrameData_O[1]
rlabel metal3 31122 62328 31122 62328 0 Tile_X0Y1_FrameData_O[20]
rlabel metal3 31122 63448 31122 63448 0 Tile_X0Y1_FrameData_O[21]
rlabel metal3 31122 64568 31122 64568 0 Tile_X0Y1_FrameData_O[22]
rlabel metal3 31122 65688 31122 65688 0 Tile_X0Y1_FrameData_O[23]
rlabel metal3 31122 66808 31122 66808 0 Tile_X0Y1_FrameData_O[24]
rlabel metal3 31122 67928 31122 67928 0 Tile_X0Y1_FrameData_O[25]
rlabel metal3 31122 69048 31122 69048 0 Tile_X0Y1_FrameData_O[26]
rlabel metal3 31122 70168 31122 70168 0 Tile_X0Y1_FrameData_O[27]
rlabel metal3 31122 71288 31122 71288 0 Tile_X0Y1_FrameData_O[28]
rlabel metal3 31122 72408 31122 72408 0 Tile_X0Y1_FrameData_O[29]
rlabel metal3 31122 42168 31122 42168 0 Tile_X0Y1_FrameData_O[2]
rlabel metal3 31122 73528 31122 73528 0 Tile_X0Y1_FrameData_O[30]
rlabel metal3 31122 74648 31122 74648 0 Tile_X0Y1_FrameData_O[31]
rlabel metal3 31122 43288 31122 43288 0 Tile_X0Y1_FrameData_O[3]
rlabel metal3 31122 44408 31122 44408 0 Tile_X0Y1_FrameData_O[4]
rlabel metal3 31122 45528 31122 45528 0 Tile_X0Y1_FrameData_O[5]
rlabel metal3 31122 46648 31122 46648 0 Tile_X0Y1_FrameData_O[6]
rlabel metal3 31122 47768 31122 47768 0 Tile_X0Y1_FrameData_O[7]
rlabel metal3 31122 48888 31122 48888 0 Tile_X0Y1_FrameData_O[8]
rlabel metal3 31122 50008 31122 50008 0 Tile_X0Y1_FrameData_O[9]
rlabel metal2 12712 1120 12712 1120 0 Tile_X0Y1_FrameStrobe[0]
rlabel metal2 27272 1960 27272 1960 0 Tile_X0Y1_FrameStrobe[10]
rlabel metal4 27048 56168 27048 56168 0 Tile_X0Y1_FrameStrobe[11]
rlabel metal2 27272 57624 27272 57624 0 Tile_X0Y1_FrameStrobe[12]
rlabel metal2 24696 350 24696 350 0 Tile_X0Y1_FrameStrobe[13]
rlabel metal2 24920 686 24920 686 0 Tile_X0Y1_FrameStrobe[14]
rlabel metal4 21336 57288 21336 57288 0 Tile_X0Y1_FrameStrobe[15]
rlabel metal3 25648 110040 25648 110040 0 Tile_X0Y1_FrameStrobe[16]
rlabel metal2 26824 109648 26824 109648 0 Tile_X0Y1_FrameStrobe[17]
rlabel metal3 26712 89096 26712 89096 0 Tile_X0Y1_FrameStrobe[18]
rlabel metal2 28392 5012 28392 5012 0 Tile_X0Y1_FrameStrobe[19]
rlabel metal2 2632 51688 2632 51688 0 Tile_X0Y1_FrameStrobe[1]
rlabel metal2 1456 55440 1456 55440 0 Tile_X0Y1_FrameStrobe[2]
rlabel metal2 2800 51352 2800 51352 0 Tile_X0Y1_FrameStrobe[3]
rlabel metal2 3416 2296 3416 2296 0 Tile_X0Y1_FrameStrobe[4]
rlabel metal2 2632 60312 2632 60312 0 Tile_X0Y1_FrameStrobe[5]
rlabel metal2 1512 48216 1512 48216 0 Tile_X0Y1_FrameStrobe[6]
rlabel metal2 2856 40656 2856 40656 0 Tile_X0Y1_FrameStrobe[7]
rlabel metal3 17360 52024 17360 52024 0 Tile_X0Y1_FrameStrobe[8]
rlabel metal2 27384 57624 27384 57624 0 Tile_X0Y1_FrameStrobe[9]
rlabel metal2 15064 9296 15064 9296 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit0.Q
rlabel metal2 16296 7728 16296 7728 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit1.Q
rlabel metal3 7112 52360 7112 52360 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit10.Q
rlabel metal2 8232 49812 8232 49812 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit11.Q
rlabel metal2 14392 33432 14392 33432 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit12.Q
rlabel metal3 12880 35000 12880 35000 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit13.Q
rlabel metal2 18200 47768 18200 47768 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit14.Q
rlabel metal3 16520 47432 16520 47432 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit15.Q
rlabel metal2 14280 2464 14280 2464 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit16.Q
rlabel metal2 11816 1792 11816 1792 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit17.Q
rlabel metal3 8624 19432 8624 19432 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit18.Q
rlabel metal3 9184 19992 9184 19992 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit19.Q
rlabel metal2 10696 46144 10696 46144 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit2.Q
rlabel metal2 14616 54768 14616 54768 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit20.Q
rlabel metal2 16072 53816 16072 53816 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit21.Q
rlabel metal2 15904 48440 15904 48440 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit22.Q
rlabel metal2 16856 50064 16856 50064 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit23.Q
rlabel metal2 15288 18928 15288 18928 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit24.Q
rlabel metal2 13944 22848 13944 22848 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit25.Q
rlabel metal2 13048 47208 13048 47208 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit26.Q
rlabel metal2 13384 48496 13384 48496 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit27.Q
rlabel metal2 8288 44520 8288 44520 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit28.Q
rlabel metal3 8680 45864 8680 45864 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit29.Q
rlabel metal2 12096 45304 12096 45304 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit3.Q
rlabel metal2 23576 22512 23576 22512 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit30.Q
rlabel metal2 23352 22064 23352 22064 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit31.Q
rlabel metal2 6776 43624 6776 43624 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit4.Q
rlabel metal2 7560 45136 7560 45136 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit5.Q
rlabel metal2 20776 7224 20776 7224 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit6.Q
rlabel metal3 22568 6664 22568 6664 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit7.Q
rlabel metal2 10584 2576 10584 2576 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit8.Q
rlabel metal2 9464 2968 9464 2968 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame0_bit9.Q
rlabel metal2 6888 37520 6888 37520 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q
rlabel metal3 7784 34328 7784 34328 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q
rlabel metal2 9912 53760 9912 53760 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit10.Q
rlabel metal2 11144 54376 11144 54376 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit11.Q
rlabel metal2 5320 52416 5320 52416 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit12.Q
rlabel metal2 6440 52024 6440 52024 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit13.Q
rlabel metal2 21448 13440 21448 13440 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit14.Q
rlabel metal3 21896 14728 21896 14728 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit15.Q
rlabel metal2 15288 4424 15288 4424 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit16.Q
rlabel metal3 15960 4536 15960 4536 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit17.Q
rlabel metal3 10080 56840 10080 56840 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit18.Q
rlabel metal2 11704 57120 11704 57120 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit19.Q
rlabel metal2 1624 41776 1624 41776 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q
rlabel metal2 6048 54488 6048 54488 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit20.Q
rlabel metal2 7448 55160 7448 55160 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit21.Q
rlabel metal2 20832 12376 20832 12376 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit22.Q
rlabel metal2 22736 15064 22736 15064 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit23.Q
rlabel metal3 13048 9016 13048 9016 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit24.Q
rlabel metal2 15176 9688 15176 9688 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit25.Q
rlabel metal2 9464 57512 9464 57512 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit26.Q
rlabel metal2 10696 57008 10696 57008 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit27.Q
rlabel metal3 4592 54712 4592 54712 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit28.Q
rlabel metal3 5600 55272 5600 55272 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit29.Q
rlabel metal2 2744 40880 2744 40880 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit3.Q
rlabel metal2 20720 8456 20720 8456 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit30.Q
rlabel metal3 22176 9240 22176 9240 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit31.Q
rlabel metal3 4256 40376 4256 40376 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q
rlabel metal2 22680 36344 22680 36344 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q
rlabel metal2 22344 35560 22344 35560 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q
rlabel metal3 24080 31864 24080 31864 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit7.Q
rlabel metal3 13664 5096 13664 5096 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit8.Q
rlabel metal3 13440 6664 13440 6664 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame1_bit9.Q
rlabel metal2 21000 29736 21000 29736 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit0.Q
rlabel metal2 18312 29680 18312 29680 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit1.Q
rlabel metal3 8176 24584 8176 24584 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit10.Q
rlabel metal3 6104 34888 6104 34888 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit11.Q
rlabel metal2 7896 36568 7896 36568 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit12.Q
rlabel metal3 8624 32760 8624 32760 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit13.Q
rlabel metal3 2240 44856 2240 44856 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit14.Q
rlabel metal2 2408 44968 2408 44968 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit15.Q
rlabel metal2 5264 40936 5264 40936 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit16.Q
rlabel metal2 22568 35952 22568 35952 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit17.Q
rlabel metal2 22456 35952 22456 35952 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit18.Q
rlabel metal2 23464 33824 23464 33824 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit19.Q
rlabel metal3 17976 30184 17976 30184 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit2.Q
rlabel metal2 20720 21000 20720 21000 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit20.Q
rlabel metal2 19936 19880 19936 19880 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit21.Q
rlabel metal3 18144 19432 18144 19432 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit22.Q
rlabel metal2 15960 20160 15960 20160 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit23.Q
rlabel metal2 16856 19404 16856 19404 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit24.Q
rlabel metal2 17248 20104 17248 20104 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit25.Q
rlabel metal3 21224 26488 21224 26488 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit26.Q
rlabel metal3 22232 25480 22232 25480 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit27.Q
rlabel metal2 9240 28112 9240 28112 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q
rlabel metal3 9856 27048 9856 27048 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q
rlabel metal3 22232 27944 22232 27944 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit3.Q
rlabel metal3 10864 23128 10864 23128 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q
rlabel metal3 6832 37128 6832 37128 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit31.Q
rlabel metal3 16632 35672 16632 35672 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit4.Q
rlabel metal2 19320 37072 19320 37072 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit5.Q
rlabel metal2 18760 33152 18760 33152 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit6.Q
rlabel metal2 20328 36624 20328 36624 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit7.Q
rlabel metal2 10360 26572 10360 26572 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit8.Q
rlabel metal2 9128 26768 9128 26768 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame2_bit9.Q
rlabel metal2 18256 12376 18256 12376 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit0.Q
rlabel metal2 19600 15064 19600 15064 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit1.Q
rlabel metal2 7224 46928 7224 46928 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit10.Q
rlabel metal2 8344 47320 8344 47320 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit11.Q
rlabel metal2 3920 50680 3920 50680 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit12.Q
rlabel metal2 5544 50904 5544 50904 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit13.Q
rlabel metal3 13776 13160 13776 13160 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit14.Q
rlabel metal2 15064 14000 15064 14000 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit15.Q
rlabel metal2 19712 17080 19712 17080 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit16.Q
rlabel metal2 20944 16296 20944 16296 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit17.Q
rlabel metal3 1456 32760 1456 32760 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit18.Q
rlabel metal2 2968 35336 2968 35336 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit19.Q
rlabel metal2 3304 31864 3304 31864 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit2.Q
rlabel metal2 5488 17864 5488 17864 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit20.Q
rlabel metal3 6832 16296 6832 16296 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit21.Q
rlabel metal3 12152 16072 12152 16072 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit22.Q
rlabel metal3 12992 14728 12992 14728 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit23.Q
rlabel metal2 18200 14224 18200 14224 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit24.Q
rlabel metal2 17472 15064 17472 15064 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit25.Q
rlabel metal2 5096 32256 5096 32256 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit26.Q
rlabel metal2 2912 32088 2912 32088 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit27.Q
rlabel metal2 8288 18424 8288 18424 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit28.Q
rlabel metal2 7728 17864 7728 17864 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit29.Q
rlabel metal2 5600 31864 5600 31864 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit3.Q
rlabel metal2 10136 15568 10136 15568 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit30.Q
rlabel metal3 8344 15288 8344 15288 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit31.Q
rlabel metal3 7000 11592 7000 11592 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit4.Q
rlabel metal3 5768 10024 5768 10024 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit5.Q
rlabel metal2 7896 13048 7896 13048 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit6.Q
rlabel metal2 10136 13048 10136 13048 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit7.Q
rlabel metal2 17864 4984 17864 4984 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit8.Q
rlabel metal2 18704 6664 18704 6664 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame3_bit9.Q
rlabel metal3 11312 15176 11312 15176 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit0.Q
rlabel metal3 6720 2184 6720 2184 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit1.Q
rlabel metal2 3696 22568 3696 22568 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit10.Q
rlabel metal2 1176 17360 1176 17360 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit11.Q
rlabel metal2 4312 24136 4312 24136 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit12.Q
rlabel metal2 3024 21784 3024 21784 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit13.Q
rlabel metal2 11928 8904 11928 8904 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit14.Q
rlabel metal3 12600 8344 12600 8344 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit15.Q
rlabel metal2 20832 6104 20832 6104 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit16.Q
rlabel metal2 22512 4536 22512 4536 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit17.Q
rlabel metal2 3192 33208 3192 33208 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit18.Q
rlabel metal2 1232 29624 1232 29624 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit19.Q
rlabel metal2 3024 19544 3024 19544 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit2.Q
rlabel metal3 3696 5880 3696 5880 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit20.Q
rlabel metal3 8176 16856 8176 16856 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit21.Q
rlabel metal2 11144 8512 11144 8512 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit22.Q
rlabel metal2 12600 10472 12600 10472 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit23.Q
rlabel metal2 18536 11088 18536 11088 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit24.Q
rlabel metal2 19768 10696 19768 10696 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit25.Q
rlabel metal2 5096 30016 5096 30016 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit26.Q
rlabel metal2 2744 24920 2744 24920 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit27.Q
rlabel metal3 7112 17080 7112 17080 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit28.Q
rlabel metal2 5096 15568 5096 15568 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit29.Q
rlabel metal3 4312 15400 4312 15400 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit3.Q
rlabel metal3 12264 10584 12264 10584 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit30.Q
rlabel metal2 10696 5376 10696 5376 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit31.Q
rlabel metal2 3472 1400 3472 1400 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit4.Q
rlabel metal2 24136 1400 24136 1400 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit5.Q
rlabel metal3 10360 5712 10360 5712 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit6.Q
rlabel metal2 23016 6160 23016 6160 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit7.Q
rlabel metal2 18200 3248 18200 3248 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit8.Q
rlabel metal2 19264 2184 19264 2184 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame4_bit9.Q
rlabel metal2 12712 4424 12712 4424 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit0.Q
rlabel metal2 11704 2408 11704 2408 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit1.Q
rlabel metal2 3752 25648 3752 25648 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit10.Q
rlabel metal2 4592 22568 4592 22568 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit11.Q
rlabel metal2 3304 19880 3304 19880 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit12.Q
rlabel metal2 1176 18760 1176 18760 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit13.Q
rlabel metal2 7336 2184 7336 2184 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit14.Q
rlabel metal2 8008 1680 8008 1680 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit15.Q
rlabel metal2 23016 4648 23016 4648 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit16.Q
rlabel metal2 21448 3920 21448 3920 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit17.Q
rlabel metal2 2856 11648 2856 11648 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit18.Q
rlabel metal2 1288 16408 1288 16408 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit19.Q
rlabel metal2 10696 18144 10696 18144 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit2.Q
rlabel metal3 4144 2968 4144 2968 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit20.Q
rlabel metal2 18312 13328 18312 13328 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit21.Q
rlabel metal4 11816 8904 11816 8904 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit22.Q
rlabel metal3 16212 9128 16212 9128 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit23.Q
rlabel metal3 17528 8008 17528 8008 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit24.Q
rlabel metal2 9184 15736 9184 15736 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit25.Q
rlabel metal3 2912 16296 2912 16296 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit26.Q
rlabel metal2 2856 17808 2856 17808 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit27.Q
rlabel metal2 3640 15512 3640 15512 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit28.Q
rlabel metal2 2856 11032 2856 11032 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit29.Q
rlabel metal2 9464 17752 9464 17752 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit3.Q
rlabel metal2 6888 5992 6888 5992 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit30.Q
rlabel metal2 4312 6720 4312 6720 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit31.Q
rlabel metal2 7224 11872 7224 11872 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit4.Q
rlabel metal2 4312 10416 4312 10416 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit5.Q
rlabel metal2 21448 4312 21448 4312 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit6.Q
rlabel metal2 19544 1400 19544 1400 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit7.Q
rlabel metal2 22960 2968 22960 2968 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit8.Q
rlabel metal4 22120 6440 22120 6440 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame5_bit9.Q
rlabel metal2 9072 40600 9072 40600 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit0.Q
rlabel metal2 10808 42448 10808 42448 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit1.Q
rlabel metal2 16016 36680 16016 36680 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit10.Q
rlabel metal2 15064 35952 15064 35952 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit11.Q
rlabel metal2 15848 28504 15848 28504 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit12.Q
rlabel metal2 14504 29288 14504 29288 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit13.Q
rlabel metal2 12152 22232 12152 22232 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit14.Q
rlabel metal3 12208 20776 12208 20776 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit15.Q
rlabel metal3 11536 19208 11536 19208 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit16.Q
rlabel metal2 13104 17864 13104 17864 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit17.Q
rlabel metal3 18816 21560 18816 21560 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit18.Q
rlabel metal2 16912 21000 16912 21000 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit19.Q
rlabel metal2 20048 22344 20048 22344 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit2.Q
rlabel metal2 15736 26992 15736 26992 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit20.Q
rlabel metal3 14000 28616 14000 28616 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit21.Q
rlabel metal2 16240 26488 16240 26488 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit22.Q
rlabel metal2 10472 35672 10472 35672 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit23.Q
rlabel metal2 11816 36792 11816 36792 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit24.Q
rlabel metal2 13048 32816 13048 32816 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit25.Q
rlabel metal2 3192 47040 3192 47040 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit26.Q
rlabel metal2 3024 49000 3024 49000 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit27.Q
rlabel metal2 1624 48776 1624 48776 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit28.Q
rlabel metal2 22120 41160 22120 41160 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit29.Q
rlabel metal2 21224 22568 21224 22568 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit3.Q
rlabel metal2 21000 42448 21000 42448 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit30.Q
rlabel metal2 21784 41552 21784 41552 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit31.Q
rlabel metal3 7280 23352 7280 23352 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit4.Q
rlabel metal3 7168 24136 7168 24136 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit5.Q
rlabel metal3 14784 43512 14784 43512 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit6.Q
rlabel metal2 15736 43792 15736 43792 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit7.Q
rlabel metal2 12376 39312 12376 39312 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit8.Q
rlabel metal3 10584 39032 10584 39032 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame6_bit9.Q
rlabel metal3 7392 24920 7392 24920 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit0.Q
rlabel metal2 7224 25704 7224 25704 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit1.Q
rlabel metal2 10584 31864 10584 31864 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q
rlabel metal2 9016 32648 9016 32648 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit11.Q
rlabel metal2 13832 42224 13832 42224 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q
rlabel metal2 14616 41664 14616 41664 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q
rlabel metal2 16520 40656 16520 40656 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit14.Q
rlabel metal2 17864 41048 17864 41048 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q
rlabel metal3 12432 29960 12432 29960 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q
rlabel metal2 12208 30744 12208 30744 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit17.Q
rlabel metal2 15736 31192 15736 31192 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit18.Q
rlabel metal2 10696 51296 10696 51296 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit19.Q
rlabel metal2 9352 43736 9352 43736 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit2.Q
rlabel metal2 9352 51408 9352 51408 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit20.Q
rlabel metal2 12040 53592 12040 53592 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit21.Q
rlabel metal2 6552 40488 6552 40488 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit22.Q
rlabel metal2 5320 41552 5320 41552 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit23.Q
rlabel metal3 8288 41832 8288 41832 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit24.Q
rlabel metal2 19432 43008 19432 43008 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit25.Q
rlabel metal2 18424 42728 18424 42728 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit26.Q
rlabel metal2 18984 45584 18984 45584 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit27.Q
rlabel metal2 13160 21840 13160 21840 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit28.Q
rlabel metal2 14280 21840 14280 21840 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit29.Q
rlabel metal2 11592 44016 11592 44016 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit3.Q
rlabel metal2 12152 50288 12152 50288 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit30.Q
rlabel metal2 13272 50288 13272 50288 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit31.Q
rlabel metal2 11480 40656 11480 40656 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit4.Q
rlabel metal3 9408 40600 9408 40600 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit5.Q
rlabel metal2 15456 38248 15456 38248 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q
rlabel metal3 13664 38808 13664 38808 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit7.Q
rlabel metal2 15624 32816 15624 32816 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit8.Q
rlabel metal3 16520 32536 16520 32536 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q
rlabel metal2 16072 23632 16072 23632 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit24.Q
rlabel metal2 16072 25312 16072 25312 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit25.Q
rlabel metal2 14280 51632 14280 51632 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit26.Q
rlabel metal2 13104 51352 13104 51352 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit27.Q
rlabel metal2 10696 48160 10696 48160 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit28.Q
rlabel metal2 9576 47712 9576 47712 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit29.Q
rlabel metal3 21840 43512 21840 43512 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit30.Q
rlabel metal2 21000 43792 21000 43792 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_ConfigMem.Inst_frame8_bit31.Q
rlabel metal2 15792 5768 15792 5768 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG4
rlabel metal3 8400 20776 8400 20776 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG5
rlabel metal2 2856 42280 2856 42280 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG6
rlabel metal2 21224 18760 21224 18760 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.J_NS4_BEG7
rlabel metal2 13496 8232 13496 8232 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S1BEG0
rlabel metal3 12544 50680 12544 50680 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S1BEG1
rlabel metal3 9576 40488 9576 40488 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S1BEG2
rlabel metal3 20048 21224 20048 21224 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S1BEG3
rlabel metal2 7392 25928 7392 25928 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG0
rlabel metal3 14728 43288 14728 43288 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG1
rlabel metal3 11480 4312 11480 4312 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG2
rlabel metal3 15344 37016 15344 37016 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG3
rlabel metal3 15960 5096 15960 5096 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG4
rlabel metal2 12880 15624 12880 15624 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG5
rlabel metal3 12936 19320 12936 19320 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG6
rlabel metal3 17024 18200 17024 18200 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S2BEG7
rlabel metal3 18312 26824 18312 26824 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S4BEG0
rlabel metal3 15568 26264 15568 26264 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S4BEG1
rlabel metal2 20216 47992 20216 47992 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S4BEG2
rlabel metal4 19880 39312 19880 39312 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.S4BEG3
rlabel metal2 7336 4480 7336 4480 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W1BEG0
rlabel metal2 10304 18200 10304 18200 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W1BEG1
rlabel metal2 5208 5768 5208 5768 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W1BEG2
rlabel metal3 19880 4312 19880 4312 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W1BEG3
rlabel metal3 5880 3752 5880 3752 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG0
rlabel metal2 12712 15512 12712 15512 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG1
rlabel metal3 2296 27384 2296 27384 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG2
rlabel metal2 1848 2352 1848 2352 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG3
rlabel metal2 9128 4424 9128 4424 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG4
rlabel metal2 896 2184 896 2184 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG5
rlabel metal4 3304 8792 3304 8792 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG6
rlabel metal2 4088 6720 4088 6720 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEG7
rlabel metal2 3864 1288 3864 1288 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb0
rlabel metal3 3752 2744 3752 2744 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb1
rlabel metal3 3976 12824 3976 12824 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb2
rlabel metal3 5880 8792 5880 8792 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb3
rlabel metal3 8400 5768 8400 5768 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb4
rlabel metal2 5712 17976 5712 17976 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb5
rlabel metal2 2408 5880 2408 5880 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb6
rlabel metal2 5432 5488 5432 5488 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W2BEGb7
rlabel metal2 19096 6720 19096 6720 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG0
rlabel metal2 1736 46984 1736 46984 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG1
rlabel metal2 8120 22232 8120 22232 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG10
rlabel metal3 8904 15176 8904 15176 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG11
rlabel metal3 3136 50792 3136 50792 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG2
rlabel metal2 15400 14896 15400 14896 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG3
rlabel metal3 19320 17752 19320 17752 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG4
rlabel metal2 2520 36960 2520 36960 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG5
rlabel metal2 5992 19656 5992 19656 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG6
rlabel metal3 12264 16184 12264 16184 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG7
rlabel metal3 17416 15624 17416 15624 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG8
rlabel metal3 2912 33432 2912 33432 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.W6BEG9
rlabel metal2 18760 4200 18760 4200 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG0
rlabel metal2 2520 27048 2520 27048 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG1
rlabel metal2 6048 15960 6048 15960 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG10
rlabel metal4 2184 8512 2184 8512 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG11
rlabel metal2 17808 16072 17808 16072 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG12
rlabel metal3 4144 35000 4144 35000 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG13
rlabel metal3 5376 15176 5376 15176 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG14
rlabel metal2 9352 14336 9352 14336 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG15
rlabel metal3 4480 25256 4480 25256 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG2
rlabel metal2 12600 8736 12600 8736 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG3
rlabel metal2 21672 8064 21672 8064 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG4
rlabel metal3 1792 33656 1792 33656 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG5
rlabel metal2 2072 13216 2072 13216 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG6
rlabel metal2 12040 10696 12040 10696 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG7
rlabel metal3 18312 11592 18312 11592 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG8
rlabel metal4 2968 21336 2968 21336 0 Tile_X0Y1_GF_SRAM_bot.Inst_GF_SRAM_bot_switch_matrix.WW4BEG9
rlabel metal2 5432 238 5432 238 0 Tile_X0Y1_N1END[0]
rlabel metal2 5656 518 5656 518 0 Tile_X0Y1_N1END[1]
rlabel metal2 5880 350 5880 350 0 Tile_X0Y1_N1END[2]
rlabel metal2 6104 854 6104 854 0 Tile_X0Y1_N1END[3]
rlabel metal2 8120 1414 8120 1414 0 Tile_X0Y1_N2END[0]
rlabel metal2 8344 854 8344 854 0 Tile_X0Y1_N2END[1]
rlabel metal2 8568 854 8568 854 0 Tile_X0Y1_N2END[2]
rlabel metal2 8792 854 8792 854 0 Tile_X0Y1_N2END[3]
rlabel metal2 9016 742 9016 742 0 Tile_X0Y1_N2END[4]
rlabel metal2 9240 910 9240 910 0 Tile_X0Y1_N2END[5]
rlabel metal2 9464 518 9464 518 0 Tile_X0Y1_N2END[6]
rlabel metal2 9688 854 9688 854 0 Tile_X0Y1_N2END[7]
rlabel metal2 6328 798 6328 798 0 Tile_X0Y1_N2MID[0]
rlabel metal2 6552 854 6552 854 0 Tile_X0Y1_N2MID[1]
rlabel metal2 6776 854 6776 854 0 Tile_X0Y1_N2MID[2]
rlabel metal2 7000 854 7000 854 0 Tile_X0Y1_N2MID[3]
rlabel metal2 7224 182 7224 182 0 Tile_X0Y1_N2MID[4]
rlabel metal2 7448 854 7448 854 0 Tile_X0Y1_N2MID[5]
rlabel metal2 7672 854 7672 854 0 Tile_X0Y1_N2MID[6]
rlabel metal2 7896 854 7896 854 0 Tile_X0Y1_N2MID[7]
rlabel metal2 9968 2408 9968 2408 0 Tile_X0Y1_N4END[0]
rlabel metal2 12152 854 12152 854 0 Tile_X0Y1_N4END[10]
rlabel metal2 12376 854 12376 854 0 Tile_X0Y1_N4END[11]
rlabel metal2 12600 854 12600 854 0 Tile_X0Y1_N4END[12]
rlabel metal2 12824 854 12824 854 0 Tile_X0Y1_N4END[13]
rlabel metal2 13048 854 13048 854 0 Tile_X0Y1_N4END[14]
rlabel metal2 13272 854 13272 854 0 Tile_X0Y1_N4END[15]
rlabel metal2 10136 854 10136 854 0 Tile_X0Y1_N4END[1]
rlabel metal2 10360 854 10360 854 0 Tile_X0Y1_N4END[2]
rlabel metal2 10584 294 10584 294 0 Tile_X0Y1_N4END[3]
rlabel metal2 10808 350 10808 350 0 Tile_X0Y1_N4END[4]
rlabel metal2 7336 87472 7336 87472 0 Tile_X0Y1_N4END[5]
rlabel metal2 11256 854 11256 854 0 Tile_X0Y1_N4END[6]
rlabel metal2 22680 60704 22680 60704 0 Tile_X0Y1_N4END[7]
rlabel metal2 11704 798 11704 798 0 Tile_X0Y1_N4END[8]
rlabel metal2 11928 854 11928 854 0 Tile_X0Y1_N4END[9]
rlabel metal2 13496 1246 13496 1246 0 Tile_X0Y1_S1BEG[0]
rlabel metal2 13720 1302 13720 1302 0 Tile_X0Y1_S1BEG[1]
rlabel metal2 13944 686 13944 686 0 Tile_X0Y1_S1BEG[2]
rlabel metal2 14168 1302 14168 1302 0 Tile_X0Y1_S1BEG[3]
rlabel metal2 14392 910 14392 910 0 Tile_X0Y1_S2BEG[0]
rlabel metal2 5208 840 5208 840 0 Tile_X0Y1_S2BEG[1]
rlabel metal2 14840 238 14840 238 0 Tile_X0Y1_S2BEG[2]
rlabel metal2 5880 896 5880 896 0 Tile_X0Y1_S2BEG[3]
rlabel metal2 8344 2240 8344 2240 0 Tile_X0Y1_S2BEG[4]
rlabel metal2 9576 1904 9576 1904 0 Tile_X0Y1_S2BEG[5]
rlabel metal2 12264 1568 12264 1568 0 Tile_X0Y1_S2BEG[6]
rlabel metal2 15960 910 15960 910 0 Tile_X0Y1_S2BEG[7]
rlabel metal2 16184 462 16184 462 0 Tile_X0Y1_S2BEGb[0]
rlabel metal2 16408 518 16408 518 0 Tile_X0Y1_S2BEGb[1]
rlabel metal2 16632 406 16632 406 0 Tile_X0Y1_S2BEGb[2]
rlabel metal2 16856 686 16856 686 0 Tile_X0Y1_S2BEGb[3]
rlabel metal2 17080 294 17080 294 0 Tile_X0Y1_S2BEGb[4]
rlabel metal2 17304 518 17304 518 0 Tile_X0Y1_S2BEGb[5]
rlabel metal2 17528 574 17528 574 0 Tile_X0Y1_S2BEGb[6]
rlabel metal2 17752 126 17752 126 0 Tile_X0Y1_S2BEGb[7]
rlabel metal2 27720 1176 27720 1176 0 Tile_X0Y1_S4BEG[0]
rlabel metal2 20216 406 20216 406 0 Tile_X0Y1_S4BEG[10]
rlabel metal2 20440 910 20440 910 0 Tile_X0Y1_S4BEG[11]
rlabel metal2 29064 616 29064 616 0 Tile_X0Y1_S4BEG[12]
rlabel metal2 27160 2240 27160 2240 0 Tile_X0Y1_S4BEG[13]
rlabel metal2 28168 1904 28168 1904 0 Tile_X0Y1_S4BEG[14]
rlabel metal2 21336 350 21336 350 0 Tile_X0Y1_S4BEG[15]
rlabel metal2 18200 462 18200 462 0 Tile_X0Y1_S4BEG[1]
rlabel metal3 27636 1064 27636 1064 0 Tile_X0Y1_S4BEG[2]
rlabel metal2 18648 1190 18648 1190 0 Tile_X0Y1_S4BEG[3]
rlabel metal3 20272 3976 20272 3976 0 Tile_X0Y1_S4BEG[4]
rlabel metal2 19096 1022 19096 1022 0 Tile_X0Y1_S4BEG[5]
rlabel metal2 19320 686 19320 686 0 Tile_X0Y1_S4BEG[6]
rlabel metal2 19544 686 19544 686 0 Tile_X0Y1_S4BEG[7]
rlabel metal2 27496 1288 27496 1288 0 Tile_X0Y1_S4BEG[8]
rlabel metal2 19992 182 19992 182 0 Tile_X0Y1_S4BEG[9]
rlabel metal3 22176 61208 22176 61208 0 Tile_X0Y1_UserCLK
rlabel metal3 854 280 854 280 0 Tile_X0Y1_W1BEG[0]
rlabel metal3 518 728 518 728 0 Tile_X0Y1_W1BEG[1]
rlabel metal3 1414 1176 1414 1176 0 Tile_X0Y1_W1BEG[2]
rlabel metal3 406 1624 406 1624 0 Tile_X0Y1_W1BEG[3]
rlabel metal3 1526 2072 1526 2072 0 Tile_X0Y1_W2BEG[0]
rlabel metal3 854 2520 854 2520 0 Tile_X0Y1_W2BEG[1]
rlabel metal3 1302 2968 1302 2968 0 Tile_X0Y1_W2BEG[2]
rlabel metal4 6328 8456 6328 8456 0 Tile_X0Y1_W2BEG[3]
rlabel metal3 910 3864 910 3864 0 Tile_X0Y1_W2BEG[4]
rlabel metal3 630 4312 630 4312 0 Tile_X0Y1_W2BEG[5]
rlabel metal3 1722 4760 1722 4760 0 Tile_X0Y1_W2BEG[6]
rlabel metal2 5880 6048 5880 6048 0 Tile_X0Y1_W2BEG[7]
rlabel metal3 182 5656 182 5656 0 Tile_X0Y1_W2BEGb[0]
rlabel metal2 8904 6440 8904 6440 0 Tile_X0Y1_W2BEGb[1]
rlabel metal3 6608 5208 6608 5208 0 Tile_X0Y1_W2BEGb[2]
rlabel metal2 2520 2240 2520 2240 0 Tile_X0Y1_W2BEGb[3]
rlabel metal2 6664 7168 6664 7168 0 Tile_X0Y1_W2BEGb[4]
rlabel metal3 1722 7896 1722 7896 0 Tile_X0Y1_W2BEGb[5]
rlabel metal3 3710 8344 3710 8344 0 Tile_X0Y1_W2BEGb[6]
rlabel metal2 6664 8232 6664 8232 0 Tile_X0Y1_W2BEGb[7]
rlabel metal3 1722 16408 1722 16408 0 Tile_X0Y1_W6BEG[0]
rlabel metal3 854 20888 854 20888 0 Tile_X0Y1_W6BEG[10]
rlabel metal3 574 21336 574 21336 0 Tile_X0Y1_W6BEG[11]
rlabel metal2 4760 16296 4760 16296 0 Tile_X0Y1_W6BEG[1]
rlabel metal3 1638 17304 1638 17304 0 Tile_X0Y1_W6BEG[2]
rlabel metal2 3976 16912 3976 16912 0 Tile_X0Y1_W6BEG[3]
rlabel metal3 2534 18200 2534 18200 0 Tile_X0Y1_W6BEG[4]
rlabel metal2 5544 18984 5544 18984 0 Tile_X0Y1_W6BEG[5]
rlabel metal2 3976 18480 3976 18480 0 Tile_X0Y1_W6BEG[6]
rlabel metal2 3304 16856 3304 16856 0 Tile_X0Y1_W6BEG[7]
rlabel metal3 1722 19992 1722 19992 0 Tile_X0Y1_W6BEG[8]
rlabel metal3 518 20440 518 20440 0 Tile_X0Y1_W6BEG[9]
rlabel metal2 1792 3752 1792 3752 0 Tile_X0Y1_WW4BEG[0]
rlabel metal3 910 13720 910 13720 0 Tile_X0Y1_WW4BEG[10]
rlabel metal2 4984 12152 4984 12152 0 Tile_X0Y1_WW4BEG[11]
rlabel metal2 1008 8344 1008 8344 0 Tile_X0Y1_WW4BEG[12]
rlabel metal2 1736 10640 1736 10640 0 Tile_X0Y1_WW4BEG[13]
rlabel metal3 574 15512 574 15512 0 Tile_X0Y1_WW4BEG[14]
rlabel metal2 4984 13944 4984 13944 0 Tile_X0Y1_WW4BEG[15]
rlabel metal2 4928 7336 4928 7336 0 Tile_X0Y1_WW4BEG[1]
rlabel metal2 1008 3752 1008 3752 0 Tile_X0Y1_WW4BEG[2]
rlabel metal2 7672 10528 7672 10528 0 Tile_X0Y1_WW4BEG[3]
rlabel metal3 2184 4200 2184 4200 0 Tile_X0Y1_WW4BEG[4]
rlabel metal3 3934 11480 3934 11480 0 Tile_X0Y1_WW4BEG[5]
rlabel metal3 728 4200 728 4200 0 Tile_X0Y1_WW4BEG[6]
rlabel metal3 2408 12488 2408 12488 0 Tile_X0Y1_WW4BEG[7]
rlabel metal3 784 5320 784 5320 0 Tile_X0Y1_WW4BEG[8]
rlabel metal2 1064 6944 1064 6944 0 Tile_X0Y1_WW4BEG[9]
rlabel metal3 31122 12824 31122 12824 0 WEN_SRAM0
rlabel metal3 31122 13720 31122 13720 0 WEN_SRAM1
rlabel metal3 31178 14616 31178 14616 0 WEN_SRAM2
rlabel metal3 31122 15512 31122 15512 0 WEN_SRAM3
rlabel metal3 31122 16408 31122 16408 0 WEN_SRAM4
rlabel metal3 31122 17304 31122 17304 0 WEN_SRAM5
rlabel metal3 31122 18200 31122 18200 0 WEN_SRAM6
rlabel metal3 31122 19096 31122 19096 0 WEN_SRAM7
rlabel metal2 3192 25368 3192 25368 0 _0000_
rlabel metal2 2632 21168 2632 21168 0 _0001_
rlabel metal3 19264 25256 19264 25256 0 _0002_
rlabel metal2 15736 29064 15736 29064 0 _0003_
rlabel metal3 2408 19208 2408 19208 0 _0004_
rlabel metal2 2968 46872 2968 46872 0 _0005_
rlabel metal2 17808 21560 17808 21560 0 _0006_
rlabel metal3 18984 98392 18984 98392 0 _0007_
rlabel metal3 17808 97496 17808 97496 0 _0008_
rlabel metal2 19152 97832 19152 97832 0 _0009_
rlabel metal2 16072 98448 16072 98448 0 _0010_
rlabel metal4 15736 66472 15736 66472 0 _0011_
rlabel metal2 15624 25760 15624 25760 0 _0012_
rlabel metal3 15176 23128 15176 23128 0 _0013_
rlabel metal2 13832 19432 13832 19432 0 _0014_
rlabel metal2 14280 22344 14280 22344 0 _0015_
rlabel metal3 14056 22568 14056 22568 0 _0016_
rlabel metal2 13496 21560 13496 21560 0 _0017_
rlabel metal2 16128 23352 16128 23352 0 _0018_
rlabel metal3 16576 25480 16576 25480 0 _0019_
rlabel metal2 17752 25984 17752 25984 0 _0020_
rlabel metal2 16968 25648 16968 25648 0 _0021_
rlabel metal2 16856 67984 16856 67984 0 _0022_
rlabel metal2 2968 74480 2968 74480 0 _0023_
rlabel metal2 11032 94248 11032 94248 0 _0024_
rlabel metal3 12488 67928 12488 67928 0 _0025_
rlabel metal2 16072 62216 16072 62216 0 _0026_
rlabel metal3 16352 61320 16352 61320 0 _0027_
rlabel metal2 15400 61768 15400 61768 0 _0028_
rlabel metal2 10696 72800 10696 72800 0 _0029_
rlabel metal3 9912 72520 9912 72520 0 _0030_
rlabel metal3 8960 74088 8960 74088 0 _0031_
rlabel metal2 11144 78848 11144 78848 0 _0032_
rlabel metal3 11872 78568 11872 78568 0 _0033_
rlabel metal2 11928 79128 11928 79128 0 _0034_
rlabel metal2 14448 79800 14448 79800 0 _0035_
rlabel metal2 14840 80528 14840 80528 0 _0036_
rlabel metal2 15344 80472 15344 80472 0 _0037_
rlabel metal2 22960 85848 22960 85848 0 _0038_
rlabel metal3 23128 86072 23128 86072 0 _0039_
rlabel metal2 13944 90160 13944 90160 0 _0040_
rlabel metal2 13944 92008 13944 92008 0 _0041_
rlabel metal2 10024 100016 10024 100016 0 _0042_
rlabel metal2 10920 99344 10920 99344 0 _0043_
rlabel metal2 3304 109368 3304 109368 0 _0044_
rlabel metal2 3304 108136 3304 108136 0 _0045_
rlabel metal3 20048 85288 20048 85288 0 _0046_
rlabel metal2 21672 84336 21672 84336 0 _0047_
rlabel metal3 17584 84168 17584 84168 0 _0048_
rlabel metal3 17080 84952 17080 84952 0 _0049_
rlabel metal2 12040 95760 12040 95760 0 _0050_
rlabel metal3 12208 96264 12208 96264 0 _0051_
rlabel metal3 5376 92904 5376 92904 0 _0052_
rlabel metal2 4872 96152 4872 96152 0 _0053_
rlabel metal2 21168 77112 21168 77112 0 _0054_
rlabel metal2 21672 78344 21672 78344 0 _0055_
rlabel metal2 18200 89768 18200 89768 0 _0056_
rlabel metal2 16632 90384 16632 90384 0 _0057_
rlabel metal2 9912 93688 9912 93688 0 _0058_
rlabel metal2 9184 92008 9184 92008 0 _0059_
rlabel metal2 2352 89768 2352 89768 0 _0060_
rlabel metal2 1624 91448 1624 91448 0 _0061_
rlabel metal2 21672 92344 21672 92344 0 _0062_
rlabel metal2 20832 94584 20832 94584 0 _0063_
rlabel metal2 20216 90608 20216 90608 0 _0064_
rlabel metal2 16632 92960 16632 92960 0 _0065_
rlabel metal2 15512 93912 15512 93912 0 _0066_
rlabel metal2 9128 94976 9128 94976 0 _0067_
rlabel metal2 3192 90104 3192 90104 0 _0068_
rlabel metal2 2072 94640 2072 94640 0 _0069_
rlabel metal2 22344 91784 22344 91784 0 _0070_
rlabel metal2 20776 91728 20776 91728 0 _0071_
rlabel metal2 18984 17808 18984 17808 0 _0072_
rlabel metal3 4144 41160 4144 41160 0 _0073_
rlabel metal2 5208 25928 5208 25928 0 _0074_
rlabel metal2 11872 25368 11872 25368 0 _0075_
rlabel metal2 22288 21000 22288 21000 0 _0076_
rlabel metal2 3080 47712 3080 47712 0 _0077_
rlabel metal3 7224 26600 7224 26600 0 _0078_
rlabel metal2 11032 22792 11032 22792 0 _0079_
rlabel metal2 21224 21392 21224 21392 0 _0080_
rlabel metal2 21784 22288 21784 22288 0 _0081_
rlabel metal3 21000 19432 21000 19432 0 _0082_
rlabel metal2 16184 21560 16184 21560 0 _0083_
rlabel metal2 18088 19544 18088 19544 0 _0084_
rlabel metal2 16968 18144 16968 18144 0 _0085_
rlabel metal2 16296 20608 16296 20608 0 _0086_
rlabel metal2 17528 20664 17528 20664 0 _0087_
rlabel metal2 17080 22680 17080 22680 0 _0088_
rlabel metal2 22232 25088 22232 25088 0 _0089_
rlabel metal3 21280 24808 21280 24808 0 _0090_
rlabel metal2 21448 25368 21448 25368 0 _0091_
rlabel metal2 15512 28280 15512 28280 0 _0092_
rlabel metal2 12824 30632 12824 30632 0 _0093_
rlabel metal2 11200 52360 11200 52360 0 _0094_
rlabel metal2 10080 51240 10080 51240 0 _0095_
rlabel metal2 5880 41720 5880 41720 0 _0096_
rlabel metal3 7784 41720 7784 41720 0 _0097_
rlabel metal2 18872 43456 18872 43456 0 _0098_
rlabel metal2 19096 42784 19096 42784 0 _0099_
rlabel metal2 17640 27888 17640 27888 0 _0100_
rlabel metal3 16072 27160 16072 27160 0 _0101_
rlabel metal3 12040 36568 12040 36568 0 _0102_
rlabel metal2 13720 33208 13720 33208 0 _0103_
rlabel metal2 3752 49056 3752 49056 0 _0104_
rlabel metal2 3304 48104 3304 48104 0 _0105_
rlabel metal3 20664 41832 20664 41832 0 _0106_
rlabel metal2 21672 40376 21672 40376 0 _0107_
rlabel metal3 18256 35000 18256 35000 0 _0108_
rlabel metal3 18200 34888 18200 34888 0 _0109_
rlabel metal2 18200 35896 18200 35896 0 _0110_
rlabel metal3 17024 33432 17024 33432 0 _0111_
rlabel metal2 19320 33488 19320 33488 0 _0112_
rlabel metal2 19656 33488 19656 33488 0 _0113_
rlabel metal2 20552 33936 20552 33936 0 _0114_
rlabel metal2 18312 32368 18312 32368 0 _0115_
rlabel metal3 18256 31528 18256 31528 0 _0116_
rlabel metal2 19544 32704 19544 32704 0 _0117_
rlabel metal2 17080 34384 17080 34384 0 _0118_
rlabel metal2 17640 32480 17640 32480 0 _0119_
rlabel metal2 18312 31640 18312 31640 0 _0120_
rlabel metal2 21224 33432 21224 33432 0 _0121_
rlabel metal2 29624 32928 29624 32928 0 _0122_
rlabel metal2 8120 25480 8120 25480 0 _0123_
rlabel metal2 7560 24640 7560 24640 0 _0124_
rlabel metal2 9800 35728 9800 35728 0 _0125_
rlabel metal3 7616 35000 7616 35000 0 _0126_
rlabel metal2 2968 45584 2968 45584 0 _0127_
rlabel metal2 2184 44520 2184 44520 0 _0128_
rlabel metal2 25480 35168 25480 35168 0 _0129_
rlabel metal2 21840 35112 21840 35112 0 _0130_
rlabel metal3 10808 27160 10808 27160 0 _0131_
rlabel metal3 10528 24920 10528 24920 0 _0132_
rlabel metal2 7448 37352 7448 37352 0 _0133_
rlabel metal3 6832 39144 6832 39144 0 _0134_
rlabel metal2 2968 42448 2968 42448 0 _0135_
rlabel metal3 3640 41720 3640 41720 0 _0136_
rlabel metal2 22008 34048 22008 34048 0 _0137_
rlabel metal2 21840 33544 21840 33544 0 _0138_
rlabel metal2 17528 33096 17528 33096 0 _0139_
rlabel metal3 16632 31752 16632 31752 0 _0140_
rlabel via2 19320 27272 19320 27272 0 _0141_
rlabel metal2 18984 33152 18984 33152 0 _0142_
rlabel metal3 22232 28056 22232 28056 0 _0143_
rlabel metal3 25368 27832 25368 27832 0 _0144_
rlabel metal2 12712 103320 12712 103320 0 _0145_
rlabel metal2 5152 92344 5152 92344 0 _0146_
rlabel metal2 23464 68824 23464 68824 0 _0147_
rlabel metal2 23744 85848 23744 85848 0 _0148_
rlabel metal3 16800 61768 16800 61768 0 _0149_
rlabel metal3 9576 73192 9576 73192 0 _0150_
rlabel metal2 12264 80248 12264 80248 0 _0151_
rlabel metal2 15176 80248 15176 80248 0 _0152_
rlabel metal4 23128 86016 23128 86016 0 _0153_
rlabel metal2 14056 25872 14056 25872 0 _0154_
rlabel metal3 19096 98168 19096 98168 0 _0155_
rlabel metal2 15064 20888 15064 20888 0 _0156_
rlabel metal3 10696 48104 10696 48104 0 _0157_
rlabel metal2 9688 44912 9688 44912 0 _0158_
rlabel metal3 23632 22904 23632 22904 0 _0159_
rlabel metal2 20664 20272 20664 20272 0 _0160_
rlabel metal2 17640 20496 17640 20496 0 _0161_
rlabel metal2 16408 20160 16408 20160 0 _0162_
rlabel metal2 22288 25704 22288 25704 0 _0163_
rlabel metal2 16072 35448 16072 35448 0 _0164_
rlabel metal2 9800 2632 9800 2632 0 _0165_
rlabel metal2 17920 29288 17920 29288 0 _0166_
rlabel metal3 16464 30408 16464 30408 0 _0167_
rlabel metal2 19208 26936 19208 26936 0 _0168_
rlabel metal3 17920 31080 17920 31080 0 _0169_
rlabel metal2 20328 30296 20328 30296 0 _0170_
rlabel metal2 20888 31024 20888 31024 0 _0171_
rlabel metal2 20888 28112 20888 28112 0 _0172_
rlabel metal2 20720 29624 20720 29624 0 _0173_
rlabel metal2 21392 27832 21392 27832 0 _0174_
rlabel metal2 18648 26880 18648 26880 0 _0175_
rlabel metal3 21952 29400 21952 29400 0 _0176_
rlabel metal2 19712 28728 19712 28728 0 _0177_
rlabel metal2 21896 29960 21896 29960 0 _0178_
rlabel metal2 21672 28280 21672 28280 0 _0179_
rlabel metal2 11592 103936 11592 103936 0 _0180_
rlabel metal2 12320 104104 12320 104104 0 _0181_
rlabel metal4 11704 104216 11704 104216 0 _0182_
rlabel metal2 10360 100800 10360 100800 0 _0183_
rlabel metal3 9688 45752 9688 45752 0 _0184_
rlabel metal3 7560 31864 7560 31864 0 _0185_
rlabel metal2 12264 48272 12264 48272 0 _0186_
rlabel metal3 12376 48104 12376 48104 0 _0187_
rlabel metal2 13496 47880 13496 47880 0 _0188_
rlabel metal2 13888 47992 13888 47992 0 _0189_
rlabel metal3 6720 92232 6720 92232 0 _0190_
rlabel metal2 7336 96264 7336 96264 0 _0191_
rlabel metal2 7784 96152 7784 96152 0 _0192_
rlabel metal2 6216 100632 6216 100632 0 _0193_
rlabel metal3 5376 44968 5376 44968 0 _0194_
rlabel metal2 7560 46816 7560 46816 0 _0195_
rlabel metal2 9744 45192 9744 45192 0 _0196_
rlabel metal2 9464 45024 9464 45024 0 _0197_
rlabel metal2 5880 45248 5880 45248 0 _0198_
rlabel metal3 9912 46088 9912 46088 0 _0199_
rlabel metal2 24808 68880 24808 68880 0 _0200_
rlabel metal2 24248 68768 24248 68768 0 _0201_
rlabel metal3 22400 68600 22400 68600 0 _0202_
rlabel metal2 24360 68768 24360 68768 0 _0203_
rlabel metal2 24248 22568 24248 22568 0 _0204_
rlabel metal2 19768 20664 19768 20664 0 _0205_
rlabel metal2 23128 23240 23128 23240 0 _0206_
rlabel metal2 23800 23128 23800 23128 0 _0207_
rlabel metal2 23464 22848 23464 22848 0 _0208_
rlabel metal2 20552 22904 20552 22904 0 _0209_
rlabel metal3 28056 55272 28056 55272 0 clknet_0_Tile_X0Y1_UserCLK
rlabel metal3 24248 55160 24248 55160 0 clknet_1_0__leaf_Tile_X0Y1_UserCLK
rlabel metal3 22624 94248 22624 94248 0 clknet_1_1__leaf_Tile_X0Y1_UserCLK
rlabel metal3 25928 20776 25928 20776 0 net1
rlabel metal3 29176 11592 29176 11592 0 net10
rlabel metal3 10416 109256 10416 109256 0 net100
rlabel metal2 10864 109928 10864 109928 0 net101
rlabel metal2 9576 108864 9576 108864 0 net102
rlabel metal2 9184 105448 9184 105448 0 net103
rlabel metal2 9912 107464 9912 107464 0 net104
rlabel metal3 6720 110376 6720 110376 0 net105
rlabel metal2 11144 110824 11144 110824 0 net106
rlabel metal2 10248 111272 10248 111272 0 net107
rlabel metal2 20944 110712 20944 110712 0 net108
rlabel metal2 22904 112616 22904 112616 0 net109
rlabel metal2 30296 36120 30296 36120 0 net11
rlabel metal2 13944 57960 13944 57960 0 net110
rlabel metal2 11592 59360 11592 59360 0 net111
rlabel metal3 1624 58968 1624 58968 0 net112
rlabel metal2 16744 58856 16744 58856 0 net113
rlabel metal3 1624 60536 1624 60536 0 net114
rlabel metal3 1624 61656 1624 61656 0 net115
rlabel metal2 1288 63616 1288 63616 0 net116
rlabel metal2 1400 58016 1400 58016 0 net117
rlabel metal2 1288 64792 1288 64792 0 net118
rlabel metal2 1736 64400 1736 64400 0 net119
rlabel metal3 24584 28728 24584 28728 0 net12
rlabel metal2 1624 65352 1624 65352 0 net120
rlabel metal3 1624 68040 1624 68040 0 net121
rlabel metal2 4984 62328 4984 62328 0 net122
rlabel metal2 5992 65632 5992 65632 0 net123
rlabel metal2 1848 67088 1848 67088 0 net124
rlabel metal3 6328 65464 6328 65464 0 net125
rlabel metal3 6664 63336 6664 63336 0 net126
rlabel metal2 4256 66472 4256 66472 0 net127
rlabel metal2 3304 70392 3304 70392 0 net128
rlabel metal3 1232 66920 1232 66920 0 net129
rlabel metal2 30240 29400 30240 29400 0 net13
rlabel metal3 12152 74312 12152 74312 0 net130
rlabel metal2 2184 84952 2184 84952 0 net131
rlabel metal2 13496 77224 13496 77224 0 net132
rlabel metal2 8120 75488 8120 75488 0 net133
rlabel metal4 1624 95032 1624 95032 0 net134
rlabel metal2 14504 71008 14504 71008 0 net135
rlabel metal4 17416 77560 17416 77560 0 net136
rlabel metal3 3920 77784 3920 77784 0 net137
rlabel metal2 1344 83720 1344 83720 0 net138
rlabel metal2 11704 76608 11704 76608 0 net139
rlabel metal2 26040 35000 26040 35000 0 net14
rlabel metal2 20104 77560 20104 77560 0 net140
rlabel metal2 8344 82208 8344 82208 0 net141
rlabel metal2 17416 63840 17416 63840 0 net142
rlabel metal3 5096 75096 5096 75096 0 net143
rlabel metal2 13888 71624 13888 71624 0 net144
rlabel metal2 20608 73192 20608 73192 0 net145
rlabel metal2 4200 78064 4200 78064 0 net146
rlabel metal2 5376 74872 5376 74872 0 net147
rlabel metal2 11872 73192 11872 73192 0 net148
rlabel metal2 1456 75656 1456 75656 0 net149
rlabel metal2 30408 31920 30408 31920 0 net15
rlabel metal2 2184 73304 2184 73304 0 net150
rlabel metal3 1344 76216 1344 76216 0 net151
rlabel metal2 15848 68824 15848 68824 0 net152
rlabel metal2 4312 70280 4312 70280 0 net153
rlabel metal2 1288 74704 1288 74704 0 net154
rlabel metal3 10080 69608 10080 69608 0 net155
rlabel metal2 19768 71988 19768 71988 0 net156
rlabel metal2 2072 75208 2072 75208 0 net157
rlabel metal2 29848 40320 29848 40320 0 net158
rlabel metal3 23800 51128 23800 51128 0 net159
rlabel metal2 30240 31976 30240 31976 0 net16
rlabel metal2 30296 52472 30296 52472 0 net160
rlabel metal2 30408 53200 30408 53200 0 net161
rlabel metal2 30184 53872 30184 53872 0 net162
rlabel metal2 21784 53760 21784 53760 0 net163
rlabel metal2 30464 55496 30464 55496 0 net164
rlabel metal2 21336 56000 21336 56000 0 net165
rlabel metal2 29904 57512 29904 57512 0 net166
rlabel metal2 29848 59080 29848 59080 0 net167
rlabel metal2 29904 60200 29904 60200 0 net168
rlabel metal2 30072 41272 30072 41272 0 net169
rlabel metal2 30464 33320 30464 33320 0 net17
rlabel metal2 29848 61096 29848 61096 0 net170
rlabel metal2 29848 62216 29848 62216 0 net171
rlabel metal2 29904 63336 29904 63336 0 net172
rlabel metal2 29848 65016 29848 65016 0 net173
rlabel metal2 30408 65912 30408 65912 0 net174
rlabel metal2 30296 67424 30296 67424 0 net175
rlabel metal2 29904 68040 29904 68040 0 net176
rlabel metal2 29848 69720 29848 69720 0 net177
rlabel metal2 30408 69468 30408 69468 0 net178
rlabel metal2 29848 71848 29848 71848 0 net179
rlabel metal2 30296 34216 30296 34216 0 net18
rlabel metal2 29848 42280 29848 42280 0 net180
rlabel metal2 23464 72856 23464 72856 0 net181
rlabel metal2 23352 73920 23352 73920 0 net182
rlabel metal2 30072 43288 30072 43288 0 net183
rlabel metal2 29904 44520 29904 44520 0 net184
rlabel metal2 29848 45416 29848 45416 0 net185
rlabel metal2 22680 46760 22680 46760 0 net186
rlabel metal2 23576 47264 23576 47264 0 net187
rlabel metal2 30296 48608 30296 48608 0 net188
rlabel metal2 30408 49840 30408 49840 0 net189
rlabel metal3 29176 35112 29176 35112 0 net19
rlabel metal2 8120 4424 8120 4424 0 net190
rlabel metal2 11928 4928 11928 4928 0 net191
rlabel metal2 10976 4200 10976 4200 0 net192
rlabel metal2 19432 6048 19432 6048 0 net193
rlabel metal2 12264 6496 12264 6496 0 net194
rlabel metal3 9576 1120 9576 1120 0 net195
rlabel metal2 9352 1848 9352 1848 0 net196
rlabel metal2 5656 1232 5656 1232 0 net197
rlabel metal2 8008 2520 8008 2520 0 net198
rlabel metal2 9240 2464 9240 2464 0 net199
rlabel metal2 30184 21000 30184 21000 0 net2
rlabel metal3 30016 25032 30016 25032 0 net20
rlabel metal2 12600 2632 12600 2632 0 net200
rlabel metal2 15848 4424 15848 4424 0 net201
rlabel metal2 15512 2408 15512 2408 0 net202
rlabel metal3 16016 952 16016 952 0 net203
rlabel metal3 16632 2072 16632 2072 0 net204
rlabel metal2 19656 2856 19656 2856 0 net205
rlabel metal2 14728 1848 14728 1848 0 net206
rlabel metal2 23352 2268 23352 2268 0 net207
rlabel metal2 16016 2632 16016 2632 0 net208
rlabel metal2 27272 952 27272 952 0 net209
rlabel metal2 29848 78344 29848 78344 0 net21
rlabel metal4 28056 55160 28056 55160 0 net210
rlabel metal3 22344 96152 22344 96152 0 net211
rlabel metal2 25088 5208 25088 5208 0 net212
rlabel metal2 29288 3416 29288 3416 0 net213
rlabel metal2 27384 3808 27384 3808 0 net214
rlabel metal2 28504 2744 28504 2744 0 net215
rlabel metal3 24920 3864 24920 3864 0 net216
rlabel metal2 21728 110712 21728 110712 0 net217
rlabel metal2 28616 1288 28616 1288 0 net218
rlabel metal2 27048 9856 27048 9856 0 net219
rlabel metal3 21448 89880 21448 89880 0 net22
rlabel metal3 23464 107576 23464 107576 0 net220
rlabel metal2 22344 110880 22344 110880 0 net221
rlabel metal4 22232 59920 22232 59920 0 net222
rlabel metal4 23296 109890 23296 109890 0 net223
rlabel metal2 27832 8680 27832 8680 0 net224
rlabel metal3 23240 94192 23240 94192 0 net225
rlabel metal2 16072 10304 16072 10304 0 net226
rlabel metal2 17080 7392 17080 7392 0 net227
rlabel metal3 5992 4200 5992 4200 0 net228
rlabel metal2 18984 4536 18984 4536 0 net229
rlabel metal2 30296 90888 30296 90888 0 net23
rlabel metal2 14952 10416 14952 10416 0 net230
rlabel metal2 12768 10472 12768 10472 0 net231
rlabel metal3 10696 12152 10696 12152 0 net232
rlabel metal2 2184 2016 2184 2016 0 net233
rlabel metal2 15512 8568 15512 8568 0 net234
rlabel metal2 1512 2772 1512 2772 0 net235
rlabel metal2 6160 4200 6160 4200 0 net236
rlabel metal2 8344 8344 8344 8344 0 net237
rlabel metal2 4200 1120 4200 1120 0 net238
rlabel metal2 4200 2856 4200 2856 0 net239
rlabel metal3 24920 91896 24920 91896 0 net24
rlabel metal3 6216 5320 6216 5320 0 net240
rlabel metal2 2576 1960 2576 1960 0 net241
rlabel metal3 7168 6776 7168 6776 0 net242
rlabel metal2 5992 7784 5992 7784 0 net243
rlabel metal3 3920 5320 3920 5320 0 net244
rlabel metal2 5992 6384 5992 6384 0 net245
rlabel metal2 15624 16604 15624 16604 0 net246
rlabel metal2 2072 22176 2072 22176 0 net247
rlabel metal2 1512 18144 1512 18144 0 net248
rlabel metal4 1960 34832 1960 34832 0 net249
rlabel metal2 30296 93296 30296 93296 0 net25
rlabel metal3 1176 50680 1176 50680 0 net250
rlabel metal2 15064 16184 15064 16184 0 net251
rlabel metal2 18312 17584 18312 17584 0 net252
rlabel metal2 1848 30520 1848 30520 0 net253
rlabel metal2 1624 18872 1624 18872 0 net254
rlabel metal3 7448 16184 7448 16184 0 net255
rlabel metal2 16688 16296 16688 16296 0 net256
rlabel metal3 1624 32200 1624 32200 0 net257
rlabel metal2 18424 4648 18424 4648 0 net258
rlabel metal2 4200 10864 4200 10864 0 net259
rlabel metal2 30408 94864 30408 94864 0 net26
rlabel metal2 2408 6720 2408 6720 0 net260
rlabel metal2 17416 15848 17416 15848 0 net261
rlabel metal2 2072 10080 2072 10080 0 net262
rlabel metal2 1400 12152 1400 12152 0 net263
rlabel metal2 5320 13832 5320 13832 0 net264
rlabel metal2 5376 7448 5376 7448 0 net265
rlabel metal2 1512 6104 1512 6104 0 net266
rlabel metal2 10360 10192 10360 10192 0 net267
rlabel metal2 2072 4368 2072 4368 0 net268
rlabel metal2 1736 6608 1736 6608 0 net269
rlabel metal2 30296 94864 30296 94864 0 net27
rlabel metal3 1680 4312 1680 4312 0 net270
rlabel metal4 2072 7448 2072 7448 0 net271
rlabel metal3 2408 12320 2408 12320 0 net272
rlabel metal2 1288 7224 1288 7224 0 net273
rlabel metal2 19208 16016 19208 16016 0 net274
rlabel metal3 19768 14952 19768 14952 0 net275
rlabel metal2 30464 25256 30464 25256 0 net276
rlabel metal3 28112 16296 28112 16296 0 net277
rlabel metal3 26488 16632 26488 16632 0 net278
rlabel metal3 29064 17864 29064 17864 0 net279
rlabel metal2 29848 96432 29848 96432 0 net28
rlabel metal3 27664 18424 27664 18424 0 net280
rlabel metal3 29120 19432 29120 19432 0 net281
rlabel metal2 30072 97720 30072 97720 0 net29
rlabel metal2 17640 22736 17640 22736 0 net3
rlabel metal3 24808 99288 24808 99288 0 net30
rlabel metal2 17640 100296 17640 100296 0 net31
rlabel metal2 30072 79352 30072 79352 0 net32
rlabel metal2 29848 100800 29848 100800 0 net33
rlabel metal3 23968 102424 23968 102424 0 net34
rlabel metal3 24920 102872 24920 102872 0 net35
rlabel metal2 30296 104272 30296 104272 0 net36
rlabel metal3 24864 105560 24864 105560 0 net37
rlabel metal2 29848 106568 29848 106568 0 net38
rlabel metal2 30408 108248 30408 108248 0 net39
rlabel metal2 30296 23240 30296 23240 0 net4
rlabel metal2 30072 108696 30072 108696 0 net40
rlabel metal2 29848 109704 29848 109704 0 net41
rlabel metal2 29848 110880 29848 110880 0 net42
rlabel metal2 29848 80752 29848 80752 0 net43
rlabel metal2 30296 111664 30296 111664 0 net44
rlabel metal2 29624 111440 29624 111440 0 net45
rlabel metal2 30072 82040 30072 82040 0 net46
rlabel metal2 30296 83048 30296 83048 0 net47
rlabel metal2 23688 83888 23688 83888 0 net48
rlabel metal3 27104 85176 27104 85176 0 net49
rlabel metal3 22848 24024 22848 24024 0 net5
rlabel metal2 30296 86184 30296 86184 0 net50
rlabel metal2 23240 87360 23240 87360 0 net51
rlabel metal2 29848 88592 29848 88592 0 net52
rlabel metal2 22064 110376 22064 110376 0 net53
rlabel metal2 24920 112112 24920 112112 0 net54
rlabel metal2 26600 112616 26600 112616 0 net55
rlabel metal2 27944 112336 27944 112336 0 net56
rlabel metal2 29512 111776 29512 111776 0 net57
rlabel metal3 27440 111832 27440 111832 0 net58
rlabel metal2 27832 111384 27832 111384 0 net59
rlabel metal3 29344 24696 29344 24696 0 net6
rlabel metal2 26824 111272 26824 111272 0 net60
rlabel metal3 28728 111944 28728 111944 0 net61
rlabel metal3 27160 110264 27160 110264 0 net62
rlabel metal2 27496 111440 27496 111440 0 net63
rlabel metal3 23128 110376 23128 110376 0 net64
rlabel metal2 22176 110264 22176 110264 0 net65
rlabel metal3 24136 109928 24136 109928 0 net66
rlabel metal2 23912 87416 23912 87416 0 net67
rlabel metal2 26320 111272 26320 111272 0 net68
rlabel metal2 23688 110936 23688 110936 0 net69
rlabel metal3 25200 25704 25200 25704 0 net7
rlabel metal2 27048 113064 27048 113064 0 net70
rlabel metal2 26936 110880 26936 110880 0 net71
rlabel metal2 28616 112392 28616 112392 0 net72
rlabel metal2 12264 110544 12264 110544 0 net73
rlabel metal2 5208 101696 5208 101696 0 net74
rlabel metal2 22960 111160 22960 111160 0 net75
rlabel metal2 21000 105280 21000 105280 0 net76
rlabel metal2 1288 107240 1288 107240 0 net77
rlabel metal3 5488 102872 5488 102872 0 net78
rlabel metal2 3752 103152 3752 103152 0 net79
rlabel metal2 30072 27272 30072 27272 0 net8
rlabel metal2 1176 110880 1176 110880 0 net80
rlabel metal2 2296 112280 2296 112280 0 net81
rlabel metal2 4088 104664 4088 104664 0 net82
rlabel metal2 3528 105896 3528 105896 0 net83
rlabel metal3 6216 109928 6216 109928 0 net84
rlabel metal2 3416 112336 3416 112336 0 net85
rlabel metal3 5264 107800 5264 107800 0 net86
rlabel metal3 24248 112504 24248 112504 0 net87
rlabel metal3 14392 107688 14392 107688 0 net88
rlabel metal2 19880 112112 19880 112112 0 net89
rlabel metal2 30296 27888 30296 27888 0 net9
rlabel metal2 22400 112280 22400 112280 0 net90
rlabel metal3 12768 109928 12768 109928 0 net91
rlabel metal2 18928 110376 18928 110376 0 net92
rlabel metal2 23184 113288 23184 113288 0 net93
rlabel metal2 15624 113064 15624 113064 0 net94
rlabel metal3 16576 46536 16576 46536 0 net95
rlabel metal2 19544 113232 19544 113232 0 net96
rlabel metal2 21560 110600 21560 110600 0 net97
rlabel metal2 10584 108864 10584 108864 0 net98
rlabel metal2 20664 111160 20664 111160 0 net99
<< properties >>
string FIXED_BBOX 0 0 31696 114912
<< end >>
