module W_IO4 (A_I_top,
    A_O_top,
    A_T_top,
    A_config_C_bit0,
    A_config_C_bit1,
    A_config_C_bit2,
    A_config_C_bit3,
    B_I_top,
    B_O_top,
    B_T_top,
    B_config_C_bit0,
    B_config_C_bit1,
    B_config_C_bit2,
    B_config_C_bit3,
    C_I_top,
    C_O_top,
    C_T_top,
    C_config_C_bit0,
    C_config_C_bit1,
    C_config_C_bit2,
    C_config_C_bit3,
    D_I_top,
    D_O_top,
    D_T_top,
    D_config_C_bit0,
    D_config_C_bit1,
    D_config_C_bit2,
    D_config_C_bit3,
    UserCLK,
    UserCLKo,
    E1BEG,
    E2BEG,
    E2BEGb,
    E6BEG,
    EE4BEG,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    W1END,
    W2END,
    W2MID,
    W6END,
    WW4END);
 output A_I_top;
 input A_O_top;
 output A_T_top;
 output A_config_C_bit0;
 output A_config_C_bit1;
 output A_config_C_bit2;
 output A_config_C_bit3;
 output B_I_top;
 input B_O_top;
 output B_T_top;
 output B_config_C_bit0;
 output B_config_C_bit1;
 output B_config_C_bit2;
 output B_config_C_bit3;
 output C_I_top;
 input C_O_top;
 output C_T_top;
 output C_config_C_bit0;
 output C_config_C_bit1;
 output C_config_C_bit2;
 output C_config_C_bit3;
 output D_I_top;
 input D_O_top;
 output D_T_top;
 output D_config_C_bit0;
 output D_config_C_bit1;
 output D_config_C_bit2;
 output D_config_C_bit3;
 input UserCLK;
 output UserCLKo;
 output [3:0] E1BEG;
 output [7:0] E2BEG;
 output [7:0] E2BEGb;
 output [11:0] E6BEG;
 output [15:0] EE4BEG;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 input [3:0] W1END;
 input [7:0] W2END;
 input [7:0] W2MID;
 input [11:0] W6END;
 input [15:0] WW4END;

 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire \Inst_A_IO_1_bidirectional_frame_config_pass.Q ;
 wire \Inst_B_IO_1_bidirectional_frame_config_pass.Q ;
 wire \Inst_C_IO_1_bidirectional_frame_config_pass.Q ;
 wire \Inst_D_IO_1_bidirectional_frame_config_pass.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame3_bit10.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame3_bit11.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame3_bit12.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame3_bit13.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame3_bit14.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame3_bit15.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame3_bit16.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame3_bit17.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame3_bit18.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame3_bit19.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame3_bit20.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame3_bit21.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame3_bit4.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame3_bit5.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame3_bit6.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame3_bit7.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame3_bit8.Q ;
 wire \Inst_W_IO4_ConfigMem.Inst_frame3_bit9.Q ;
 wire \Inst_W_IO4_switch_matrix.E1BEG0 ;
 wire \Inst_W_IO4_switch_matrix.E1BEG1 ;
 wire \Inst_W_IO4_switch_matrix.E1BEG2 ;
 wire \Inst_W_IO4_switch_matrix.E1BEG3 ;
 wire \Inst_W_IO4_switch_matrix.E2BEG0 ;
 wire \Inst_W_IO4_switch_matrix.E2BEG1 ;
 wire \Inst_W_IO4_switch_matrix.E2BEG2 ;
 wire \Inst_W_IO4_switch_matrix.E2BEG3 ;
 wire \Inst_W_IO4_switch_matrix.E2BEG4 ;
 wire \Inst_W_IO4_switch_matrix.E2BEG5 ;
 wire \Inst_W_IO4_switch_matrix.E2BEG6 ;
 wire \Inst_W_IO4_switch_matrix.E2BEG7 ;
 wire \Inst_W_IO4_switch_matrix.E2BEGb0 ;
 wire \Inst_W_IO4_switch_matrix.E2BEGb1 ;
 wire \Inst_W_IO4_switch_matrix.E2BEGb2 ;
 wire \Inst_W_IO4_switch_matrix.E2BEGb3 ;
 wire \Inst_W_IO4_switch_matrix.E2BEGb4 ;
 wire \Inst_W_IO4_switch_matrix.E2BEGb5 ;
 wire \Inst_W_IO4_switch_matrix.E2BEGb6 ;
 wire \Inst_W_IO4_switch_matrix.E2BEGb7 ;
 wire \Inst_W_IO4_switch_matrix.E6BEG0 ;
 wire \Inst_W_IO4_switch_matrix.E6BEG1 ;
 wire \Inst_W_IO4_switch_matrix.E6BEG10 ;
 wire \Inst_W_IO4_switch_matrix.E6BEG11 ;
 wire \Inst_W_IO4_switch_matrix.E6BEG2 ;
 wire \Inst_W_IO4_switch_matrix.E6BEG3 ;
 wire \Inst_W_IO4_switch_matrix.E6BEG4 ;
 wire \Inst_W_IO4_switch_matrix.E6BEG5 ;
 wire \Inst_W_IO4_switch_matrix.E6BEG6 ;
 wire \Inst_W_IO4_switch_matrix.E6BEG7 ;
 wire \Inst_W_IO4_switch_matrix.E6BEG8 ;
 wire \Inst_W_IO4_switch_matrix.E6BEG9 ;
 wire \Inst_W_IO4_switch_matrix.EE4BEG0 ;
 wire \Inst_W_IO4_switch_matrix.EE4BEG1 ;
 wire \Inst_W_IO4_switch_matrix.EE4BEG10 ;
 wire \Inst_W_IO4_switch_matrix.EE4BEG11 ;
 wire \Inst_W_IO4_switch_matrix.EE4BEG12 ;
 wire \Inst_W_IO4_switch_matrix.EE4BEG13 ;
 wire \Inst_W_IO4_switch_matrix.EE4BEG14 ;
 wire \Inst_W_IO4_switch_matrix.EE4BEG15 ;
 wire \Inst_W_IO4_switch_matrix.EE4BEG2 ;
 wire \Inst_W_IO4_switch_matrix.EE4BEG3 ;
 wire \Inst_W_IO4_switch_matrix.EE4BEG4 ;
 wire \Inst_W_IO4_switch_matrix.EE4BEG5 ;
 wire \Inst_W_IO4_switch_matrix.EE4BEG6 ;
 wire \Inst_W_IO4_switch_matrix.EE4BEG7 ;
 wire \Inst_W_IO4_switch_matrix.EE4BEG8 ;
 wire \Inst_W_IO4_switch_matrix.EE4BEG9 ;
 wire net143;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net144;
 wire net145;
 wire UserCLK_regs;
 wire clknet_0_UserCLK;
 wire clknet_1_0__leaf_UserCLK;
 wire clknet_0_UserCLK_regs;
 wire clknet_1_0__leaf_UserCLK_regs;
 wire clknet_1_1__leaf_UserCLK_regs;

 gf180mcu_fd_sc_mcu7t5v0__inv_1 _078_ (.I(W2MID[5]),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _079_ (.I(W2MID[7]),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _080_ (.I(W2END[0]),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _081_ (.I(W2END[1]),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _082_ (.I(\Inst_W_IO4_ConfigMem.Inst_frame0_bit9.Q ),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _083_ (.I(\Inst_W_IO4_ConfigMem.Inst_frame0_bit16.Q ),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _084_ (.I(\Inst_W_IO4_ConfigMem.Inst_frame0_bit23.Q ),
    .ZN(_006_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _085_ (.I(\Inst_W_IO4_ConfigMem.Inst_frame0_bit30.Q ),
    .ZN(_007_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _086_ (.I(\Inst_W_IO4_ConfigMem.Inst_frame0_bit27.Q ),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _087_ (.I(\Inst_W_IO4_ConfigMem.Inst_frame0_bit20.Q ),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _088_ (.I(\Inst_W_IO4_ConfigMem.Inst_frame0_bit13.Q ),
    .ZN(_010_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _089_ (.I(\Inst_W_IO4_ConfigMem.Inst_frame0_bit6.Q ),
    .ZN(_011_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _090_ (.I0(W2MID[5]),
    .I1(WW4END[5]),
    .I2(WW4END[13]),
    .I3(W6END[5]),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame3_bit16.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame3_bit17.Q ),
    .Z(\Inst_W_IO4_switch_matrix.E2BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _091_ (.I0(W2MID[6]),
    .I1(WW4END[6]),
    .I2(WW4END[14]),
    .I3(W6END[6]),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame3_bit14.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame3_bit15.Q ),
    .Z(\Inst_W_IO4_switch_matrix.E2BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _092_ (.I0(W2MID[7]),
    .I1(WW4END[7]),
    .I2(WW4END[15]),
    .I3(W6END[7]),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame3_bit12.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame3_bit13.Q ),
    .Z(\Inst_W_IO4_switch_matrix.E2BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _093_ (.I0(W1END[0]),
    .I1(W1END[3]),
    .I2(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .I3(\Inst_D_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame3_bit10.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame3_bit11.Q ),
    .Z(\Inst_W_IO4_switch_matrix.E1BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _094_ (.I0(W1END[0]),
    .I1(W1END[1]),
    .I2(B_O_top),
    .I3(D_O_top),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame3_bit8.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame3_bit9.Q ),
    .Z(\Inst_W_IO4_switch_matrix.E1BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _095_ (.I0(W1END[1]),
    .I1(W1END[2]),
    .I2(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .I3(\Inst_C_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame3_bit6.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame3_bit7.Q ),
    .Z(\Inst_W_IO4_switch_matrix.E1BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _096_ (.I0(W1END[2]),
    .I1(A_O_top),
    .I2(W1END[3]),
    .I3(C_O_top),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame3_bit5.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame3_bit4.Q ),
    .Z(\Inst_W_IO4_switch_matrix.E1BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _097_ (.A1(W2MID[7]),
    .A2(\Inst_W_IO4_ConfigMem.Inst_frame0_bit9.Q ),
    .ZN(_012_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _098_ (.A1(_003_),
    .A2(\Inst_W_IO4_ConfigMem.Inst_frame0_bit9.Q ),
    .B(\Inst_W_IO4_ConfigMem.Inst_frame0_bit10.Q ),
    .C(_012_),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _099_ (.A1(_004_),
    .A2(W2END[3]),
    .A3(\Inst_W_IO4_ConfigMem.Inst_frame0_bit10.Q ),
    .Z(_014_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _100_ (.A1(_002_),
    .A2(\Inst_W_IO4_ConfigMem.Inst_frame0_bit9.Q ),
    .A3(\Inst_W_IO4_ConfigMem.Inst_frame0_bit10.Q ),
    .ZN(_015_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _101_ (.A1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit9.Q ),
    .A2(W2END[4]),
    .B(\Inst_W_IO4_ConfigMem.Inst_frame0_bit10.Q ),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _102_ (.A1(W2END[2]),
    .A2(\Inst_W_IO4_ConfigMem.Inst_frame0_bit9.Q ),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _103_ (.A1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit8.Q ),
    .A2(_016_),
    .A3(_017_),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _104_ (.A1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit8.Q ),
    .A2(_013_),
    .A3(_014_),
    .B1(_015_),
    .B2(_018_),
    .ZN(net2));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _105_ (.A1(W2MID[6]),
    .A2(\Inst_W_IO4_ConfigMem.Inst_frame0_bit16.Q ),
    .ZN(_019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _106_ (.A1(_002_),
    .A2(\Inst_W_IO4_ConfigMem.Inst_frame0_bit16.Q ),
    .B(\Inst_W_IO4_ConfigMem.Inst_frame0_bit17.Q ),
    .C(_019_),
    .ZN(_020_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _107_ (.A1(_005_),
    .A2(W2END[5]),
    .A3(\Inst_W_IO4_ConfigMem.Inst_frame0_bit17.Q ),
    .Z(_021_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _108_ (.A1(_001_),
    .A2(\Inst_W_IO4_ConfigMem.Inst_frame0_bit16.Q ),
    .A3(\Inst_W_IO4_ConfigMem.Inst_frame0_bit17.Q ),
    .ZN(_022_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _109_ (.A1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit16.Q ),
    .A2(W2END[6]),
    .B(\Inst_W_IO4_ConfigMem.Inst_frame0_bit17.Q ),
    .ZN(_023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _110_ (.A1(W2END[4]),
    .A2(\Inst_W_IO4_ConfigMem.Inst_frame0_bit16.Q ),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _111_ (.A1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit15.Q ),
    .A2(_023_),
    .A3(_024_),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _112_ (.A1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit15.Q ),
    .A2(_020_),
    .A3(_021_),
    .B1(_022_),
    .B2(_025_),
    .ZN(net8));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _113_ (.A1(W2MID[7]),
    .A2(\Inst_W_IO4_ConfigMem.Inst_frame0_bit23.Q ),
    .ZN(_026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _114_ (.A1(_003_),
    .A2(\Inst_W_IO4_ConfigMem.Inst_frame0_bit23.Q ),
    .B(\Inst_W_IO4_ConfigMem.Inst_frame0_bit24.Q ),
    .C(_026_),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _115_ (.A1(W2END[3]),
    .A2(_006_),
    .A3(\Inst_W_IO4_ConfigMem.Inst_frame0_bit24.Q ),
    .Z(_028_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _116_ (.A1(_002_),
    .A2(\Inst_W_IO4_ConfigMem.Inst_frame0_bit23.Q ),
    .A3(\Inst_W_IO4_ConfigMem.Inst_frame0_bit24.Q ),
    .ZN(_029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _117_ (.A1(W2END[4]),
    .A2(\Inst_W_IO4_ConfigMem.Inst_frame0_bit23.Q ),
    .B(\Inst_W_IO4_ConfigMem.Inst_frame0_bit24.Q ),
    .ZN(_030_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _118_ (.A1(W2END[2]),
    .A2(\Inst_W_IO4_ConfigMem.Inst_frame0_bit23.Q ),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _119_ (.A1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit22.Q ),
    .A2(_030_),
    .A3(_031_),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _120_ (.A1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit22.Q ),
    .A2(_027_),
    .A3(_028_),
    .B1(_029_),
    .B2(_032_),
    .ZN(net14));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _121_ (.A1(W2MID[6]),
    .A2(\Inst_W_IO4_ConfigMem.Inst_frame0_bit30.Q ),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _122_ (.A1(_002_),
    .A2(\Inst_W_IO4_ConfigMem.Inst_frame0_bit30.Q ),
    .B(\Inst_W_IO4_ConfigMem.Inst_frame0_bit31.Q ),
    .C(_033_),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _123_ (.A1(W2END[5]),
    .A2(_007_),
    .A3(\Inst_W_IO4_ConfigMem.Inst_frame0_bit31.Q ),
    .Z(_035_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _124_ (.A1(_001_),
    .A2(\Inst_W_IO4_ConfigMem.Inst_frame0_bit30.Q ),
    .A3(\Inst_W_IO4_ConfigMem.Inst_frame0_bit31.Q ),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _125_ (.A1(W2END[6]),
    .A2(\Inst_W_IO4_ConfigMem.Inst_frame0_bit30.Q ),
    .B(\Inst_W_IO4_ConfigMem.Inst_frame0_bit31.Q ),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _126_ (.A1(W2END[4]),
    .A2(\Inst_W_IO4_ConfigMem.Inst_frame0_bit30.Q ),
    .ZN(_038_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _127_ (.A1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit29.Q ),
    .A2(_037_),
    .A3(_038_),
    .ZN(_039_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _128_ (.A1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit29.Q ),
    .A2(_034_),
    .A3(_035_),
    .B1(_036_),
    .B2(_039_),
    .ZN(net20));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _129_ (.I0(W2END[0]),
    .I1(W2END[2]),
    .I2(W2END[1]),
    .I3(W2END[3]),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame0_bit26.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit25.Q ),
    .Z(_040_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _130_ (.A1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit27.Q ),
    .A2(_040_),
    .ZN(_041_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _131_ (.I0(W2END[4]),
    .I1(W2END[5]),
    .I2(W2END[6]),
    .I3(W2END[7]),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame0_bit25.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit26.Q ),
    .Z(_042_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _132_ (.A1(_008_),
    .A2(_042_),
    .B(\Inst_W_IO4_ConfigMem.Inst_frame0_bit28.Q ),
    .ZN(_043_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _133_ (.I0(W2MID[0]),
    .I1(W2MID[1]),
    .I2(W2MID[2]),
    .I3(W2MID[3]),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame0_bit25.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit26.Q ),
    .Z(_044_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _134_ (.A1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit27.Q ),
    .A2(_044_),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _135_ (.I0(W2MID[6]),
    .I1(W2MID[7]),
    .S(\Inst_W_IO4_ConfigMem.Inst_frame0_bit25.Q ),
    .Z(_046_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _136_ (.A1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit25.Q ),
    .A2(W2MID[4]),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _137_ (.A1(_000_),
    .A2(\Inst_W_IO4_ConfigMem.Inst_frame0_bit25.Q ),
    .B(\Inst_W_IO4_ConfigMem.Inst_frame0_bit26.Q ),
    .C(_047_),
    .ZN(_048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _138_ (.A1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit26.Q ),
    .A2(_046_),
    .B(_048_),
    .C(_008_),
    .ZN(_049_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _139_ (.A1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit28.Q ),
    .A2(_045_),
    .A3(_049_),
    .B1(_041_),
    .B2(_043_),
    .ZN(net19));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _140_ (.I0(W2END[0]),
    .I1(W2END[2]),
    .I2(W2END[1]),
    .I3(W2END[3]),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame0_bit19.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit18.Q ),
    .Z(_050_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _141_ (.A1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit20.Q ),
    .A2(_050_),
    .ZN(_051_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _142_ (.I0(W2END[4]),
    .I1(W2END[5]),
    .I2(W2END[6]),
    .I3(W2END[7]),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame0_bit18.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit19.Q ),
    .Z(_052_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _143_ (.A1(_009_),
    .A2(_052_),
    .B(\Inst_W_IO4_ConfigMem.Inst_frame0_bit21.Q ),
    .ZN(_053_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _144_ (.I0(W2MID[4]),
    .I1(W2MID[6]),
    .I2(W2MID[5]),
    .I3(W2MID[7]),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame0_bit19.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit18.Q ),
    .Z(_054_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _145_ (.A1(_009_),
    .A2(_054_),
    .ZN(_055_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _146_ (.I0(W2MID[0]),
    .I1(W2MID[1]),
    .I2(W2MID[2]),
    .I3(W2MID[3]),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame0_bit18.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit19.Q ),
    .Z(_056_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _147_ (.A1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit20.Q ),
    .A2(_056_),
    .ZN(_057_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _148_ (.A1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit21.Q ),
    .A2(_055_),
    .A3(_057_),
    .B1(_051_),
    .B2(_053_),
    .ZN(net13));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _149_ (.I0(W2END[0]),
    .I1(W2END[2]),
    .I2(W2END[1]),
    .I3(W2END[3]),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame0_bit12.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit11.Q ),
    .Z(_058_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _150_ (.A1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit13.Q ),
    .A2(_058_),
    .ZN(_059_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _151_ (.I0(W2END[4]),
    .I1(W2END[5]),
    .I2(W2END[6]),
    .I3(W2END[7]),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame0_bit11.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit12.Q ),
    .Z(_060_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _152_ (.A1(_010_),
    .A2(_060_),
    .B(\Inst_W_IO4_ConfigMem.Inst_frame0_bit14.Q ),
    .ZN(_061_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _153_ (.I0(W2MID[0]),
    .I1(W2MID[1]),
    .I2(W2MID[2]),
    .I3(W2MID[3]),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame0_bit11.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit12.Q ),
    .Z(_062_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _154_ (.A1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit13.Q ),
    .A2(_062_),
    .ZN(_063_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _155_ (.I0(W2MID[6]),
    .I1(W2MID[7]),
    .S(\Inst_W_IO4_ConfigMem.Inst_frame0_bit11.Q ),
    .Z(_064_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _156_ (.A1(W2MID[4]),
    .A2(\Inst_W_IO4_ConfigMem.Inst_frame0_bit11.Q ),
    .ZN(_065_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _157_ (.A1(_000_),
    .A2(\Inst_W_IO4_ConfigMem.Inst_frame0_bit11.Q ),
    .B(\Inst_W_IO4_ConfigMem.Inst_frame0_bit12.Q ),
    .C(_065_),
    .ZN(_066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _158_ (.A1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit12.Q ),
    .A2(_064_),
    .B(_066_),
    .C(_010_),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _159_ (.A1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit14.Q ),
    .A2(_063_),
    .A3(_067_),
    .B1(_059_),
    .B2(_061_),
    .ZN(net7));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _160_ (.I0(W2END[0]),
    .I1(W2END[2]),
    .I2(W2END[1]),
    .I3(W2END[3]),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame0_bit5.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit4.Q ),
    .Z(_068_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _161_ (.A1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit6.Q ),
    .A2(_068_),
    .ZN(_069_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _162_ (.I0(W2END[4]),
    .I1(W2END[5]),
    .I2(W2END[6]),
    .I3(W2END[7]),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame0_bit4.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit5.Q ),
    .Z(_070_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _163_ (.A1(_011_),
    .A2(_070_),
    .B(\Inst_W_IO4_ConfigMem.Inst_frame0_bit7.Q ),
    .ZN(_071_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _164_ (.I0(W2MID[0]),
    .I1(W2MID[1]),
    .I2(W2MID[2]),
    .I3(W2MID[3]),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame0_bit4.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit5.Q ),
    .Z(_072_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _165_ (.A1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit6.Q ),
    .A2(_072_),
    .ZN(_073_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _166_ (.I0(W2MID[6]),
    .I1(W2MID[7]),
    .S(\Inst_W_IO4_ConfigMem.Inst_frame0_bit4.Q ),
    .Z(_074_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _167_ (.A1(W2MID[4]),
    .A2(\Inst_W_IO4_ConfigMem.Inst_frame0_bit4.Q ),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _168_ (.A1(_000_),
    .A2(\Inst_W_IO4_ConfigMem.Inst_frame0_bit4.Q ),
    .B(\Inst_W_IO4_ConfigMem.Inst_frame0_bit5.Q ),
    .C(_075_),
    .ZN(_076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _169_ (.A1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit5.Q ),
    .A2(_074_),
    .B(_076_),
    .C(_011_),
    .ZN(_077_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _170_ (.A1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit7.Q ),
    .A2(_073_),
    .A3(_077_),
    .B1(_069_),
    .B2(_071_),
    .ZN(net1));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _171_ (.I0(W1END[0]),
    .I1(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .I2(WW4END[0]),
    .I3(\Inst_D_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame0_bit3.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit2.Q ),
    .Z(\Inst_W_IO4_switch_matrix.E6BEG11 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _172_ (.I0(W1END[1]),
    .I1(B_O_top),
    .I2(WW4END[1]),
    .I3(D_O_top),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame0_bit1.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame0_bit0.Q ),
    .Z(\Inst_W_IO4_switch_matrix.E6BEG10 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _173_ (.I0(WW4END[4]),
    .I1(WW4END[12]),
    .I2(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .I3(\Inst_D_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame1_bit30.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame1_bit31.Q ),
    .Z(\Inst_W_IO4_switch_matrix.E6BEG9 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _174_ (.I0(WW4END[5]),
    .I1(WW4END[13]),
    .I2(B_O_top),
    .I3(D_O_top),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame1_bit28.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame1_bit29.Q ),
    .Z(\Inst_W_IO4_switch_matrix.E6BEG8 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _175_ (.I0(W1END[0]),
    .I1(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .I2(WW4END[8]),
    .I3(\Inst_D_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame1_bit27.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame1_bit26.Q ),
    .Z(\Inst_W_IO4_switch_matrix.E6BEG7 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _176_ (.I0(W1END[1]),
    .I1(B_O_top),
    .I2(WW4END[9]),
    .I3(D_O_top),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame1_bit25.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame1_bit24.Q ),
    .Z(\Inst_W_IO4_switch_matrix.E6BEG6 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _177_ (.I0(W1END[3]),
    .I1(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .I2(WW4END[2]),
    .I3(\Inst_C_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame1_bit23.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame1_bit22.Q ),
    .Z(\Inst_W_IO4_switch_matrix.E6BEG5 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _178_ (.I0(W1END[2]),
    .I1(A_O_top),
    .I2(WW4END[3]),
    .I3(C_O_top),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame1_bit21.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame1_bit20.Q ),
    .Z(\Inst_W_IO4_switch_matrix.E6BEG4 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _179_ (.I0(WW4END[6]),
    .I1(WW4END[14]),
    .I2(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .I3(\Inst_C_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame1_bit18.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame1_bit19.Q ),
    .Z(\Inst_W_IO4_switch_matrix.E6BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _180_ (.I0(WW4END[7]),
    .I1(WW4END[15]),
    .I2(A_O_top),
    .I3(C_O_top),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame1_bit16.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame1_bit17.Q ),
    .Z(\Inst_W_IO4_switch_matrix.E6BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _181_ (.I0(W1END[3]),
    .I1(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .I2(WW4END[10]),
    .I3(\Inst_C_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame1_bit15.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame1_bit14.Q ),
    .Z(\Inst_W_IO4_switch_matrix.E6BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _182_ (.I0(W1END[2]),
    .I1(A_O_top),
    .I2(WW4END[11]),
    .I3(C_O_top),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame1_bit13.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame1_bit12.Q ),
    .Z(\Inst_W_IO4_switch_matrix.E6BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _183_ (.I0(W2MID[3]),
    .I1(W2MID[7]),
    .I2(W2MID[5]),
    .I3(\Inst_D_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame1_bit11.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame1_bit10.Q ),
    .Z(\Inst_W_IO4_switch_matrix.EE4BEG15 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _184_ (.I0(W2MID[2]),
    .I1(W2MID[4]),
    .I2(W2MID[6]),
    .I3(\Inst_C_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame1_bit8.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame1_bit9.Q ),
    .Z(\Inst_W_IO4_switch_matrix.EE4BEG14 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _185_ (.I0(W6END[7]),
    .I1(W6END[9]),
    .I2(W6END[11]),
    .I3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame1_bit6.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame1_bit7.Q ),
    .Z(\Inst_W_IO4_switch_matrix.EE4BEG13 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _186_ (.I0(W6END[1]),
    .I1(W6END[3]),
    .I2(W6END[5]),
    .I3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame1_bit4.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame1_bit5.Q ),
    .Z(\Inst_W_IO4_switch_matrix.EE4BEG12 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _187_ (.I0(W6END[6]),
    .I1(W6END[8]),
    .I2(W6END[10]),
    .I3(B_O_top),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame1_bit2.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame1_bit3.Q ),
    .Z(\Inst_W_IO4_switch_matrix.EE4BEG11 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _188_ (.I0(W6END[0]),
    .I1(W6END[2]),
    .I2(W6END[4]),
    .I3(A_O_top),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame1_bit0.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame1_bit1.Q ),
    .Z(\Inst_W_IO4_switch_matrix.EE4BEG10 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _189_ (.I0(W6END[3]),
    .I1(W6END[7]),
    .I2(W6END[5]),
    .I3(D_O_top),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame2_bit31.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame2_bit30.Q ),
    .Z(\Inst_W_IO4_switch_matrix.EE4BEG9 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _190_ (.I0(W6END[6]),
    .I1(W6END[8]),
    .I2(W6END[10]),
    .I3(C_O_top),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame2_bit28.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame2_bit29.Q ),
    .Z(\Inst_W_IO4_switch_matrix.EE4BEG8 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _191_ (.I0(W2MID[3]),
    .I1(W2MID[7]),
    .I2(W2MID[5]),
    .I3(\Inst_D_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame2_bit27.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame2_bit26.Q ),
    .Z(\Inst_W_IO4_switch_matrix.EE4BEG7 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _192_ (.I0(W2MID[2]),
    .I1(W2MID[4]),
    .I2(W2MID[6]),
    .I3(\Inst_C_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame2_bit24.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame2_bit25.Q ),
    .Z(\Inst_W_IO4_switch_matrix.EE4BEG6 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _193_ (.I0(W2END[3]),
    .I1(W2END[5]),
    .I2(W2END[7]),
    .I3(D_O_top),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame2_bit22.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame2_bit23.Q ),
    .Z(\Inst_W_IO4_switch_matrix.EE4BEG5 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _194_ (.I0(W2END[2]),
    .I1(W2END[4]),
    .I2(W2END[6]),
    .I3(C_O_top),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame2_bit20.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame2_bit21.Q ),
    .Z(\Inst_W_IO4_switch_matrix.EE4BEG4 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _195_ (.I0(W6END[7]),
    .I1(W6END[9]),
    .I2(W6END[11]),
    .I3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame2_bit18.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame2_bit19.Q ),
    .Z(\Inst_W_IO4_switch_matrix.EE4BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _196_ (.I0(W6END[1]),
    .I1(W6END[3]),
    .I2(W6END[5]),
    .I3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame2_bit16.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame2_bit17.Q ),
    .Z(\Inst_W_IO4_switch_matrix.EE4BEG2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _197_ (.I0(W6END[6]),
    .I1(W6END[8]),
    .I2(W6END[10]),
    .I3(B_O_top),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame2_bit14.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame2_bit15.Q ),
    .Z(\Inst_W_IO4_switch_matrix.EE4BEG1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _198_ (.I0(W6END[0]),
    .I1(W6END[2]),
    .I2(W6END[4]),
    .I3(A_O_top),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame2_bit12.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame2_bit13.Q ),
    .Z(\Inst_W_IO4_switch_matrix.EE4BEG0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _199_ (.I0(W2END[0]),
    .I1(WW4END[0]),
    .I2(WW4END[8]),
    .I3(W6END[0]),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame2_bit10.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame2_bit11.Q ),
    .Z(\Inst_W_IO4_switch_matrix.E2BEGb7 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _200_ (.I0(W2END[1]),
    .I1(WW4END[1]),
    .I2(WW4END[9]),
    .I3(W6END[1]),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame2_bit8.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame2_bit9.Q ),
    .Z(\Inst_W_IO4_switch_matrix.E2BEGb6 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _201_ (.I0(W2END[2]),
    .I1(WW4END[2]),
    .I2(WW4END[10]),
    .I3(W6END[2]),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame2_bit6.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame2_bit7.Q ),
    .Z(\Inst_W_IO4_switch_matrix.E2BEGb5 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _202_ (.I0(W2END[3]),
    .I1(WW4END[3]),
    .I2(WW4END[11]),
    .I3(W6END[3]),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame2_bit4.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame2_bit5.Q ),
    .Z(\Inst_W_IO4_switch_matrix.E2BEGb4 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _203_ (.I0(W2END[4]),
    .I1(WW4END[4]),
    .I2(WW4END[12]),
    .I3(W6END[4]),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame2_bit2.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame2_bit3.Q ),
    .Z(\Inst_W_IO4_switch_matrix.E2BEGb3 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _204_ (.I0(W2END[5]),
    .I1(WW4END[13]),
    .I2(WW4END[5]),
    .I3(W6END[5]),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame2_bit1.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame2_bit0.Q ),
    .Z(\Inst_W_IO4_switch_matrix.E2BEGb2 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _205_ (.I0(W2END[6]),
    .I1(WW4END[14]),
    .I2(WW4END[6]),
    .I3(W6END[6]),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame3_bit31.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame3_bit30.Q ),
    .Z(\Inst_W_IO4_switch_matrix.E2BEGb1 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _206_ (.I0(W2END[7]),
    .I1(WW4END[15]),
    .I2(WW4END[7]),
    .I3(W6END[7]),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame3_bit29.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame3_bit28.Q ),
    .Z(\Inst_W_IO4_switch_matrix.E2BEGb0 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _207_ (.I0(W2MID[0]),
    .I1(WW4END[0]),
    .I2(WW4END[8]),
    .I3(W6END[0]),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame3_bit26.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame3_bit27.Q ),
    .Z(\Inst_W_IO4_switch_matrix.E2BEG7 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _208_ (.I0(W2MID[1]),
    .I1(WW4END[1]),
    .I2(WW4END[9]),
    .I3(W6END[1]),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame3_bit24.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame3_bit25.Q ),
    .Z(\Inst_W_IO4_switch_matrix.E2BEG6 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _209_ (.I0(W2MID[2]),
    .I1(WW4END[2]),
    .I2(WW4END[10]),
    .I3(W6END[2]),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame3_bit22.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame3_bit23.Q ),
    .Z(\Inst_W_IO4_switch_matrix.E2BEG5 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _210_ (.I0(W2MID[3]),
    .I1(WW4END[3]),
    .I2(WW4END[11]),
    .I3(W6END[3]),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame3_bit20.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame3_bit21.Q ),
    .Z(\Inst_W_IO4_switch_matrix.E2BEG4 ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _211_ (.I0(W2MID[4]),
    .I1(WW4END[4]),
    .I2(WW4END[12]),
    .I3(W6END[4]),
    .S0(\Inst_W_IO4_ConfigMem.Inst_frame3_bit18.Q ),
    .S1(\Inst_W_IO4_ConfigMem.Inst_frame3_bit19.Q ),
    .Z(\Inst_W_IO4_switch_matrix.E2BEG3 ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _212_ (.D(FrameData[20]),
    .E(net38),
    .Q(net3));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _213_ (.D(FrameData[21]),
    .E(net38),
    .Q(net4));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _214_ (.D(FrameData[22]),
    .E(net38),
    .Q(net5));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _215_ (.D(FrameData[23]),
    .E(net38),
    .Q(net6));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _216_ (.D(FrameData[24]),
    .E(net38),
    .Q(net9));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _217_ (.D(FrameData[25]),
    .E(net38),
    .Q(net10));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _218_ (.D(FrameData[26]),
    .E(net38),
    .Q(net11));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _219_ (.D(FrameData[27]),
    .E(net38),
    .Q(net12));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _220_ (.D(FrameData[28]),
    .E(FrameStrobe[4]),
    .Q(net15));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _221_ (.D(FrameData[29]),
    .E(FrameStrobe[4]),
    .Q(net16));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _222_ (.D(FrameData[30]),
    .E(FrameStrobe[4]),
    .Q(net17));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _223_ (.D(FrameData[31]),
    .E(net38),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _224_ (.D(FrameData[0]),
    .E(net41),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _225_ (.D(FrameData[1]),
    .E(net41),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _226_ (.D(FrameData[2]),
    .E(net41),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _227_ (.D(FrameData[3]),
    .E(net41),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _228_ (.D(FrameData[4]),
    .E(net42),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame3_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _229_ (.D(FrameData[5]),
    .E(net41),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame3_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _230_ (.D(FrameData[6]),
    .E(net42),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame3_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _231_ (.D(FrameData[7]),
    .E(net42),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame3_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _232_ (.D(FrameData[8]),
    .E(net41),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame3_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _233_ (.D(FrameData[9]),
    .E(net42),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame3_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _234_ (.D(FrameData[10]),
    .E(net41),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame3_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _235_ (.D(FrameData[11]),
    .E(net42),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame3_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _236_ (.D(FrameData[12]),
    .E(net39),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame3_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _237_ (.D(FrameData[13]),
    .E(net39),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame3_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _238_ (.D(FrameData[14]),
    .E(net39),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame3_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _239_ (.D(FrameData[15]),
    .E(net40),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame3_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _240_ (.D(FrameData[16]),
    .E(net40),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame3_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _241_ (.D(FrameData[17]),
    .E(net40),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame3_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _242_ (.D(FrameData[18]),
    .E(net39),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame3_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _243_ (.D(FrameData[19]),
    .E(net39),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame3_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _244_ (.D(FrameData[20]),
    .E(net40),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame3_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _245_ (.D(FrameData[21]),
    .E(net40),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame3_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _246_ (.D(FrameData[22]),
    .E(net39),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame3_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _247_ (.D(FrameData[23]),
    .E(net40),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame3_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _248_ (.D(FrameData[24]),
    .E(net39),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame3_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _249_ (.D(FrameData[25]),
    .E(net39),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame3_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _250_ (.D(FrameData[26]),
    .E(net39),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame3_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _251_ (.D(FrameData[27]),
    .E(net39),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame3_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _252_ (.D(FrameData[28]),
    .E(net40),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame3_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _253_ (.D(FrameData[29]),
    .E(net40),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame3_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _254_ (.D(FrameData[30]),
    .E(net41),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame3_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _255_ (.D(FrameData[31]),
    .E(net41),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame3_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _256_ (.D(FrameData[0]),
    .E(net46),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame2_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _257_ (.D(FrameData[1]),
    .E(net43),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame2_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _258_ (.D(FrameData[2]),
    .E(net44),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame2_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _259_ (.D(FrameData[3]),
    .E(net45),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame2_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _260_ (.D(FrameData[4]),
    .E(net46),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame2_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _261_ (.D(FrameData[5]),
    .E(net46),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame2_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _262_ (.D(FrameData[6]),
    .E(net45),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame2_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _263_ (.D(FrameData[7]),
    .E(net44),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame2_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _264_ (.D(FrameData[8]),
    .E(net43),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame2_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _265_ (.D(FrameData[9]),
    .E(net43),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame2_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _266_ (.D(FrameData[10]),
    .E(net43),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame2_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _267_ (.D(FrameData[11]),
    .E(net43),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame2_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _268_ (.D(FrameData[12]),
    .E(net44),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame2_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _269_ (.D(FrameData[13]),
    .E(net44),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame2_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _270_ (.D(FrameData[14]),
    .E(net44),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame2_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _271_ (.D(FrameData[15]),
    .E(net44),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame2_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _272_ (.D(FrameData[16]),
    .E(net45),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame2_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _273_ (.D(FrameData[17]),
    .E(net45),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame2_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _274_ (.D(FrameData[18]),
    .E(net45),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame2_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _275_ (.D(FrameData[19]),
    .E(net45),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame2_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _276_ (.D(FrameData[20]),
    .E(net44),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame2_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _277_ (.D(FrameData[21]),
    .E(net44),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame2_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _278_ (.D(FrameData[22]),
    .E(net43),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame2_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _279_ (.D(FrameData[23]),
    .E(net46),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame2_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _280_ (.D(FrameData[24]),
    .E(net43),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame2_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _281_ (.D(FrameData[25]),
    .E(net43),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame2_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _282_ (.D(FrameData[26]),
    .E(net43),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame2_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _283_ (.D(FrameData[27]),
    .E(net43),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame2_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _284_ (.D(FrameData[28]),
    .E(net44),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame2_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _285_ (.D(FrameData[29]),
    .E(net44),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame2_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _286_ (.D(FrameData[30]),
    .E(net45),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame2_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _287_ (.D(FrameData[31]),
    .E(net45),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame2_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _288_ (.D(FrameData[0]),
    .E(net48),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame1_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _289_ (.D(FrameData[1]),
    .E(net48),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame1_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _290_ (.D(FrameData[2]),
    .E(net49),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame1_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _291_ (.D(FrameData[3]),
    .E(net49),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame1_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _292_ (.D(FrameData[4]),
    .E(net49),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame1_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _293_ (.D(FrameData[5]),
    .E(net49),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame1_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _294_ (.D(FrameData[6]),
    .E(net49),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame1_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _295_ (.D(FrameData[7]),
    .E(net49),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame1_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _296_ (.D(FrameData[8]),
    .E(net47),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame1_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _297_ (.D(FrameData[9]),
    .E(net47),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame1_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _298_ (.D(FrameData[10]),
    .E(net47),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame1_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _299_ (.D(FrameData[11]),
    .E(net47),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame1_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _300_ (.D(FrameData[12]),
    .E(net50),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame1_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _301_ (.D(FrameData[13]),
    .E(net47),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame1_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _302_ (.D(FrameData[14]),
    .E(net48),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame1_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _303_ (.D(FrameData[15]),
    .E(net48),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame1_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _304_ (.D(FrameData[16]),
    .E(net47),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame1_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _305_ (.D(FrameData[17]),
    .E(net47),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame1_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _306_ (.D(FrameData[18]),
    .E(net48),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame1_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _307_ (.D(FrameData[19]),
    .E(net48),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame1_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _308_ (.D(FrameData[20]),
    .E(net50),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame1_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _309_ (.D(FrameData[21]),
    .E(net47),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame1_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _310_ (.D(FrameData[22]),
    .E(net48),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame1_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _311_ (.D(FrameData[23]),
    .E(net48),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame1_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _312_ (.D(FrameData[24]),
    .E(net49),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame1_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _313_ (.D(FrameData[25]),
    .E(net49),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame1_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _314_ (.D(FrameData[26]),
    .E(net49),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame1_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _315_ (.D(FrameData[27]),
    .E(net49),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame1_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _316_ (.D(FrameData[28]),
    .E(net47),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame1_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _317_ (.D(FrameData[29]),
    .E(net47),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame1_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _318_ (.D(FrameData[30]),
    .E(net48),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame1_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _319_ (.D(FrameData[31]),
    .E(net48),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame1_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _320_ (.D(FrameData[0]),
    .E(net55),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame0_bit0.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _321_ (.D(FrameData[1]),
    .E(net55),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame0_bit1.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _322_ (.D(FrameData[2]),
    .E(net55),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame0_bit2.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _323_ (.D(FrameData[3]),
    .E(net55),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame0_bit3.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _324_ (.D(FrameData[4]),
    .E(net51),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame0_bit4.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _325_ (.D(FrameData[5]),
    .E(net51),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame0_bit5.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _326_ (.D(FrameData[6]),
    .E(net54),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame0_bit6.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _327_ (.D(FrameData[7]),
    .E(net54),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame0_bit7.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _328_ (.D(FrameData[8]),
    .E(net52),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame0_bit8.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _329_ (.D(FrameData[9]),
    .E(net53),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame0_bit9.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _330_ (.D(FrameData[10]),
    .E(net53),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame0_bit10.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _331_ (.D(FrameData[11]),
    .E(net52),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame0_bit11.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _332_ (.D(FrameData[12]),
    .E(net52),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame0_bit12.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _333_ (.D(FrameData[13]),
    .E(net52),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame0_bit13.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _334_ (.D(FrameData[14]),
    .E(net52),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame0_bit14.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _335_ (.D(FrameData[15]),
    .E(net51),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame0_bit15.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _336_ (.D(FrameData[16]),
    .E(net51),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame0_bit16.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _337_ (.D(FrameData[17]),
    .E(net51),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame0_bit17.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _338_ (.D(FrameData[18]),
    .E(net51),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame0_bit18.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _339_ (.D(FrameData[19]),
    .E(net52),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame0_bit19.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _340_ (.D(FrameData[20]),
    .E(net51),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame0_bit20.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _341_ (.D(FrameData[21]),
    .E(net51),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame0_bit21.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _342_ (.D(FrameData[22]),
    .E(net51),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame0_bit22.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _343_ (.D(FrameData[23]),
    .E(net53),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame0_bit23.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _344_ (.D(FrameData[24]),
    .E(net53),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame0_bit24.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _345_ (.D(FrameData[25]),
    .E(net52),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame0_bit25.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _346_ (.D(FrameData[26]),
    .E(net52),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame0_bit26.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _347_ (.D(FrameData[27]),
    .E(net52),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame0_bit27.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _348_ (.D(FrameData[28]),
    .E(net51),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame0_bit28.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _349_ (.D(FrameData[29]),
    .E(net54),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame0_bit29.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _350_ (.D(FrameData[30]),
    .E(net54),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame0_bit30.Q ));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _351_ (.D(FrameData[31]),
    .E(net54),
    .Q(\Inst_W_IO4_ConfigMem.Inst_frame0_bit31.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _352_ (.D(A_O_top),
    .CLK(clknet_1_0__leaf_UserCLK_regs),
    .Q(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _353_ (.D(B_O_top),
    .CLK(clknet_1_1__leaf_UserCLK_regs),
    .Q(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _354_ (.D(C_O_top),
    .CLK(clknet_1_0__leaf_UserCLK_regs),
    .Q(\Inst_C_IO_1_bidirectional_frame_config_pass.Q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _355_ (.D(D_O_top),
    .CLK(clknet_1_1__leaf_UserCLK_regs),
    .Q(\Inst_D_IO_1_bidirectional_frame_config_pass.Q ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _356_ (.I(\Inst_W_IO4_switch_matrix.E1BEG0 ),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _357_ (.I(\Inst_W_IO4_switch_matrix.E1BEG1 ),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _358_ (.I(\Inst_W_IO4_switch_matrix.E1BEG2 ),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _359_ (.I(\Inst_W_IO4_switch_matrix.E1BEG3 ),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _360_ (.I(\Inst_W_IO4_switch_matrix.E2BEG0 ),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _361_ (.I(\Inst_W_IO4_switch_matrix.E2BEG1 ),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _362_ (.I(\Inst_W_IO4_switch_matrix.E2BEG2 ),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _363_ (.I(\Inst_W_IO4_switch_matrix.E2BEG3 ),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _364_ (.I(\Inst_W_IO4_switch_matrix.E2BEG4 ),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _365_ (.I(\Inst_W_IO4_switch_matrix.E2BEG5 ),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _366_ (.I(\Inst_W_IO4_switch_matrix.E2BEG6 ),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _367_ (.I(\Inst_W_IO4_switch_matrix.E2BEG7 ),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _368_ (.I(\Inst_W_IO4_switch_matrix.E2BEGb0 ),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _369_ (.I(\Inst_W_IO4_switch_matrix.E2BEGb1 ),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _370_ (.I(\Inst_W_IO4_switch_matrix.E2BEGb2 ),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _371_ (.I(\Inst_W_IO4_switch_matrix.E2BEGb3 ),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _372_ (.I(\Inst_W_IO4_switch_matrix.E2BEGb4 ),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _373_ (.I(\Inst_W_IO4_switch_matrix.E2BEGb5 ),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _374_ (.I(\Inst_W_IO4_switch_matrix.E2BEGb6 ),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _375_ (.I(\Inst_W_IO4_switch_matrix.E2BEGb7 ),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _376_ (.I(\Inst_W_IO4_switch_matrix.E6BEG0 ),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _377_ (.I(\Inst_W_IO4_switch_matrix.E6BEG1 ),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _378_ (.I(\Inst_W_IO4_switch_matrix.E6BEG2 ),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _379_ (.I(\Inst_W_IO4_switch_matrix.E6BEG3 ),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _380_ (.I(\Inst_W_IO4_switch_matrix.E6BEG4 ),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _381_ (.I(\Inst_W_IO4_switch_matrix.E6BEG5 ),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _382_ (.I(\Inst_W_IO4_switch_matrix.E6BEG6 ),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _383_ (.I(\Inst_W_IO4_switch_matrix.E6BEG7 ),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _384_ (.I(\Inst_W_IO4_switch_matrix.E6BEG8 ),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _385_ (.I(\Inst_W_IO4_switch_matrix.E6BEG9 ),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _386_ (.I(\Inst_W_IO4_switch_matrix.E6BEG10 ),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _387_ (.I(\Inst_W_IO4_switch_matrix.E6BEG11 ),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _388_ (.I(\Inst_W_IO4_switch_matrix.EE4BEG0 ),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _389_ (.I(\Inst_W_IO4_switch_matrix.EE4BEG1 ),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _390_ (.I(\Inst_W_IO4_switch_matrix.EE4BEG2 ),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _391_ (.I(\Inst_W_IO4_switch_matrix.EE4BEG3 ),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _392_ (.I(\Inst_W_IO4_switch_matrix.EE4BEG4 ),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _393_ (.I(\Inst_W_IO4_switch_matrix.EE4BEG5 ),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _394_ (.I(\Inst_W_IO4_switch_matrix.EE4BEG6 ),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _395_ (.I(\Inst_W_IO4_switch_matrix.EE4BEG7 ),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _396_ (.I(\Inst_W_IO4_switch_matrix.EE4BEG8 ),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _397_ (.I(\Inst_W_IO4_switch_matrix.EE4BEG9 ),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _398_ (.I(\Inst_W_IO4_switch_matrix.EE4BEG10 ),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _399_ (.I(\Inst_W_IO4_switch_matrix.EE4BEG11 ),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _400_ (.I(\Inst_W_IO4_switch_matrix.EE4BEG12 ),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _401_ (.I(\Inst_W_IO4_switch_matrix.EE4BEG13 ),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _402_ (.I(\Inst_W_IO4_switch_matrix.EE4BEG14 ),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _403_ (.I(\Inst_W_IO4_switch_matrix.EE4BEG15 ),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _404_ (.I(FrameData[0]),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _405_ (.I(FrameData[1]),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _406_ (.I(FrameData[2]),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _407_ (.I(FrameData[3]),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _408_ (.I(FrameData[4]),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _409_ (.I(FrameData[5]),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _410_ (.I(FrameData[6]),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _411_ (.I(FrameData[7]),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _412_ (.I(FrameData[8]),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _413_ (.I(FrameData[9]),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _414_ (.I(FrameData[10]),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _415_ (.I(FrameData[11]),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _416_ (.I(FrameData[12]),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _417_ (.I(FrameData[13]),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _418_ (.I(FrameData[14]),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _419_ (.I(FrameData[15]),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _420_ (.I(FrameData[16]),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _421_ (.I(FrameData[17]),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _422_ (.I(FrameData[18]),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _423_ (.I(FrameData[19]),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _424_ (.I(FrameData[20]),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _425_ (.I(FrameData[21]),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _426_ (.I(FrameData[22]),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _427_ (.I(FrameData[23]),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _428_ (.I(FrameData[24]),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _429_ (.I(FrameData[25]),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _430_ (.I(FrameData[26]),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _431_ (.I(FrameData[27]),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _432_ (.I(FrameData[28]),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _433_ (.I(FrameData[29]),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _434_ (.I(FrameData[30]),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _435_ (.I(FrameData[31]),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _436_ (.I(net55),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _437_ (.I(net50),
    .Z(net134));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _438_ (.I(net45),
    .Z(net135));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _439_ (.I(net41),
    .Z(net136));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _440_ (.I(net38),
    .Z(net137));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _441_ (.I(FrameStrobe[5]),
    .Z(net138));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _442_ (.I(FrameStrobe[6]),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _443_ (.I(FrameStrobe[7]),
    .Z(net140));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _444_ (.I(FrameStrobe[8]),
    .Z(net141));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _445_ (.I(FrameStrobe[9]),
    .Z(net142));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _446_ (.I(FrameStrobe[10]),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _447_ (.I(FrameStrobe[11]),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _448_ (.I(FrameStrobe[12]),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _449_ (.I(FrameStrobe[13]),
    .Z(net127));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _450_ (.I(FrameStrobe[14]),
    .Z(net128));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _451_ (.I(FrameStrobe[15]),
    .Z(net129));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _452_ (.I(FrameStrobe[16]),
    .Z(net130));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _453_ (.I(FrameStrobe[17]),
    .Z(net131));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _454_ (.I(FrameStrobe[18]),
    .Z(net132));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _455_ (.I(FrameStrobe[19]),
    .Z(net133));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _456_ (.I(clknet_1_0__leaf_UserCLK),
    .Z(net143));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Left_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Left_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Left_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Left_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Left_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Left_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Left_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Left_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Left_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_362 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout38 (.I(FrameStrobe[4]),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout39 (.I(net40),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout40 (.I(FrameStrobe[3]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout41 (.I(FrameStrobe[3]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout42 (.I(FrameStrobe[3]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout43 (.I(net46),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout44 (.I(net45),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout45 (.I(net46),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout46 (.I(FrameStrobe[2]),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout47 (.I(net50),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout48 (.I(net50),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout49 (.I(net50),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout50 (.I(FrameStrobe[1]),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout51 (.I(net52),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout52 (.I(net53),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout53 (.I(net54),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout54 (.I(net55),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout55 (.I(FrameStrobe[0]),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output1 (.I(net1),
    .Z(A_I_top));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output2 (.I(net2),
    .Z(A_T_top));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output3 (.I(net3),
    .Z(A_config_C_bit0));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output4 (.I(net4),
    .Z(A_config_C_bit1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output5 (.I(net5),
    .Z(A_config_C_bit2));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output6 (.I(net6),
    .Z(A_config_C_bit3));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output7 (.I(net144),
    .Z(B_I_top));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output8 (.I(net8),
    .Z(B_T_top));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output9 (.I(net9),
    .Z(B_config_C_bit0));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output10 (.I(net10),
    .Z(B_config_C_bit1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output11 (.I(net11),
    .Z(B_config_C_bit2));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output12 (.I(net12),
    .Z(B_config_C_bit3));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output13 (.I(net145),
    .Z(C_I_top));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output14 (.I(net14),
    .Z(C_T_top));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output15 (.I(net15),
    .Z(C_config_C_bit0));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output16 (.I(net16),
    .Z(C_config_C_bit1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output17 (.I(net17),
    .Z(C_config_C_bit2));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output18 (.I(net18),
    .Z(C_config_C_bit3));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output19 (.I(net19),
    .Z(D_I_top));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output20 (.I(net20),
    .Z(D_T_top));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output21 (.I(net21),
    .Z(D_config_C_bit0));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output22 (.I(net22),
    .Z(D_config_C_bit1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output23 (.I(net23),
    .Z(D_config_C_bit2));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output24 (.I(net24),
    .Z(D_config_C_bit3));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output25 (.I(net25),
    .Z(E1BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output26 (.I(net26),
    .Z(E1BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output27 (.I(net27),
    .Z(E1BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output28 (.I(net28),
    .Z(E1BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output29 (.I(net29),
    .Z(E2BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output30 (.I(net30),
    .Z(E2BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output31 (.I(net31),
    .Z(E2BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output32 (.I(net32),
    .Z(E2BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output33 (.I(net33),
    .Z(E2BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output34 (.I(net34),
    .Z(E2BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output35 (.I(net35),
    .Z(E2BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output36 (.I(net36),
    .Z(E2BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output37 (.I(net37),
    .Z(E2BEGb[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output38 (.I(net56),
    .Z(E2BEGb[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output39 (.I(net57),
    .Z(E2BEGb[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output40 (.I(net58),
    .Z(E2BEGb[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output41 (.I(net59),
    .Z(E2BEGb[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output42 (.I(net60),
    .Z(E2BEGb[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output43 (.I(net61),
    .Z(E2BEGb[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output44 (.I(net62),
    .Z(E2BEGb[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output45 (.I(net63),
    .Z(E6BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output46 (.I(net64),
    .Z(E6BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output47 (.I(net65),
    .Z(E6BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output48 (.I(net66),
    .Z(E6BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output49 (.I(net67),
    .Z(E6BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output50 (.I(net68),
    .Z(E6BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output51 (.I(net69),
    .Z(E6BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output52 (.I(net70),
    .Z(E6BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output53 (.I(net71),
    .Z(E6BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output54 (.I(net72),
    .Z(E6BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output55 (.I(net73),
    .Z(E6BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output56 (.I(net74),
    .Z(E6BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output57 (.I(net75),
    .Z(EE4BEG[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output58 (.I(net76),
    .Z(EE4BEG[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output59 (.I(net77),
    .Z(EE4BEG[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output60 (.I(net78),
    .Z(EE4BEG[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output61 (.I(net79),
    .Z(EE4BEG[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output62 (.I(net80),
    .Z(EE4BEG[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output63 (.I(net81),
    .Z(EE4BEG[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output64 (.I(net82),
    .Z(EE4BEG[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output65 (.I(net83),
    .Z(EE4BEG[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output66 (.I(net84),
    .Z(EE4BEG[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output67 (.I(net85),
    .Z(EE4BEG[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output68 (.I(net86),
    .Z(EE4BEG[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output69 (.I(net87),
    .Z(EE4BEG[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output70 (.I(net88),
    .Z(EE4BEG[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output71 (.I(net89),
    .Z(EE4BEG[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output72 (.I(net90),
    .Z(EE4BEG[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output73 (.I(net91),
    .Z(FrameData_O[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output74 (.I(net92),
    .Z(FrameData_O[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output75 (.I(net93),
    .Z(FrameData_O[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output76 (.I(net94),
    .Z(FrameData_O[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output77 (.I(net95),
    .Z(FrameData_O[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output78 (.I(net96),
    .Z(FrameData_O[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output79 (.I(net97),
    .Z(FrameData_O[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output80 (.I(net98),
    .Z(FrameData_O[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output81 (.I(net99),
    .Z(FrameData_O[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output82 (.I(net100),
    .Z(FrameData_O[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output83 (.I(net101),
    .Z(FrameData_O[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output84 (.I(net102),
    .Z(FrameData_O[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output85 (.I(net103),
    .Z(FrameData_O[20]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output86 (.I(net104),
    .Z(FrameData_O[21]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output87 (.I(net105),
    .Z(FrameData_O[22]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output88 (.I(net106),
    .Z(FrameData_O[23]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output89 (.I(net107),
    .Z(FrameData_O[24]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output90 (.I(net108),
    .Z(FrameData_O[25]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output91 (.I(net109),
    .Z(FrameData_O[26]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output92 (.I(net110),
    .Z(FrameData_O[27]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output93 (.I(net111),
    .Z(FrameData_O[28]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output94 (.I(net112),
    .Z(FrameData_O[29]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output95 (.I(net113),
    .Z(FrameData_O[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output96 (.I(net114),
    .Z(FrameData_O[30]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output97 (.I(net115),
    .Z(FrameData_O[31]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output98 (.I(net116),
    .Z(FrameData_O[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output99 (.I(net117),
    .Z(FrameData_O[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output100 (.I(net118),
    .Z(FrameData_O[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output101 (.I(net119),
    .Z(FrameData_O[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output102 (.I(net120),
    .Z(FrameData_O[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output103 (.I(net121),
    .Z(FrameData_O[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output104 (.I(net122),
    .Z(FrameData_O[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output105 (.I(net123),
    .Z(FrameStrobe_O[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output106 (.I(net124),
    .Z(FrameStrobe_O[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output107 (.I(net125),
    .Z(FrameStrobe_O[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output108 (.I(net126),
    .Z(FrameStrobe_O[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output109 (.I(net127),
    .Z(FrameStrobe_O[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output110 (.I(net128),
    .Z(FrameStrobe_O[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output111 (.I(net129),
    .Z(FrameStrobe_O[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output112 (.I(net130),
    .Z(FrameStrobe_O[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output113 (.I(net131),
    .Z(FrameStrobe_O[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output114 (.I(net132),
    .Z(FrameStrobe_O[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output115 (.I(net133),
    .Z(FrameStrobe_O[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output116 (.I(net134),
    .Z(FrameStrobe_O[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output117 (.I(net135),
    .Z(FrameStrobe_O[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output118 (.I(net136),
    .Z(FrameStrobe_O[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output119 (.I(net137),
    .Z(FrameStrobe_O[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output120 (.I(net138),
    .Z(FrameStrobe_O[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output121 (.I(net139),
    .Z(FrameStrobe_O[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output122 (.I(net140),
    .Z(FrameStrobe_O[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output123 (.I(net141),
    .Z(FrameStrobe_O[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 output124 (.I(net142),
    .Z(FrameStrobe_O[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output125 (.I(net143),
    .Z(UserCLKo));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 wire126 (.I(net7),
    .Z(net144));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 wire127 (.I(net13),
    .Z(net145));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_regs_0_UserCLK (.I(UserCLK),
    .Z(UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_UserCLK (.I(UserCLK),
    .Z(clknet_0_UserCLK));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_0__f_UserCLK (.I(clknet_0_UserCLK),
    .Z(clknet_1_0__leaf_UserCLK));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_UserCLK_regs (.I(UserCLK_regs),
    .Z(clknet_0_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_0__f_UserCLK_regs (.I(clknet_0_UserCLK_regs),
    .Z(clknet_1_0__leaf_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_1__f_UserCLK_regs (.I(clknet_0_UserCLK_regs),
    .Z(clknet_1_1__leaf_UserCLK_regs));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_240 ();
endmodule
