magic
tech gf180mcuD
magscale 1 10
timestamp 1764971362
<< metal1 >>
rect 672 56474 27888 56508
rect 672 56422 3806 56474
rect 3858 56422 3910 56474
rect 3962 56422 4014 56474
rect 4066 56422 23806 56474
rect 23858 56422 23910 56474
rect 23962 56422 24014 56474
rect 24066 56422 27888 56474
rect 672 56388 27888 56422
rect 3614 56306 3666 56318
rect 3614 56242 3666 56254
rect 5518 56306 5570 56318
rect 5518 56242 5570 56254
rect 8990 56306 9042 56318
rect 8990 56242 9042 56254
rect 10558 56306 10610 56318
rect 10558 56242 10610 56254
rect 13022 56306 13074 56318
rect 13022 56242 13074 56254
rect 14590 56306 14642 56318
rect 14590 56242 14642 56254
rect 16494 56306 16546 56318
rect 16494 56242 16546 56254
rect 18510 56306 18562 56318
rect 18510 56242 18562 56254
rect 20638 56306 20690 56318
rect 20638 56242 20690 56254
rect 21870 56306 21922 56318
rect 21870 56242 21922 56254
rect 24446 56306 24498 56318
rect 24446 56242 24498 56254
rect 26014 56306 26066 56318
rect 26014 56242 26066 56254
rect 7410 56142 7422 56194
rect 7474 56142 7486 56194
rect 5170 56030 5182 56082
rect 5234 56030 5246 56082
rect 20178 56030 20190 56082
rect 20242 56030 20254 56082
rect 25666 56030 25678 56082
rect 25730 56030 25742 56082
rect 1026 55918 1038 55970
rect 1090 55918 1102 55970
rect 3042 55918 3054 55970
rect 3106 55918 3118 55970
rect 8082 55918 8094 55970
rect 8146 55918 8158 55970
rect 9986 55918 9998 55970
rect 10050 55918 10062 55970
rect 11554 55918 11566 55970
rect 11618 55918 11630 55970
rect 14018 55918 14030 55970
rect 14082 55918 14094 55970
rect 15586 55918 15598 55970
rect 15650 55918 15662 55970
rect 17490 55918 17502 55970
rect 17554 55918 17566 55970
rect 19506 55918 19518 55970
rect 19570 55918 19582 55970
rect 22866 55918 22878 55970
rect 22930 55918 22942 55970
rect 23874 55918 23886 55970
rect 23938 55918 23950 55970
rect 1374 55858 1426 55870
rect 1374 55794 1426 55806
rect 672 55690 27888 55724
rect 672 55638 4466 55690
rect 4518 55638 4570 55690
rect 4622 55638 4674 55690
rect 4726 55638 24466 55690
rect 24518 55638 24570 55690
rect 24622 55638 24674 55690
rect 24726 55638 27888 55690
rect 672 55604 27888 55638
rect 18846 55410 18898 55422
rect 21634 55358 21646 55410
rect 21698 55358 21710 55410
rect 18846 55346 18898 55358
rect 20526 55298 20578 55310
rect 3490 55246 3502 55298
rect 3554 55246 3566 55298
rect 7522 55246 7534 55298
rect 7586 55246 7598 55298
rect 12898 55246 12910 55298
rect 12962 55246 12974 55298
rect 18274 55246 18286 55298
rect 18338 55246 18350 55298
rect 19282 55246 19294 55298
rect 19346 55246 19358 55298
rect 20066 55246 20078 55298
rect 20130 55246 20142 55298
rect 20850 55246 20862 55298
rect 20914 55246 20926 55298
rect 23650 55246 23662 55298
rect 23714 55246 23726 55298
rect 24658 55246 24670 55298
rect 24722 55246 24734 55298
rect 26226 55246 26238 55298
rect 26290 55246 26302 55298
rect 20526 55234 20578 55246
rect 2494 55186 2546 55198
rect 2494 55122 2546 55134
rect 6526 55186 6578 55198
rect 6526 55122 6578 55134
rect 11902 55186 11954 55198
rect 11902 55122 11954 55134
rect 17278 55186 17330 55198
rect 17278 55122 17330 55134
rect 22654 55186 22706 55198
rect 25554 55134 25566 55186
rect 25618 55134 25630 55186
rect 22654 55122 22706 55134
rect 27246 55074 27298 55086
rect 27246 55010 27298 55022
rect 672 54906 27888 54940
rect 672 54854 3806 54906
rect 3858 54854 3910 54906
rect 3962 54854 4014 54906
rect 4066 54854 23806 54906
rect 23858 54854 23910 54906
rect 23962 54854 24014 54906
rect 24066 54854 27888 54906
rect 672 54820 27888 54854
rect 22542 54738 22594 54750
rect 22542 54674 22594 54686
rect 24110 54738 24162 54750
rect 24110 54674 24162 54686
rect 19394 54574 19406 54626
rect 19458 54574 19470 54626
rect 21074 54574 21086 54626
rect 21138 54574 21150 54626
rect 25442 54574 25454 54626
rect 25506 54574 25518 54626
rect 19058 54462 19070 54514
rect 19122 54462 19134 54514
rect 24658 54462 24670 54514
rect 24722 54462 24734 54514
rect 21522 54350 21534 54402
rect 21586 54350 21598 54402
rect 23090 54350 23102 54402
rect 23154 54350 23166 54402
rect 26226 54350 26238 54402
rect 26290 54350 26302 54402
rect 27010 54350 27022 54402
rect 27074 54350 27086 54402
rect 20638 54290 20690 54302
rect 20638 54226 20690 54238
rect 672 54122 27888 54156
rect 672 54070 4466 54122
rect 4518 54070 4570 54122
rect 4622 54070 4674 54122
rect 4726 54070 24466 54122
rect 24518 54070 24570 54122
rect 24622 54070 24674 54122
rect 24726 54070 27888 54122
rect 672 54036 27888 54070
rect 20526 53730 20578 53742
rect 20526 53666 20578 53678
rect 20862 53730 20914 53742
rect 22318 53730 22370 53742
rect 21858 53678 21870 53730
rect 21922 53678 21934 53730
rect 22866 53678 22878 53730
rect 22930 53678 22942 53730
rect 24882 53678 24894 53730
rect 24946 53678 24958 53730
rect 26226 53678 26238 53730
rect 26290 53678 26302 53730
rect 20862 53666 20914 53678
rect 22318 53666 22370 53678
rect 19966 53618 20018 53630
rect 23774 53618 23826 53630
rect 21298 53566 21310 53618
rect 21362 53566 21374 53618
rect 25554 53566 25566 53618
rect 25618 53566 25630 53618
rect 19966 53554 20018 53566
rect 23774 53554 23826 53566
rect 27246 53506 27298 53518
rect 27246 53442 27298 53454
rect 672 53338 27888 53372
rect 672 53286 3806 53338
rect 3858 53286 3910 53338
rect 3962 53286 4014 53338
rect 4066 53286 23806 53338
rect 23858 53286 23910 53338
rect 23962 53286 24014 53338
rect 24066 53286 27888 53338
rect 672 53252 27888 53286
rect 24110 53170 24162 53182
rect 24110 53106 24162 53118
rect 21746 53006 21758 53058
rect 21810 53006 21822 53058
rect 22642 53006 22654 53058
rect 22706 53006 22718 53058
rect 27122 53006 27134 53058
rect 27186 53006 27198 53058
rect 21410 52894 21422 52946
rect 21474 52894 21486 52946
rect 23202 52894 23214 52946
rect 23266 52894 23278 52946
rect 24658 52894 24670 52946
rect 24722 52894 24734 52946
rect 25442 52782 25454 52834
rect 25506 52782 25518 52834
rect 26226 52782 26238 52834
rect 26290 52782 26302 52834
rect 22206 52722 22258 52734
rect 22206 52658 22258 52670
rect 672 52554 27888 52588
rect 672 52502 4466 52554
rect 4518 52502 4570 52554
rect 4622 52502 4674 52554
rect 4726 52502 24466 52554
rect 24518 52502 24570 52554
rect 24622 52502 24674 52554
rect 24726 52502 27888 52554
rect 672 52468 27888 52502
rect 21870 52274 21922 52286
rect 22754 52222 22766 52274
rect 22818 52222 22830 52274
rect 23538 52222 23550 52274
rect 23602 52222 23614 52274
rect 24658 52222 24670 52274
rect 24722 52222 24734 52274
rect 21870 52210 21922 52222
rect 22430 52162 22482 52174
rect 26226 52110 26238 52162
rect 26290 52110 26302 52162
rect 22430 52098 22482 52110
rect 25554 51998 25566 52050
rect 25618 51998 25630 52050
rect 27246 51938 27298 51950
rect 27246 51874 27298 51886
rect 672 51770 27888 51804
rect 672 51718 3806 51770
rect 3858 51718 3910 51770
rect 3962 51718 4014 51770
rect 4066 51718 23806 51770
rect 23858 51718 23910 51770
rect 23962 51718 24014 51770
rect 24066 51718 27888 51770
rect 672 51684 27888 51718
rect 23326 51490 23378 51502
rect 23326 51426 23378 51438
rect 24334 51490 24386 51502
rect 25330 51438 25342 51490
rect 25394 51438 25406 51490
rect 24334 51426 24386 51438
rect 24658 51214 24670 51266
rect 24722 51214 24734 51266
rect 26226 51214 26238 51266
rect 26290 51214 26302 51266
rect 27010 51214 27022 51266
rect 27074 51214 27086 51266
rect 22766 51154 22818 51166
rect 22766 51090 22818 51102
rect 23774 51154 23826 51166
rect 23774 51090 23826 51102
rect 672 50986 27888 51020
rect 672 50934 4466 50986
rect 4518 50934 4570 50986
rect 4622 50934 4674 50986
rect 4726 50934 24466 50986
rect 24518 50934 24570 50986
rect 24622 50934 24674 50986
rect 24726 50934 27888 50986
rect 672 50900 27888 50934
rect 23438 50706 23490 50718
rect 23438 50642 23490 50654
rect 23874 50542 23886 50594
rect 23938 50542 23950 50594
rect 24882 50542 24894 50594
rect 24946 50542 24958 50594
rect 26338 50542 26350 50594
rect 26402 50542 26414 50594
rect 25554 50430 25566 50482
rect 25618 50430 25630 50482
rect 27246 50370 27298 50382
rect 27246 50306 27298 50318
rect 672 50202 27888 50236
rect 672 50150 3806 50202
rect 3858 50150 3910 50202
rect 3962 50150 4014 50202
rect 4066 50150 23806 50202
rect 23858 50150 23910 50202
rect 23962 50150 24014 50202
rect 24066 50150 27888 50202
rect 672 50116 27888 50150
rect 25678 49922 25730 49934
rect 24210 49870 24222 49922
rect 24274 49870 24286 49922
rect 27122 49870 27134 49922
rect 27186 49870 27198 49922
rect 25678 49858 25730 49870
rect 26338 49758 26350 49810
rect 26402 49758 26414 49810
rect 24658 49646 24670 49698
rect 24722 49646 24734 49698
rect 23774 49586 23826 49598
rect 23774 49522 23826 49534
rect 672 49418 27888 49452
rect 672 49366 4466 49418
rect 4518 49366 4570 49418
rect 4622 49366 4674 49418
rect 4726 49366 24466 49418
rect 24518 49366 24570 49418
rect 24622 49366 24674 49418
rect 24726 49366 27888 49418
rect 672 49332 27888 49366
rect 24658 48974 24670 49026
rect 24722 48974 24734 49026
rect 26226 48974 26238 49026
rect 26290 48974 26302 49026
rect 25678 48802 25730 48814
rect 25678 48738 25730 48750
rect 27246 48802 27298 48814
rect 27246 48738 27298 48750
rect 672 48634 27888 48668
rect 672 48582 3806 48634
rect 3858 48582 3910 48634
rect 3962 48582 4014 48634
rect 4066 48582 23806 48634
rect 23858 48582 23910 48634
rect 23962 48582 24014 48634
rect 24066 48582 27888 48634
rect 672 48548 27888 48582
rect 25006 48354 25058 48366
rect 25778 48302 25790 48354
rect 25842 48302 25854 48354
rect 25006 48290 25058 48302
rect 26226 48078 26238 48130
rect 26290 48078 26302 48130
rect 27010 48078 27022 48130
rect 27074 48078 27086 48130
rect 24446 48018 24498 48030
rect 24446 47954 24498 47966
rect 25342 48018 25394 48030
rect 25342 47954 25394 47966
rect 672 47850 27888 47884
rect 672 47798 4466 47850
rect 4518 47798 4570 47850
rect 4622 47798 4674 47850
rect 4726 47798 24466 47850
rect 24518 47798 24570 47850
rect 24622 47798 24674 47850
rect 24726 47798 27888 47850
rect 672 47764 27888 47798
rect 24658 47406 24670 47458
rect 24722 47406 24734 47458
rect 26450 47406 26462 47458
rect 26514 47406 26526 47458
rect 25678 47346 25730 47358
rect 25678 47282 25730 47294
rect 27246 47234 27298 47246
rect 27246 47170 27298 47182
rect 672 47066 27888 47100
rect 672 47014 3806 47066
rect 3858 47014 3910 47066
rect 3962 47014 4014 47066
rect 4066 47014 23806 47066
rect 23858 47014 23910 47066
rect 23962 47014 24014 47066
rect 24066 47014 27888 47066
rect 672 46980 27888 47014
rect 25678 46786 25730 46798
rect 27122 46734 27134 46786
rect 27186 46734 27198 46786
rect 25678 46722 25730 46734
rect 24882 46622 24894 46674
rect 24946 46622 24958 46674
rect 26338 46622 26350 46674
rect 26402 46622 26414 46674
rect 672 46282 27888 46316
rect 672 46230 4466 46282
rect 4518 46230 4570 46282
rect 4622 46230 4674 46282
rect 4726 46230 24466 46282
rect 24518 46230 24570 46282
rect 24622 46230 24674 46282
rect 24726 46230 27888 46282
rect 672 46196 27888 46230
rect 24658 45838 24670 45890
rect 24722 45838 24734 45890
rect 26226 45838 26238 45890
rect 26290 45838 26302 45890
rect 25678 45666 25730 45678
rect 25678 45602 25730 45614
rect 27246 45666 27298 45678
rect 27246 45602 27298 45614
rect 672 45498 27888 45532
rect 672 45446 3806 45498
rect 3858 45446 3910 45498
rect 3962 45446 4014 45498
rect 4066 45446 23806 45498
rect 23858 45446 23910 45498
rect 23962 45446 24014 45498
rect 24066 45446 27888 45498
rect 672 45412 27888 45446
rect 26226 44942 26238 44994
rect 26290 44942 26302 44994
rect 27010 44942 27022 44994
rect 27074 44942 27086 44994
rect 672 44714 27888 44748
rect 672 44662 4466 44714
rect 4518 44662 4570 44714
rect 4622 44662 4674 44714
rect 4726 44662 24466 44714
rect 24518 44662 24570 44714
rect 24622 44662 24674 44714
rect 24726 44662 27888 44714
rect 672 44628 27888 44662
rect 24658 44270 24670 44322
rect 24722 44270 24734 44322
rect 26226 44270 26238 44322
rect 26290 44270 26302 44322
rect 25678 44210 25730 44222
rect 25678 44146 25730 44158
rect 27246 44098 27298 44110
rect 27246 44034 27298 44046
rect 672 43930 27888 43964
rect 672 43878 3806 43930
rect 3858 43878 3910 43930
rect 3962 43878 4014 43930
rect 4066 43878 23806 43930
rect 23858 43878 23910 43930
rect 23962 43878 24014 43930
rect 24066 43878 27888 43930
rect 672 43844 27888 43878
rect 25678 43650 25730 43662
rect 25678 43586 25730 43598
rect 24882 43486 24894 43538
rect 24946 43486 24958 43538
rect 26226 43374 26238 43426
rect 26290 43374 26302 43426
rect 26798 43314 26850 43326
rect 26798 43250 26850 43262
rect 672 43146 27888 43180
rect 672 43094 4466 43146
rect 4518 43094 4570 43146
rect 4622 43094 4674 43146
rect 4726 43094 24466 43146
rect 24518 43094 24570 43146
rect 24622 43094 24674 43146
rect 24726 43094 27888 43146
rect 672 43060 27888 43094
rect 24658 42702 24670 42754
rect 24722 42702 24734 42754
rect 26226 42702 26238 42754
rect 26290 42702 26302 42754
rect 25678 42530 25730 42542
rect 25678 42466 25730 42478
rect 27246 42530 27298 42542
rect 27246 42466 27298 42478
rect 672 42362 27888 42396
rect 672 42310 3806 42362
rect 3858 42310 3910 42362
rect 3962 42310 4014 42362
rect 4066 42310 23806 42362
rect 23858 42310 23910 42362
rect 23962 42310 24014 42362
rect 24066 42310 27888 42362
rect 672 42276 27888 42310
rect 4174 41970 4226 41982
rect 16258 41918 16270 41970
rect 16322 41918 16334 41970
rect 4174 41906 4226 41918
rect 18386 41806 18398 41858
rect 18450 41806 18462 41858
rect 26226 41806 26238 41858
rect 26290 41806 26302 41858
rect 3614 41746 3666 41758
rect 3614 41682 3666 41694
rect 26798 41746 26850 41758
rect 26798 41682 26850 41694
rect 672 41578 27888 41612
rect 672 41526 4466 41578
rect 4518 41526 4570 41578
rect 4622 41526 4674 41578
rect 4726 41526 24466 41578
rect 24518 41526 24570 41578
rect 24622 41526 24674 41578
rect 24726 41526 27888 41578
rect 672 41492 27888 41526
rect 6078 41410 6130 41422
rect 6078 41346 6130 41358
rect 6638 41298 6690 41310
rect 4274 41246 4286 41298
rect 4338 41246 4350 41298
rect 10546 41246 10558 41298
rect 10610 41246 10622 41298
rect 6638 41234 6690 41246
rect 8878 41186 8930 41198
rect 3826 41134 3838 41186
rect 3890 41134 3902 41186
rect 24770 41134 24782 41186
rect 24834 41134 24846 41186
rect 26226 41134 26238 41186
rect 26290 41134 26302 41186
rect 8878 41122 8930 41134
rect 9438 41074 9490 41086
rect 25678 41074 25730 41086
rect 10210 41022 10222 41074
rect 10274 41022 10286 41074
rect 9438 41010 9490 41022
rect 25678 41010 25730 41022
rect 5518 40962 5570 40974
rect 5518 40898 5570 40910
rect 11790 40962 11842 40974
rect 11790 40898 11842 40910
rect 27246 40962 27298 40974
rect 27246 40898 27298 40910
rect 672 40794 27888 40828
rect 672 40742 3806 40794
rect 3858 40742 3910 40794
rect 3962 40742 4014 40794
rect 4066 40742 23806 40794
rect 23858 40742 23910 40794
rect 23962 40742 24014 40794
rect 24066 40742 27888 40794
rect 672 40708 27888 40742
rect 2158 40514 2210 40526
rect 25678 40514 25730 40526
rect 13346 40462 13358 40514
rect 13410 40462 13422 40514
rect 15474 40462 15486 40514
rect 15538 40462 15550 40514
rect 2158 40450 2210 40462
rect 25678 40450 25730 40462
rect 4286 40402 4338 40414
rect 8766 40402 8818 40414
rect 1698 40350 1710 40402
rect 1762 40350 1774 40402
rect 2594 40350 2606 40402
rect 2658 40350 2670 40402
rect 7634 40350 7646 40402
rect 7698 40350 7710 40402
rect 8082 40350 8094 40402
rect 8146 40350 8158 40402
rect 9314 40350 9326 40402
rect 9378 40350 9390 40402
rect 10434 40350 10446 40402
rect 10498 40350 10510 40402
rect 17714 40350 17726 40402
rect 17778 40350 17790 40402
rect 18386 40350 18398 40402
rect 18450 40350 18462 40402
rect 24658 40350 24670 40402
rect 24722 40350 24734 40402
rect 26226 40350 26238 40402
rect 26290 40350 26302 40402
rect 4286 40338 4338 40350
rect 8766 40338 8818 40350
rect 6974 40290 7026 40302
rect 3042 40238 3054 40290
rect 3106 40238 3118 40290
rect 6974 40226 7026 40238
rect 7310 40290 7362 40302
rect 8306 40238 8318 40290
rect 8370 40238 8382 40290
rect 7310 40226 7362 40238
rect 6414 40178 6466 40190
rect 6414 40114 6466 40126
rect 12910 40178 12962 40190
rect 12910 40114 12962 40126
rect 26798 40178 26850 40190
rect 26798 40114 26850 40126
rect 672 40010 27888 40044
rect 672 39958 4466 40010
rect 4518 39958 4570 40010
rect 4622 39958 4674 40010
rect 4726 39958 24466 40010
rect 24518 39958 24570 40010
rect 24622 39958 24674 40010
rect 24726 39958 27888 40010
rect 672 39924 27888 39958
rect 6066 39790 6078 39842
rect 6130 39790 6142 39842
rect 9874 39790 9886 39842
rect 9938 39790 9950 39842
rect 12450 39790 12462 39842
rect 12514 39790 12526 39842
rect 2270 39730 2322 39742
rect 2270 39666 2322 39678
rect 3166 39730 3218 39742
rect 3166 39666 3218 39678
rect 5070 39730 5122 39742
rect 5070 39666 5122 39678
rect 12910 39730 12962 39742
rect 24658 39678 24670 39730
rect 24722 39678 24734 39730
rect 12910 39666 12962 39678
rect 1710 39618 1762 39630
rect 1710 39554 1762 39566
rect 2606 39618 2658 39630
rect 6750 39618 6802 39630
rect 5506 39566 5518 39618
rect 5570 39566 5582 39618
rect 5842 39566 5854 39618
rect 5906 39566 5918 39618
rect 7074 39566 7086 39618
rect 7138 39566 7150 39618
rect 7298 39566 7310 39618
rect 7362 39566 7374 39618
rect 8194 39566 8206 39618
rect 8258 39566 8270 39618
rect 9426 39566 9438 39618
rect 9490 39566 9502 39618
rect 11778 39566 11790 39618
rect 11842 39566 11854 39618
rect 12338 39566 12350 39618
rect 12402 39566 12414 39618
rect 13570 39566 13582 39618
rect 13634 39566 13646 39618
rect 14578 39566 14590 39618
rect 14642 39566 14654 39618
rect 16706 39566 16718 39618
rect 16770 39566 16782 39618
rect 26226 39566 26238 39618
rect 26290 39566 26302 39618
rect 2606 39554 2658 39566
rect 6750 39554 6802 39566
rect 11006 39506 11058 39518
rect 11006 39442 11058 39454
rect 11454 39506 11506 39518
rect 18722 39454 18734 39506
rect 18786 39454 18798 39506
rect 11454 39442 11506 39454
rect 25678 39394 25730 39406
rect 25678 39330 25730 39342
rect 27246 39394 27298 39406
rect 27246 39330 27298 39342
rect 672 39226 27888 39260
rect 672 39174 3806 39226
rect 3858 39174 3910 39226
rect 3962 39174 4014 39226
rect 4066 39174 23806 39226
rect 23858 39174 23910 39226
rect 23962 39174 24014 39226
rect 24066 39174 27888 39226
rect 672 39140 27888 39174
rect 7198 39058 7250 39070
rect 7198 38994 7250 39006
rect 2034 38894 2046 38946
rect 2098 38894 2110 38946
rect 2706 38894 2718 38946
rect 2770 38894 2782 38946
rect 5618 38894 5630 38946
rect 5682 38894 5694 38946
rect 13346 38894 13358 38946
rect 13410 38894 13422 38946
rect 26898 38894 26910 38946
rect 26962 38894 26974 38946
rect 4286 38834 4338 38846
rect 10546 38782 10558 38834
rect 10610 38782 10622 38834
rect 15810 38782 15822 38834
rect 15874 38782 15886 38834
rect 26226 38782 26238 38834
rect 26290 38782 26302 38834
rect 4286 38770 4338 38782
rect 3042 38670 3054 38722
rect 3106 38670 3118 38722
rect 5954 38670 5966 38722
rect 6018 38670 6030 38722
rect 10994 38670 11006 38722
rect 11058 38670 11070 38722
rect 18610 38670 18622 38722
rect 18674 38670 18686 38722
rect 1598 38610 1650 38622
rect 1598 38546 1650 38558
rect 12126 38610 12178 38622
rect 12126 38546 12178 38558
rect 12910 38610 12962 38622
rect 12910 38546 12962 38558
rect 672 38442 27888 38476
rect 672 38390 4466 38442
rect 4518 38390 4570 38442
rect 4622 38390 4674 38442
rect 4726 38390 24466 38442
rect 24518 38390 24570 38442
rect 24622 38390 24674 38442
rect 24726 38390 27888 38442
rect 672 38356 27888 38390
rect 6302 38274 6354 38286
rect 12562 38222 12574 38274
rect 12626 38222 12638 38274
rect 15138 38222 15150 38274
rect 15202 38222 15214 38274
rect 6302 38210 6354 38222
rect 7310 38162 7362 38174
rect 2370 38110 2382 38162
rect 2434 38110 2446 38162
rect 5058 38110 5070 38162
rect 5122 38110 5134 38162
rect 7310 38098 7362 38110
rect 7758 38162 7810 38174
rect 9986 38110 9998 38162
rect 10050 38110 10062 38162
rect 7758 38098 7810 38110
rect 6750 38050 6802 38062
rect 4610 37998 4622 38050
rect 4674 37998 4686 38050
rect 6750 37986 6802 37998
rect 8318 38050 8370 38062
rect 11118 38050 11170 38062
rect 9538 37998 9550 38050
rect 9602 37998 9614 38050
rect 11890 37998 11902 38050
rect 11954 37998 11966 38050
rect 12450 38004 12462 38056
rect 12514 38004 12526 38056
rect 15486 38050 15538 38062
rect 13122 37998 13134 38050
rect 13186 37998 13198 38050
rect 13570 37998 13582 38050
rect 13634 37998 13646 38050
rect 14690 37998 14702 38050
rect 14754 37998 14766 38050
rect 16706 37998 16718 38050
rect 16770 37998 16782 38050
rect 24882 37998 24894 38050
rect 24946 37998 24958 38050
rect 26226 37998 26238 38050
rect 26290 37998 26302 38050
rect 8318 37986 8370 37998
rect 11118 37986 11170 37998
rect 15486 37986 15538 37998
rect 11566 37938 11618 37950
rect 25678 37938 25730 37950
rect 2706 37886 2718 37938
rect 2770 37886 2782 37938
rect 17490 37886 17502 37938
rect 17554 37886 17566 37938
rect 19730 37886 19742 37938
rect 19794 37886 19806 37938
rect 11566 37874 11618 37886
rect 25678 37874 25730 37886
rect 1150 37826 1202 37838
rect 1150 37762 1202 37774
rect 27246 37826 27298 37838
rect 27246 37762 27298 37774
rect 672 37658 27888 37692
rect 672 37606 3806 37658
rect 3858 37606 3910 37658
rect 3962 37606 4014 37658
rect 4066 37606 23806 37658
rect 23858 37606 23910 37658
rect 23962 37606 24014 37658
rect 24066 37606 27888 37658
rect 672 37572 27888 37606
rect 6750 37490 6802 37502
rect 6750 37426 6802 37438
rect 2494 37378 2546 37390
rect 1474 37326 1486 37378
rect 1538 37326 1550 37378
rect 16482 37326 16494 37378
rect 16546 37326 16558 37378
rect 2494 37314 2546 37326
rect 8990 37266 9042 37278
rect 2034 37214 2046 37266
rect 2098 37214 2110 37266
rect 5170 37214 5182 37266
rect 5234 37214 5246 37266
rect 7858 37214 7870 37266
rect 7922 37214 7934 37266
rect 8306 37214 8318 37266
rect 8370 37214 8382 37266
rect 9538 37214 9550 37266
rect 9602 37214 9614 37266
rect 10658 37214 10670 37266
rect 10722 37214 10734 37266
rect 18610 37214 18622 37266
rect 18674 37214 18686 37266
rect 26226 37214 26238 37266
rect 26290 37214 26302 37266
rect 8990 37202 9042 37214
rect 7534 37154 7586 37166
rect 8530 37102 8542 37154
rect 8594 37102 8606 37154
rect 16594 37102 16606 37154
rect 16658 37102 16670 37154
rect 24658 37102 24670 37154
rect 24722 37102 24734 37154
rect 25442 37102 25454 37154
rect 25506 37102 25518 37154
rect 7534 37090 7586 37102
rect 1038 37042 1090 37054
rect 1038 36978 1090 36990
rect 1934 37042 1986 37054
rect 26798 37042 26850 37054
rect 5618 36990 5630 37042
rect 5682 36990 5694 37042
rect 1934 36978 1986 36990
rect 26798 36978 26850 36990
rect 672 36874 27888 36908
rect 672 36822 4466 36874
rect 4518 36822 4570 36874
rect 4622 36822 4674 36874
rect 4726 36822 24466 36874
rect 24518 36822 24570 36874
rect 24622 36822 24674 36874
rect 24726 36822 27888 36874
rect 672 36788 27888 36822
rect 10098 36654 10110 36706
rect 10162 36654 10174 36706
rect 18846 36594 18898 36606
rect 1586 36542 1598 36594
rect 1650 36542 1662 36594
rect 3938 36542 3950 36594
rect 4002 36542 4014 36594
rect 12114 36542 12126 36594
rect 12178 36542 12190 36594
rect 15698 36542 15710 36594
rect 15762 36542 15774 36594
rect 18846 36530 18898 36542
rect 6190 36482 6242 36494
rect 1250 36430 1262 36482
rect 1314 36430 1326 36482
rect 3378 36430 3390 36482
rect 3442 36430 3454 36482
rect 6190 36418 6242 36430
rect 8318 36482 8370 36494
rect 8318 36418 8370 36430
rect 14366 36482 14418 36494
rect 14366 36418 14418 36430
rect 14814 36482 14866 36494
rect 18286 36482 18338 36494
rect 15922 36430 15934 36482
rect 15986 36430 15998 36482
rect 17826 36430 17838 36482
rect 17890 36430 17902 36482
rect 24882 36430 24894 36482
rect 24946 36430 24958 36482
rect 26338 36430 26350 36482
rect 26402 36430 26414 36482
rect 14814 36418 14866 36430
rect 18286 36418 18338 36430
rect 6750 36370 6802 36382
rect 7858 36318 7870 36370
rect 7922 36318 7934 36370
rect 10546 36318 10558 36370
rect 10610 36318 10622 36370
rect 11778 36318 11790 36370
rect 11842 36318 11854 36370
rect 13906 36318 13918 36370
rect 13970 36318 13982 36370
rect 6750 36306 6802 36318
rect 2830 36258 2882 36270
rect 2830 36194 2882 36206
rect 5070 36258 5122 36270
rect 5070 36194 5122 36206
rect 8990 36258 9042 36270
rect 8990 36194 9042 36206
rect 13358 36258 13410 36270
rect 13358 36194 13410 36206
rect 15150 36258 15202 36270
rect 15150 36194 15202 36206
rect 17390 36258 17442 36270
rect 17390 36194 17442 36206
rect 25678 36258 25730 36270
rect 25678 36194 25730 36206
rect 27246 36258 27298 36270
rect 27246 36194 27298 36206
rect 672 36090 27888 36124
rect 672 36038 3806 36090
rect 3858 36038 3910 36090
rect 3962 36038 4014 36090
rect 4066 36038 23806 36090
rect 23858 36038 23910 36090
rect 23962 36038 24014 36090
rect 24066 36038 27888 36090
rect 672 36004 27888 36038
rect 7422 35810 7474 35822
rect 5842 35758 5854 35810
rect 5906 35758 5918 35810
rect 7422 35746 7474 35758
rect 11454 35810 11506 35822
rect 12898 35758 12910 35810
rect 12962 35758 12974 35810
rect 15474 35758 15486 35810
rect 15538 35758 15550 35810
rect 26898 35758 26910 35810
rect 26962 35758 26974 35810
rect 11454 35746 11506 35758
rect 9326 35698 9378 35710
rect 2594 35646 2606 35698
rect 2658 35646 2670 35698
rect 8306 35646 8318 35698
rect 8370 35646 8382 35698
rect 8642 35646 8654 35698
rect 8706 35646 8718 35698
rect 9986 35646 9998 35698
rect 10050 35646 10062 35698
rect 10882 35646 10894 35698
rect 10946 35646 10958 35698
rect 11890 35646 11902 35698
rect 11954 35646 11966 35698
rect 18386 35646 18398 35698
rect 18450 35646 18462 35698
rect 9326 35634 9378 35646
rect 7870 35586 7922 35598
rect 26226 35534 26238 35586
rect 26290 35534 26302 35586
rect 7870 35522 7922 35534
rect 4286 35474 4338 35486
rect 13358 35474 13410 35486
rect 3154 35422 3166 35474
rect 3218 35422 3230 35474
rect 6290 35422 6302 35474
rect 6354 35422 6366 35474
rect 8866 35422 8878 35474
rect 8930 35422 8942 35474
rect 4286 35410 4338 35422
rect 13358 35410 13410 35422
rect 672 35306 27888 35340
rect 672 35254 4466 35306
rect 4518 35254 4570 35306
rect 4622 35254 4674 35306
rect 4726 35254 24466 35306
rect 24518 35254 24570 35306
rect 24622 35254 24674 35306
rect 24726 35254 27888 35306
rect 672 35220 27888 35254
rect 16830 35138 16882 35150
rect 6066 35086 6078 35138
rect 6130 35086 6142 35138
rect 10994 35086 11006 35138
rect 11058 35086 11070 35138
rect 13570 35086 13582 35138
rect 13634 35086 13646 35138
rect 16830 35074 16882 35086
rect 14030 35026 14082 35038
rect 19854 35026 19906 35038
rect 3042 34974 3054 35026
rect 3106 34974 3118 35026
rect 17938 34974 17950 35026
rect 18002 34974 18014 35026
rect 14030 34962 14082 34974
rect 19854 34962 19906 34974
rect 20414 35026 20466 35038
rect 20414 34962 20466 34974
rect 2158 34914 2210 34926
rect 4286 34914 4338 34926
rect 6750 34914 6802 34926
rect 12126 34914 12178 34926
rect 18958 34914 19010 34926
rect 2594 34862 2606 34914
rect 2658 34862 2670 34914
rect 5394 34862 5406 34914
rect 5458 34862 5470 34914
rect 5954 34862 5966 34914
rect 6018 34862 6030 34914
rect 7186 34862 7198 34914
rect 7250 34862 7262 34914
rect 8082 34862 8094 34914
rect 8146 34862 8158 34914
rect 12898 34862 12910 34914
rect 12962 34862 12974 34914
rect 13346 34862 13358 34914
rect 13410 34862 13422 34914
rect 14578 34862 14590 34914
rect 14642 34862 14654 34914
rect 15698 34862 15710 34914
rect 15762 34862 15774 34914
rect 24658 34862 24670 34914
rect 24722 34862 24734 34914
rect 26226 34862 26238 34914
rect 26290 34862 26302 34914
rect 2158 34850 2210 34862
rect 4286 34850 4338 34862
rect 6750 34850 6802 34862
rect 12126 34850 12178 34862
rect 18958 34850 19010 34862
rect 5070 34802 5122 34814
rect 12574 34802 12626 34814
rect 25678 34802 25730 34814
rect 1698 34750 1710 34802
rect 1762 34750 1774 34802
rect 10546 34750 10558 34802
rect 10610 34750 10622 34802
rect 18386 34750 18398 34802
rect 18450 34750 18462 34802
rect 19394 34750 19406 34802
rect 19458 34750 19470 34802
rect 5070 34738 5122 34750
rect 12574 34738 12626 34750
rect 25678 34738 25730 34750
rect 27246 34690 27298 34702
rect 27246 34626 27298 34638
rect 672 34522 27888 34556
rect 672 34470 3806 34522
rect 3858 34470 3910 34522
rect 3962 34470 4014 34522
rect 4066 34470 23806 34522
rect 23858 34470 23910 34522
rect 23962 34470 24014 34522
rect 24066 34470 27888 34522
rect 672 34436 27888 34470
rect 6750 34354 6802 34366
rect 6750 34290 6802 34302
rect 25678 34242 25730 34254
rect 16706 34190 16718 34242
rect 16770 34190 16782 34242
rect 25678 34178 25730 34190
rect 2830 34130 2882 34142
rect 1474 34078 1486 34130
rect 1538 34078 1550 34130
rect 1922 34078 1934 34130
rect 1986 34078 1998 34130
rect 3266 34078 3278 34130
rect 3330 34078 3342 34130
rect 4274 34078 4286 34130
rect 4338 34078 4350 34130
rect 5170 34078 5182 34130
rect 5234 34078 5246 34130
rect 9202 34078 9214 34130
rect 9266 34078 9278 34130
rect 18498 34078 18510 34130
rect 18562 34078 18574 34130
rect 2830 34066 2882 34078
rect 1150 34018 1202 34030
rect 2146 33966 2158 34018
rect 2210 33966 2222 34018
rect 24658 33966 24670 34018
rect 24722 33966 24734 34018
rect 26226 33966 26238 34018
rect 26290 33966 26302 34018
rect 1150 33954 1202 33966
rect 7534 33906 7586 33918
rect 26798 33906 26850 33918
rect 5618 33854 5630 33906
rect 5682 33854 5694 33906
rect 8642 33854 8654 33906
rect 8706 33854 8718 33906
rect 7534 33842 7586 33854
rect 26798 33842 26850 33854
rect 672 33738 27888 33772
rect 672 33686 4466 33738
rect 4518 33686 4570 33738
rect 4622 33686 4674 33738
rect 4726 33686 24466 33738
rect 24518 33686 24570 33738
rect 24622 33686 24674 33738
rect 24726 33686 27888 33738
rect 672 33652 27888 33686
rect 6066 33518 6078 33570
rect 6130 33518 6142 33570
rect 9986 33518 9998 33570
rect 10050 33518 10062 33570
rect 18386 33518 18398 33570
rect 18450 33518 18462 33570
rect 8206 33458 8258 33470
rect 14590 33458 14642 33470
rect 1586 33406 1598 33458
rect 1650 33406 1662 33458
rect 12338 33406 12350 33458
rect 12402 33406 12414 33458
rect 8206 33394 8258 33406
rect 14590 33394 14642 33406
rect 7646 33346 7698 33358
rect 17390 33346 17442 33358
rect 9538 33294 9550 33346
rect 9602 33294 9614 33346
rect 11778 33294 11790 33346
rect 11842 33294 11854 33346
rect 17826 33294 17838 33346
rect 17890 33294 17902 33346
rect 24658 33294 24670 33346
rect 24722 33294 24734 33346
rect 26338 33294 26350 33346
rect 26402 33294 26414 33346
rect 7646 33282 7698 33294
rect 17390 33282 17442 33294
rect 1250 33182 1262 33234
rect 1314 33182 1326 33234
rect 5618 33182 5630 33234
rect 5682 33182 5694 33234
rect 15026 33182 15038 33234
rect 15090 33182 15102 33234
rect 16930 33182 16942 33234
rect 16994 33182 17006 33234
rect 17938 33182 17950 33234
rect 18002 33182 18014 33234
rect 2830 33122 2882 33134
rect 2830 33058 2882 33070
rect 7198 33122 7250 33134
rect 7198 33058 7250 33070
rect 11118 33122 11170 33134
rect 11118 33058 11170 33070
rect 13470 33122 13522 33134
rect 13470 33058 13522 33070
rect 19518 33122 19570 33134
rect 19518 33058 19570 33070
rect 25678 33122 25730 33134
rect 25678 33058 25730 33070
rect 27246 33122 27298 33134
rect 27246 33058 27298 33070
rect 672 32954 27888 32988
rect 672 32902 3806 32954
rect 3858 32902 3910 32954
rect 3962 32902 4014 32954
rect 4066 32902 23806 32954
rect 23858 32902 23910 32954
rect 23962 32902 24014 32954
rect 24066 32902 27888 32954
rect 672 32868 27888 32902
rect 18286 32786 18338 32798
rect 18286 32722 18338 32734
rect 14366 32674 14418 32686
rect 13346 32622 13358 32674
rect 13410 32622 13422 32674
rect 14366 32610 14418 32622
rect 17278 32674 17330 32686
rect 17278 32610 17330 32622
rect 18622 32674 18674 32686
rect 26898 32622 26910 32674
rect 26962 32622 26974 32674
rect 18622 32610 18674 32622
rect 7758 32562 7810 32574
rect 1586 32510 1598 32562
rect 1650 32510 1662 32562
rect 6738 32510 6750 32562
rect 6802 32510 6814 32562
rect 7074 32510 7086 32562
rect 7138 32510 7150 32562
rect 8418 32510 8430 32562
rect 8482 32510 8494 32562
rect 9314 32510 9326 32562
rect 9378 32510 9390 32562
rect 10434 32510 10446 32562
rect 10498 32510 10510 32562
rect 13010 32510 13022 32562
rect 13074 32510 13086 32562
rect 15138 32510 15150 32562
rect 15202 32510 15214 32562
rect 19058 32510 19070 32562
rect 19122 32510 19134 32562
rect 26226 32510 26238 32562
rect 26290 32510 26302 32562
rect 7758 32498 7810 32510
rect 4286 32450 4338 32462
rect 2146 32398 2158 32450
rect 2210 32398 2222 32450
rect 4286 32386 4338 32398
rect 6302 32450 6354 32462
rect 7298 32398 7310 32450
rect 7362 32398 7374 32450
rect 15586 32398 15598 32450
rect 15650 32398 15662 32450
rect 19170 32398 19182 32450
rect 19234 32398 19246 32450
rect 6302 32386 6354 32398
rect 3278 32338 3330 32350
rect 3278 32274 3330 32286
rect 3726 32338 3778 32350
rect 12126 32338 12178 32350
rect 10994 32286 11006 32338
rect 11058 32286 11070 32338
rect 3726 32274 3778 32286
rect 12126 32274 12178 32286
rect 13806 32338 13858 32350
rect 13806 32274 13858 32286
rect 16830 32338 16882 32350
rect 16830 32274 16882 32286
rect 17838 32338 17890 32350
rect 17838 32274 17890 32286
rect 672 32170 27888 32204
rect 672 32118 4466 32170
rect 4518 32118 4570 32170
rect 4622 32118 4674 32170
rect 4726 32118 24466 32170
rect 24518 32118 24570 32170
rect 24622 32118 24674 32170
rect 24726 32118 27888 32170
rect 672 32084 27888 32118
rect 13010 31950 13022 32002
rect 13074 31950 13086 32002
rect 17714 31950 17726 32002
rect 17778 31950 17790 32002
rect 3278 31890 3330 31902
rect 2818 31838 2830 31890
rect 2882 31838 2894 31890
rect 3278 31826 3330 31838
rect 18174 31890 18226 31902
rect 18174 31826 18226 31838
rect 8878 31778 8930 31790
rect 2258 31726 2270 31778
rect 2322 31726 2334 31778
rect 2706 31726 2718 31778
rect 2770 31726 2782 31778
rect 4050 31726 4062 31778
rect 4114 31726 4126 31778
rect 4834 31726 4846 31778
rect 4898 31726 4910 31778
rect 7298 31726 7310 31778
rect 7362 31726 7374 31778
rect 12338 31726 12350 31778
rect 12402 31726 12414 31778
rect 12786 31726 12798 31778
rect 12850 31726 12862 31778
rect 13570 31726 13582 31778
rect 13634 31726 13646 31778
rect 14242 31726 14254 31778
rect 14306 31726 14318 31778
rect 15026 31726 15038 31778
rect 15090 31726 15102 31778
rect 17042 31726 17054 31778
rect 17106 31726 17118 31778
rect 17490 31726 17502 31778
rect 17554 31726 17566 31778
rect 18946 31726 18958 31778
rect 19010 31726 19022 31778
rect 19842 31726 19854 31778
rect 19906 31726 19918 31778
rect 24658 31726 24670 31778
rect 24722 31726 24734 31778
rect 26338 31726 26350 31778
rect 26402 31726 26414 31778
rect 8878 31714 8930 31726
rect 1822 31666 1874 31678
rect 12014 31666 12066 31678
rect 7970 31614 7982 31666
rect 8034 31614 8046 31666
rect 9314 31614 9326 31666
rect 9378 31614 9390 31666
rect 1822 31602 1874 31614
rect 12014 31602 12066 31614
rect 16718 31666 16770 31678
rect 16718 31602 16770 31614
rect 25678 31666 25730 31678
rect 26898 31614 26910 31666
rect 26962 31614 26974 31666
rect 25678 31602 25730 31614
rect 672 31386 27888 31420
rect 672 31334 3806 31386
rect 3858 31334 3910 31386
rect 3962 31334 4014 31386
rect 4066 31334 23806 31386
rect 23858 31334 23910 31386
rect 23962 31334 24014 31386
rect 24066 31334 27888 31386
rect 672 31300 27888 31334
rect 15822 31218 15874 31230
rect 15822 31154 15874 31166
rect 4398 31106 4450 31118
rect 11902 31106 11954 31118
rect 6626 31054 6638 31106
rect 6690 31054 6702 31106
rect 7186 31054 7198 31106
rect 7250 31054 7262 31106
rect 4398 31042 4450 31054
rect 11902 31042 11954 31054
rect 27246 31106 27298 31118
rect 27246 31042 27298 31054
rect 11342 30994 11394 31006
rect 18398 30994 18450 31006
rect 1250 30942 1262 30994
rect 1314 30942 1326 30994
rect 2370 30942 2382 30994
rect 2434 30942 2446 30994
rect 3490 30942 3502 30994
rect 3554 30942 3566 30994
rect 3938 30942 3950 30994
rect 4002 30942 4014 30994
rect 8082 30942 8094 30994
rect 8146 30942 8158 30994
rect 10434 30942 10446 30994
rect 10498 30942 10510 30994
rect 14242 30942 14254 30994
rect 14306 30942 14318 30994
rect 17154 30942 17166 30994
rect 17218 30942 17230 30994
rect 17490 30942 17502 30994
rect 17554 30942 17566 30994
rect 18722 30942 18734 30994
rect 18786 30942 18798 30994
rect 19842 30942 19854 30994
rect 19906 30942 19918 30994
rect 24882 30942 24894 30994
rect 24946 30942 24958 30994
rect 11342 30930 11394 30942
rect 18398 30930 18450 30942
rect 2942 30882 2994 30894
rect 10894 30882 10946 30894
rect 8642 30830 8654 30882
rect 8706 30830 8718 30882
rect 2942 30818 2994 30830
rect 10894 30818 10946 30830
rect 16718 30882 16770 30894
rect 17714 30830 17726 30882
rect 17778 30830 17790 30882
rect 25442 30830 25454 30882
rect 25506 30830 25518 30882
rect 26226 30830 26238 30882
rect 26290 30830 26302 30882
rect 16718 30818 16770 30830
rect 6190 30770 6242 30782
rect 3378 30718 3390 30770
rect 3442 30718 3454 30770
rect 6190 30706 6242 30718
rect 7646 30770 7698 30782
rect 7646 30706 7698 30718
rect 9774 30770 9826 30782
rect 14690 30718 14702 30770
rect 14754 30718 14766 30770
rect 9774 30706 9826 30718
rect 672 30602 27888 30636
rect 672 30550 4466 30602
rect 4518 30550 4570 30602
rect 4622 30550 4674 30602
rect 4726 30550 24466 30602
rect 24518 30550 24570 30602
rect 24622 30550 24674 30602
rect 24726 30550 27888 30602
rect 672 30516 27888 30550
rect 3166 30434 3218 30446
rect 6066 30382 6078 30434
rect 6130 30382 6142 30434
rect 10434 30382 10446 30434
rect 10498 30382 10510 30434
rect 3166 30370 3218 30382
rect 16158 30322 16210 30334
rect 17266 30270 17278 30322
rect 17330 30270 17342 30322
rect 16158 30258 16210 30270
rect 6750 30210 6802 30222
rect 9438 30210 9490 30222
rect 11118 30210 11170 30222
rect 14142 30210 14194 30222
rect 1026 30158 1038 30210
rect 1090 30158 1102 30210
rect 5394 30158 5406 30210
rect 5458 30158 5470 30210
rect 5842 30158 5854 30210
rect 5906 30158 5918 30210
rect 7074 30158 7086 30210
rect 7138 30158 7150 30210
rect 8194 30158 8206 30210
rect 8258 30158 8270 30210
rect 9762 30158 9774 30210
rect 9826 30158 9838 30210
rect 10210 30158 10222 30210
rect 10274 30158 10286 30210
rect 11442 30158 11454 30210
rect 11506 30158 11518 30210
rect 12562 30158 12574 30210
rect 12626 30158 12638 30210
rect 15698 30158 15710 30210
rect 15762 30158 15774 30210
rect 16818 30158 16830 30210
rect 16882 30158 16894 30210
rect 26226 30158 26238 30210
rect 26290 30158 26302 30210
rect 6750 30146 6802 30158
rect 9438 30146 9490 30158
rect 11118 30146 11170 30158
rect 14142 30146 14194 30158
rect 5070 30098 5122 30110
rect 2706 30046 2718 30098
rect 2770 30046 2782 30098
rect 5070 30034 5122 30046
rect 14702 30098 14754 30110
rect 14702 30034 14754 30046
rect 18510 30098 18562 30110
rect 26898 30046 26910 30098
rect 26962 30046 26974 30098
rect 18510 30034 18562 30046
rect 2046 29986 2098 29998
rect 2046 29922 2098 29934
rect 672 29818 27888 29852
rect 672 29766 3806 29818
rect 3858 29766 3910 29818
rect 3962 29766 4014 29818
rect 4066 29766 23806 29818
rect 23858 29766 23910 29818
rect 23962 29766 24014 29818
rect 24066 29766 27888 29818
rect 672 29732 27888 29766
rect 2830 29650 2882 29662
rect 2830 29586 2882 29598
rect 6750 29650 6802 29662
rect 6750 29586 6802 29598
rect 17502 29650 17554 29662
rect 17502 29586 17554 29598
rect 27246 29538 27298 29550
rect 1250 29486 1262 29538
rect 1314 29486 1326 29538
rect 5170 29486 5182 29538
rect 5234 29486 5246 29538
rect 12114 29486 12126 29538
rect 12178 29486 12190 29538
rect 15922 29486 15934 29538
rect 15986 29486 15998 29538
rect 27246 29474 27298 29486
rect 19742 29426 19794 29438
rect 8530 29374 8542 29426
rect 8594 29374 8606 29426
rect 11778 29374 11790 29426
rect 11842 29374 11854 29426
rect 13570 29374 13582 29426
rect 13634 29374 13646 29426
rect 18162 29374 18174 29426
rect 18226 29374 18238 29426
rect 19742 29362 19794 29374
rect 1586 29262 1598 29314
rect 1650 29262 1662 29314
rect 5506 29262 5518 29314
rect 5570 29262 5582 29314
rect 14130 29262 14142 29314
rect 14194 29262 14206 29314
rect 18610 29262 18622 29314
rect 18674 29262 18686 29314
rect 26226 29262 26238 29314
rect 26290 29262 26302 29314
rect 10110 29202 10162 29214
rect 8978 29150 8990 29202
rect 9042 29150 9054 29202
rect 10110 29138 10162 29150
rect 15262 29202 15314 29214
rect 16370 29150 16382 29202
rect 16434 29150 16446 29202
rect 15262 29138 15314 29150
rect 672 29034 27888 29068
rect 672 28982 4466 29034
rect 4518 28982 4570 29034
rect 4622 28982 4674 29034
rect 4726 28982 24466 29034
rect 24518 28982 24570 29034
rect 24622 28982 24674 29034
rect 24726 28982 27888 29034
rect 672 28948 27888 28982
rect 2830 28866 2882 28878
rect 2830 28802 2882 28814
rect 5070 28866 5122 28878
rect 11330 28814 11342 28866
rect 11394 28814 11406 28866
rect 13906 28814 13918 28866
rect 13970 28814 13982 28866
rect 5070 28802 5122 28814
rect 5518 28754 5570 28766
rect 12910 28754 12962 28766
rect 1586 28702 1598 28754
rect 1650 28702 1662 28754
rect 3826 28702 3838 28754
rect 3890 28702 3902 28754
rect 6962 28702 6974 28754
rect 7026 28702 7038 28754
rect 5518 28690 5570 28702
rect 12910 28690 12962 28702
rect 18398 28754 18450 28766
rect 19394 28702 19406 28754
rect 19458 28702 19470 28754
rect 26226 28702 26238 28754
rect 26290 28702 26302 28754
rect 18398 28690 18450 28702
rect 12462 28642 12514 28654
rect 14366 28642 14418 28654
rect 20078 28642 20130 28654
rect 1250 28590 1262 28642
rect 1314 28590 1326 28642
rect 5954 28590 5966 28642
rect 6018 28590 6030 28642
rect 13234 28590 13246 28642
rect 13298 28590 13310 28642
rect 13682 28590 13694 28642
rect 13746 28590 13758 28642
rect 14914 28590 14926 28642
rect 14978 28590 14990 28642
rect 15922 28590 15934 28642
rect 15986 28590 15998 28642
rect 18834 28590 18846 28642
rect 18898 28590 18910 28642
rect 19170 28590 19182 28642
rect 19234 28590 19246 28642
rect 20402 28590 20414 28642
rect 20466 28590 20478 28642
rect 20626 28590 20638 28642
rect 20690 28590 20702 28642
rect 21410 28590 21422 28642
rect 21474 28590 21486 28642
rect 12462 28578 12514 28590
rect 14366 28578 14418 28590
rect 20078 28578 20130 28590
rect 27246 28530 27298 28542
rect 3490 28478 3502 28530
rect 3554 28478 3566 28530
rect 6626 28478 6638 28530
rect 6690 28478 6702 28530
rect 10882 28478 10894 28530
rect 10946 28478 10958 28530
rect 27246 28466 27298 28478
rect 8206 28418 8258 28430
rect 8206 28354 8258 28366
rect 672 28250 27888 28284
rect 672 28198 3806 28250
rect 3858 28198 3910 28250
rect 3962 28198 4014 28250
rect 4066 28198 23806 28250
rect 23858 28198 23910 28250
rect 23962 28198 24014 28250
rect 24066 28198 27888 28250
rect 672 28164 27888 28198
rect 19070 28082 19122 28094
rect 19070 28018 19122 28030
rect 27246 28082 27298 28094
rect 27246 28018 27298 28030
rect 4958 27970 5010 27982
rect 1474 27918 1486 27970
rect 1538 27918 1550 27970
rect 4958 27906 5010 27918
rect 8990 27970 9042 27982
rect 8990 27906 9042 27918
rect 13582 27970 13634 27982
rect 20078 27970 20130 27982
rect 17490 27918 17502 27970
rect 17554 27918 17566 27970
rect 13582 27906 13634 27918
rect 20078 27906 20130 27918
rect 25678 27970 25730 27982
rect 25678 27906 25730 27918
rect 1038 27858 1090 27870
rect 4286 27858 4338 27870
rect 10446 27858 10498 27870
rect 15262 27858 15314 27870
rect 2594 27806 2606 27858
rect 2658 27806 2670 27858
rect 5282 27806 5294 27858
rect 5346 27806 5358 27858
rect 5730 27806 5742 27858
rect 5794 27806 5806 27858
rect 6514 27806 6526 27858
rect 6578 27806 6590 27858
rect 7186 27806 7198 27858
rect 7250 27806 7262 27858
rect 8082 27806 8094 27858
rect 8146 27806 8158 27858
rect 9314 27806 9326 27858
rect 9378 27806 9390 27858
rect 9762 27806 9774 27858
rect 9826 27806 9838 27858
rect 11218 27806 11230 27858
rect 11282 27806 11294 27858
rect 12002 27806 12014 27858
rect 12066 27806 12078 27858
rect 14018 27806 14030 27858
rect 14082 27806 14094 27858
rect 14466 27806 14478 27858
rect 14530 27806 14542 27858
rect 15586 27806 15598 27858
rect 15650 27806 15662 27858
rect 16594 27806 16606 27858
rect 16658 27806 16670 27858
rect 26338 27806 26350 27858
rect 26402 27806 26414 27858
rect 1038 27794 1090 27806
rect 4286 27794 4338 27806
rect 10446 27794 10498 27806
rect 15262 27794 15314 27806
rect 19518 27746 19570 27758
rect 3042 27694 3054 27746
rect 3106 27694 3118 27746
rect 5954 27694 5966 27746
rect 6018 27694 6030 27746
rect 17826 27694 17838 27746
rect 17890 27694 17902 27746
rect 24658 27694 24670 27746
rect 24722 27694 24734 27746
rect 19518 27682 19570 27694
rect 9986 27582 9998 27634
rect 10050 27582 10062 27634
rect 14578 27582 14590 27634
rect 14642 27582 14654 27634
rect 672 27466 27888 27500
rect 672 27414 4466 27466
rect 4518 27414 4570 27466
rect 4622 27414 4674 27466
rect 4726 27414 24466 27466
rect 24518 27414 24570 27466
rect 24622 27414 24674 27466
rect 24726 27414 27888 27466
rect 672 27380 27888 27414
rect 6526 27298 6578 27310
rect 5394 27246 5406 27298
rect 5458 27246 5470 27298
rect 6526 27234 6578 27246
rect 10222 27298 10274 27310
rect 10222 27234 10274 27246
rect 12910 27298 12962 27310
rect 12910 27234 12962 27246
rect 15150 27298 15202 27310
rect 15150 27234 15202 27246
rect 15598 27298 15650 27310
rect 15598 27234 15650 27246
rect 10782 27186 10834 27198
rect 16158 27186 16210 27198
rect 1586 27134 1598 27186
rect 1650 27134 1662 27186
rect 11666 27134 11678 27186
rect 11730 27134 11742 27186
rect 13906 27134 13918 27186
rect 13970 27134 13982 27186
rect 18162 27134 18174 27186
rect 18226 27134 18238 27186
rect 24658 27134 24670 27186
rect 24722 27134 24734 27186
rect 10782 27122 10834 27134
rect 16158 27122 16210 27134
rect 1250 27022 1262 27074
rect 1314 27022 1326 27074
rect 4834 27022 4846 27074
rect 4898 27022 4910 27074
rect 11330 27022 11342 27074
rect 11394 27022 11406 27074
rect 13458 27022 13470 27074
rect 13522 27022 13534 27074
rect 17714 27022 17726 27074
rect 17778 27022 17790 27074
rect 26226 27022 26238 27074
rect 26290 27022 26302 27074
rect 27246 26962 27298 26974
rect 27246 26898 27298 26910
rect 2830 26850 2882 26862
rect 2830 26786 2882 26798
rect 19406 26850 19458 26862
rect 19406 26786 19458 26798
rect 25678 26850 25730 26862
rect 25678 26786 25730 26798
rect 672 26682 27888 26716
rect 672 26630 3806 26682
rect 3858 26630 3910 26682
rect 3962 26630 4014 26682
rect 4066 26630 23806 26682
rect 23858 26630 23910 26682
rect 23962 26630 24014 26682
rect 24066 26630 27888 26682
rect 672 26596 27888 26630
rect 27246 26514 27298 26526
rect 27246 26450 27298 26462
rect 13358 26402 13410 26414
rect 1698 26350 1710 26402
rect 1762 26350 1774 26402
rect 4162 26350 4174 26402
rect 4226 26350 4238 26402
rect 7634 26350 7646 26402
rect 7698 26350 7710 26402
rect 13358 26338 13410 26350
rect 14590 26402 14642 26414
rect 16482 26350 16494 26402
rect 16546 26350 16558 26402
rect 19618 26350 19630 26402
rect 19682 26350 19694 26402
rect 14590 26338 14642 26350
rect 12898 26238 12910 26290
rect 12962 26238 12974 26290
rect 2034 26126 2046 26178
rect 2098 26126 2110 26178
rect 26226 26126 26238 26178
rect 26290 26126 26302 26178
rect 3278 26066 3330 26078
rect 3278 26002 3330 26014
rect 3726 26066 3778 26078
rect 9214 26066 9266 26078
rect 8082 26014 8094 26066
rect 8146 26014 8158 26066
rect 3726 26002 3778 26014
rect 9214 26002 9266 26014
rect 14030 26066 14082 26078
rect 18062 26066 18114 26078
rect 16930 26014 16942 26066
rect 16994 26014 17006 26066
rect 14030 26002 14082 26014
rect 18062 26002 18114 26014
rect 19182 26066 19234 26078
rect 19182 26002 19234 26014
rect 672 25898 27888 25932
rect 672 25846 4466 25898
rect 4518 25846 4570 25898
rect 4622 25846 4674 25898
rect 4726 25846 24466 25898
rect 24518 25846 24570 25898
rect 24622 25846 24674 25898
rect 24726 25846 27888 25898
rect 672 25812 27888 25846
rect 3042 25678 3054 25730
rect 3106 25678 3118 25730
rect 3502 25618 3554 25630
rect 9438 25618 9490 25630
rect 15262 25618 15314 25630
rect 6626 25566 6638 25618
rect 6690 25566 6702 25618
rect 10882 25566 10894 25618
rect 10946 25566 10958 25618
rect 13122 25566 13134 25618
rect 13186 25566 13198 25618
rect 3502 25554 3554 25566
rect 9438 25554 9490 25566
rect 15262 25554 15314 25566
rect 17502 25618 17554 25630
rect 18498 25566 18510 25618
rect 18562 25566 18574 25618
rect 24658 25566 24670 25618
rect 24722 25566 24734 25618
rect 17502 25554 17554 25566
rect 8878 25506 8930 25518
rect 2482 25454 2494 25506
rect 2546 25454 2558 25506
rect 2818 25454 2830 25506
rect 2882 25454 2894 25506
rect 4274 25454 4286 25506
rect 4338 25454 4350 25506
rect 5058 25454 5070 25506
rect 5122 25454 5134 25506
rect 6290 25454 6302 25506
rect 6354 25454 6366 25506
rect 8878 25442 8930 25454
rect 14702 25506 14754 25518
rect 19182 25506 19234 25518
rect 17938 25454 17950 25506
rect 18002 25454 18014 25506
rect 18386 25454 18398 25506
rect 18450 25454 18462 25506
rect 19730 25454 19742 25506
rect 19794 25454 19806 25506
rect 20514 25454 20526 25506
rect 20578 25454 20590 25506
rect 26226 25454 26238 25506
rect 26290 25454 26302 25506
rect 14702 25442 14754 25454
rect 19182 25442 19234 25454
rect 2046 25394 2098 25406
rect 27246 25394 27298 25406
rect 10434 25342 10446 25394
rect 10498 25342 10510 25394
rect 12674 25342 12686 25394
rect 12738 25342 12750 25394
rect 2046 25330 2098 25342
rect 27246 25330 27298 25342
rect 7870 25282 7922 25294
rect 7870 25218 7922 25230
rect 12014 25282 12066 25294
rect 12014 25218 12066 25230
rect 14254 25282 14306 25294
rect 14254 25218 14306 25230
rect 25678 25282 25730 25294
rect 25678 25218 25730 25230
rect 672 25114 27888 25148
rect 672 25062 3806 25114
rect 3858 25062 3910 25114
rect 3962 25062 4014 25114
rect 4066 25062 23806 25114
rect 23858 25062 23910 25114
rect 23962 25062 24014 25114
rect 24066 25062 27888 25114
rect 672 25028 27888 25062
rect 27246 24946 27298 24958
rect 27246 24882 27298 24894
rect 6190 24834 6242 24846
rect 6190 24770 6242 24782
rect 7534 24834 7586 24846
rect 19518 24834 19570 24846
rect 18162 24782 18174 24834
rect 18226 24782 18238 24834
rect 7534 24770 7586 24782
rect 19518 24770 19570 24782
rect 2718 24722 2770 24734
rect 9214 24722 9266 24734
rect 14366 24722 14418 24734
rect 18958 24722 19010 24734
rect 1250 24670 1262 24722
rect 1314 24670 1326 24722
rect 2258 24670 2270 24722
rect 2322 24670 2334 24722
rect 3490 24670 3502 24722
rect 3554 24670 3566 24722
rect 4050 24670 4062 24722
rect 4114 24670 4126 24722
rect 7858 24670 7870 24722
rect 7922 24670 7934 24722
rect 8306 24670 8318 24722
rect 8370 24670 8382 24722
rect 9762 24670 9774 24722
rect 9826 24670 9838 24722
rect 10658 24670 10670 24722
rect 10722 24670 10734 24722
rect 13346 24670 13358 24722
rect 13410 24670 13422 24722
rect 13794 24670 13806 24722
rect 13858 24670 13870 24722
rect 14914 24670 14926 24722
rect 14978 24670 14990 24722
rect 15922 24670 15934 24722
rect 15986 24670 15998 24722
rect 24882 24670 24894 24722
rect 24946 24670 24958 24722
rect 26226 24670 26238 24722
rect 26290 24670 26302 24722
rect 2718 24658 2770 24670
rect 9214 24658 9266 24670
rect 14366 24658 14418 24670
rect 18958 24658 19010 24670
rect 4398 24610 4450 24622
rect 12238 24610 12290 24622
rect 8530 24558 8542 24610
rect 8594 24558 8606 24610
rect 4398 24546 4450 24558
rect 12238 24546 12290 24558
rect 12910 24610 12962 24622
rect 13906 24558 13918 24610
rect 13970 24558 13982 24610
rect 25442 24558 25454 24610
rect 25506 24558 25518 24610
rect 12910 24546 12962 24558
rect 5630 24498 5682 24510
rect 3378 24446 3390 24498
rect 3442 24446 3454 24498
rect 5630 24434 5682 24446
rect 12014 24498 12066 24510
rect 12014 24434 12066 24446
rect 12126 24498 12178 24510
rect 12126 24434 12178 24446
rect 16606 24498 16658 24510
rect 17714 24446 17726 24498
rect 17778 24446 17790 24498
rect 16606 24434 16658 24446
rect 672 24330 27888 24364
rect 672 24278 4466 24330
rect 4518 24278 4570 24330
rect 4622 24278 4674 24330
rect 4726 24278 24466 24330
rect 24518 24278 24570 24330
rect 24622 24278 24674 24330
rect 24726 24278 27888 24330
rect 672 24244 27888 24278
rect 1486 24162 1538 24174
rect 1486 24098 1538 24110
rect 2494 24162 2546 24174
rect 5618 24110 5630 24162
rect 5682 24110 5694 24162
rect 13794 24110 13806 24162
rect 13858 24110 13870 24162
rect 2494 24098 2546 24110
rect 6078 24050 6130 24062
rect 3602 23998 3614 24050
rect 3666 23998 3678 24050
rect 6078 23986 6130 23998
rect 9326 24050 9378 24062
rect 11218 23998 11230 24050
rect 11282 23998 11294 24050
rect 17938 23998 17950 24050
rect 18002 23998 18014 24050
rect 24658 23998 24670 24050
rect 24722 23998 24734 24050
rect 9326 23986 9378 23998
rect 2046 23938 2098 23950
rect 9886 23938 9938 23950
rect 5058 23886 5070 23938
rect 5122 23886 5134 23938
rect 5394 23886 5406 23938
rect 5458 23886 5470 23938
rect 6626 23886 6638 23938
rect 6690 23886 6702 23938
rect 7746 23886 7758 23938
rect 7810 23886 7822 23938
rect 2046 23874 2098 23886
rect 9886 23874 9938 23886
rect 12350 23938 12402 23950
rect 14254 23938 14306 23950
rect 19406 23938 19458 23950
rect 13122 23886 13134 23938
rect 13186 23886 13198 23938
rect 13682 23886 13694 23938
rect 13746 23886 13758 23938
rect 14914 23886 14926 23938
rect 14978 23886 14990 23938
rect 15922 23886 15934 23938
rect 15986 23886 15998 23938
rect 18386 23886 18398 23938
rect 18450 23886 18462 23938
rect 26226 23886 26238 23938
rect 26290 23886 26302 23938
rect 12350 23874 12402 23886
rect 14254 23874 14306 23886
rect 19406 23874 19458 23886
rect 4622 23826 4674 23838
rect 12798 23826 12850 23838
rect 27246 23826 27298 23838
rect 4050 23774 4062 23826
rect 4114 23774 4126 23826
rect 10770 23774 10782 23826
rect 10834 23774 10846 23826
rect 19842 23774 19854 23826
rect 19906 23774 19918 23826
rect 4622 23762 4674 23774
rect 12798 23762 12850 23774
rect 27246 23762 27298 23774
rect 16830 23714 16882 23726
rect 16830 23650 16882 23662
rect 25678 23714 25730 23726
rect 25678 23650 25730 23662
rect 672 23546 27888 23580
rect 672 23494 3806 23546
rect 3858 23494 3910 23546
rect 3962 23494 4014 23546
rect 4066 23494 23806 23546
rect 23858 23494 23910 23546
rect 23962 23494 24014 23546
rect 24066 23494 27888 23546
rect 672 23460 27888 23494
rect 3838 23378 3890 23390
rect 27246 23378 27298 23390
rect 11666 23326 11678 23378
rect 11730 23326 11742 23378
rect 3838 23314 3890 23326
rect 27246 23314 27298 23326
rect 1150 23266 1202 23278
rect 1150 23202 1202 23214
rect 6190 23266 6242 23278
rect 16942 23266 16994 23278
rect 6738 23214 6750 23266
rect 6802 23214 6814 23266
rect 18946 23214 18958 23266
rect 19010 23214 19022 23266
rect 6190 23202 6242 23214
rect 16942 23202 16994 23214
rect 1586 23102 1598 23154
rect 1650 23102 1662 23154
rect 2146 23102 2158 23154
rect 2210 23102 2222 23154
rect 8978 23102 8990 23154
rect 9042 23102 9054 23154
rect 11442 23102 11454 23154
rect 11506 23102 11518 23154
rect 13122 23102 13134 23154
rect 13186 23102 13198 23154
rect 13682 23102 13694 23154
rect 13746 23102 13758 23154
rect 14354 23102 14366 23154
rect 14418 23102 14430 23154
rect 14802 23102 14814 23154
rect 14866 23102 14878 23154
rect 15922 23102 15934 23154
rect 15986 23102 15998 23154
rect 26338 23102 26350 23154
rect 26402 23102 26414 23154
rect 5630 23042 5682 23054
rect 10558 23042 10610 23054
rect 12238 23042 12290 23054
rect 2706 22990 2718 23042
rect 2770 22990 2782 23042
rect 9426 22990 9438 23042
rect 9490 22990 9502 23042
rect 12002 22990 12014 23042
rect 12066 22990 12078 23042
rect 5630 22978 5682 22990
rect 10558 22978 10610 22990
rect 12238 22978 12290 22990
rect 12798 23042 12850 23054
rect 13794 22990 13806 23042
rect 13858 22990 13870 23042
rect 18498 22990 18510 23042
rect 18562 22990 18574 23042
rect 12798 22978 12850 22990
rect 8318 22930 8370 22942
rect 16382 22930 16434 22942
rect 7186 22878 7198 22930
rect 7250 22878 7262 22930
rect 11778 22878 11790 22930
rect 11842 22878 11854 22930
rect 8318 22866 8370 22878
rect 16382 22866 16434 22878
rect 17390 22930 17442 22942
rect 17390 22866 17442 22878
rect 672 22762 27888 22796
rect 672 22710 4466 22762
rect 4518 22710 4570 22762
rect 4622 22710 4674 22762
rect 4726 22710 24466 22762
rect 24518 22710 24570 22762
rect 24622 22710 24674 22762
rect 24726 22710 27888 22762
rect 672 22676 27888 22710
rect 1150 22594 1202 22606
rect 2706 22542 2718 22594
rect 2770 22542 2782 22594
rect 5954 22542 5966 22594
rect 6018 22542 6030 22594
rect 9874 22542 9886 22594
rect 9938 22542 9950 22594
rect 15138 22542 15150 22594
rect 15202 22542 15214 22594
rect 1150 22530 1202 22542
rect 10334 22482 10386 22494
rect 10334 22418 10386 22430
rect 14702 22482 14754 22494
rect 18610 22430 18622 22482
rect 18674 22430 18686 22482
rect 26226 22430 26238 22482
rect 26290 22430 26302 22482
rect 14702 22418 14754 22430
rect 6414 22370 6466 22382
rect 16830 22370 16882 22382
rect 2258 22318 2270 22370
rect 2322 22318 2334 22370
rect 5282 22318 5294 22370
rect 5346 22318 5358 22370
rect 5842 22318 5854 22370
rect 5906 22318 5918 22370
rect 6962 22318 6974 22370
rect 7026 22318 7038 22370
rect 8082 22318 8094 22370
rect 8146 22318 8158 22370
rect 9202 22318 9214 22370
rect 9266 22318 9278 22370
rect 9650 22318 9662 22370
rect 9714 22318 9726 22370
rect 11106 22318 11118 22370
rect 11170 22318 11182 22370
rect 11890 22318 11902 22370
rect 11954 22318 11966 22370
rect 13010 22318 13022 22370
rect 13074 22318 13086 22370
rect 13906 22318 13918 22370
rect 13970 22318 13982 22370
rect 15250 22318 15262 22370
rect 15314 22318 15326 22370
rect 15810 22318 15822 22370
rect 15874 22318 15886 22370
rect 24882 22318 24894 22370
rect 24946 22318 24958 22370
rect 6414 22306 6466 22318
rect 16830 22306 16882 22318
rect 4958 22258 5010 22270
rect 1586 22206 1598 22258
rect 1650 22206 1662 22258
rect 4958 22194 5010 22206
rect 8878 22258 8930 22270
rect 8878 22194 8930 22206
rect 16158 22258 16210 22270
rect 27246 22258 27298 22270
rect 18946 22206 18958 22258
rect 19010 22206 19022 22258
rect 16158 22194 16210 22206
rect 27246 22194 27298 22206
rect 3838 22146 3890 22158
rect 3838 22082 3890 22094
rect 16718 22146 16770 22158
rect 16718 22082 16770 22094
rect 17390 22146 17442 22158
rect 17390 22082 17442 22094
rect 25678 22146 25730 22158
rect 25678 22082 25730 22094
rect 672 21978 27888 22012
rect 672 21926 3806 21978
rect 3858 21926 3910 21978
rect 3962 21926 4014 21978
rect 4066 21926 23806 21978
rect 23858 21926 23910 21978
rect 23962 21926 24014 21978
rect 24066 21926 27888 21978
rect 672 21892 27888 21926
rect 4286 21810 4338 21822
rect 4286 21746 4338 21758
rect 11678 21810 11730 21822
rect 11678 21746 11730 21758
rect 12798 21810 12850 21822
rect 12798 21746 12850 21758
rect 13134 21810 13186 21822
rect 13134 21746 13186 21758
rect 27246 21810 27298 21822
rect 27246 21746 27298 21758
rect 1698 21646 1710 21698
rect 1762 21646 1774 21698
rect 5506 21646 5518 21698
rect 5570 21646 5582 21698
rect 18722 21646 18734 21698
rect 18786 21646 18798 21698
rect 2706 21534 2718 21586
rect 2770 21534 2782 21586
rect 6738 21534 6750 21586
rect 6802 21534 6814 21586
rect 7074 21534 7086 21586
rect 7138 21534 7150 21586
rect 7858 21534 7870 21586
rect 7922 21534 7934 21586
rect 8530 21534 8542 21586
rect 8594 21534 8606 21586
rect 9426 21534 9438 21586
rect 9490 21534 9502 21586
rect 10098 21534 10110 21586
rect 10162 21534 10174 21586
rect 13570 21534 13582 21586
rect 13634 21534 13646 21586
rect 14466 21534 14478 21586
rect 14530 21534 14542 21586
rect 15810 21534 15822 21586
rect 15874 21534 15886 21586
rect 16370 21534 16382 21586
rect 16434 21534 16446 21586
rect 6302 21474 6354 21486
rect 12238 21474 12290 21486
rect 3042 21422 3054 21474
rect 3106 21422 3118 21474
rect 10434 21422 10446 21474
rect 10498 21422 10510 21474
rect 6302 21410 6354 21422
rect 12238 21410 12290 21422
rect 15262 21474 15314 21486
rect 15262 21410 15314 21422
rect 16718 21474 16770 21486
rect 16718 21410 16770 21422
rect 17166 21474 17218 21486
rect 19294 21474 19346 21486
rect 18274 21422 18286 21474
rect 18338 21422 18350 21474
rect 26226 21422 26238 21474
rect 26290 21422 26302 21474
rect 17166 21410 17218 21422
rect 19294 21410 19346 21422
rect 2158 21362 2210 21374
rect 2158 21298 2210 21310
rect 5966 21362 6018 21374
rect 12126 21362 12178 21374
rect 7298 21310 7310 21362
rect 7362 21310 7374 21362
rect 5966 21298 6018 21310
rect 12126 21298 12178 21310
rect 12910 21362 12962 21374
rect 19854 21362 19906 21374
rect 15698 21310 15710 21362
rect 15762 21310 15774 21362
rect 12910 21298 12962 21310
rect 19854 21298 19906 21310
rect 672 21194 27888 21228
rect 672 21142 4466 21194
rect 4518 21142 4570 21194
rect 4622 21142 4674 21194
rect 4726 21142 24466 21194
rect 24518 21142 24570 21194
rect 24622 21142 24674 21194
rect 24726 21142 27888 21194
rect 672 21108 27888 21142
rect 1374 21026 1426 21038
rect 7870 21026 7922 21038
rect 3266 20974 3278 21026
rect 3330 20974 3342 21026
rect 1374 20962 1426 20974
rect 7870 20962 7922 20974
rect 9774 21026 9826 21038
rect 9774 20962 9826 20974
rect 17614 21026 17666 21038
rect 19854 21026 19906 21038
rect 18722 20974 18734 21026
rect 18786 20974 18798 21026
rect 17614 20962 17666 20974
rect 19854 20962 19906 20974
rect 1934 20914 1986 20926
rect 1934 20850 1986 20862
rect 2270 20914 2322 20926
rect 2270 20850 2322 20862
rect 3726 20914 3778 20926
rect 9550 20914 9602 20926
rect 6738 20862 6750 20914
rect 6802 20862 6814 20914
rect 13906 20862 13918 20914
rect 13970 20862 13982 20914
rect 20402 20862 20414 20914
rect 20466 20862 20478 20914
rect 20738 20862 20750 20914
rect 20802 20862 20814 20914
rect 3726 20850 3778 20862
rect 9550 20850 9602 20862
rect 9886 20802 9938 20814
rect 2594 20750 2606 20802
rect 2658 20750 2670 20802
rect 3042 20750 3054 20802
rect 3106 20750 3118 20802
rect 4498 20750 4510 20802
rect 4562 20750 4574 20802
rect 5282 20750 5294 20802
rect 5346 20750 5358 20802
rect 9886 20738 9938 20750
rect 9998 20802 10050 20814
rect 9998 20738 10050 20750
rect 10446 20802 10498 20814
rect 14590 20802 14642 20814
rect 20190 20802 20242 20814
rect 10994 20750 11006 20802
rect 11058 20750 11070 20802
rect 11554 20750 11566 20802
rect 11618 20750 11630 20802
rect 11890 20750 11902 20802
rect 11954 20750 11966 20802
rect 13346 20750 13358 20802
rect 13410 20750 13422 20802
rect 13794 20750 13806 20802
rect 13858 20750 13870 20802
rect 14914 20750 14926 20802
rect 14978 20750 14990 20802
rect 15922 20750 15934 20802
rect 15986 20750 15998 20802
rect 16706 20750 16718 20802
rect 16770 20750 16782 20802
rect 19170 20750 19182 20802
rect 19234 20750 19246 20802
rect 10446 20738 10498 20750
rect 14590 20738 14642 20750
rect 20190 20738 20242 20750
rect 12910 20690 12962 20702
rect 6290 20638 6302 20690
rect 6354 20638 6366 20690
rect 11778 20638 11790 20690
rect 11842 20638 11854 20690
rect 12910 20626 12962 20638
rect 16718 20578 16770 20590
rect 10770 20526 10782 20578
rect 10834 20526 10846 20578
rect 16718 20514 16770 20526
rect 17054 20578 17106 20590
rect 17054 20514 17106 20526
rect 672 20410 27888 20444
rect 672 20358 3806 20410
rect 3858 20358 3910 20410
rect 3962 20358 4014 20410
rect 4066 20358 23806 20410
rect 23858 20358 23910 20410
rect 23962 20358 24014 20410
rect 24066 20358 27888 20410
rect 672 20324 27888 20358
rect 2830 20242 2882 20254
rect 2830 20178 2882 20190
rect 12910 20242 12962 20254
rect 16034 20190 16046 20242
rect 16098 20190 16110 20242
rect 12910 20178 12962 20190
rect 8318 20130 8370 20142
rect 10558 20130 10610 20142
rect 6738 20078 6750 20130
rect 6802 20078 6814 20130
rect 8978 20078 8990 20130
rect 9042 20078 9054 20130
rect 8318 20066 8370 20078
rect 10558 20066 10610 20078
rect 13246 20130 13298 20142
rect 19742 20130 19794 20142
rect 15026 20078 15038 20130
rect 15090 20078 15102 20130
rect 18162 20078 18174 20130
rect 18226 20078 18238 20130
rect 13246 20066 13298 20078
rect 19742 20066 19794 20078
rect 11454 20018 11506 20030
rect 1250 19966 1262 20018
rect 1314 19966 1326 20018
rect 3602 19966 3614 20018
rect 3666 19966 3678 20018
rect 8866 19966 8878 20018
rect 8930 19966 8942 20018
rect 11454 19954 11506 19966
rect 11902 20018 11954 20030
rect 15486 20018 15538 20030
rect 12226 19966 12238 20018
rect 12290 19966 12302 20018
rect 14690 19966 14702 20018
rect 14754 19966 14766 20018
rect 11902 19954 11954 19966
rect 15486 19954 15538 19966
rect 15822 20018 15874 20030
rect 16258 19966 16270 20018
rect 16322 19966 16334 20018
rect 15822 19954 15874 19966
rect 6190 19906 6242 19918
rect 1026 19854 1038 19906
rect 1090 19854 1102 19906
rect 9314 19854 9326 19906
rect 9378 19854 9390 19906
rect 11666 19854 11678 19906
rect 11730 19854 11742 19906
rect 13458 19854 13470 19906
rect 13522 19854 13534 19906
rect 13794 19854 13806 19906
rect 13858 19854 13870 19906
rect 18498 19854 18510 19906
rect 18562 19854 18574 19906
rect 6190 19842 6242 19854
rect 1598 19794 1650 19806
rect 1598 19730 1650 19742
rect 5630 19794 5682 19806
rect 15598 19794 15650 19806
rect 7186 19742 7198 19794
rect 7250 19742 7262 19794
rect 11778 19742 11790 19794
rect 11842 19742 11854 19794
rect 5630 19730 5682 19742
rect 15598 19730 15650 19742
rect 672 19626 27888 19660
rect 672 19574 4466 19626
rect 4518 19574 4570 19626
rect 4622 19574 4674 19626
rect 4726 19574 24466 19626
rect 24518 19574 24570 19626
rect 24622 19574 24674 19626
rect 24726 19574 27888 19626
rect 672 19540 27888 19574
rect 1598 19458 1650 19470
rect 1598 19394 1650 19406
rect 5742 19458 5794 19470
rect 5742 19394 5794 19406
rect 8206 19458 8258 19470
rect 11554 19406 11566 19458
rect 11618 19406 11630 19458
rect 8206 19394 8258 19406
rect 11118 19346 11170 19358
rect 2706 19294 2718 19346
rect 2770 19294 2782 19346
rect 4498 19294 4510 19346
rect 4562 19294 4574 19346
rect 6962 19294 6974 19346
rect 7026 19294 7038 19346
rect 11118 19282 11170 19294
rect 12574 19346 12626 19358
rect 14366 19346 14418 19358
rect 13906 19294 13918 19346
rect 13970 19294 13982 19346
rect 12574 19282 12626 19294
rect 14366 19282 14418 19294
rect 16718 19346 16770 19358
rect 16718 19282 16770 19294
rect 16942 19346 16994 19358
rect 16942 19282 16994 19294
rect 12910 19234 12962 19246
rect 6626 19182 6638 19234
rect 6690 19182 6702 19234
rect 9538 19182 9550 19234
rect 9602 19182 9614 19234
rect 10322 19182 10334 19234
rect 10386 19182 10398 19234
rect 11778 19182 11790 19234
rect 11842 19182 11854 19234
rect 12114 19182 12126 19234
rect 12178 19182 12190 19234
rect 13346 19182 13358 19234
rect 13410 19182 13422 19234
rect 13794 19182 13806 19234
rect 13858 19182 13870 19234
rect 14914 19182 14926 19234
rect 14978 19182 14990 19234
rect 16034 19182 16046 19234
rect 16098 19182 16110 19234
rect 12910 19170 12962 19182
rect 16830 19122 16882 19134
rect 3154 19070 3166 19122
rect 3218 19070 3230 19122
rect 4162 19070 4174 19122
rect 4226 19070 4238 19122
rect 16830 19058 16882 19070
rect 672 18842 27888 18876
rect 672 18790 3806 18842
rect 3858 18790 3910 18842
rect 3962 18790 4014 18842
rect 4066 18790 23806 18842
rect 23858 18790 23910 18842
rect 23962 18790 24014 18842
rect 24066 18790 27888 18842
rect 672 18756 27888 18790
rect 7198 18674 7250 18686
rect 7198 18610 7250 18622
rect 13806 18674 13858 18686
rect 13806 18610 13858 18622
rect 15822 18674 15874 18686
rect 15822 18610 15874 18622
rect 3166 18562 3218 18574
rect 16046 18562 16098 18574
rect 4274 18510 4286 18562
rect 4338 18510 4350 18562
rect 10322 18510 10334 18562
rect 10386 18510 10398 18562
rect 16258 18510 16270 18562
rect 16322 18510 16334 18562
rect 3166 18498 3218 18510
rect 16046 18498 16098 18510
rect 15598 18450 15650 18462
rect 1474 18398 1486 18450
rect 1538 18398 1550 18450
rect 2258 18398 2270 18450
rect 2322 18398 2334 18450
rect 2706 18398 2718 18450
rect 2770 18398 2782 18450
rect 3938 18398 3950 18450
rect 4002 18398 4014 18450
rect 5618 18398 5630 18450
rect 5682 18398 5694 18450
rect 8082 18398 8094 18450
rect 8146 18398 8158 18450
rect 14578 18398 14590 18450
rect 14642 18398 14654 18450
rect 15598 18386 15650 18398
rect 19518 18450 19570 18462
rect 19518 18386 19570 18398
rect 15262 18338 15314 18350
rect 5954 18286 5966 18338
rect 6018 18286 6030 18338
rect 8418 18286 8430 18338
rect 8482 18286 8494 18338
rect 14354 18286 14366 18338
rect 14418 18286 14430 18338
rect 15262 18274 15314 18286
rect 1710 18226 1762 18238
rect 1710 18162 1762 18174
rect 9662 18226 9714 18238
rect 11902 18226 11954 18238
rect 10770 18174 10782 18226
rect 10834 18174 10846 18226
rect 9662 18162 9714 18174
rect 11902 18162 11954 18174
rect 13470 18226 13522 18238
rect 13470 18162 13522 18174
rect 15150 18226 15202 18238
rect 15150 18162 15202 18174
rect 16270 18226 16322 18238
rect 16270 18162 16322 18174
rect 16494 18226 16546 18238
rect 16494 18162 16546 18174
rect 16942 18226 16994 18238
rect 16942 18162 16994 18174
rect 17054 18226 17106 18238
rect 17054 18162 17106 18174
rect 17166 18226 17218 18238
rect 17166 18162 17218 18174
rect 17390 18226 17442 18238
rect 17390 18162 17442 18174
rect 18958 18226 19010 18238
rect 18958 18162 19010 18174
rect 672 18058 27888 18092
rect 672 18006 4466 18058
rect 4518 18006 4570 18058
rect 4622 18006 4674 18058
rect 4726 18006 24466 18058
rect 24518 18006 24570 18058
rect 24622 18006 24674 18058
rect 24726 18006 27888 18058
rect 672 17972 27888 18006
rect 1038 17890 1090 17902
rect 11230 17890 11282 17902
rect 16046 17890 16098 17902
rect 4834 17838 4846 17890
rect 4898 17838 4910 17890
rect 14466 17838 14478 17890
rect 14530 17838 14542 17890
rect 1038 17826 1090 17838
rect 11230 17826 11282 17838
rect 16046 17826 16098 17838
rect 2594 17726 2606 17778
rect 2658 17726 2670 17778
rect 6962 17726 6974 17778
rect 7026 17726 7038 17778
rect 9986 17726 9998 17778
rect 10050 17726 10062 17778
rect 3726 17666 3778 17678
rect 13806 17666 13858 17678
rect 2034 17614 2046 17666
rect 2098 17614 2110 17666
rect 4274 17614 4286 17666
rect 4338 17614 4350 17666
rect 6626 17614 6638 17666
rect 6690 17614 6702 17666
rect 9538 17614 9550 17666
rect 9602 17614 9614 17666
rect 12338 17614 12350 17666
rect 12402 17614 12414 17666
rect 13234 17614 13246 17666
rect 13298 17614 13310 17666
rect 3726 17602 3778 17614
rect 13806 17602 13858 17614
rect 14030 17666 14082 17678
rect 14690 17614 14702 17666
rect 14754 17614 14766 17666
rect 15026 17614 15038 17666
rect 15090 17614 15102 17666
rect 14030 17602 14082 17614
rect 1598 17554 1650 17566
rect 15486 17554 15538 17566
rect 4386 17502 4398 17554
rect 4450 17502 4462 17554
rect 9650 17502 9662 17554
rect 9714 17502 9726 17554
rect 16146 17502 16158 17554
rect 16210 17502 16222 17554
rect 1598 17490 1650 17502
rect 15486 17490 15538 17502
rect 5966 17442 6018 17454
rect 5966 17378 6018 17390
rect 8206 17442 8258 17454
rect 8206 17378 8258 17390
rect 15822 17442 15874 17454
rect 15822 17378 15874 17390
rect 672 17274 27888 17308
rect 672 17222 3806 17274
rect 3858 17222 3910 17274
rect 3962 17222 4014 17274
rect 4066 17222 23806 17274
rect 23858 17222 23910 17274
rect 23962 17222 24014 17274
rect 24066 17222 27888 17274
rect 672 17188 27888 17222
rect 12798 17106 12850 17118
rect 12798 17042 12850 17054
rect 13134 17106 13186 17118
rect 13134 17042 13186 17054
rect 14254 17106 14306 17118
rect 14254 17042 14306 17054
rect 1038 16994 1090 17006
rect 1038 16930 1090 16942
rect 2494 16994 2546 17006
rect 2494 16930 2546 16942
rect 8318 16994 8370 17006
rect 14926 16994 14978 17006
rect 10210 16942 10222 16994
rect 10274 16942 10286 16994
rect 12114 16942 12126 16994
rect 12178 16942 12190 16994
rect 8318 16930 8370 16942
rect 14926 16930 14978 16942
rect 3838 16882 3890 16894
rect 10894 16882 10946 16894
rect 1474 16830 1486 16882
rect 1538 16830 1550 16882
rect 4946 16830 4958 16882
rect 5010 16830 5022 16882
rect 6626 16830 6638 16882
rect 6690 16830 6702 16882
rect 10546 16830 10558 16882
rect 10610 16830 10622 16882
rect 3838 16818 3890 16830
rect 10894 16818 10946 16830
rect 11006 16882 11058 16894
rect 13806 16882 13858 16894
rect 16382 16882 16434 16894
rect 11778 16830 11790 16882
rect 11842 16830 11854 16882
rect 14018 16830 14030 16882
rect 14082 16830 14094 16882
rect 14354 16830 14366 16882
rect 14418 16830 14430 16882
rect 15250 16830 15262 16882
rect 15314 16830 15326 16882
rect 15698 16830 15710 16882
rect 15762 16830 15774 16882
rect 16930 16830 16942 16882
rect 16994 16830 17006 16882
rect 17938 16830 17950 16882
rect 18002 16830 18014 16882
rect 11006 16818 11058 16830
rect 13806 16818 13858 16830
rect 16382 16818 16434 16830
rect 9886 16770 9938 16782
rect 7074 16718 7086 16770
rect 7138 16718 7150 16770
rect 9886 16706 9938 16718
rect 10110 16770 10162 16782
rect 10110 16706 10162 16718
rect 11342 16770 11394 16782
rect 11342 16706 11394 16718
rect 12910 16770 12962 16782
rect 15922 16718 15934 16770
rect 15986 16718 15998 16770
rect 12910 16706 12962 16718
rect 1934 16658 1986 16670
rect 1934 16594 1986 16606
rect 4398 16658 4450 16670
rect 4398 16594 4450 16606
rect 5518 16658 5570 16670
rect 5518 16594 5570 16606
rect 11230 16658 11282 16670
rect 11230 16594 11282 16606
rect 14590 16658 14642 16670
rect 14590 16594 14642 16606
rect 672 16490 27888 16524
rect 672 16438 4466 16490
rect 4518 16438 4570 16490
rect 4622 16438 4674 16490
rect 4726 16438 24466 16490
rect 24518 16438 24570 16490
rect 24622 16438 24674 16490
rect 24726 16438 27888 16490
rect 672 16404 27888 16438
rect 10110 16322 10162 16334
rect 3042 16270 3054 16322
rect 3106 16270 3118 16322
rect 4722 16270 4734 16322
rect 4786 16270 4798 16322
rect 11778 16270 11790 16322
rect 11842 16270 11854 16322
rect 17938 16270 17950 16322
rect 18002 16270 18014 16322
rect 10110 16258 10162 16270
rect 9550 16210 9602 16222
rect 6850 16158 6862 16210
rect 6914 16158 6926 16210
rect 9550 16146 9602 16158
rect 10334 16210 10386 16222
rect 10334 16146 10386 16158
rect 12238 16210 12290 16222
rect 12238 16146 12290 16158
rect 15262 16210 15314 16222
rect 15262 16146 15314 16158
rect 15710 16210 15762 16222
rect 15710 16146 15762 16158
rect 9886 16098 9938 16110
rect 3602 16046 3614 16098
rect 3666 16046 3678 16098
rect 4162 16046 4174 16098
rect 4226 16046 4238 16098
rect 6514 16046 6526 16098
rect 6578 16046 6590 16098
rect 9090 16046 9102 16098
rect 9154 16046 9166 16098
rect 9314 16046 9326 16098
rect 9378 16046 9390 16098
rect 9886 16034 9938 16046
rect 9998 16098 10050 16110
rect 16270 16098 16322 16110
rect 11106 16046 11118 16098
rect 11170 16046 11182 16098
rect 11666 16046 11678 16098
rect 11730 16046 11742 16098
rect 13010 16046 13022 16098
rect 13074 16046 13086 16098
rect 13906 16046 13918 16098
rect 13970 16046 13982 16098
rect 15922 16046 15934 16098
rect 15986 16046 15998 16098
rect 18386 16046 18398 16098
rect 18450 16046 18462 16098
rect 9998 16034 10050 16046
rect 16270 16034 16322 16046
rect 8094 15986 8146 15998
rect 8094 15922 8146 15934
rect 10782 15986 10834 15998
rect 10782 15922 10834 15934
rect 1934 15874 1986 15886
rect 1934 15810 1986 15822
rect 5854 15874 5906 15886
rect 5854 15810 5906 15822
rect 9662 15874 9714 15886
rect 9662 15810 9714 15822
rect 15374 15874 15426 15886
rect 15374 15810 15426 15822
rect 16046 15874 16098 15886
rect 16046 15810 16098 15822
rect 16830 15874 16882 15886
rect 16830 15810 16882 15822
rect 672 15706 27888 15740
rect 672 15654 3806 15706
rect 3858 15654 3910 15706
rect 3962 15654 4014 15706
rect 4066 15654 23806 15706
rect 23858 15654 23910 15706
rect 23962 15654 24014 15706
rect 24066 15654 27888 15706
rect 672 15620 27888 15654
rect 11230 15538 11282 15550
rect 11230 15474 11282 15486
rect 11902 15538 11954 15550
rect 11902 15474 11954 15486
rect 9550 15426 9602 15438
rect 3490 15374 3502 15426
rect 3554 15374 3566 15426
rect 5730 15374 5742 15426
rect 5794 15374 5806 15426
rect 9550 15362 9602 15374
rect 11006 15426 11058 15438
rect 11006 15362 11058 15374
rect 15262 15426 15314 15438
rect 16482 15374 16494 15426
rect 16546 15374 16558 15426
rect 18498 15374 18510 15426
rect 18562 15374 18574 15426
rect 15262 15362 15314 15374
rect 10110 15314 10162 15326
rect 7858 15262 7870 15314
rect 7922 15262 7934 15314
rect 10110 15250 10162 15262
rect 10558 15314 10610 15326
rect 10558 15250 10610 15262
rect 11454 15314 11506 15326
rect 11454 15250 11506 15262
rect 11790 15314 11842 15326
rect 11790 15250 11842 15262
rect 13694 15314 13746 15326
rect 13694 15250 13746 15262
rect 15150 15314 15202 15326
rect 15150 15250 15202 15262
rect 15822 15314 15874 15326
rect 15822 15250 15874 15262
rect 16046 15314 16098 15326
rect 16046 15250 16098 15262
rect 10782 15202 10834 15214
rect 3154 15150 3166 15202
rect 3218 15150 3230 15202
rect 6066 15150 6078 15202
rect 6130 15150 6142 15202
rect 8306 15150 8318 15202
rect 8370 15150 8382 15202
rect 10782 15138 10834 15150
rect 11902 15202 11954 15214
rect 11902 15138 11954 15150
rect 14926 15202 14978 15214
rect 14926 15138 14978 15150
rect 15934 15202 15986 15214
rect 15934 15138 15986 15150
rect 16942 15202 16994 15214
rect 18050 15150 18062 15202
rect 18114 15150 18126 15202
rect 16942 15138 16994 15150
rect 1934 15090 1986 15102
rect 1934 15026 1986 15038
rect 7310 15090 7362 15102
rect 7310 15026 7362 15038
rect 9998 15090 10050 15102
rect 9998 15026 10050 15038
rect 10670 15090 10722 15102
rect 10670 15026 10722 15038
rect 13358 15090 13410 15102
rect 13358 15026 13410 15038
rect 15374 15090 15426 15102
rect 15374 15026 15426 15038
rect 672 14922 27888 14956
rect 672 14870 4466 14922
rect 4518 14870 4570 14922
rect 4622 14870 4674 14922
rect 4726 14870 24466 14922
rect 24518 14870 24570 14922
rect 24622 14870 24674 14922
rect 24726 14870 27888 14922
rect 672 14836 27888 14870
rect 1934 14754 1986 14766
rect 1934 14690 1986 14702
rect 2830 14754 2882 14766
rect 2830 14690 2882 14702
rect 9438 14754 9490 14766
rect 9438 14690 9490 14702
rect 11118 14754 11170 14766
rect 11118 14690 11170 14702
rect 11230 14754 11282 14766
rect 15486 14754 15538 14766
rect 14354 14702 14366 14754
rect 14418 14702 14430 14754
rect 11230 14690 11282 14702
rect 15486 14690 15538 14702
rect 16270 14754 16322 14766
rect 16270 14690 16322 14702
rect 17614 14754 17666 14766
rect 17614 14690 17666 14702
rect 4510 14642 4562 14654
rect 5966 14642 6018 14654
rect 5506 14590 5518 14642
rect 5570 14590 5582 14642
rect 4510 14578 4562 14590
rect 5966 14578 6018 14590
rect 9550 14642 9602 14654
rect 9550 14578 9602 14590
rect 10110 14642 10162 14654
rect 10110 14578 10162 14590
rect 10222 14642 10274 14654
rect 10222 14578 10274 14590
rect 15934 14642 15986 14654
rect 15934 14578 15986 14590
rect 16046 14642 16098 14654
rect 16046 14578 16098 14590
rect 9998 14530 10050 14542
rect 16718 14530 16770 14542
rect 4834 14478 4846 14530
rect 4898 14478 4910 14530
rect 5282 14478 5294 14530
rect 5346 14478 5358 14530
rect 6514 14478 6526 14530
rect 6578 14478 6590 14530
rect 7634 14478 7646 14530
rect 7698 14478 7710 14530
rect 10658 14478 10670 14530
rect 10722 14478 10734 14530
rect 9998 14466 10050 14478
rect 16718 14466 16770 14478
rect 17166 14530 17218 14542
rect 17166 14466 17218 14478
rect 17390 14530 17442 14542
rect 17390 14466 17442 14478
rect 2494 14418 2546 14430
rect 3266 14366 3278 14418
rect 3330 14366 3342 14418
rect 13906 14366 13918 14418
rect 13970 14366 13982 14418
rect 17490 14366 17502 14418
rect 17554 14366 17566 14418
rect 2494 14354 2546 14366
rect 9438 14306 9490 14318
rect 9438 14242 9490 14254
rect 11006 14306 11058 14318
rect 11006 14242 11058 14254
rect 16942 14306 16994 14318
rect 16942 14242 16994 14254
rect 672 14138 27888 14172
rect 672 14086 3806 14138
rect 3858 14086 3910 14138
rect 3962 14086 4014 14138
rect 4066 14086 23806 14138
rect 23858 14086 23910 14138
rect 23962 14086 24014 14138
rect 24066 14086 27888 14138
rect 672 14052 27888 14086
rect 7422 13970 7474 13982
rect 7422 13906 7474 13918
rect 16942 13970 16994 13982
rect 16942 13906 16994 13918
rect 17278 13970 17330 13982
rect 17278 13906 17330 13918
rect 17390 13970 17442 13982
rect 17390 13906 17442 13918
rect 1150 13858 1202 13870
rect 1150 13794 1202 13806
rect 16382 13858 16434 13870
rect 16382 13794 16434 13806
rect 2606 13746 2658 13758
rect 16046 13746 16098 13758
rect 1586 13694 1598 13746
rect 1650 13694 1662 13746
rect 1922 13694 1934 13746
rect 1986 13694 1998 13746
rect 3378 13694 3390 13746
rect 3442 13694 3454 13746
rect 4274 13694 4286 13746
rect 4338 13694 4350 13746
rect 5170 13694 5182 13746
rect 5234 13694 5246 13746
rect 8194 13694 8206 13746
rect 8258 13694 8270 13746
rect 9314 13694 9326 13746
rect 9378 13694 9390 13746
rect 13122 13694 13134 13746
rect 13186 13694 13198 13746
rect 15698 13694 15710 13746
rect 15762 13694 15774 13746
rect 2606 13682 2658 13694
rect 16046 13682 16098 13694
rect 16158 13746 16210 13758
rect 16158 13682 16210 13694
rect 16494 13746 16546 13758
rect 16494 13682 16546 13694
rect 17054 13746 17106 13758
rect 17054 13682 17106 13694
rect 15262 13634 15314 13646
rect 5618 13582 5630 13634
rect 5682 13582 5694 13634
rect 9762 13582 9774 13634
rect 9826 13582 9838 13634
rect 13682 13582 13694 13634
rect 13746 13582 13758 13634
rect 15262 13570 15314 13582
rect 15374 13634 15426 13646
rect 15374 13570 15426 13582
rect 6750 13522 6802 13534
rect 2146 13470 2158 13522
rect 2210 13470 2222 13522
rect 6750 13458 6802 13470
rect 11006 13522 11058 13534
rect 11006 13458 11058 13470
rect 14814 13522 14866 13534
rect 14814 13458 14866 13470
rect 672 13354 27888 13388
rect 672 13302 4466 13354
rect 4518 13302 4570 13354
rect 4622 13302 4674 13354
rect 4726 13302 24466 13354
rect 24518 13302 24570 13354
rect 24622 13302 24674 13354
rect 24726 13302 27888 13354
rect 672 13268 27888 13302
rect 7758 13186 7810 13198
rect 2594 13134 2606 13186
rect 2658 13134 2670 13186
rect 7758 13122 7810 13134
rect 15374 13186 15426 13198
rect 15374 13122 15426 13134
rect 16046 13186 16098 13198
rect 16046 13122 16098 13134
rect 3726 13074 3778 13086
rect 11902 13074 11954 13086
rect 5170 13022 5182 13074
rect 5234 13022 5246 13074
rect 9426 13022 9438 13074
rect 9490 13022 9502 13074
rect 3726 13010 3778 13022
rect 11902 13010 11954 13022
rect 14478 13074 14530 13086
rect 14478 13010 14530 13022
rect 14814 13074 14866 13086
rect 14814 13010 14866 13022
rect 15262 13074 15314 13086
rect 15262 13010 15314 13022
rect 16158 13074 16210 13086
rect 16158 13010 16210 13022
rect 5854 12962 5906 12974
rect 11342 12962 11394 12974
rect 2146 12910 2158 12962
rect 2210 12910 2222 12962
rect 4498 12910 4510 12962
rect 4562 12910 4574 12962
rect 4946 12910 4958 12962
rect 5010 12910 5022 12962
rect 6402 12910 6414 12962
rect 6466 12910 6478 12962
rect 7186 12910 7198 12962
rect 7250 12910 7262 12962
rect 5854 12898 5906 12910
rect 11342 12898 11394 12910
rect 12238 12962 12290 12974
rect 12238 12898 12290 12910
rect 12798 12962 12850 12974
rect 12798 12898 12850 12910
rect 4174 12850 4226 12862
rect 15486 12850 15538 12862
rect 8194 12798 8206 12850
rect 8258 12798 8270 12850
rect 9090 12798 9102 12850
rect 9154 12798 9166 12850
rect 4174 12786 4226 12798
rect 15486 12786 15538 12798
rect 10670 12738 10722 12750
rect 10670 12674 10722 12686
rect 672 12570 27888 12604
rect 672 12518 3806 12570
rect 3858 12518 3910 12570
rect 3962 12518 4014 12570
rect 4066 12518 23806 12570
rect 23858 12518 23910 12570
rect 23962 12518 24014 12570
rect 24066 12518 27888 12570
rect 672 12484 27888 12518
rect 1598 12290 1650 12302
rect 1598 12226 1650 12238
rect 2494 12290 2546 12302
rect 5966 12290 6018 12302
rect 3266 12238 3278 12290
rect 3330 12238 3342 12290
rect 2494 12226 2546 12238
rect 5966 12226 6018 12238
rect 12798 12290 12850 12302
rect 12798 12226 12850 12238
rect 2830 12178 2882 12190
rect 8542 12178 8594 12190
rect 10670 12178 10722 12190
rect 1138 12126 1150 12178
rect 1202 12126 1214 12178
rect 2034 12126 2046 12178
rect 2098 12126 2110 12178
rect 5506 12126 5518 12178
rect 5570 12126 5582 12178
rect 6850 12126 6862 12178
rect 6914 12126 6926 12178
rect 9314 12126 9326 12178
rect 9378 12126 9390 12178
rect 9874 12126 9886 12178
rect 9938 12126 9950 12178
rect 11218 12126 11230 12178
rect 11282 12126 11294 12178
rect 12114 12126 12126 12178
rect 12178 12126 12190 12178
rect 13122 12126 13134 12178
rect 13186 12126 13198 12178
rect 13570 12126 13582 12178
rect 13634 12126 13646 12178
rect 15026 12126 15038 12178
rect 15090 12126 15102 12178
rect 15922 12126 15934 12178
rect 15986 12126 15998 12178
rect 2830 12114 2882 12126
rect 8542 12114 8594 12126
rect 10670 12114 10722 12126
rect 8990 12066 9042 12078
rect 14254 12066 14306 12078
rect 7298 12014 7310 12066
rect 7362 12014 7374 12066
rect 9986 12014 9998 12066
rect 10050 12014 10062 12066
rect 8990 12002 9042 12014
rect 14254 12002 14306 12014
rect 13794 11902 13806 11954
rect 13858 11902 13870 11954
rect 672 11786 27888 11820
rect 672 11734 4466 11786
rect 4518 11734 4570 11786
rect 4622 11734 4674 11786
rect 4726 11734 24466 11786
rect 24518 11734 24570 11786
rect 24622 11734 24674 11786
rect 24726 11734 27888 11786
rect 672 11700 27888 11734
rect 10882 11566 10894 11618
rect 10946 11566 10958 11618
rect 2606 11506 2658 11518
rect 2258 11454 2270 11506
rect 2322 11454 2334 11506
rect 2606 11442 2658 11454
rect 3166 11506 3218 11518
rect 9886 11506 9938 11518
rect 4834 11454 4846 11506
rect 4898 11454 4910 11506
rect 6962 11454 6974 11506
rect 7026 11454 7038 11506
rect 14690 11454 14702 11506
rect 14754 11454 14766 11506
rect 15138 11454 15150 11506
rect 15202 11454 15214 11506
rect 3166 11442 3218 11454
rect 9886 11442 9938 11454
rect 8206 11394 8258 11406
rect 4274 11342 4286 11394
rect 4338 11342 4350 11394
rect 6626 11342 6638 11394
rect 6690 11342 6702 11394
rect 10210 11342 10222 11394
rect 10274 11342 10286 11394
rect 10770 11342 10782 11394
rect 10834 11342 10846 11394
rect 11442 11342 11454 11394
rect 11506 11342 11518 11394
rect 12002 11342 12014 11394
rect 12066 11342 12078 11394
rect 13010 11342 13022 11394
rect 13074 11342 13086 11394
rect 8206 11330 8258 11342
rect 1262 11170 1314 11182
rect 1262 11106 1314 11118
rect 5966 11170 6018 11182
rect 5966 11106 6018 11118
rect 14142 11170 14194 11182
rect 14142 11106 14194 11118
rect 14478 11170 14530 11182
rect 14478 11106 14530 11118
rect 672 11002 27888 11036
rect 672 10950 3806 11002
rect 3858 10950 3910 11002
rect 3962 10950 4014 11002
rect 4066 10950 23806 11002
rect 23858 10950 23910 11002
rect 23962 10950 24014 11002
rect 24066 10950 27888 11002
rect 672 10916 27888 10950
rect 12126 10834 12178 10846
rect 12126 10770 12178 10782
rect 5854 10722 5906 10734
rect 5854 10658 5906 10670
rect 6750 10722 6802 10734
rect 6750 10658 6802 10670
rect 14030 10722 14082 10734
rect 14030 10658 14082 10670
rect 14926 10722 14978 10734
rect 14926 10658 14978 10670
rect 14366 10610 14418 10622
rect 5394 10558 5406 10610
rect 5458 10558 5470 10610
rect 7074 10558 7086 10610
rect 7138 10558 7150 10610
rect 7522 10558 7534 10610
rect 7586 10558 7598 10610
rect 8306 10558 8318 10610
rect 8370 10558 8382 10610
rect 8978 10558 8990 10610
rect 9042 10558 9054 10610
rect 9874 10558 9886 10610
rect 9938 10558 9950 10610
rect 10434 10558 10446 10610
rect 10498 10558 10510 10610
rect 13570 10558 13582 10610
rect 13634 10558 13646 10610
rect 14366 10546 14418 10558
rect 10882 10446 10894 10498
rect 10946 10446 10958 10498
rect 7746 10334 7758 10386
rect 7810 10334 7822 10386
rect 672 10218 27888 10252
rect 672 10166 4466 10218
rect 4518 10166 4570 10218
rect 4622 10166 4674 10218
rect 4726 10166 24466 10218
rect 24518 10166 24570 10218
rect 24622 10166 24674 10218
rect 24726 10166 27888 10218
rect 672 10132 27888 10166
rect 7534 10050 7586 10062
rect 7534 9986 7586 9998
rect 4734 9938 4786 9950
rect 4734 9874 4786 9886
rect 10110 9938 10162 9950
rect 11106 9886 11118 9938
rect 11170 9886 11182 9938
rect 10110 9874 10162 9886
rect 11566 9826 11618 9838
rect 2146 9774 2158 9826
rect 2210 9774 2222 9826
rect 5170 9774 5182 9826
rect 5234 9774 5246 9826
rect 10434 9774 10446 9826
rect 10498 9774 10510 9826
rect 10882 9774 10894 9826
rect 10946 9774 10958 9826
rect 12114 9774 12126 9826
rect 12178 9774 12190 9826
rect 13122 9774 13134 9826
rect 13186 9774 13198 9826
rect 11566 9762 11618 9774
rect 6974 9714 7026 9726
rect 6974 9650 7026 9662
rect 1262 9602 1314 9614
rect 1262 9538 1314 9550
rect 672 9434 27888 9468
rect 672 9382 3806 9434
rect 3858 9382 3910 9434
rect 3962 9382 4014 9434
rect 4066 9382 23806 9434
rect 23858 9382 23910 9434
rect 23962 9382 24014 9434
rect 24066 9382 27888 9434
rect 672 9348 27888 9382
rect 8878 9266 8930 9278
rect 8878 9202 8930 9214
rect 11118 9266 11170 9278
rect 11118 9202 11170 9214
rect 7298 9102 7310 9154
rect 7362 9102 7374 9154
rect 9538 9102 9550 9154
rect 9602 9102 9614 9154
rect 7634 8878 7646 8930
rect 7698 8878 7710 8930
rect 9874 8878 9886 8930
rect 9938 8878 9950 8930
rect 672 8650 27888 8684
rect 672 8598 4466 8650
rect 4518 8598 4570 8650
rect 4622 8598 4674 8650
rect 4726 8598 24466 8650
rect 24518 8598 24570 8650
rect 24622 8598 24674 8650
rect 24726 8598 27888 8650
rect 672 8564 27888 8598
rect 7758 8482 7810 8494
rect 7758 8418 7810 8430
rect 11342 8482 11394 8494
rect 11342 8418 11394 8430
rect 10210 8318 10222 8370
rect 10274 8318 10286 8370
rect 9650 8206 9662 8258
rect 9714 8206 9726 8258
rect 8318 8146 8370 8158
rect 8318 8082 8370 8094
rect 672 7866 27888 7900
rect 672 7814 3806 7866
rect 3858 7814 3910 7866
rect 3962 7814 4014 7866
rect 4066 7814 23806 7866
rect 23858 7814 23910 7866
rect 23962 7814 24014 7866
rect 24066 7814 27888 7866
rect 672 7780 27888 7814
rect 11566 7586 11618 7598
rect 11566 7522 11618 7534
rect 11006 7474 11058 7486
rect 10210 7422 10222 7474
rect 10274 7422 10286 7474
rect 11006 7410 11058 7422
rect 10670 7362 10722 7374
rect 10670 7298 10722 7310
rect 672 7082 27888 7116
rect 672 7030 4466 7082
rect 4518 7030 4570 7082
rect 4622 7030 4674 7082
rect 4726 7030 24466 7082
rect 24518 7030 24570 7082
rect 24622 7030 24674 7082
rect 24726 7030 27888 7082
rect 672 6996 27888 7030
rect 2258 6750 2270 6802
rect 2322 6750 2334 6802
rect 1262 6578 1314 6590
rect 1262 6514 1314 6526
rect 672 6298 27888 6332
rect 672 6246 3806 6298
rect 3858 6246 3910 6298
rect 3962 6246 4014 6298
rect 4066 6246 23806 6298
rect 23858 6246 23910 6298
rect 23962 6246 24014 6298
rect 24066 6246 27888 6298
rect 672 6212 27888 6246
rect 1262 6018 1314 6030
rect 1262 5954 1314 5966
rect 2258 5854 2270 5906
rect 2322 5854 2334 5906
rect 672 5514 27888 5548
rect 672 5462 4466 5514
rect 4518 5462 4570 5514
rect 4622 5462 4674 5514
rect 4726 5462 24466 5514
rect 24518 5462 24570 5514
rect 24622 5462 24674 5514
rect 24726 5462 27888 5514
rect 672 5428 27888 5462
rect 672 4730 27888 4764
rect 672 4678 3806 4730
rect 3858 4678 3910 4730
rect 3962 4678 4014 4730
rect 4066 4678 23806 4730
rect 23858 4678 23910 4730
rect 23962 4678 24014 4730
rect 24066 4678 27888 4730
rect 672 4644 27888 4678
rect 672 3946 27888 3980
rect 672 3894 4466 3946
rect 4518 3894 4570 3946
rect 4622 3894 4674 3946
rect 4726 3894 24466 3946
rect 24518 3894 24570 3946
rect 24622 3894 24674 3946
rect 24726 3894 27888 3946
rect 672 3860 27888 3894
rect 672 3162 27888 3196
rect 672 3110 3806 3162
rect 3858 3110 3910 3162
rect 3962 3110 4014 3162
rect 4066 3110 23806 3162
rect 23858 3110 23910 3162
rect 23962 3110 24014 3162
rect 24066 3110 27888 3162
rect 672 3076 27888 3110
rect 672 2378 27888 2412
rect 672 2326 4466 2378
rect 4518 2326 4570 2378
rect 4622 2326 4674 2378
rect 4726 2326 24466 2378
rect 24518 2326 24570 2378
rect 24622 2326 24674 2378
rect 24726 2326 27888 2378
rect 672 2292 27888 2326
rect 672 1594 27888 1628
rect 672 1542 3806 1594
rect 3858 1542 3910 1594
rect 3962 1542 4014 1594
rect 4066 1542 23806 1594
rect 23858 1542 23910 1594
rect 23962 1542 24014 1594
rect 24066 1542 27888 1594
rect 672 1508 27888 1542
rect 672 810 27888 844
rect 672 758 4466 810
rect 4518 758 4570 810
rect 4622 758 4674 810
rect 4726 758 24466 810
rect 24518 758 24570 810
rect 24622 758 24674 810
rect 24726 758 27888 810
rect 672 724 27888 758
<< via1 >>
rect 3806 56422 3858 56474
rect 3910 56422 3962 56474
rect 4014 56422 4066 56474
rect 23806 56422 23858 56474
rect 23910 56422 23962 56474
rect 24014 56422 24066 56474
rect 3614 56254 3666 56306
rect 5518 56254 5570 56306
rect 8990 56254 9042 56306
rect 10558 56254 10610 56306
rect 13022 56254 13074 56306
rect 14590 56254 14642 56306
rect 16494 56254 16546 56306
rect 18510 56254 18562 56306
rect 20638 56254 20690 56306
rect 21870 56254 21922 56306
rect 24446 56254 24498 56306
rect 26014 56254 26066 56306
rect 7422 56142 7474 56194
rect 5182 56030 5234 56082
rect 20190 56030 20242 56082
rect 25678 56030 25730 56082
rect 1038 55918 1090 55970
rect 3054 55918 3106 55970
rect 8094 55918 8146 55970
rect 9998 55918 10050 55970
rect 11566 55918 11618 55970
rect 14030 55918 14082 55970
rect 15598 55918 15650 55970
rect 17502 55918 17554 55970
rect 19518 55918 19570 55970
rect 22878 55918 22930 55970
rect 23886 55918 23938 55970
rect 1374 55806 1426 55858
rect 4466 55638 4518 55690
rect 4570 55638 4622 55690
rect 4674 55638 4726 55690
rect 24466 55638 24518 55690
rect 24570 55638 24622 55690
rect 24674 55638 24726 55690
rect 18846 55358 18898 55410
rect 21646 55358 21698 55410
rect 3502 55246 3554 55298
rect 7534 55246 7586 55298
rect 12910 55246 12962 55298
rect 18286 55246 18338 55298
rect 19294 55246 19346 55298
rect 20078 55246 20130 55298
rect 20526 55246 20578 55298
rect 20862 55246 20914 55298
rect 23662 55246 23714 55298
rect 24670 55246 24722 55298
rect 26238 55246 26290 55298
rect 2494 55134 2546 55186
rect 6526 55134 6578 55186
rect 11902 55134 11954 55186
rect 17278 55134 17330 55186
rect 22654 55134 22706 55186
rect 25566 55134 25618 55186
rect 27246 55022 27298 55074
rect 3806 54854 3858 54906
rect 3910 54854 3962 54906
rect 4014 54854 4066 54906
rect 23806 54854 23858 54906
rect 23910 54854 23962 54906
rect 24014 54854 24066 54906
rect 22542 54686 22594 54738
rect 24110 54686 24162 54738
rect 19406 54574 19458 54626
rect 21086 54574 21138 54626
rect 25454 54574 25506 54626
rect 19070 54462 19122 54514
rect 24670 54462 24722 54514
rect 21534 54350 21586 54402
rect 23102 54350 23154 54402
rect 26238 54350 26290 54402
rect 27022 54350 27074 54402
rect 20638 54238 20690 54290
rect 4466 54070 4518 54122
rect 4570 54070 4622 54122
rect 4674 54070 4726 54122
rect 24466 54070 24518 54122
rect 24570 54070 24622 54122
rect 24674 54070 24726 54122
rect 20526 53678 20578 53730
rect 20862 53678 20914 53730
rect 21870 53678 21922 53730
rect 22318 53678 22370 53730
rect 22878 53678 22930 53730
rect 24894 53678 24946 53730
rect 26238 53678 26290 53730
rect 19966 53566 20018 53618
rect 21310 53566 21362 53618
rect 23774 53566 23826 53618
rect 25566 53566 25618 53618
rect 27246 53454 27298 53506
rect 3806 53286 3858 53338
rect 3910 53286 3962 53338
rect 4014 53286 4066 53338
rect 23806 53286 23858 53338
rect 23910 53286 23962 53338
rect 24014 53286 24066 53338
rect 24110 53118 24162 53170
rect 21758 53006 21810 53058
rect 22654 53006 22706 53058
rect 27134 53006 27186 53058
rect 21422 52894 21474 52946
rect 23214 52894 23266 52946
rect 24670 52894 24722 52946
rect 25454 52782 25506 52834
rect 26238 52782 26290 52834
rect 22206 52670 22258 52722
rect 4466 52502 4518 52554
rect 4570 52502 4622 52554
rect 4674 52502 4726 52554
rect 24466 52502 24518 52554
rect 24570 52502 24622 52554
rect 24674 52502 24726 52554
rect 21870 52222 21922 52274
rect 22766 52222 22818 52274
rect 23550 52222 23602 52274
rect 24670 52222 24722 52274
rect 22430 52110 22482 52162
rect 26238 52110 26290 52162
rect 25566 51998 25618 52050
rect 27246 51886 27298 51938
rect 3806 51718 3858 51770
rect 3910 51718 3962 51770
rect 4014 51718 4066 51770
rect 23806 51718 23858 51770
rect 23910 51718 23962 51770
rect 24014 51718 24066 51770
rect 23326 51438 23378 51490
rect 24334 51438 24386 51490
rect 25342 51438 25394 51490
rect 24670 51214 24722 51266
rect 26238 51214 26290 51266
rect 27022 51214 27074 51266
rect 22766 51102 22818 51154
rect 23774 51102 23826 51154
rect 4466 50934 4518 50986
rect 4570 50934 4622 50986
rect 4674 50934 4726 50986
rect 24466 50934 24518 50986
rect 24570 50934 24622 50986
rect 24674 50934 24726 50986
rect 23438 50654 23490 50706
rect 23886 50542 23938 50594
rect 24894 50542 24946 50594
rect 26350 50542 26402 50594
rect 25566 50430 25618 50482
rect 27246 50318 27298 50370
rect 3806 50150 3858 50202
rect 3910 50150 3962 50202
rect 4014 50150 4066 50202
rect 23806 50150 23858 50202
rect 23910 50150 23962 50202
rect 24014 50150 24066 50202
rect 24222 49870 24274 49922
rect 25678 49870 25730 49922
rect 27134 49870 27186 49922
rect 26350 49758 26402 49810
rect 24670 49646 24722 49698
rect 23774 49534 23826 49586
rect 4466 49366 4518 49418
rect 4570 49366 4622 49418
rect 4674 49366 4726 49418
rect 24466 49366 24518 49418
rect 24570 49366 24622 49418
rect 24674 49366 24726 49418
rect 24670 48974 24722 49026
rect 26238 48974 26290 49026
rect 25678 48750 25730 48802
rect 27246 48750 27298 48802
rect 3806 48582 3858 48634
rect 3910 48582 3962 48634
rect 4014 48582 4066 48634
rect 23806 48582 23858 48634
rect 23910 48582 23962 48634
rect 24014 48582 24066 48634
rect 25006 48302 25058 48354
rect 25790 48302 25842 48354
rect 26238 48078 26290 48130
rect 27022 48078 27074 48130
rect 24446 47966 24498 48018
rect 25342 47966 25394 48018
rect 4466 47798 4518 47850
rect 4570 47798 4622 47850
rect 4674 47798 4726 47850
rect 24466 47798 24518 47850
rect 24570 47798 24622 47850
rect 24674 47798 24726 47850
rect 24670 47406 24722 47458
rect 26462 47406 26514 47458
rect 25678 47294 25730 47346
rect 27246 47182 27298 47234
rect 3806 47014 3858 47066
rect 3910 47014 3962 47066
rect 4014 47014 4066 47066
rect 23806 47014 23858 47066
rect 23910 47014 23962 47066
rect 24014 47014 24066 47066
rect 25678 46734 25730 46786
rect 27134 46734 27186 46786
rect 24894 46622 24946 46674
rect 26350 46622 26402 46674
rect 4466 46230 4518 46282
rect 4570 46230 4622 46282
rect 4674 46230 4726 46282
rect 24466 46230 24518 46282
rect 24570 46230 24622 46282
rect 24674 46230 24726 46282
rect 24670 45838 24722 45890
rect 26238 45838 26290 45890
rect 25678 45614 25730 45666
rect 27246 45614 27298 45666
rect 3806 45446 3858 45498
rect 3910 45446 3962 45498
rect 4014 45446 4066 45498
rect 23806 45446 23858 45498
rect 23910 45446 23962 45498
rect 24014 45446 24066 45498
rect 26238 44942 26290 44994
rect 27022 44942 27074 44994
rect 4466 44662 4518 44714
rect 4570 44662 4622 44714
rect 4674 44662 4726 44714
rect 24466 44662 24518 44714
rect 24570 44662 24622 44714
rect 24674 44662 24726 44714
rect 24670 44270 24722 44322
rect 26238 44270 26290 44322
rect 25678 44158 25730 44210
rect 27246 44046 27298 44098
rect 3806 43878 3858 43930
rect 3910 43878 3962 43930
rect 4014 43878 4066 43930
rect 23806 43878 23858 43930
rect 23910 43878 23962 43930
rect 24014 43878 24066 43930
rect 25678 43598 25730 43650
rect 24894 43486 24946 43538
rect 26238 43374 26290 43426
rect 26798 43262 26850 43314
rect 4466 43094 4518 43146
rect 4570 43094 4622 43146
rect 4674 43094 4726 43146
rect 24466 43094 24518 43146
rect 24570 43094 24622 43146
rect 24674 43094 24726 43146
rect 24670 42702 24722 42754
rect 26238 42702 26290 42754
rect 25678 42478 25730 42530
rect 27246 42478 27298 42530
rect 3806 42310 3858 42362
rect 3910 42310 3962 42362
rect 4014 42310 4066 42362
rect 23806 42310 23858 42362
rect 23910 42310 23962 42362
rect 24014 42310 24066 42362
rect 4174 41918 4226 41970
rect 16270 41918 16322 41970
rect 18398 41806 18450 41858
rect 26238 41806 26290 41858
rect 3614 41694 3666 41746
rect 26798 41694 26850 41746
rect 4466 41526 4518 41578
rect 4570 41526 4622 41578
rect 4674 41526 4726 41578
rect 24466 41526 24518 41578
rect 24570 41526 24622 41578
rect 24674 41526 24726 41578
rect 6078 41358 6130 41410
rect 4286 41246 4338 41298
rect 6638 41246 6690 41298
rect 10558 41246 10610 41298
rect 3838 41134 3890 41186
rect 8878 41134 8930 41186
rect 24782 41134 24834 41186
rect 26238 41134 26290 41186
rect 9438 41022 9490 41074
rect 10222 41022 10274 41074
rect 25678 41022 25730 41074
rect 5518 40910 5570 40962
rect 11790 40910 11842 40962
rect 27246 40910 27298 40962
rect 3806 40742 3858 40794
rect 3910 40742 3962 40794
rect 4014 40742 4066 40794
rect 23806 40742 23858 40794
rect 23910 40742 23962 40794
rect 24014 40742 24066 40794
rect 2158 40462 2210 40514
rect 13358 40462 13410 40514
rect 15486 40462 15538 40514
rect 25678 40462 25730 40514
rect 1710 40350 1762 40402
rect 2606 40350 2658 40402
rect 4286 40350 4338 40402
rect 7646 40350 7698 40402
rect 8094 40350 8146 40402
rect 8766 40350 8818 40402
rect 9326 40350 9378 40402
rect 10446 40350 10498 40402
rect 17726 40350 17778 40402
rect 18398 40350 18450 40402
rect 24670 40350 24722 40402
rect 26238 40350 26290 40402
rect 3054 40238 3106 40290
rect 6974 40238 7026 40290
rect 7310 40238 7362 40290
rect 8318 40238 8370 40290
rect 6414 40126 6466 40178
rect 12910 40126 12962 40178
rect 26798 40126 26850 40178
rect 4466 39958 4518 40010
rect 4570 39958 4622 40010
rect 4674 39958 4726 40010
rect 24466 39958 24518 40010
rect 24570 39958 24622 40010
rect 24674 39958 24726 40010
rect 6078 39790 6130 39842
rect 9886 39790 9938 39842
rect 12462 39790 12514 39842
rect 2270 39678 2322 39730
rect 3166 39678 3218 39730
rect 5070 39678 5122 39730
rect 12910 39678 12962 39730
rect 24670 39678 24722 39730
rect 1710 39566 1762 39618
rect 2606 39566 2658 39618
rect 5518 39566 5570 39618
rect 5854 39566 5906 39618
rect 6750 39566 6802 39618
rect 7086 39566 7138 39618
rect 7310 39566 7362 39618
rect 8206 39566 8258 39618
rect 9438 39566 9490 39618
rect 11790 39566 11842 39618
rect 12350 39566 12402 39618
rect 13582 39566 13634 39618
rect 14590 39566 14642 39618
rect 16718 39566 16770 39618
rect 26238 39566 26290 39618
rect 11006 39454 11058 39506
rect 11454 39454 11506 39506
rect 18734 39454 18786 39506
rect 25678 39342 25730 39394
rect 27246 39342 27298 39394
rect 3806 39174 3858 39226
rect 3910 39174 3962 39226
rect 4014 39174 4066 39226
rect 23806 39174 23858 39226
rect 23910 39174 23962 39226
rect 24014 39174 24066 39226
rect 7198 39006 7250 39058
rect 2046 38894 2098 38946
rect 2718 38894 2770 38946
rect 5630 38894 5682 38946
rect 13358 38894 13410 38946
rect 26910 38894 26962 38946
rect 4286 38782 4338 38834
rect 10558 38782 10610 38834
rect 15822 38782 15874 38834
rect 26238 38782 26290 38834
rect 3054 38670 3106 38722
rect 5966 38670 6018 38722
rect 11006 38670 11058 38722
rect 18622 38670 18674 38722
rect 1598 38558 1650 38610
rect 12126 38558 12178 38610
rect 12910 38558 12962 38610
rect 4466 38390 4518 38442
rect 4570 38390 4622 38442
rect 4674 38390 4726 38442
rect 24466 38390 24518 38442
rect 24570 38390 24622 38442
rect 24674 38390 24726 38442
rect 6302 38222 6354 38274
rect 12574 38222 12626 38274
rect 15150 38222 15202 38274
rect 2382 38110 2434 38162
rect 5070 38110 5122 38162
rect 7310 38110 7362 38162
rect 7758 38110 7810 38162
rect 9998 38110 10050 38162
rect 4622 37998 4674 38050
rect 6750 37998 6802 38050
rect 8318 37998 8370 38050
rect 9550 37998 9602 38050
rect 11118 37998 11170 38050
rect 11902 37998 11954 38050
rect 12462 38004 12514 38056
rect 13134 37998 13186 38050
rect 13582 37998 13634 38050
rect 14702 37998 14754 38050
rect 15486 37998 15538 38050
rect 16718 37998 16770 38050
rect 24894 37998 24946 38050
rect 26238 37998 26290 38050
rect 2718 37886 2770 37938
rect 11566 37886 11618 37938
rect 17502 37886 17554 37938
rect 19742 37886 19794 37938
rect 25678 37886 25730 37938
rect 1150 37774 1202 37826
rect 27246 37774 27298 37826
rect 3806 37606 3858 37658
rect 3910 37606 3962 37658
rect 4014 37606 4066 37658
rect 23806 37606 23858 37658
rect 23910 37606 23962 37658
rect 24014 37606 24066 37658
rect 6750 37438 6802 37490
rect 1486 37326 1538 37378
rect 2494 37326 2546 37378
rect 16494 37326 16546 37378
rect 2046 37214 2098 37266
rect 5182 37214 5234 37266
rect 7870 37214 7922 37266
rect 8318 37214 8370 37266
rect 8990 37214 9042 37266
rect 9550 37214 9602 37266
rect 10670 37214 10722 37266
rect 18622 37214 18674 37266
rect 26238 37214 26290 37266
rect 7534 37102 7586 37154
rect 8542 37102 8594 37154
rect 16606 37102 16658 37154
rect 24670 37102 24722 37154
rect 25454 37102 25506 37154
rect 1038 36990 1090 37042
rect 1934 36990 1986 37042
rect 5630 36990 5682 37042
rect 26798 36990 26850 37042
rect 4466 36822 4518 36874
rect 4570 36822 4622 36874
rect 4674 36822 4726 36874
rect 24466 36822 24518 36874
rect 24570 36822 24622 36874
rect 24674 36822 24726 36874
rect 10110 36654 10162 36706
rect 1598 36542 1650 36594
rect 3950 36542 4002 36594
rect 12126 36542 12178 36594
rect 15710 36542 15762 36594
rect 18846 36542 18898 36594
rect 1262 36430 1314 36482
rect 3390 36430 3442 36482
rect 6190 36430 6242 36482
rect 8318 36430 8370 36482
rect 14366 36430 14418 36482
rect 14814 36430 14866 36482
rect 15934 36430 15986 36482
rect 17838 36430 17890 36482
rect 18286 36430 18338 36482
rect 24894 36430 24946 36482
rect 26350 36430 26402 36482
rect 6750 36318 6802 36370
rect 7870 36318 7922 36370
rect 10558 36318 10610 36370
rect 11790 36318 11842 36370
rect 13918 36318 13970 36370
rect 2830 36206 2882 36258
rect 5070 36206 5122 36258
rect 8990 36206 9042 36258
rect 13358 36206 13410 36258
rect 15150 36206 15202 36258
rect 17390 36206 17442 36258
rect 25678 36206 25730 36258
rect 27246 36206 27298 36258
rect 3806 36038 3858 36090
rect 3910 36038 3962 36090
rect 4014 36038 4066 36090
rect 23806 36038 23858 36090
rect 23910 36038 23962 36090
rect 24014 36038 24066 36090
rect 5854 35758 5906 35810
rect 7422 35758 7474 35810
rect 11454 35758 11506 35810
rect 12910 35758 12962 35810
rect 15486 35758 15538 35810
rect 26910 35758 26962 35810
rect 2606 35646 2658 35698
rect 8318 35646 8370 35698
rect 8654 35646 8706 35698
rect 9326 35646 9378 35698
rect 9998 35646 10050 35698
rect 10894 35646 10946 35698
rect 11902 35646 11954 35698
rect 18398 35646 18450 35698
rect 7870 35534 7922 35586
rect 26238 35534 26290 35586
rect 3166 35422 3218 35474
rect 4286 35422 4338 35474
rect 6302 35422 6354 35474
rect 8878 35422 8930 35474
rect 13358 35422 13410 35474
rect 4466 35254 4518 35306
rect 4570 35254 4622 35306
rect 4674 35254 4726 35306
rect 24466 35254 24518 35306
rect 24570 35254 24622 35306
rect 24674 35254 24726 35306
rect 6078 35086 6130 35138
rect 11006 35086 11058 35138
rect 13582 35086 13634 35138
rect 16830 35086 16882 35138
rect 3054 34974 3106 35026
rect 14030 34974 14082 35026
rect 17950 34974 18002 35026
rect 19854 34974 19906 35026
rect 20414 34974 20466 35026
rect 2158 34862 2210 34914
rect 2606 34862 2658 34914
rect 4286 34862 4338 34914
rect 5406 34862 5458 34914
rect 5966 34862 6018 34914
rect 6750 34862 6802 34914
rect 7198 34862 7250 34914
rect 8094 34862 8146 34914
rect 12126 34862 12178 34914
rect 12910 34862 12962 34914
rect 13358 34862 13410 34914
rect 14590 34862 14642 34914
rect 15710 34862 15762 34914
rect 18958 34862 19010 34914
rect 24670 34862 24722 34914
rect 26238 34862 26290 34914
rect 1710 34750 1762 34802
rect 5070 34750 5122 34802
rect 10558 34750 10610 34802
rect 12574 34750 12626 34802
rect 18398 34750 18450 34802
rect 19406 34750 19458 34802
rect 25678 34750 25730 34802
rect 27246 34638 27298 34690
rect 3806 34470 3858 34522
rect 3910 34470 3962 34522
rect 4014 34470 4066 34522
rect 23806 34470 23858 34522
rect 23910 34470 23962 34522
rect 24014 34470 24066 34522
rect 6750 34302 6802 34354
rect 16718 34190 16770 34242
rect 25678 34190 25730 34242
rect 1486 34078 1538 34130
rect 1934 34078 1986 34130
rect 2830 34078 2882 34130
rect 3278 34078 3330 34130
rect 4286 34078 4338 34130
rect 5182 34078 5234 34130
rect 9214 34078 9266 34130
rect 18510 34078 18562 34130
rect 1150 33966 1202 34018
rect 2158 33966 2210 34018
rect 24670 33966 24722 34018
rect 26238 33966 26290 34018
rect 5630 33854 5682 33906
rect 7534 33854 7586 33906
rect 8654 33854 8706 33906
rect 26798 33854 26850 33906
rect 4466 33686 4518 33738
rect 4570 33686 4622 33738
rect 4674 33686 4726 33738
rect 24466 33686 24518 33738
rect 24570 33686 24622 33738
rect 24674 33686 24726 33738
rect 6078 33518 6130 33570
rect 9998 33518 10050 33570
rect 18398 33518 18450 33570
rect 1598 33406 1650 33458
rect 8206 33406 8258 33458
rect 12350 33406 12402 33458
rect 14590 33406 14642 33458
rect 7646 33294 7698 33346
rect 9550 33294 9602 33346
rect 11790 33294 11842 33346
rect 17390 33294 17442 33346
rect 17838 33294 17890 33346
rect 24670 33294 24722 33346
rect 26350 33294 26402 33346
rect 1262 33182 1314 33234
rect 5630 33182 5682 33234
rect 15038 33182 15090 33234
rect 16942 33182 16994 33234
rect 17950 33182 18002 33234
rect 2830 33070 2882 33122
rect 7198 33070 7250 33122
rect 11118 33070 11170 33122
rect 13470 33070 13522 33122
rect 19518 33070 19570 33122
rect 25678 33070 25730 33122
rect 27246 33070 27298 33122
rect 3806 32902 3858 32954
rect 3910 32902 3962 32954
rect 4014 32902 4066 32954
rect 23806 32902 23858 32954
rect 23910 32902 23962 32954
rect 24014 32902 24066 32954
rect 18286 32734 18338 32786
rect 13358 32622 13410 32674
rect 14366 32622 14418 32674
rect 17278 32622 17330 32674
rect 18622 32622 18674 32674
rect 26910 32622 26962 32674
rect 1598 32510 1650 32562
rect 6750 32510 6802 32562
rect 7086 32510 7138 32562
rect 7758 32510 7810 32562
rect 8430 32510 8482 32562
rect 9326 32510 9378 32562
rect 10446 32510 10498 32562
rect 13022 32510 13074 32562
rect 15150 32510 15202 32562
rect 19070 32510 19122 32562
rect 26238 32510 26290 32562
rect 2158 32398 2210 32450
rect 4286 32398 4338 32450
rect 6302 32398 6354 32450
rect 7310 32398 7362 32450
rect 15598 32398 15650 32450
rect 19182 32398 19234 32450
rect 3278 32286 3330 32338
rect 3726 32286 3778 32338
rect 11006 32286 11058 32338
rect 12126 32286 12178 32338
rect 13806 32286 13858 32338
rect 16830 32286 16882 32338
rect 17838 32286 17890 32338
rect 4466 32118 4518 32170
rect 4570 32118 4622 32170
rect 4674 32118 4726 32170
rect 24466 32118 24518 32170
rect 24570 32118 24622 32170
rect 24674 32118 24726 32170
rect 13022 31950 13074 32002
rect 17726 31950 17778 32002
rect 2830 31838 2882 31890
rect 3278 31838 3330 31890
rect 18174 31838 18226 31890
rect 2270 31726 2322 31778
rect 2718 31726 2770 31778
rect 4062 31726 4114 31778
rect 4846 31726 4898 31778
rect 7310 31726 7362 31778
rect 8878 31726 8930 31778
rect 12350 31726 12402 31778
rect 12798 31726 12850 31778
rect 13582 31726 13634 31778
rect 14254 31726 14306 31778
rect 15038 31726 15090 31778
rect 17054 31726 17106 31778
rect 17502 31726 17554 31778
rect 18958 31726 19010 31778
rect 19854 31726 19906 31778
rect 24670 31726 24722 31778
rect 26350 31726 26402 31778
rect 1822 31614 1874 31666
rect 7982 31614 8034 31666
rect 9326 31614 9378 31666
rect 12014 31614 12066 31666
rect 16718 31614 16770 31666
rect 25678 31614 25730 31666
rect 26910 31614 26962 31666
rect 3806 31334 3858 31386
rect 3910 31334 3962 31386
rect 4014 31334 4066 31386
rect 23806 31334 23858 31386
rect 23910 31334 23962 31386
rect 24014 31334 24066 31386
rect 15822 31166 15874 31218
rect 4398 31054 4450 31106
rect 6638 31054 6690 31106
rect 7198 31054 7250 31106
rect 11902 31054 11954 31106
rect 27246 31054 27298 31106
rect 1262 30942 1314 30994
rect 2382 30942 2434 30994
rect 3502 30942 3554 30994
rect 3950 30942 4002 30994
rect 8094 30942 8146 30994
rect 10446 30942 10498 30994
rect 11342 30942 11394 30994
rect 14254 30942 14306 30994
rect 17166 30942 17218 30994
rect 17502 30942 17554 30994
rect 18398 30942 18450 30994
rect 18734 30942 18786 30994
rect 19854 30942 19906 30994
rect 24894 30942 24946 30994
rect 2942 30830 2994 30882
rect 8654 30830 8706 30882
rect 10894 30830 10946 30882
rect 16718 30830 16770 30882
rect 17726 30830 17778 30882
rect 25454 30830 25506 30882
rect 26238 30830 26290 30882
rect 3390 30718 3442 30770
rect 6190 30718 6242 30770
rect 7646 30718 7698 30770
rect 9774 30718 9826 30770
rect 14702 30718 14754 30770
rect 4466 30550 4518 30602
rect 4570 30550 4622 30602
rect 4674 30550 4726 30602
rect 24466 30550 24518 30602
rect 24570 30550 24622 30602
rect 24674 30550 24726 30602
rect 3166 30382 3218 30434
rect 6078 30382 6130 30434
rect 10446 30382 10498 30434
rect 16158 30270 16210 30322
rect 17278 30270 17330 30322
rect 1038 30158 1090 30210
rect 5406 30158 5458 30210
rect 5854 30158 5906 30210
rect 6750 30158 6802 30210
rect 7086 30158 7138 30210
rect 8206 30158 8258 30210
rect 9438 30158 9490 30210
rect 9774 30158 9826 30210
rect 10222 30158 10274 30210
rect 11118 30158 11170 30210
rect 11454 30158 11506 30210
rect 12574 30158 12626 30210
rect 14142 30158 14194 30210
rect 15710 30158 15762 30210
rect 16830 30158 16882 30210
rect 26238 30158 26290 30210
rect 2718 30046 2770 30098
rect 5070 30046 5122 30098
rect 14702 30046 14754 30098
rect 18510 30046 18562 30098
rect 26910 30046 26962 30098
rect 2046 29934 2098 29986
rect 3806 29766 3858 29818
rect 3910 29766 3962 29818
rect 4014 29766 4066 29818
rect 23806 29766 23858 29818
rect 23910 29766 23962 29818
rect 24014 29766 24066 29818
rect 2830 29598 2882 29650
rect 6750 29598 6802 29650
rect 17502 29598 17554 29650
rect 1262 29486 1314 29538
rect 5182 29486 5234 29538
rect 12126 29486 12178 29538
rect 15934 29486 15986 29538
rect 27246 29486 27298 29538
rect 8542 29374 8594 29426
rect 11790 29374 11842 29426
rect 13582 29374 13634 29426
rect 18174 29374 18226 29426
rect 19742 29374 19794 29426
rect 1598 29262 1650 29314
rect 5518 29262 5570 29314
rect 14142 29262 14194 29314
rect 18622 29262 18674 29314
rect 26238 29262 26290 29314
rect 8990 29150 9042 29202
rect 10110 29150 10162 29202
rect 15262 29150 15314 29202
rect 16382 29150 16434 29202
rect 4466 28982 4518 29034
rect 4570 28982 4622 29034
rect 4674 28982 4726 29034
rect 24466 28982 24518 29034
rect 24570 28982 24622 29034
rect 24674 28982 24726 29034
rect 2830 28814 2882 28866
rect 5070 28814 5122 28866
rect 11342 28814 11394 28866
rect 13918 28814 13970 28866
rect 1598 28702 1650 28754
rect 3838 28702 3890 28754
rect 5518 28702 5570 28754
rect 6974 28702 7026 28754
rect 12910 28702 12962 28754
rect 18398 28702 18450 28754
rect 19406 28702 19458 28754
rect 26238 28702 26290 28754
rect 1262 28590 1314 28642
rect 5966 28590 6018 28642
rect 12462 28590 12514 28642
rect 13246 28590 13298 28642
rect 13694 28590 13746 28642
rect 14366 28590 14418 28642
rect 14926 28590 14978 28642
rect 15934 28590 15986 28642
rect 18846 28590 18898 28642
rect 19182 28590 19234 28642
rect 20078 28590 20130 28642
rect 20414 28590 20466 28642
rect 20638 28590 20690 28642
rect 21422 28590 21474 28642
rect 3502 28478 3554 28530
rect 6638 28478 6690 28530
rect 10894 28478 10946 28530
rect 27246 28478 27298 28530
rect 8206 28366 8258 28418
rect 3806 28198 3858 28250
rect 3910 28198 3962 28250
rect 4014 28198 4066 28250
rect 23806 28198 23858 28250
rect 23910 28198 23962 28250
rect 24014 28198 24066 28250
rect 19070 28030 19122 28082
rect 27246 28030 27298 28082
rect 1486 27918 1538 27970
rect 4958 27918 5010 27970
rect 8990 27918 9042 27970
rect 13582 27918 13634 27970
rect 17502 27918 17554 27970
rect 20078 27918 20130 27970
rect 25678 27918 25730 27970
rect 1038 27806 1090 27858
rect 2606 27806 2658 27858
rect 4286 27806 4338 27858
rect 5294 27806 5346 27858
rect 5742 27806 5794 27858
rect 6526 27806 6578 27858
rect 7198 27806 7250 27858
rect 8094 27806 8146 27858
rect 9326 27806 9378 27858
rect 9774 27806 9826 27858
rect 10446 27806 10498 27858
rect 11230 27806 11282 27858
rect 12014 27806 12066 27858
rect 14030 27806 14082 27858
rect 14478 27806 14530 27858
rect 15262 27806 15314 27858
rect 15598 27806 15650 27858
rect 16606 27806 16658 27858
rect 26350 27806 26402 27858
rect 3054 27694 3106 27746
rect 5966 27694 6018 27746
rect 17838 27694 17890 27746
rect 19518 27694 19570 27746
rect 24670 27694 24722 27746
rect 9998 27582 10050 27634
rect 14590 27582 14642 27634
rect 4466 27414 4518 27466
rect 4570 27414 4622 27466
rect 4674 27414 4726 27466
rect 24466 27414 24518 27466
rect 24570 27414 24622 27466
rect 24674 27414 24726 27466
rect 5406 27246 5458 27298
rect 6526 27246 6578 27298
rect 10222 27246 10274 27298
rect 12910 27246 12962 27298
rect 15150 27246 15202 27298
rect 15598 27246 15650 27298
rect 1598 27134 1650 27186
rect 10782 27134 10834 27186
rect 11678 27134 11730 27186
rect 13918 27134 13970 27186
rect 16158 27134 16210 27186
rect 18174 27134 18226 27186
rect 24670 27134 24722 27186
rect 1262 27022 1314 27074
rect 4846 27022 4898 27074
rect 11342 27022 11394 27074
rect 13470 27022 13522 27074
rect 17726 27022 17778 27074
rect 26238 27022 26290 27074
rect 27246 26910 27298 26962
rect 2830 26798 2882 26850
rect 19406 26798 19458 26850
rect 25678 26798 25730 26850
rect 3806 26630 3858 26682
rect 3910 26630 3962 26682
rect 4014 26630 4066 26682
rect 23806 26630 23858 26682
rect 23910 26630 23962 26682
rect 24014 26630 24066 26682
rect 27246 26462 27298 26514
rect 1710 26350 1762 26402
rect 4174 26350 4226 26402
rect 7646 26350 7698 26402
rect 13358 26350 13410 26402
rect 14590 26350 14642 26402
rect 16494 26350 16546 26402
rect 19630 26350 19682 26402
rect 12910 26238 12962 26290
rect 2046 26126 2098 26178
rect 26238 26126 26290 26178
rect 3278 26014 3330 26066
rect 3726 26014 3778 26066
rect 8094 26014 8146 26066
rect 9214 26014 9266 26066
rect 14030 26014 14082 26066
rect 16942 26014 16994 26066
rect 18062 26014 18114 26066
rect 19182 26014 19234 26066
rect 4466 25846 4518 25898
rect 4570 25846 4622 25898
rect 4674 25846 4726 25898
rect 24466 25846 24518 25898
rect 24570 25846 24622 25898
rect 24674 25846 24726 25898
rect 3054 25678 3106 25730
rect 3502 25566 3554 25618
rect 6638 25566 6690 25618
rect 9438 25566 9490 25618
rect 10894 25566 10946 25618
rect 13134 25566 13186 25618
rect 15262 25566 15314 25618
rect 17502 25566 17554 25618
rect 18510 25566 18562 25618
rect 24670 25566 24722 25618
rect 2494 25454 2546 25506
rect 2830 25454 2882 25506
rect 4286 25454 4338 25506
rect 5070 25454 5122 25506
rect 6302 25454 6354 25506
rect 8878 25454 8930 25506
rect 14702 25454 14754 25506
rect 17950 25454 18002 25506
rect 18398 25454 18450 25506
rect 19182 25454 19234 25506
rect 19742 25454 19794 25506
rect 20526 25454 20578 25506
rect 26238 25454 26290 25506
rect 2046 25342 2098 25394
rect 10446 25342 10498 25394
rect 12686 25342 12738 25394
rect 27246 25342 27298 25394
rect 7870 25230 7922 25282
rect 12014 25230 12066 25282
rect 14254 25230 14306 25282
rect 25678 25230 25730 25282
rect 3806 25062 3858 25114
rect 3910 25062 3962 25114
rect 4014 25062 4066 25114
rect 23806 25062 23858 25114
rect 23910 25062 23962 25114
rect 24014 25062 24066 25114
rect 27246 24894 27298 24946
rect 6190 24782 6242 24834
rect 7534 24782 7586 24834
rect 18174 24782 18226 24834
rect 19518 24782 19570 24834
rect 1262 24670 1314 24722
rect 2270 24670 2322 24722
rect 2718 24670 2770 24722
rect 3502 24670 3554 24722
rect 4062 24670 4114 24722
rect 7870 24670 7922 24722
rect 8318 24670 8370 24722
rect 9214 24670 9266 24722
rect 9774 24670 9826 24722
rect 10670 24670 10722 24722
rect 13358 24670 13410 24722
rect 13806 24670 13858 24722
rect 14366 24670 14418 24722
rect 14926 24670 14978 24722
rect 15934 24670 15986 24722
rect 18958 24670 19010 24722
rect 24894 24670 24946 24722
rect 26238 24670 26290 24722
rect 4398 24558 4450 24610
rect 8542 24558 8594 24610
rect 12238 24558 12290 24610
rect 12910 24558 12962 24610
rect 13918 24558 13970 24610
rect 25454 24558 25506 24610
rect 3390 24446 3442 24498
rect 5630 24446 5682 24498
rect 12014 24446 12066 24498
rect 12126 24446 12178 24498
rect 16606 24446 16658 24498
rect 17726 24446 17778 24498
rect 4466 24278 4518 24330
rect 4570 24278 4622 24330
rect 4674 24278 4726 24330
rect 24466 24278 24518 24330
rect 24570 24278 24622 24330
rect 24674 24278 24726 24330
rect 1486 24110 1538 24162
rect 2494 24110 2546 24162
rect 5630 24110 5682 24162
rect 13806 24110 13858 24162
rect 3614 23998 3666 24050
rect 6078 23998 6130 24050
rect 9326 23998 9378 24050
rect 11230 23998 11282 24050
rect 17950 23998 18002 24050
rect 24670 23998 24722 24050
rect 2046 23886 2098 23938
rect 5070 23886 5122 23938
rect 5406 23886 5458 23938
rect 6638 23886 6690 23938
rect 7758 23886 7810 23938
rect 9886 23886 9938 23938
rect 12350 23886 12402 23938
rect 13134 23886 13186 23938
rect 13694 23886 13746 23938
rect 14254 23886 14306 23938
rect 14926 23886 14978 23938
rect 15934 23886 15986 23938
rect 18398 23886 18450 23938
rect 19406 23886 19458 23938
rect 26238 23886 26290 23938
rect 4062 23774 4114 23826
rect 4622 23774 4674 23826
rect 10782 23774 10834 23826
rect 12798 23774 12850 23826
rect 19854 23774 19906 23826
rect 27246 23774 27298 23826
rect 16830 23662 16882 23714
rect 25678 23662 25730 23714
rect 3806 23494 3858 23546
rect 3910 23494 3962 23546
rect 4014 23494 4066 23546
rect 23806 23494 23858 23546
rect 23910 23494 23962 23546
rect 24014 23494 24066 23546
rect 3838 23326 3890 23378
rect 11678 23326 11730 23378
rect 27246 23326 27298 23378
rect 1150 23214 1202 23266
rect 6190 23214 6242 23266
rect 6750 23214 6802 23266
rect 16942 23214 16994 23266
rect 18958 23214 19010 23266
rect 1598 23102 1650 23154
rect 2158 23102 2210 23154
rect 8990 23102 9042 23154
rect 11454 23102 11506 23154
rect 13134 23102 13186 23154
rect 13694 23102 13746 23154
rect 14366 23102 14418 23154
rect 14814 23102 14866 23154
rect 15934 23102 15986 23154
rect 26350 23102 26402 23154
rect 2718 22990 2770 23042
rect 5630 22990 5682 23042
rect 9438 22990 9490 23042
rect 10558 22990 10610 23042
rect 12014 22990 12066 23042
rect 12238 22990 12290 23042
rect 12798 22990 12850 23042
rect 13806 22990 13858 23042
rect 18510 22990 18562 23042
rect 7198 22878 7250 22930
rect 8318 22878 8370 22930
rect 11790 22878 11842 22930
rect 16382 22878 16434 22930
rect 17390 22878 17442 22930
rect 4466 22710 4518 22762
rect 4570 22710 4622 22762
rect 4674 22710 4726 22762
rect 24466 22710 24518 22762
rect 24570 22710 24622 22762
rect 24674 22710 24726 22762
rect 1150 22542 1202 22594
rect 2718 22542 2770 22594
rect 5966 22542 6018 22594
rect 9886 22542 9938 22594
rect 15150 22542 15202 22594
rect 10334 22430 10386 22482
rect 14702 22430 14754 22482
rect 18622 22430 18674 22482
rect 26238 22430 26290 22482
rect 2270 22318 2322 22370
rect 5294 22318 5346 22370
rect 5854 22318 5906 22370
rect 6414 22318 6466 22370
rect 6974 22318 7026 22370
rect 8094 22318 8146 22370
rect 9214 22318 9266 22370
rect 9662 22318 9714 22370
rect 11118 22318 11170 22370
rect 11902 22318 11954 22370
rect 13022 22318 13074 22370
rect 13918 22318 13970 22370
rect 15262 22318 15314 22370
rect 15822 22318 15874 22370
rect 16830 22318 16882 22370
rect 24894 22318 24946 22370
rect 1598 22206 1650 22258
rect 4958 22206 5010 22258
rect 8878 22206 8930 22258
rect 16158 22206 16210 22258
rect 18958 22206 19010 22258
rect 27246 22206 27298 22258
rect 3838 22094 3890 22146
rect 16718 22094 16770 22146
rect 17390 22094 17442 22146
rect 25678 22094 25730 22146
rect 3806 21926 3858 21978
rect 3910 21926 3962 21978
rect 4014 21926 4066 21978
rect 23806 21926 23858 21978
rect 23910 21926 23962 21978
rect 24014 21926 24066 21978
rect 4286 21758 4338 21810
rect 11678 21758 11730 21810
rect 12798 21758 12850 21810
rect 13134 21758 13186 21810
rect 27246 21758 27298 21810
rect 1710 21646 1762 21698
rect 5518 21646 5570 21698
rect 18734 21646 18786 21698
rect 2718 21534 2770 21586
rect 6750 21534 6802 21586
rect 7086 21534 7138 21586
rect 7870 21534 7922 21586
rect 8542 21534 8594 21586
rect 9438 21534 9490 21586
rect 10110 21534 10162 21586
rect 13582 21534 13634 21586
rect 14478 21534 14530 21586
rect 15822 21534 15874 21586
rect 16382 21534 16434 21586
rect 3054 21422 3106 21474
rect 6302 21422 6354 21474
rect 10446 21422 10498 21474
rect 12238 21422 12290 21474
rect 15262 21422 15314 21474
rect 16718 21422 16770 21474
rect 17166 21422 17218 21474
rect 18286 21422 18338 21474
rect 19294 21422 19346 21474
rect 26238 21422 26290 21474
rect 2158 21310 2210 21362
rect 5966 21310 6018 21362
rect 7310 21310 7362 21362
rect 12126 21310 12178 21362
rect 12910 21310 12962 21362
rect 15710 21310 15762 21362
rect 19854 21310 19906 21362
rect 4466 21142 4518 21194
rect 4570 21142 4622 21194
rect 4674 21142 4726 21194
rect 24466 21142 24518 21194
rect 24570 21142 24622 21194
rect 24674 21142 24726 21194
rect 1374 20974 1426 21026
rect 3278 20974 3330 21026
rect 7870 20974 7922 21026
rect 9774 20974 9826 21026
rect 17614 20974 17666 21026
rect 18734 20974 18786 21026
rect 19854 20974 19906 21026
rect 1934 20862 1986 20914
rect 2270 20862 2322 20914
rect 3726 20862 3778 20914
rect 6750 20862 6802 20914
rect 9550 20862 9602 20914
rect 13918 20862 13970 20914
rect 20414 20862 20466 20914
rect 20750 20862 20802 20914
rect 2606 20750 2658 20802
rect 3054 20750 3106 20802
rect 4510 20750 4562 20802
rect 5294 20750 5346 20802
rect 9886 20750 9938 20802
rect 9998 20750 10050 20802
rect 10446 20750 10498 20802
rect 11006 20750 11058 20802
rect 11566 20750 11618 20802
rect 11902 20750 11954 20802
rect 13358 20750 13410 20802
rect 13806 20750 13858 20802
rect 14590 20750 14642 20802
rect 14926 20750 14978 20802
rect 15934 20750 15986 20802
rect 16718 20750 16770 20802
rect 19182 20750 19234 20802
rect 20190 20750 20242 20802
rect 6302 20638 6354 20690
rect 11790 20638 11842 20690
rect 12910 20638 12962 20690
rect 10782 20526 10834 20578
rect 16718 20526 16770 20578
rect 17054 20526 17106 20578
rect 3806 20358 3858 20410
rect 3910 20358 3962 20410
rect 4014 20358 4066 20410
rect 23806 20358 23858 20410
rect 23910 20358 23962 20410
rect 24014 20358 24066 20410
rect 2830 20190 2882 20242
rect 12910 20190 12962 20242
rect 16046 20190 16098 20242
rect 6750 20078 6802 20130
rect 8318 20078 8370 20130
rect 8990 20078 9042 20130
rect 10558 20078 10610 20130
rect 13246 20078 13298 20130
rect 15038 20078 15090 20130
rect 18174 20078 18226 20130
rect 19742 20078 19794 20130
rect 1262 19966 1314 20018
rect 3614 19966 3666 20018
rect 8878 19966 8930 20018
rect 11454 19966 11506 20018
rect 11902 19966 11954 20018
rect 12238 19966 12290 20018
rect 14702 19966 14754 20018
rect 15486 19966 15538 20018
rect 15822 19966 15874 20018
rect 16270 19966 16322 20018
rect 1038 19854 1090 19906
rect 6190 19854 6242 19906
rect 9326 19854 9378 19906
rect 11678 19854 11730 19906
rect 13470 19854 13522 19906
rect 13806 19854 13858 19906
rect 18510 19854 18562 19906
rect 1598 19742 1650 19794
rect 5630 19742 5682 19794
rect 7198 19742 7250 19794
rect 11790 19742 11842 19794
rect 15598 19742 15650 19794
rect 4466 19574 4518 19626
rect 4570 19574 4622 19626
rect 4674 19574 4726 19626
rect 24466 19574 24518 19626
rect 24570 19574 24622 19626
rect 24674 19574 24726 19626
rect 1598 19406 1650 19458
rect 5742 19406 5794 19458
rect 8206 19406 8258 19458
rect 11566 19406 11618 19458
rect 2718 19294 2770 19346
rect 4510 19294 4562 19346
rect 6974 19294 7026 19346
rect 11118 19294 11170 19346
rect 12574 19294 12626 19346
rect 13918 19294 13970 19346
rect 14366 19294 14418 19346
rect 16718 19294 16770 19346
rect 16942 19294 16994 19346
rect 6638 19182 6690 19234
rect 9550 19182 9602 19234
rect 10334 19182 10386 19234
rect 11790 19182 11842 19234
rect 12126 19182 12178 19234
rect 12910 19182 12962 19234
rect 13358 19182 13410 19234
rect 13806 19182 13858 19234
rect 14926 19182 14978 19234
rect 16046 19182 16098 19234
rect 3166 19070 3218 19122
rect 4174 19070 4226 19122
rect 16830 19070 16882 19122
rect 3806 18790 3858 18842
rect 3910 18790 3962 18842
rect 4014 18790 4066 18842
rect 23806 18790 23858 18842
rect 23910 18790 23962 18842
rect 24014 18790 24066 18842
rect 7198 18622 7250 18674
rect 13806 18622 13858 18674
rect 15822 18622 15874 18674
rect 3166 18510 3218 18562
rect 4286 18510 4338 18562
rect 10334 18510 10386 18562
rect 16046 18510 16098 18562
rect 16270 18510 16322 18562
rect 1486 18398 1538 18450
rect 2270 18398 2322 18450
rect 2718 18398 2770 18450
rect 3950 18398 4002 18450
rect 5630 18398 5682 18450
rect 8094 18398 8146 18450
rect 14590 18398 14642 18450
rect 15598 18398 15650 18450
rect 19518 18398 19570 18450
rect 5966 18286 6018 18338
rect 8430 18286 8482 18338
rect 14366 18286 14418 18338
rect 15262 18286 15314 18338
rect 1710 18174 1762 18226
rect 9662 18174 9714 18226
rect 10782 18174 10834 18226
rect 11902 18174 11954 18226
rect 13470 18174 13522 18226
rect 15150 18174 15202 18226
rect 16270 18174 16322 18226
rect 16494 18174 16546 18226
rect 16942 18174 16994 18226
rect 17054 18174 17106 18226
rect 17166 18174 17218 18226
rect 17390 18174 17442 18226
rect 18958 18174 19010 18226
rect 4466 18006 4518 18058
rect 4570 18006 4622 18058
rect 4674 18006 4726 18058
rect 24466 18006 24518 18058
rect 24570 18006 24622 18058
rect 24674 18006 24726 18058
rect 1038 17838 1090 17890
rect 4846 17838 4898 17890
rect 11230 17838 11282 17890
rect 14478 17838 14530 17890
rect 16046 17838 16098 17890
rect 2606 17726 2658 17778
rect 6974 17726 7026 17778
rect 9998 17726 10050 17778
rect 2046 17614 2098 17666
rect 3726 17614 3778 17666
rect 4286 17614 4338 17666
rect 6638 17614 6690 17666
rect 9550 17614 9602 17666
rect 12350 17614 12402 17666
rect 13246 17614 13298 17666
rect 13806 17614 13858 17666
rect 14030 17614 14082 17666
rect 14702 17614 14754 17666
rect 15038 17614 15090 17666
rect 1598 17502 1650 17554
rect 4398 17502 4450 17554
rect 9662 17502 9714 17554
rect 15486 17502 15538 17554
rect 16158 17502 16210 17554
rect 5966 17390 6018 17442
rect 8206 17390 8258 17442
rect 15822 17390 15874 17442
rect 3806 17222 3858 17274
rect 3910 17222 3962 17274
rect 4014 17222 4066 17274
rect 23806 17222 23858 17274
rect 23910 17222 23962 17274
rect 24014 17222 24066 17274
rect 12798 17054 12850 17106
rect 13134 17054 13186 17106
rect 14254 17054 14306 17106
rect 1038 16942 1090 16994
rect 2494 16942 2546 16994
rect 8318 16942 8370 16994
rect 10222 16942 10274 16994
rect 12126 16942 12178 16994
rect 14926 16942 14978 16994
rect 1486 16830 1538 16882
rect 3838 16830 3890 16882
rect 4958 16830 5010 16882
rect 6638 16830 6690 16882
rect 10558 16830 10610 16882
rect 10894 16830 10946 16882
rect 11006 16830 11058 16882
rect 11790 16830 11842 16882
rect 13806 16830 13858 16882
rect 14030 16830 14082 16882
rect 14366 16830 14418 16882
rect 15262 16830 15314 16882
rect 15710 16830 15762 16882
rect 16382 16830 16434 16882
rect 16942 16830 16994 16882
rect 17950 16830 18002 16882
rect 7086 16718 7138 16770
rect 9886 16718 9938 16770
rect 10110 16718 10162 16770
rect 11342 16718 11394 16770
rect 12910 16718 12962 16770
rect 15934 16718 15986 16770
rect 1934 16606 1986 16658
rect 4398 16606 4450 16658
rect 5518 16606 5570 16658
rect 11230 16606 11282 16658
rect 14590 16606 14642 16658
rect 4466 16438 4518 16490
rect 4570 16438 4622 16490
rect 4674 16438 4726 16490
rect 24466 16438 24518 16490
rect 24570 16438 24622 16490
rect 24674 16438 24726 16490
rect 3054 16270 3106 16322
rect 4734 16270 4786 16322
rect 10110 16270 10162 16322
rect 11790 16270 11842 16322
rect 17950 16270 18002 16322
rect 6862 16158 6914 16210
rect 9550 16158 9602 16210
rect 10334 16158 10386 16210
rect 12238 16158 12290 16210
rect 15262 16158 15314 16210
rect 15710 16158 15762 16210
rect 3614 16046 3666 16098
rect 4174 16046 4226 16098
rect 6526 16046 6578 16098
rect 9102 16046 9154 16098
rect 9326 16046 9378 16098
rect 9886 16046 9938 16098
rect 9998 16046 10050 16098
rect 11118 16046 11170 16098
rect 11678 16046 11730 16098
rect 13022 16046 13074 16098
rect 13918 16046 13970 16098
rect 15934 16046 15986 16098
rect 16270 16046 16322 16098
rect 18398 16046 18450 16098
rect 8094 15934 8146 15986
rect 10782 15934 10834 15986
rect 1934 15822 1986 15874
rect 5854 15822 5906 15874
rect 9662 15822 9714 15874
rect 15374 15822 15426 15874
rect 16046 15822 16098 15874
rect 16830 15822 16882 15874
rect 3806 15654 3858 15706
rect 3910 15654 3962 15706
rect 4014 15654 4066 15706
rect 23806 15654 23858 15706
rect 23910 15654 23962 15706
rect 24014 15654 24066 15706
rect 11230 15486 11282 15538
rect 11902 15486 11954 15538
rect 3502 15374 3554 15426
rect 5742 15374 5794 15426
rect 9550 15374 9602 15426
rect 11006 15374 11058 15426
rect 15262 15374 15314 15426
rect 16494 15374 16546 15426
rect 18510 15374 18562 15426
rect 7870 15262 7922 15314
rect 10110 15262 10162 15314
rect 10558 15262 10610 15314
rect 11454 15262 11506 15314
rect 11790 15262 11842 15314
rect 13694 15262 13746 15314
rect 15150 15262 15202 15314
rect 15822 15262 15874 15314
rect 16046 15262 16098 15314
rect 3166 15150 3218 15202
rect 6078 15150 6130 15202
rect 8318 15150 8370 15202
rect 10782 15150 10834 15202
rect 11902 15150 11954 15202
rect 14926 15150 14978 15202
rect 15934 15150 15986 15202
rect 16942 15150 16994 15202
rect 18062 15150 18114 15202
rect 1934 15038 1986 15090
rect 7310 15038 7362 15090
rect 9998 15038 10050 15090
rect 10670 15038 10722 15090
rect 13358 15038 13410 15090
rect 15374 15038 15426 15090
rect 4466 14870 4518 14922
rect 4570 14870 4622 14922
rect 4674 14870 4726 14922
rect 24466 14870 24518 14922
rect 24570 14870 24622 14922
rect 24674 14870 24726 14922
rect 1934 14702 1986 14754
rect 2830 14702 2882 14754
rect 9438 14702 9490 14754
rect 11118 14702 11170 14754
rect 11230 14702 11282 14754
rect 14366 14702 14418 14754
rect 15486 14702 15538 14754
rect 16270 14702 16322 14754
rect 17614 14702 17666 14754
rect 4510 14590 4562 14642
rect 5518 14590 5570 14642
rect 5966 14590 6018 14642
rect 9550 14590 9602 14642
rect 10110 14590 10162 14642
rect 10222 14590 10274 14642
rect 15934 14590 15986 14642
rect 16046 14590 16098 14642
rect 4846 14478 4898 14530
rect 5294 14478 5346 14530
rect 6526 14478 6578 14530
rect 7646 14478 7698 14530
rect 9998 14478 10050 14530
rect 10670 14478 10722 14530
rect 16718 14478 16770 14530
rect 17166 14478 17218 14530
rect 17390 14478 17442 14530
rect 2494 14366 2546 14418
rect 3278 14366 3330 14418
rect 13918 14366 13970 14418
rect 17502 14366 17554 14418
rect 9438 14254 9490 14306
rect 11006 14254 11058 14306
rect 16942 14254 16994 14306
rect 3806 14086 3858 14138
rect 3910 14086 3962 14138
rect 4014 14086 4066 14138
rect 23806 14086 23858 14138
rect 23910 14086 23962 14138
rect 24014 14086 24066 14138
rect 7422 13918 7474 13970
rect 16942 13918 16994 13970
rect 17278 13918 17330 13970
rect 17390 13918 17442 13970
rect 1150 13806 1202 13858
rect 16382 13806 16434 13858
rect 1598 13694 1650 13746
rect 1934 13694 1986 13746
rect 2606 13694 2658 13746
rect 3390 13694 3442 13746
rect 4286 13694 4338 13746
rect 5182 13694 5234 13746
rect 8206 13694 8258 13746
rect 9326 13694 9378 13746
rect 13134 13694 13186 13746
rect 15710 13694 15762 13746
rect 16046 13694 16098 13746
rect 16158 13694 16210 13746
rect 16494 13694 16546 13746
rect 17054 13694 17106 13746
rect 5630 13582 5682 13634
rect 9774 13582 9826 13634
rect 13694 13582 13746 13634
rect 15262 13582 15314 13634
rect 15374 13582 15426 13634
rect 2158 13470 2210 13522
rect 6750 13470 6802 13522
rect 11006 13470 11058 13522
rect 14814 13470 14866 13522
rect 4466 13302 4518 13354
rect 4570 13302 4622 13354
rect 4674 13302 4726 13354
rect 24466 13302 24518 13354
rect 24570 13302 24622 13354
rect 24674 13302 24726 13354
rect 2606 13134 2658 13186
rect 7758 13134 7810 13186
rect 15374 13134 15426 13186
rect 16046 13134 16098 13186
rect 3726 13022 3778 13074
rect 5182 13022 5234 13074
rect 9438 13022 9490 13074
rect 11902 13022 11954 13074
rect 14478 13022 14530 13074
rect 14814 13022 14866 13074
rect 15262 13022 15314 13074
rect 16158 13022 16210 13074
rect 2158 12910 2210 12962
rect 4510 12910 4562 12962
rect 4958 12910 5010 12962
rect 5854 12910 5906 12962
rect 6414 12910 6466 12962
rect 7198 12910 7250 12962
rect 11342 12910 11394 12962
rect 12238 12910 12290 12962
rect 12798 12910 12850 12962
rect 4174 12798 4226 12850
rect 8206 12798 8258 12850
rect 9102 12798 9154 12850
rect 15486 12798 15538 12850
rect 10670 12686 10722 12738
rect 3806 12518 3858 12570
rect 3910 12518 3962 12570
rect 4014 12518 4066 12570
rect 23806 12518 23858 12570
rect 23910 12518 23962 12570
rect 24014 12518 24066 12570
rect 1598 12238 1650 12290
rect 2494 12238 2546 12290
rect 3278 12238 3330 12290
rect 5966 12238 6018 12290
rect 12798 12238 12850 12290
rect 1150 12126 1202 12178
rect 2046 12126 2098 12178
rect 2830 12126 2882 12178
rect 5518 12126 5570 12178
rect 6862 12126 6914 12178
rect 8542 12126 8594 12178
rect 9326 12126 9378 12178
rect 9886 12126 9938 12178
rect 10670 12126 10722 12178
rect 11230 12126 11282 12178
rect 12126 12126 12178 12178
rect 13134 12126 13186 12178
rect 13582 12126 13634 12178
rect 15038 12126 15090 12178
rect 15934 12126 15986 12178
rect 7310 12014 7362 12066
rect 8990 12014 9042 12066
rect 9998 12014 10050 12066
rect 14254 12014 14306 12066
rect 13806 11902 13858 11954
rect 4466 11734 4518 11786
rect 4570 11734 4622 11786
rect 4674 11734 4726 11786
rect 24466 11734 24518 11786
rect 24570 11734 24622 11786
rect 24674 11734 24726 11786
rect 10894 11566 10946 11618
rect 2270 11454 2322 11506
rect 2606 11454 2658 11506
rect 3166 11454 3218 11506
rect 4846 11454 4898 11506
rect 6974 11454 7026 11506
rect 9886 11454 9938 11506
rect 14702 11454 14754 11506
rect 15150 11454 15202 11506
rect 4286 11342 4338 11394
rect 6638 11342 6690 11394
rect 8206 11342 8258 11394
rect 10222 11342 10274 11394
rect 10782 11342 10834 11394
rect 11454 11342 11506 11394
rect 12014 11342 12066 11394
rect 13022 11342 13074 11394
rect 1262 11118 1314 11170
rect 5966 11118 6018 11170
rect 14142 11118 14194 11170
rect 14478 11118 14530 11170
rect 3806 10950 3858 11002
rect 3910 10950 3962 11002
rect 4014 10950 4066 11002
rect 23806 10950 23858 11002
rect 23910 10950 23962 11002
rect 24014 10950 24066 11002
rect 12126 10782 12178 10834
rect 5854 10670 5906 10722
rect 6750 10670 6802 10722
rect 14030 10670 14082 10722
rect 14926 10670 14978 10722
rect 5406 10558 5458 10610
rect 7086 10558 7138 10610
rect 7534 10558 7586 10610
rect 8318 10558 8370 10610
rect 8990 10558 9042 10610
rect 9886 10558 9938 10610
rect 10446 10558 10498 10610
rect 13582 10558 13634 10610
rect 14366 10558 14418 10610
rect 10894 10446 10946 10498
rect 7758 10334 7810 10386
rect 4466 10166 4518 10218
rect 4570 10166 4622 10218
rect 4674 10166 4726 10218
rect 24466 10166 24518 10218
rect 24570 10166 24622 10218
rect 24674 10166 24726 10218
rect 7534 9998 7586 10050
rect 4734 9886 4786 9938
rect 10110 9886 10162 9938
rect 11118 9886 11170 9938
rect 2158 9774 2210 9826
rect 5182 9774 5234 9826
rect 10446 9774 10498 9826
rect 10894 9774 10946 9826
rect 11566 9774 11618 9826
rect 12126 9774 12178 9826
rect 13134 9774 13186 9826
rect 6974 9662 7026 9714
rect 1262 9550 1314 9602
rect 3806 9382 3858 9434
rect 3910 9382 3962 9434
rect 4014 9382 4066 9434
rect 23806 9382 23858 9434
rect 23910 9382 23962 9434
rect 24014 9382 24066 9434
rect 8878 9214 8930 9266
rect 11118 9214 11170 9266
rect 7310 9102 7362 9154
rect 9550 9102 9602 9154
rect 7646 8878 7698 8930
rect 9886 8878 9938 8930
rect 4466 8598 4518 8650
rect 4570 8598 4622 8650
rect 4674 8598 4726 8650
rect 24466 8598 24518 8650
rect 24570 8598 24622 8650
rect 24674 8598 24726 8650
rect 7758 8430 7810 8482
rect 11342 8430 11394 8482
rect 10222 8318 10274 8370
rect 9662 8206 9714 8258
rect 8318 8094 8370 8146
rect 3806 7814 3858 7866
rect 3910 7814 3962 7866
rect 4014 7814 4066 7866
rect 23806 7814 23858 7866
rect 23910 7814 23962 7866
rect 24014 7814 24066 7866
rect 11566 7534 11618 7586
rect 10222 7422 10274 7474
rect 11006 7422 11058 7474
rect 10670 7310 10722 7362
rect 4466 7030 4518 7082
rect 4570 7030 4622 7082
rect 4674 7030 4726 7082
rect 24466 7030 24518 7082
rect 24570 7030 24622 7082
rect 24674 7030 24726 7082
rect 2270 6750 2322 6802
rect 1262 6526 1314 6578
rect 3806 6246 3858 6298
rect 3910 6246 3962 6298
rect 4014 6246 4066 6298
rect 23806 6246 23858 6298
rect 23910 6246 23962 6298
rect 24014 6246 24066 6298
rect 1262 5966 1314 6018
rect 2270 5854 2322 5906
rect 4466 5462 4518 5514
rect 4570 5462 4622 5514
rect 4674 5462 4726 5514
rect 24466 5462 24518 5514
rect 24570 5462 24622 5514
rect 24674 5462 24726 5514
rect 3806 4678 3858 4730
rect 3910 4678 3962 4730
rect 4014 4678 4066 4730
rect 23806 4678 23858 4730
rect 23910 4678 23962 4730
rect 24014 4678 24066 4730
rect 4466 3894 4518 3946
rect 4570 3894 4622 3946
rect 4674 3894 4726 3946
rect 24466 3894 24518 3946
rect 24570 3894 24622 3946
rect 24674 3894 24726 3946
rect 3806 3110 3858 3162
rect 3910 3110 3962 3162
rect 4014 3110 4066 3162
rect 23806 3110 23858 3162
rect 23910 3110 23962 3162
rect 24014 3110 24066 3162
rect 4466 2326 4518 2378
rect 4570 2326 4622 2378
rect 4674 2326 4726 2378
rect 24466 2326 24518 2378
rect 24570 2326 24622 2378
rect 24674 2326 24726 2378
rect 3806 1542 3858 1594
rect 3910 1542 3962 1594
rect 4014 1542 4066 1594
rect 23806 1542 23858 1594
rect 23910 1542 23962 1594
rect 24014 1542 24066 1594
rect 4466 758 4518 810
rect 4570 758 4622 810
rect 4674 758 4726 810
rect 24466 758 24518 810
rect 24570 758 24622 810
rect 24674 758 24726 810
<< metal2 >>
rect 672 57344 784 57456
rect 2016 57344 2128 57456
rect 3360 57344 3472 57456
rect 4704 57344 4816 57456
rect 6048 57344 6160 57456
rect 7392 57344 7504 57456
rect 8736 57344 8848 57456
rect 10080 57344 10192 57456
rect 11424 57344 11536 57456
rect 12768 57344 12880 57456
rect 14112 57344 14224 57456
rect 15456 57344 15568 57456
rect 16800 57344 16912 57456
rect 18144 57344 18256 57456
rect 19488 57344 19600 57456
rect 20832 57344 20944 57456
rect 22176 57344 22288 57456
rect 23520 57344 23632 57456
rect 24864 57344 24976 57456
rect 26208 57344 26320 57456
rect 27552 57344 27664 57456
rect 700 55972 756 57344
rect 1036 55972 1092 55982
rect 700 55970 1092 55972
rect 700 55918 1038 55970
rect 1090 55918 1092 55970
rect 700 55916 1092 55918
rect 1036 55906 1092 55916
rect 1372 55858 1428 55870
rect 1372 55806 1374 55858
rect 1426 55806 1428 55858
rect 364 53620 420 53630
rect 252 36148 308 36158
rect 140 29204 196 29214
rect 140 13300 196 29148
rect 252 26180 308 36092
rect 252 26114 308 26124
rect 364 19348 420 53564
rect 1372 52948 1428 55806
rect 2044 55468 2100 57344
rect 3388 56308 3444 57344
rect 4732 57316 4788 57344
rect 4732 57250 4788 57260
rect 5516 57316 5572 57326
rect 3804 56476 4068 56486
rect 3860 56420 3908 56476
rect 3964 56420 4012 56476
rect 3804 56410 4068 56420
rect 3612 56308 3668 56318
rect 3388 56306 3668 56308
rect 3388 56254 3614 56306
rect 3666 56254 3668 56306
rect 3388 56252 3668 56254
rect 3612 56242 3668 56252
rect 5516 56306 5572 57260
rect 6076 57204 6132 57344
rect 6076 57148 6580 57204
rect 5516 56254 5518 56306
rect 5570 56254 5572 56306
rect 5516 56242 5572 56254
rect 5180 56082 5236 56094
rect 5180 56030 5182 56082
rect 5234 56030 5236 56082
rect 3052 55972 3108 55982
rect 3052 55878 3108 55916
rect 4464 55692 4728 55702
rect 4520 55636 4568 55692
rect 4624 55636 4672 55692
rect 4464 55626 4728 55636
rect 5180 55468 5236 56030
rect 2044 55412 2548 55468
rect 5180 55412 6468 55468
rect 2492 55186 2548 55412
rect 2492 55134 2494 55186
rect 2546 55134 2548 55186
rect 2492 55122 2548 55134
rect 3500 55298 3556 55310
rect 3500 55246 3502 55298
rect 3554 55246 3556 55298
rect 1372 52882 1428 52892
rect 1820 52276 1876 52286
rect 1484 42980 1540 42990
rect 812 40180 868 40190
rect 588 38836 644 38846
rect 476 37044 532 37054
rect 476 28084 532 36988
rect 476 28018 532 28028
rect 588 28756 644 38780
rect 588 19796 644 28700
rect 588 19730 644 19740
rect 700 30996 756 31006
rect 364 19282 420 19292
rect 700 13860 756 30940
rect 812 29316 868 40124
rect 1148 37828 1204 37838
rect 1148 37826 1428 37828
rect 1148 37774 1150 37826
rect 1202 37774 1428 37826
rect 1148 37772 1428 37774
rect 1148 37762 1204 37772
rect 1260 37604 1316 37614
rect 812 20580 868 29260
rect 924 37492 980 37502
rect 924 27748 980 37436
rect 1036 37044 1092 37054
rect 1036 36950 1092 36988
rect 1260 36482 1316 37548
rect 1260 36430 1262 36482
rect 1314 36430 1316 36482
rect 1260 36418 1316 36430
rect 1372 34132 1428 37772
rect 1484 37378 1540 42924
rect 1708 41300 1764 41310
rect 1708 40404 1764 41244
rect 1708 40310 1764 40348
rect 1708 39618 1764 39630
rect 1708 39566 1710 39618
rect 1762 39566 1764 39618
rect 1708 38724 1764 39566
rect 1596 38610 1652 38622
rect 1596 38558 1598 38610
rect 1650 38558 1652 38610
rect 1596 38276 1652 38558
rect 1708 38612 1764 38668
rect 1708 38546 1764 38556
rect 1596 38220 1764 38276
rect 1484 37326 1486 37378
rect 1538 37326 1540 37378
rect 1484 37314 1540 37326
rect 1596 38052 1652 38062
rect 1596 37156 1652 37996
rect 1484 37100 1652 37156
rect 1484 36372 1540 37100
rect 1596 36932 1652 36942
rect 1596 36594 1652 36876
rect 1596 36542 1598 36594
rect 1650 36542 1652 36594
rect 1596 36530 1652 36542
rect 1708 36596 1764 38220
rect 1708 36530 1764 36540
rect 1484 36316 1652 36372
rect 1484 34132 1540 34142
rect 1372 34130 1540 34132
rect 1372 34078 1486 34130
rect 1538 34078 1540 34130
rect 1372 34076 1540 34078
rect 1484 34066 1540 34076
rect 1148 34018 1204 34030
rect 1148 33966 1150 34018
rect 1202 33966 1204 34018
rect 924 27682 980 27692
rect 1036 30210 1092 30222
rect 1036 30158 1038 30210
rect 1090 30158 1092 30210
rect 1036 27858 1092 30158
rect 1148 30212 1204 33966
rect 1596 33458 1652 36316
rect 1708 34802 1764 34814
rect 1708 34750 1710 34802
rect 1762 34750 1764 34802
rect 1708 34356 1764 34750
rect 1708 34290 1764 34300
rect 1596 33406 1598 33458
rect 1650 33406 1652 33458
rect 1260 33234 1316 33246
rect 1260 33182 1262 33234
rect 1314 33182 1316 33234
rect 1260 32564 1316 33182
rect 1596 32788 1652 33406
rect 1484 32732 1652 32788
rect 1708 33236 1764 33246
rect 1316 32508 1428 32564
rect 1260 32498 1316 32508
rect 1260 31668 1316 31678
rect 1260 30996 1316 31612
rect 1260 30902 1316 30940
rect 1148 30146 1204 30156
rect 1036 27806 1038 27858
rect 1090 27806 1092 27858
rect 812 20514 868 20524
rect 924 26964 980 26974
rect 700 13794 756 13804
rect 140 13234 196 13244
rect 924 12292 980 26908
rect 1036 26908 1092 27806
rect 1260 29540 1316 29550
rect 1372 29540 1428 32508
rect 1260 29538 1428 29540
rect 1260 29486 1262 29538
rect 1314 29486 1428 29538
rect 1260 29484 1428 29486
rect 1260 28644 1316 29484
rect 1484 29204 1540 32732
rect 1596 32564 1652 32574
rect 1596 32470 1652 32508
rect 1708 31668 1764 33180
rect 1820 32788 1876 52220
rect 1932 50932 1988 50942
rect 1932 40628 1988 50876
rect 3276 46900 3332 46910
rect 2268 44996 2324 45006
rect 1932 40562 1988 40572
rect 2044 42084 2100 42094
rect 1932 40404 1988 40414
rect 1932 37268 1988 40348
rect 2044 38946 2100 42028
rect 2156 40628 2212 40638
rect 2156 40514 2212 40572
rect 2156 40462 2158 40514
rect 2210 40462 2212 40514
rect 2156 40450 2212 40462
rect 2044 38894 2046 38946
rect 2098 38894 2100 38946
rect 2044 38882 2100 38894
rect 2156 40292 2212 40302
rect 2156 38668 2212 40236
rect 2268 39730 2324 44940
rect 3276 41748 3332 46844
rect 3500 43652 3556 55246
rect 3804 54908 4068 54918
rect 3860 54852 3908 54908
rect 3964 54852 4012 54908
rect 3804 54842 4068 54852
rect 4464 54124 4728 54134
rect 4520 54068 4568 54124
rect 4624 54068 4672 54124
rect 4464 54058 4728 54068
rect 3804 53340 4068 53350
rect 3860 53284 3908 53340
rect 3964 53284 4012 53340
rect 3804 53274 4068 53284
rect 6300 53060 6356 53070
rect 4464 52556 4728 52566
rect 4520 52500 4568 52556
rect 4624 52500 4672 52556
rect 4464 52490 4728 52500
rect 5964 51940 6020 51950
rect 3804 51772 4068 51782
rect 3860 51716 3908 51772
rect 3964 51716 4012 51772
rect 3804 51706 4068 51716
rect 4172 51380 4228 51390
rect 3804 50204 4068 50214
rect 3860 50148 3908 50204
rect 3964 50148 4012 50204
rect 3804 50138 4068 50148
rect 3804 48636 4068 48646
rect 3860 48580 3908 48636
rect 3964 48580 4012 48636
rect 3804 48570 4068 48580
rect 3804 47068 4068 47078
rect 3860 47012 3908 47068
rect 3964 47012 4012 47068
rect 3804 47002 4068 47012
rect 3804 45500 4068 45510
rect 3860 45444 3908 45500
rect 3964 45444 4012 45500
rect 3804 45434 4068 45444
rect 3804 43932 4068 43942
rect 3860 43876 3908 43932
rect 3964 43876 4012 43932
rect 3804 43866 4068 43876
rect 3500 43586 3556 43596
rect 3804 42364 4068 42374
rect 3860 42308 3908 42364
rect 3964 42308 4012 42364
rect 3804 42298 4068 42308
rect 4172 41970 4228 51324
rect 4464 50988 4728 50998
rect 4520 50932 4568 50988
rect 4624 50932 4672 50988
rect 4464 50922 4728 50932
rect 5740 49588 5796 49598
rect 4464 49420 4728 49430
rect 4520 49364 4568 49420
rect 4624 49364 4672 49420
rect 4464 49354 4728 49364
rect 4464 47852 4728 47862
rect 4520 47796 4568 47852
rect 4624 47796 4672 47852
rect 4464 47786 4728 47796
rect 4464 46284 4728 46294
rect 4520 46228 4568 46284
rect 4624 46228 4672 46284
rect 4464 46218 4728 46228
rect 4464 44716 4728 44726
rect 4520 44660 4568 44716
rect 4624 44660 4672 44716
rect 4464 44650 4728 44660
rect 4464 43148 4728 43158
rect 4520 43092 4568 43148
rect 4624 43092 4672 43148
rect 4464 43082 4728 43092
rect 4172 41918 4174 41970
rect 4226 41918 4228 41970
rect 4172 41906 4228 41918
rect 3612 41748 3668 41758
rect 3276 41746 3668 41748
rect 3276 41694 3614 41746
rect 3666 41694 3668 41746
rect 3276 41692 3668 41694
rect 3276 41188 3332 41692
rect 3612 41682 3668 41692
rect 4464 41580 4728 41590
rect 4520 41524 4568 41580
rect 4624 41524 4672 41580
rect 4464 41514 4728 41524
rect 5292 41412 5348 41422
rect 4284 41300 4340 41310
rect 4284 41206 4340 41244
rect 3836 41188 3892 41198
rect 2604 40404 2660 40414
rect 2268 39678 2270 39730
rect 2322 39678 2324 39730
rect 2268 39666 2324 39678
rect 2492 40402 2660 40404
rect 2492 40350 2606 40402
rect 2658 40350 2660 40402
rect 2492 40348 2660 40350
rect 1932 37202 1988 37212
rect 2044 38612 2212 38668
rect 2044 37266 2100 38612
rect 2380 38164 2436 38174
rect 2044 37214 2046 37266
rect 2098 37214 2100 37266
rect 2044 37202 2100 37214
rect 2268 37268 2324 37278
rect 1932 37042 1988 37054
rect 1932 36990 1934 37042
rect 1986 36990 1988 37042
rect 1932 36708 1988 36990
rect 1932 36642 1988 36652
rect 2044 36596 2100 36606
rect 1932 34130 1988 34142
rect 1932 34078 1934 34130
rect 1986 34078 1988 34130
rect 1932 33236 1988 34078
rect 1932 33170 1988 33180
rect 1820 32732 1988 32788
rect 1708 31602 1764 31612
rect 1820 31666 1876 31678
rect 1820 31614 1822 31666
rect 1874 31614 1876 31666
rect 1820 31220 1876 31614
rect 1820 31154 1876 31164
rect 1596 29316 1652 29326
rect 1596 29222 1652 29260
rect 1484 29138 1540 29148
rect 1596 28756 1652 28766
rect 1596 28662 1652 28700
rect 1820 28644 1876 28654
rect 1260 28642 1540 28644
rect 1260 28590 1262 28642
rect 1314 28590 1540 28642
rect 1260 28588 1540 28590
rect 1260 27076 1316 28588
rect 1484 27970 1540 28588
rect 1484 27918 1486 27970
rect 1538 27918 1540 27970
rect 1484 27906 1540 27918
rect 1260 26982 1316 27020
rect 1484 27748 1540 27758
rect 1484 27188 1540 27692
rect 1596 27188 1652 27198
rect 1484 27186 1652 27188
rect 1484 27134 1598 27186
rect 1650 27134 1652 27186
rect 1484 27132 1652 27134
rect 1036 26852 1204 26908
rect 1036 26180 1092 26190
rect 1036 22596 1092 26124
rect 1148 25172 1204 26852
rect 1484 26068 1540 27132
rect 1596 27122 1652 27132
rect 1708 27076 1764 27086
rect 1708 26402 1764 27020
rect 1708 26350 1710 26402
rect 1762 26350 1764 26402
rect 1708 26338 1764 26350
rect 1148 25116 1428 25172
rect 1148 24948 1204 24958
rect 1148 23266 1204 24892
rect 1260 24724 1316 24734
rect 1260 24630 1316 24668
rect 1148 23214 1150 23266
rect 1202 23214 1204 23266
rect 1148 23202 1204 23214
rect 1148 22596 1204 22606
rect 1036 22594 1204 22596
rect 1036 22542 1150 22594
rect 1202 22542 1204 22594
rect 1036 22540 1204 22542
rect 1148 22530 1204 22540
rect 1372 21026 1428 25116
rect 1484 24162 1540 26012
rect 1484 24110 1486 24162
rect 1538 24110 1540 24162
rect 1484 24098 1540 24110
rect 1708 25508 1764 25518
rect 1708 23492 1764 25452
rect 1596 23436 1764 23492
rect 1596 23380 1652 23436
rect 1484 23324 1652 23380
rect 1484 21476 1540 23324
rect 1708 23268 1764 23278
rect 1596 23156 1652 23166
rect 1596 23062 1652 23100
rect 1596 22484 1652 22494
rect 1596 22258 1652 22428
rect 1596 22206 1598 22258
rect 1650 22206 1652 22258
rect 1596 22194 1652 22206
rect 1708 21698 1764 23212
rect 1820 22372 1876 28588
rect 1932 22596 1988 32732
rect 2044 32116 2100 36540
rect 2156 34914 2212 34926
rect 2156 34862 2158 34914
rect 2210 34862 2212 34914
rect 2156 34018 2212 34862
rect 2156 33966 2158 34018
rect 2210 33966 2212 34018
rect 2156 33954 2212 33966
rect 2156 32452 2212 32462
rect 2268 32452 2324 37212
rect 2156 32450 2268 32452
rect 2156 32398 2158 32450
rect 2210 32398 2268 32450
rect 2156 32396 2268 32398
rect 2156 32386 2212 32396
rect 2268 32358 2324 32396
rect 2044 32050 2100 32060
rect 2268 32116 2324 32126
rect 2268 31778 2324 32060
rect 2268 31726 2270 31778
rect 2322 31726 2324 31778
rect 2268 31714 2324 31726
rect 2380 31556 2436 38108
rect 2492 37604 2548 40348
rect 2604 40338 2660 40348
rect 3052 40290 3108 40302
rect 3052 40238 3054 40290
rect 3106 40238 3108 40290
rect 2604 39618 2660 39630
rect 2604 39566 2606 39618
rect 2658 39566 2660 39618
rect 2604 38668 2660 39566
rect 2716 38948 2772 38958
rect 2716 38854 2772 38892
rect 3052 38722 3108 40238
rect 3164 39732 3220 39742
rect 3164 39638 3220 39676
rect 3052 38670 3054 38722
rect 3106 38670 3108 38722
rect 3052 38668 3108 38670
rect 2604 38612 3108 38668
rect 2604 38164 2660 38612
rect 2604 38098 2660 38108
rect 2716 37938 2772 37950
rect 2716 37886 2718 37938
rect 2770 37886 2772 37938
rect 2716 37828 2772 37886
rect 2716 37604 2772 37772
rect 2492 37548 2660 37604
rect 2492 37380 2548 37390
rect 2492 37286 2548 37324
rect 2604 36484 2660 37548
rect 2716 37538 2772 37548
rect 3164 37940 3220 37950
rect 2604 35698 2660 36428
rect 3052 36708 3108 36718
rect 2604 35646 2606 35698
rect 2658 35646 2660 35698
rect 2604 34916 2660 35646
rect 2268 31500 2436 31556
rect 2492 34914 2660 34916
rect 2492 34862 2606 34914
rect 2658 34862 2660 34914
rect 2492 34860 2660 34862
rect 2492 34244 2548 34860
rect 2604 34850 2660 34860
rect 2828 36258 2884 36270
rect 2828 36206 2830 36258
rect 2882 36206 2884 36258
rect 2156 30212 2212 30222
rect 2044 29986 2100 29998
rect 2044 29934 2046 29986
rect 2098 29934 2100 29986
rect 2044 29540 2100 29934
rect 2044 29474 2100 29484
rect 2044 26180 2100 26190
rect 2044 25620 2100 26124
rect 2044 25554 2100 25564
rect 2044 25396 2100 25406
rect 2156 25396 2212 30156
rect 2268 29876 2324 31500
rect 2380 30994 2436 31006
rect 2380 30942 2382 30994
rect 2434 30942 2436 30994
rect 2380 30772 2436 30942
rect 2380 30706 2436 30716
rect 2492 30548 2548 34188
rect 2828 34130 2884 36206
rect 3052 35026 3108 36652
rect 3052 34974 3054 35026
rect 3106 34974 3108 35026
rect 3052 34962 3108 34974
rect 3164 35474 3220 37884
rect 3164 35422 3166 35474
rect 3218 35422 3220 35474
rect 3164 34692 3220 35422
rect 2828 34078 2830 34130
rect 2882 34078 2884 34130
rect 2828 34066 2884 34078
rect 2940 34636 3220 34692
rect 2828 33122 2884 33134
rect 2828 33070 2830 33122
rect 2882 33070 2884 33122
rect 2268 29810 2324 29820
rect 2380 30492 2548 30548
rect 2604 32452 2660 32462
rect 2044 25394 2212 25396
rect 2044 25342 2046 25394
rect 2098 25342 2212 25394
rect 2044 25340 2212 25342
rect 2268 29652 2324 29662
rect 2044 24164 2100 25340
rect 2268 25284 2324 29596
rect 2044 24098 2100 24108
rect 2156 25228 2324 25284
rect 2044 23940 2100 23950
rect 2156 23940 2212 25228
rect 2044 23938 2212 23940
rect 2044 23886 2046 23938
rect 2098 23886 2212 23938
rect 2044 23884 2212 23886
rect 2268 24722 2324 24734
rect 2268 24670 2270 24722
rect 2322 24670 2324 24722
rect 2044 23874 2100 23884
rect 2268 23828 2324 24670
rect 2268 23762 2324 23772
rect 2156 23716 2212 23726
rect 1932 22530 1988 22540
rect 2044 23604 2100 23614
rect 2044 22484 2100 23548
rect 2156 23154 2212 23660
rect 2156 23102 2158 23154
rect 2210 23102 2212 23154
rect 2156 23090 2212 23102
rect 2044 22428 2212 22484
rect 1820 22316 2100 22372
rect 1708 21646 1710 21698
rect 1762 21646 1764 21698
rect 1708 21634 1764 21646
rect 1484 21420 1764 21476
rect 1372 20974 1374 21026
rect 1426 20974 1428 21026
rect 1260 20020 1316 20030
rect 1372 20020 1428 20974
rect 1708 20132 1764 21420
rect 1932 20916 1988 20926
rect 1932 20822 1988 20860
rect 2044 20188 2100 22316
rect 2156 22148 2212 22428
rect 2268 22372 2324 22382
rect 2380 22372 2436 30492
rect 2604 29764 2660 32396
rect 2828 32116 2884 33070
rect 2828 32050 2884 32060
rect 2828 31892 2884 31902
rect 2828 31798 2884 31836
rect 2716 31780 2772 31790
rect 2716 31686 2772 31724
rect 2940 31668 2996 34636
rect 3276 34356 3332 41132
rect 3612 41186 3892 41188
rect 3612 41134 3838 41186
rect 3890 41134 3892 41186
rect 3612 41132 3892 41134
rect 3612 38948 3668 41132
rect 3836 41122 3892 41132
rect 3804 40796 4068 40806
rect 3860 40740 3908 40796
rect 3964 40740 4012 40796
rect 3804 40730 4068 40740
rect 4284 40404 4340 40414
rect 4284 40310 4340 40348
rect 5068 40180 5124 40190
rect 4464 40012 4728 40022
rect 4520 39956 4568 40012
rect 4624 39956 4672 40012
rect 4464 39946 4728 39956
rect 5068 39730 5124 40124
rect 5068 39678 5070 39730
rect 5122 39678 5124 39730
rect 5068 39666 5124 39678
rect 5292 39956 5348 41356
rect 3804 39228 4068 39238
rect 3860 39172 3908 39228
rect 3964 39172 4012 39228
rect 3804 39162 4068 39172
rect 3612 38882 3668 38892
rect 5180 38948 5236 38958
rect 4284 38836 4340 38846
rect 4284 38742 4340 38780
rect 4464 38444 4728 38454
rect 4520 38388 4568 38444
rect 4624 38388 4672 38444
rect 4464 38378 4728 38388
rect 5068 38162 5124 38174
rect 5068 38110 5070 38162
rect 5122 38110 5124 38162
rect 4620 38052 4676 38062
rect 3612 38050 4676 38052
rect 3612 37998 4622 38050
rect 4674 37998 4676 38050
rect 3612 37996 4676 37998
rect 3500 37268 3556 37278
rect 3388 36484 3444 36494
rect 3388 36390 3444 36428
rect 2828 31612 2996 31668
rect 3052 34300 3332 34356
rect 2828 30884 2884 31612
rect 2828 30818 2884 30828
rect 2940 30882 2996 30894
rect 2940 30830 2942 30882
rect 2994 30830 2996 30882
rect 2492 29708 2660 29764
rect 2716 30098 2772 30110
rect 2716 30046 2718 30098
rect 2770 30046 2772 30098
rect 2492 28644 2548 29708
rect 2492 28578 2548 28588
rect 2604 29540 2660 29550
rect 2604 27972 2660 29484
rect 2716 28756 2772 30046
rect 2828 30100 2884 30110
rect 2828 29650 2884 30044
rect 2828 29598 2830 29650
rect 2882 29598 2884 29650
rect 2828 29586 2884 29598
rect 2828 28868 2884 28878
rect 2940 28868 2996 30830
rect 2828 28866 2996 28868
rect 2828 28814 2830 28866
rect 2882 28814 2996 28866
rect 2828 28812 2996 28814
rect 2828 28802 2884 28812
rect 2716 28690 2772 28700
rect 2604 27858 2660 27916
rect 2604 27806 2606 27858
rect 2658 27806 2660 27858
rect 2604 27794 2660 27806
rect 3052 27746 3108 34300
rect 3276 34130 3332 34142
rect 3276 34078 3278 34130
rect 3330 34078 3332 34130
rect 3276 33572 3332 34078
rect 3276 33506 3332 33516
rect 3276 32338 3332 32350
rect 3276 32286 3278 32338
rect 3330 32286 3332 32338
rect 3276 31890 3332 32286
rect 3276 31838 3278 31890
rect 3330 31838 3332 31890
rect 3276 31826 3332 31838
rect 3500 31780 3556 37212
rect 3500 30994 3556 31724
rect 3500 30942 3502 30994
rect 3554 30942 3556 30994
rect 3500 30930 3556 30942
rect 3388 30772 3444 30782
rect 3612 30772 3668 37996
rect 4620 37986 4676 37996
rect 3804 37660 4068 37670
rect 3860 37604 3908 37660
rect 3964 37604 4012 37660
rect 3804 37594 4068 37604
rect 5068 37044 5124 38110
rect 5068 36978 5124 36988
rect 5180 37266 5236 38892
rect 5292 38668 5348 39900
rect 5516 40962 5572 40974
rect 5516 40910 5518 40962
rect 5570 40910 5572 40962
rect 5516 39618 5572 40910
rect 5516 39566 5518 39618
rect 5570 39566 5572 39618
rect 5516 39554 5572 39566
rect 5628 38948 5684 38958
rect 5628 38854 5684 38892
rect 5292 38612 5572 38668
rect 5180 37214 5182 37266
rect 5234 37214 5236 37266
rect 4464 36876 4728 36886
rect 4520 36820 4568 36876
rect 4624 36820 4672 36876
rect 4464 36810 4728 36820
rect 3948 36596 4004 36606
rect 3948 36502 4004 36540
rect 5180 36372 5236 37214
rect 5180 36316 5460 36372
rect 5068 36260 5124 36270
rect 5068 36258 5348 36260
rect 5068 36206 5070 36258
rect 5122 36206 5348 36258
rect 5068 36204 5348 36206
rect 5068 36194 5124 36204
rect 3804 36092 4068 36102
rect 3860 36036 3908 36092
rect 3964 36036 4012 36092
rect 3804 36026 4068 36036
rect 4284 35476 4340 35486
rect 4284 35474 5012 35476
rect 4284 35422 4286 35474
rect 4338 35422 5012 35474
rect 4284 35420 5012 35422
rect 4284 35410 4340 35420
rect 4464 35308 4728 35318
rect 4520 35252 4568 35308
rect 4624 35252 4672 35308
rect 4464 35242 4728 35252
rect 4284 34916 4340 34926
rect 4284 34822 4340 34860
rect 3804 34524 4068 34534
rect 3860 34468 3908 34524
rect 3964 34468 4012 34524
rect 3804 34458 4068 34468
rect 4284 34132 4340 34142
rect 4284 34038 4340 34076
rect 4464 33740 4728 33750
rect 4520 33684 4568 33740
rect 4624 33684 4672 33740
rect 4464 33674 4728 33684
rect 4172 33572 4228 33582
rect 3804 32956 4068 32966
rect 3860 32900 3908 32956
rect 3964 32900 4012 32956
rect 3804 32890 4068 32900
rect 3724 32338 3780 32350
rect 3724 32286 3726 32338
rect 3778 32286 3780 32338
rect 3724 31892 3780 32286
rect 3724 31826 3780 31836
rect 4060 31780 4116 31790
rect 4060 31686 4116 31724
rect 3804 31388 4068 31398
rect 3860 31332 3908 31388
rect 3964 31332 4012 31388
rect 3804 31322 4068 31332
rect 3164 30770 3444 30772
rect 3164 30718 3390 30770
rect 3442 30718 3444 30770
rect 3164 30716 3444 30718
rect 3164 30434 3220 30716
rect 3388 30706 3444 30716
rect 3500 30716 3668 30772
rect 3948 30994 4004 31006
rect 3948 30942 3950 30994
rect 4002 30942 4004 30994
rect 3164 30382 3166 30434
rect 3218 30382 3220 30434
rect 3164 30370 3220 30382
rect 3500 28756 3556 30716
rect 3948 30100 4004 30942
rect 3948 30034 4004 30044
rect 3804 29820 4068 29830
rect 3860 29764 3908 29820
rect 3964 29764 4012 29820
rect 3804 29754 4068 29764
rect 4060 29540 4116 29550
rect 3836 28756 3892 28766
rect 3388 28700 3556 28756
rect 3612 28754 3892 28756
rect 3612 28702 3838 28754
rect 3890 28702 3892 28754
rect 3612 28700 3892 28702
rect 3388 28308 3444 28700
rect 3500 28532 3556 28542
rect 3500 28438 3556 28476
rect 3388 28252 3556 28308
rect 3052 27694 3054 27746
rect 3106 27694 3108 27746
rect 3052 26908 3108 27694
rect 2492 26852 2548 26862
rect 2492 25506 2548 26796
rect 2828 26852 2884 26862
rect 2828 26758 2884 26796
rect 2940 26852 3108 26908
rect 3388 28084 3444 28094
rect 2492 25454 2494 25506
rect 2546 25454 2548 25506
rect 2492 25442 2548 25454
rect 2828 26180 2884 26190
rect 2828 25506 2884 26124
rect 2828 25454 2830 25506
rect 2882 25454 2884 25506
rect 2716 25396 2772 25406
rect 2716 24948 2772 25340
rect 2828 25284 2884 25454
rect 2828 25218 2884 25228
rect 2716 24892 2884 24948
rect 2716 24724 2772 24734
rect 2492 24722 2772 24724
rect 2492 24670 2718 24722
rect 2770 24670 2772 24722
rect 2492 24668 2772 24670
rect 2492 24162 2548 24668
rect 2716 24658 2772 24668
rect 2492 24110 2494 24162
rect 2546 24110 2548 24162
rect 2492 24098 2548 24110
rect 2716 23044 2772 23054
rect 2828 23044 2884 24892
rect 2268 22370 2436 22372
rect 2268 22318 2270 22370
rect 2322 22318 2436 22370
rect 2268 22316 2436 22318
rect 2268 22306 2324 22316
rect 2156 22092 2324 22148
rect 2268 21700 2324 22092
rect 2156 21362 2212 21374
rect 2156 21310 2158 21362
rect 2210 21310 2212 21362
rect 2156 21028 2212 21310
rect 2156 20962 2212 20972
rect 2268 20914 2324 21644
rect 2268 20862 2270 20914
rect 2322 20862 2324 20914
rect 2268 20850 2324 20862
rect 1260 20018 1428 20020
rect 1260 19966 1262 20018
rect 1314 19966 1428 20018
rect 1260 19964 1428 19966
rect 1484 20076 1764 20132
rect 1820 20132 2100 20188
rect 2156 20804 2212 20814
rect 1260 19954 1316 19964
rect 1036 19906 1092 19918
rect 1036 19854 1038 19906
rect 1090 19854 1092 19906
rect 1036 17890 1092 19854
rect 1484 18450 1540 20076
rect 1708 19908 1764 19918
rect 1596 19796 1652 19806
rect 1708 19796 1764 19852
rect 1596 19794 1764 19796
rect 1596 19742 1598 19794
rect 1650 19742 1764 19794
rect 1596 19740 1764 19742
rect 1596 19730 1652 19740
rect 1596 19460 1652 19470
rect 1596 19366 1652 19404
rect 1484 18398 1486 18450
rect 1538 18398 1540 18450
rect 1484 18386 1540 18398
rect 1036 17838 1038 17890
rect 1090 17838 1092 17890
rect 1036 16994 1092 17838
rect 1708 18226 1764 18238
rect 1708 18174 1710 18226
rect 1762 18174 1764 18226
rect 1596 17554 1652 17566
rect 1596 17502 1598 17554
rect 1650 17502 1652 17554
rect 1596 17108 1652 17502
rect 1596 17042 1652 17052
rect 1036 16942 1038 16994
rect 1090 16942 1092 16994
rect 1036 16930 1092 16942
rect 1484 16882 1540 16894
rect 1484 16830 1486 16882
rect 1538 16830 1540 16882
rect 1148 13860 1204 13870
rect 1148 13766 1204 13804
rect 924 12226 980 12236
rect 1148 13188 1204 13198
rect 1148 12178 1204 13132
rect 1148 12126 1150 12178
rect 1202 12126 1204 12178
rect 1148 12114 1204 12126
rect 1260 11170 1316 11182
rect 1260 11118 1262 11170
rect 1314 11118 1316 11170
rect 1260 10612 1316 11118
rect 1260 10546 1316 10556
rect 1260 9602 1316 9614
rect 1260 9550 1262 9602
rect 1314 9550 1316 9602
rect 1260 9268 1316 9550
rect 1260 9202 1316 9212
rect 1484 8428 1540 16830
rect 1596 15092 1652 15102
rect 1596 13746 1652 15036
rect 1596 13694 1598 13746
rect 1650 13694 1652 13746
rect 1596 13682 1652 13694
rect 1708 12964 1764 18174
rect 1820 15316 1876 20132
rect 2044 17892 2100 17902
rect 2044 17666 2100 17836
rect 2156 17780 2212 20748
rect 2380 20244 2436 22316
rect 2380 20178 2436 20188
rect 2492 23042 2884 23044
rect 2492 22990 2718 23042
rect 2770 22990 2884 23042
rect 2492 22988 2884 22990
rect 2268 18788 2324 18798
rect 2268 18450 2324 18732
rect 2492 18676 2548 22988
rect 2716 22978 2772 22988
rect 2716 22596 2772 22606
rect 2716 22502 2772 22540
rect 2716 21586 2772 21598
rect 2716 21534 2718 21586
rect 2770 21534 2772 21586
rect 2604 20802 2660 20814
rect 2604 20750 2606 20802
rect 2658 20750 2660 20802
rect 2604 19460 2660 20750
rect 2716 19572 2772 21534
rect 2940 20804 2996 26852
rect 3276 26066 3332 26078
rect 3276 26014 3278 26066
rect 3330 26014 3332 26066
rect 3276 25844 3332 26014
rect 3276 25778 3332 25788
rect 3052 25732 3108 25742
rect 3052 25638 3108 25676
rect 3388 25060 3444 28028
rect 3500 26516 3556 28252
rect 3500 26450 3556 26460
rect 3612 26740 3668 28700
rect 3836 28690 3892 28700
rect 4060 28420 4116 29484
rect 4172 28868 4228 33516
rect 4284 32452 4340 32462
rect 4284 32358 4340 32396
rect 4464 32172 4728 32182
rect 4520 32116 4568 32172
rect 4624 32116 4672 32172
rect 4464 32106 4728 32116
rect 4284 31780 4340 31790
rect 4284 30772 4340 31724
rect 4844 31778 4900 31790
rect 4844 31726 4846 31778
rect 4898 31726 4900 31778
rect 4844 31668 4900 31726
rect 4844 31602 4900 31612
rect 4396 31556 4452 31566
rect 4396 31220 4452 31500
rect 4396 31106 4452 31164
rect 4396 31054 4398 31106
rect 4450 31054 4452 31106
rect 4396 31042 4452 31054
rect 4284 30706 4340 30716
rect 4844 30772 4900 30782
rect 4464 30604 4728 30614
rect 4520 30548 4568 30604
rect 4624 30548 4672 30604
rect 4464 30538 4728 30548
rect 4464 29036 4728 29046
rect 4520 28980 4568 29036
rect 4624 28980 4672 29036
rect 4464 28970 4728 28980
rect 4172 28812 4452 28868
rect 4060 28364 4228 28420
rect 3804 28252 4068 28262
rect 3860 28196 3908 28252
rect 3964 28196 4012 28252
rect 3804 28186 4068 28196
rect 3500 25844 3556 25854
rect 3500 25618 3556 25788
rect 3500 25566 3502 25618
rect 3554 25566 3556 25618
rect 3500 25554 3556 25566
rect 3052 25004 3444 25060
rect 3500 25284 3556 25294
rect 3052 23716 3108 25004
rect 3500 24724 3556 25228
rect 3052 23650 3108 23660
rect 3164 24722 3556 24724
rect 3164 24670 3502 24722
rect 3554 24670 3556 24722
rect 3164 24668 3556 24670
rect 3052 22596 3108 22606
rect 3052 21476 3108 22540
rect 3164 21588 3220 24668
rect 3500 24658 3556 24668
rect 3388 24500 3444 24510
rect 3276 24498 3444 24500
rect 3276 24446 3390 24498
rect 3442 24446 3444 24498
rect 3276 24444 3444 24446
rect 3276 23156 3332 24444
rect 3388 24434 3444 24444
rect 3612 24052 3668 26684
rect 3804 26684 4068 26694
rect 3860 26628 3908 26684
rect 3964 26628 4012 26684
rect 3804 26618 4068 26628
rect 3836 26516 3892 26526
rect 3724 26066 3780 26078
rect 3724 26014 3726 26066
rect 3778 26014 3780 26066
rect 3724 25732 3780 26014
rect 3724 25666 3780 25676
rect 3836 25508 3892 26460
rect 4172 26402 4228 28364
rect 4284 27860 4340 27870
rect 4284 27766 4340 27804
rect 4396 27636 4452 28812
rect 4844 28532 4900 30716
rect 4956 28644 5012 35420
rect 5068 34802 5124 34814
rect 5068 34750 5070 34802
rect 5122 34750 5124 34802
rect 5068 31892 5124 34750
rect 5180 34244 5236 34254
rect 5180 34130 5236 34188
rect 5180 34078 5182 34130
rect 5234 34078 5236 34130
rect 5180 33684 5236 34078
rect 5180 33618 5236 33628
rect 5068 31826 5124 31836
rect 5180 33236 5236 33246
rect 5068 30098 5124 30110
rect 5068 30046 5070 30098
rect 5122 30046 5124 30098
rect 5068 29876 5124 30046
rect 5068 29810 5124 29820
rect 5180 29652 5236 33180
rect 5292 31668 5348 36204
rect 5404 35588 5460 36316
rect 5404 35522 5460 35532
rect 5404 34916 5460 34926
rect 5404 34822 5460 34860
rect 5292 31602 5348 31612
rect 5404 34132 5460 34142
rect 5404 30436 5460 34076
rect 5404 30370 5460 30380
rect 5404 30212 5460 30222
rect 5180 29538 5236 29596
rect 5180 29486 5182 29538
rect 5234 29486 5236 29538
rect 5180 29474 5236 29486
rect 5292 30210 5460 30212
rect 5292 30158 5406 30210
rect 5458 30158 5460 30210
rect 5292 30156 5460 30158
rect 5292 29204 5348 30156
rect 5404 30146 5460 30156
rect 5516 29652 5572 38612
rect 5628 37044 5684 37054
rect 5628 36950 5684 36988
rect 5740 35476 5796 49532
rect 5964 39732 6020 51884
rect 6076 48244 6132 48254
rect 6076 41412 6132 48188
rect 6076 41318 6132 41356
rect 6300 40852 6356 53004
rect 6412 41076 6468 55412
rect 6524 55186 6580 57148
rect 7420 56194 7476 57344
rect 8764 56644 8820 57344
rect 10108 56756 10164 57344
rect 10108 56700 10612 56756
rect 8764 56588 9044 56644
rect 8988 56306 9044 56588
rect 8988 56254 8990 56306
rect 9042 56254 9044 56306
rect 8988 56242 9044 56254
rect 10556 56306 10612 56700
rect 10556 56254 10558 56306
rect 10610 56254 10612 56306
rect 10556 56242 10612 56254
rect 7420 56142 7422 56194
rect 7474 56142 7476 56194
rect 7420 56130 7476 56142
rect 8092 55972 8148 55982
rect 8092 55878 8148 55916
rect 9996 55970 10052 55982
rect 9996 55918 9998 55970
rect 10050 55918 10052 55970
rect 6524 55134 6526 55186
rect 6578 55134 6580 55186
rect 6524 55122 6580 55134
rect 7532 55298 7588 55310
rect 7532 55246 7534 55298
rect 7586 55246 7588 55298
rect 6636 51492 6692 51502
rect 6636 41298 6692 51436
rect 7420 49588 7476 49598
rect 6636 41246 6638 41298
rect 6690 41246 6692 41298
rect 6636 41234 6692 41246
rect 7196 49028 7252 49038
rect 6412 41020 6692 41076
rect 6300 40796 6580 40852
rect 6412 40180 6468 40190
rect 6076 40178 6468 40180
rect 6076 40126 6414 40178
rect 6466 40126 6468 40178
rect 6076 40124 6468 40126
rect 6076 39842 6132 40124
rect 6412 40114 6468 40124
rect 6524 39956 6580 40796
rect 6076 39790 6078 39842
rect 6130 39790 6132 39842
rect 6076 39778 6132 39790
rect 6412 39900 6580 39956
rect 5964 39666 6020 39676
rect 5852 39618 5908 39630
rect 5852 39566 5854 39618
rect 5906 39566 5908 39618
rect 5852 36036 5908 39566
rect 6188 38948 6244 38958
rect 5964 38724 6020 38762
rect 5964 38658 6020 38668
rect 6188 38276 6244 38892
rect 6300 38276 6356 38286
rect 6188 38274 6356 38276
rect 6188 38222 6302 38274
rect 6354 38222 6356 38274
rect 6188 38220 6356 38222
rect 6300 38210 6356 38220
rect 6188 36482 6244 36494
rect 6188 36430 6190 36482
rect 6242 36430 6244 36482
rect 5852 35980 6020 36036
rect 5852 35812 5908 35822
rect 5852 35718 5908 35756
rect 5628 33908 5684 33918
rect 5740 33908 5796 35420
rect 5628 33906 5796 33908
rect 5628 33854 5630 33906
rect 5682 33854 5796 33906
rect 5628 33852 5796 33854
rect 5628 33842 5684 33852
rect 5628 33236 5684 33246
rect 5628 33142 5684 33180
rect 5628 30436 5684 30446
rect 5628 29764 5684 30380
rect 5740 29988 5796 33852
rect 5852 35588 5908 35598
rect 5852 30436 5908 35532
rect 5964 34914 6020 35980
rect 6076 35140 6132 35150
rect 6188 35140 6244 36430
rect 6300 35476 6356 35486
rect 6300 35382 6356 35420
rect 6076 35138 6244 35140
rect 6076 35086 6078 35138
rect 6130 35086 6244 35138
rect 6076 35084 6244 35086
rect 6076 35074 6132 35084
rect 5964 34862 5966 34914
rect 6018 34862 6020 34914
rect 5964 34468 6020 34862
rect 5964 34402 6020 34412
rect 6076 34804 6132 34814
rect 6076 33572 6132 34748
rect 6076 33478 6132 33516
rect 6300 32450 6356 32462
rect 6300 32398 6302 32450
rect 6354 32398 6356 32450
rect 6300 31892 6356 32398
rect 5852 30370 5908 30380
rect 5964 31668 6020 31678
rect 5852 30212 5908 30222
rect 5964 30212 6020 31612
rect 6188 30770 6244 30782
rect 6188 30718 6190 30770
rect 6242 30718 6244 30770
rect 6076 30436 6132 30446
rect 6188 30436 6244 30718
rect 6300 30660 6356 31836
rect 6300 30594 6356 30604
rect 6076 30434 6244 30436
rect 6076 30382 6078 30434
rect 6130 30382 6244 30434
rect 6076 30380 6244 30382
rect 6076 30370 6132 30380
rect 5964 30156 6132 30212
rect 5852 30118 5908 30156
rect 5740 29932 5908 29988
rect 5628 29708 5796 29764
rect 5516 29596 5684 29652
rect 5516 29316 5572 29326
rect 5068 29148 5348 29204
rect 5404 29314 5572 29316
rect 5404 29262 5518 29314
rect 5570 29262 5572 29314
rect 5404 29260 5572 29262
rect 5068 28866 5124 29148
rect 5068 28814 5070 28866
rect 5122 28814 5124 28866
rect 5068 28802 5124 28814
rect 4956 28588 5236 28644
rect 4844 28476 5012 28532
rect 4956 28084 5012 28476
rect 4172 26350 4174 26402
rect 4226 26350 4228 26402
rect 4172 26338 4228 26350
rect 4284 27580 4452 27636
rect 4844 27972 4900 27982
rect 3836 25442 3892 25452
rect 4284 25506 4340 27580
rect 4464 27468 4728 27478
rect 4520 27412 4568 27468
rect 4624 27412 4672 27468
rect 4464 27402 4728 27412
rect 4844 27074 4900 27916
rect 4956 27970 5012 28028
rect 4956 27918 4958 27970
rect 5010 27918 5012 27970
rect 4956 27906 5012 27918
rect 5068 28420 5124 28430
rect 4844 27022 4846 27074
rect 4898 27022 4900 27074
rect 4844 27010 4900 27022
rect 4464 25900 4728 25910
rect 4520 25844 4568 25900
rect 4624 25844 4672 25900
rect 4464 25834 4728 25844
rect 4284 25454 4286 25506
rect 4338 25454 4340 25506
rect 3804 25116 4068 25126
rect 3860 25060 3908 25116
rect 3964 25060 4012 25116
rect 3804 25050 4068 25060
rect 4060 24724 4116 24734
rect 4060 24722 4228 24724
rect 4060 24670 4062 24722
rect 4114 24670 4228 24722
rect 4060 24668 4228 24670
rect 4060 24658 4116 24668
rect 3276 23090 3332 23100
rect 3388 24050 3668 24052
rect 3388 23998 3614 24050
rect 3666 23998 3668 24050
rect 3388 23996 3668 23998
rect 3164 21532 3332 21588
rect 3052 21474 3220 21476
rect 3052 21422 3054 21474
rect 3106 21422 3220 21474
rect 3052 21420 3220 21422
rect 3052 21410 3108 21420
rect 2940 20738 2996 20748
rect 3052 21252 3108 21262
rect 3052 20802 3108 21196
rect 3052 20750 3054 20802
rect 3106 20750 3108 20802
rect 3052 20738 3108 20750
rect 2828 20244 2884 20282
rect 2828 20178 2884 20188
rect 3164 20188 3220 21420
rect 3276 21252 3332 21532
rect 3276 21186 3332 21196
rect 3276 21028 3332 21038
rect 3276 20934 3332 20972
rect 3164 20132 3332 20188
rect 2716 19516 2884 19572
rect 2604 19394 2660 19404
rect 2716 19348 2772 19358
rect 2716 19254 2772 19292
rect 2716 18788 2772 18798
rect 2492 18620 2660 18676
rect 2268 18398 2270 18450
rect 2322 18398 2324 18450
rect 2268 18386 2324 18398
rect 2492 18452 2548 18462
rect 2156 17714 2212 17724
rect 2044 17614 2046 17666
rect 2098 17614 2100 17666
rect 2044 17602 2100 17614
rect 2492 16994 2548 18396
rect 2604 18004 2660 18620
rect 2716 18450 2772 18732
rect 2716 18398 2718 18450
rect 2770 18398 2772 18450
rect 2716 18386 2772 18398
rect 2604 17948 2772 18004
rect 2604 17780 2660 17790
rect 2604 17556 2660 17724
rect 2604 17490 2660 17500
rect 2492 16942 2494 16994
rect 2546 16942 2548 16994
rect 2492 16930 2548 16942
rect 1932 16658 1988 16670
rect 1932 16606 1934 16658
rect 1986 16606 1988 16658
rect 1932 16212 1988 16606
rect 1932 16146 1988 16156
rect 1932 15876 1988 15886
rect 1932 15874 2660 15876
rect 1932 15822 1934 15874
rect 1986 15822 2660 15874
rect 1932 15820 2660 15822
rect 1932 15810 1988 15820
rect 1820 15260 2100 15316
rect 1932 15092 1988 15130
rect 1932 15026 1988 15036
rect 1932 14868 1988 14878
rect 1932 14754 1988 14812
rect 1932 14702 1934 14754
rect 1986 14702 1988 14754
rect 1932 14690 1988 14702
rect 1932 13746 1988 13758
rect 1932 13694 1934 13746
rect 1986 13694 1988 13746
rect 1932 13524 1988 13694
rect 1932 13458 1988 13468
rect 2044 13300 2100 15260
rect 2492 14418 2548 14430
rect 2492 14366 2494 14418
rect 2546 14366 2548 14418
rect 2492 13972 2548 14366
rect 2492 13906 2548 13916
rect 2604 13746 2660 15820
rect 2604 13694 2606 13746
rect 2658 13694 2660 13746
rect 2604 13682 2660 13694
rect 2156 13524 2212 13534
rect 2156 13522 2548 13524
rect 2156 13470 2158 13522
rect 2210 13470 2548 13522
rect 2156 13468 2548 13470
rect 2156 13458 2212 13468
rect 1708 12898 1764 12908
rect 1932 13244 2100 13300
rect 1596 12292 1652 12302
rect 1596 12198 1652 12236
rect 1932 11956 1988 13244
rect 2044 13076 2100 13086
rect 2044 12178 2100 13020
rect 2156 12964 2212 12974
rect 2156 12870 2212 12908
rect 2492 12740 2548 13468
rect 2604 13188 2660 13198
rect 2716 13188 2772 17948
rect 2828 17892 2884 19516
rect 2828 17826 2884 17836
rect 2940 19460 2996 19470
rect 2828 14756 2884 14766
rect 2828 14662 2884 14700
rect 2940 14532 2996 19404
rect 3052 19348 3108 19358
rect 3052 16322 3108 19292
rect 3164 19122 3220 19134
rect 3164 19070 3166 19122
rect 3218 19070 3220 19122
rect 3164 18788 3220 19070
rect 3164 18722 3220 18732
rect 3164 18564 3220 18574
rect 3164 18470 3220 18508
rect 3052 16270 3054 16322
rect 3106 16270 3108 16322
rect 3052 15204 3108 16270
rect 3052 14868 3108 15148
rect 3164 16212 3220 16222
rect 3276 16212 3332 20132
rect 3220 16156 3332 16212
rect 3164 15202 3220 16156
rect 3164 15150 3166 15202
rect 3218 15150 3220 15202
rect 3164 15138 3220 15150
rect 3052 14802 3108 14812
rect 3388 14868 3444 23996
rect 3612 23986 3668 23996
rect 4060 23826 4116 23838
rect 4060 23774 4062 23826
rect 4114 23774 4116 23826
rect 4060 23716 4116 23774
rect 4060 23650 4116 23660
rect 3804 23548 4068 23558
rect 3860 23492 3908 23548
rect 3964 23492 4012 23548
rect 3804 23482 4068 23492
rect 3836 23380 3892 23390
rect 4172 23380 4228 24668
rect 4284 24612 4340 25454
rect 5068 25506 5124 28364
rect 5068 25454 5070 25506
rect 5122 25454 5124 25506
rect 4396 24612 4452 24622
rect 4284 24610 4452 24612
rect 4284 24558 4398 24610
rect 4450 24558 4452 24610
rect 4284 24556 4452 24558
rect 4396 24500 4452 24556
rect 4396 24444 4900 24500
rect 4464 24332 4728 24342
rect 4520 24276 4568 24332
rect 4624 24276 4672 24332
rect 4464 24266 4728 24276
rect 4844 23940 4900 24444
rect 5068 24164 5124 25454
rect 4844 23874 4900 23884
rect 4956 24108 5124 24164
rect 4620 23828 4676 23838
rect 3836 23378 4228 23380
rect 3836 23326 3838 23378
rect 3890 23326 4228 23378
rect 3836 23324 4228 23326
rect 4284 23716 4340 23726
rect 3836 23314 3892 23324
rect 4284 23268 4340 23660
rect 4172 23212 4340 23268
rect 3836 22148 3892 22158
rect 3612 22146 3892 22148
rect 3612 22094 3838 22146
rect 3890 22094 3892 22146
rect 3612 22092 3892 22094
rect 3612 20916 3668 22092
rect 3836 22082 3892 22092
rect 3804 21980 4068 21990
rect 3860 21924 3908 21980
rect 3964 21924 4012 21980
rect 3804 21914 4068 21924
rect 3724 20916 3780 20926
rect 3612 20914 3780 20916
rect 3612 20862 3726 20914
rect 3778 20862 3780 20914
rect 3612 20860 3780 20862
rect 3724 20850 3780 20860
rect 3804 20412 4068 20422
rect 3860 20356 3908 20412
rect 3964 20356 4012 20412
rect 3804 20346 4068 20356
rect 3612 20018 3668 20030
rect 3612 19966 3614 20018
rect 3666 19966 3668 20018
rect 3500 19908 3556 19918
rect 3500 16100 3556 19852
rect 3612 18788 3668 19966
rect 4172 19908 4228 23212
rect 4620 22932 4676 23772
rect 4956 23716 5012 24108
rect 5068 23940 5124 23950
rect 5180 23940 5236 28588
rect 5292 27860 5348 27870
rect 5292 27766 5348 27804
rect 5404 27636 5460 29260
rect 5516 29250 5572 29260
rect 5516 29092 5572 29102
rect 5516 28754 5572 29036
rect 5516 28702 5518 28754
rect 5570 28702 5572 28754
rect 5516 28690 5572 28702
rect 5292 27580 5460 27636
rect 5292 25396 5348 27580
rect 5628 27524 5684 29596
rect 5740 28420 5796 29708
rect 5740 28354 5796 28364
rect 5740 27860 5796 27870
rect 5740 27766 5796 27804
rect 5404 27468 5684 27524
rect 5404 27298 5460 27468
rect 5404 27246 5406 27298
rect 5458 27246 5460 27298
rect 5404 27234 5460 27246
rect 5516 27300 5572 27310
rect 5292 25330 5348 25340
rect 5068 23938 5236 23940
rect 5068 23886 5070 23938
rect 5122 23886 5236 23938
rect 5068 23884 5236 23886
rect 5404 23940 5460 23950
rect 5068 23874 5124 23884
rect 4956 23660 5236 23716
rect 5068 23380 5124 23390
rect 4620 22876 4900 22932
rect 4464 22764 4728 22774
rect 4520 22708 4568 22764
rect 4624 22708 4672 22764
rect 4464 22698 4728 22708
rect 4284 22372 4340 22382
rect 4284 21810 4340 22316
rect 4844 22260 4900 22876
rect 4956 22260 5012 22270
rect 4844 22258 5012 22260
rect 4844 22206 4958 22258
rect 5010 22206 5012 22258
rect 4844 22204 5012 22206
rect 4284 21758 4286 21810
rect 4338 21758 4340 21810
rect 4284 21746 4340 21758
rect 4956 21252 5012 22204
rect 4464 21196 4728 21206
rect 4520 21140 4568 21196
rect 4624 21140 4672 21196
rect 4956 21186 5012 21196
rect 4464 21130 4728 21140
rect 4508 20802 4564 20814
rect 4508 20750 4510 20802
rect 4562 20750 4564 20802
rect 4508 20468 4564 20750
rect 4508 20402 4564 20412
rect 4172 19842 4228 19852
rect 4956 20020 5012 20030
rect 4464 19628 4728 19638
rect 4520 19572 4568 19628
rect 4624 19572 4672 19628
rect 4464 19562 4728 19572
rect 4508 19348 4564 19358
rect 4508 19254 4564 19292
rect 4172 19124 4228 19134
rect 4172 19122 4452 19124
rect 4172 19070 4174 19122
rect 4226 19070 4452 19122
rect 4172 19068 4452 19070
rect 4172 19058 4228 19068
rect 3804 18844 4068 18854
rect 3860 18788 3908 18844
rect 3964 18788 4012 18844
rect 3804 18778 4068 18788
rect 4284 18788 4340 18798
rect 3612 17332 3668 18732
rect 4284 18562 4340 18732
rect 4284 18510 4286 18562
rect 4338 18510 4340 18562
rect 4284 18498 4340 18510
rect 3948 18450 4004 18462
rect 3948 18398 3950 18450
rect 4002 18398 4004 18450
rect 3948 18340 4004 18398
rect 4396 18340 4452 19068
rect 4956 18788 5012 19964
rect 4956 18722 5012 18732
rect 3948 17780 4004 18284
rect 4284 18284 4452 18340
rect 4284 17892 4340 18284
rect 4464 18060 4728 18070
rect 4520 18004 4568 18060
rect 4624 18004 4672 18060
rect 4464 17994 4728 18004
rect 3948 17724 4228 17780
rect 3724 17668 3780 17678
rect 3724 17574 3780 17612
rect 3612 17266 3668 17276
rect 3804 17276 4068 17286
rect 3860 17220 3908 17276
rect 3964 17220 4012 17276
rect 3804 17210 4068 17220
rect 3836 16884 3892 16894
rect 3836 16790 3892 16828
rect 4172 16324 4228 17724
rect 4284 17666 4340 17836
rect 4844 17892 4900 17930
rect 4844 17826 4900 17836
rect 4284 17614 4286 17666
rect 4338 17614 4340 17666
rect 4284 17602 4340 17614
rect 4844 17668 4900 17678
rect 4396 17556 4452 17566
rect 4396 17554 4564 17556
rect 4396 17502 4398 17554
rect 4450 17502 4564 17554
rect 4396 17500 4564 17502
rect 4396 17490 4452 17500
rect 4508 17332 4564 17500
rect 4508 17266 4564 17276
rect 4396 16660 4452 16698
rect 4396 16594 4452 16604
rect 4464 16492 4728 16502
rect 4520 16436 4568 16492
rect 4624 16436 4672 16492
rect 4464 16426 4728 16436
rect 4732 16324 4788 16334
rect 4172 16268 4452 16324
rect 3612 16100 3668 16110
rect 4172 16100 4228 16110
rect 3500 16098 4228 16100
rect 3500 16046 3614 16098
rect 3666 16046 4174 16098
rect 4226 16046 4228 16098
rect 3500 16044 4228 16046
rect 3612 16034 3668 16044
rect 4172 16034 4228 16044
rect 3388 14802 3444 14812
rect 3500 15764 3556 15774
rect 3500 15426 3556 15708
rect 3804 15708 4068 15718
rect 3500 15374 3502 15426
rect 3554 15374 3556 15426
rect 3388 14644 3444 14654
rect 2940 14476 3220 14532
rect 2660 13132 2772 13188
rect 2940 14308 2996 14318
rect 2604 13094 2660 13132
rect 2492 12684 2884 12740
rect 2044 12126 2046 12178
rect 2098 12126 2100 12178
rect 2044 12114 2100 12126
rect 2156 12404 2212 12414
rect 1932 11890 1988 11900
rect 2156 9826 2212 12348
rect 2492 12292 2548 12302
rect 2492 12198 2548 12236
rect 2828 12178 2884 12684
rect 2828 12126 2830 12178
rect 2882 12126 2884 12178
rect 2828 12114 2884 12126
rect 2380 11956 2436 11966
rect 2268 11620 2324 11630
rect 2268 11506 2324 11564
rect 2268 11454 2270 11506
rect 2322 11454 2324 11506
rect 2268 11442 2324 11454
rect 2156 9774 2158 9826
rect 2210 9774 2212 9826
rect 2156 9762 2212 9774
rect 2380 8428 2436 11900
rect 2604 11508 2660 11518
rect 2604 11414 2660 11452
rect 2940 8428 2996 14252
rect 3164 14196 3220 14476
rect 3276 14420 3332 14430
rect 3276 14326 3332 14364
rect 3164 14140 3332 14196
rect 1372 8372 1540 8428
rect 2268 8372 2436 8428
rect 2716 8372 2996 8428
rect 3052 13524 3108 13534
rect 1260 6580 1316 6590
rect 1260 6486 1316 6524
rect 1260 6018 1316 6030
rect 1260 5966 1262 6018
rect 1314 5966 1316 6018
rect 1260 5236 1316 5966
rect 1260 5170 1316 5180
rect 1372 2436 1428 8372
rect 2268 6802 2324 8372
rect 2268 6750 2270 6802
rect 2322 6750 2324 6802
rect 2268 6738 2324 6750
rect 2268 5908 2324 5918
rect 2716 5908 2772 8372
rect 2268 5906 2772 5908
rect 2268 5854 2270 5906
rect 2322 5854 2772 5906
rect 2268 5852 2772 5854
rect 2268 5842 2324 5852
rect 3052 3892 3108 13468
rect 3164 12740 3220 12750
rect 3164 11506 3220 12684
rect 3276 12290 3332 14140
rect 3388 13746 3444 14588
rect 3388 13694 3390 13746
rect 3442 13694 3444 13746
rect 3388 12852 3444 13694
rect 3388 12786 3444 12796
rect 3276 12238 3278 12290
rect 3330 12238 3332 12290
rect 3276 12226 3332 12238
rect 3164 11454 3166 11506
rect 3218 11454 3220 11506
rect 3164 11442 3220 11454
rect 3500 11396 3556 15374
rect 3500 11330 3556 11340
rect 3612 15652 3668 15662
rect 3860 15652 3908 15708
rect 3964 15652 4012 15708
rect 3804 15642 4068 15652
rect 3052 3826 3108 3836
rect 1372 2370 1428 2380
rect 3388 2436 3444 2446
rect 700 1652 756 1662
rect 700 112 756 1596
rect 2044 1428 2100 1438
rect 2044 112 2100 1372
rect 3388 112 3444 2380
rect 3612 196 3668 15596
rect 4396 15092 4452 16268
rect 4732 16230 4788 16268
rect 4396 15026 4452 15036
rect 4464 14924 4728 14934
rect 4520 14868 4568 14924
rect 4624 14868 4672 14924
rect 4464 14858 4728 14868
rect 4508 14644 4564 14654
rect 4508 14550 4564 14588
rect 4844 14530 4900 17612
rect 4956 16884 5012 16894
rect 4956 16790 5012 16828
rect 4956 15764 5012 15774
rect 4956 14644 5012 15708
rect 4956 14578 5012 14588
rect 4844 14478 4846 14530
rect 4898 14478 4900 14530
rect 4844 14466 4900 14478
rect 3804 14140 4068 14150
rect 3860 14084 3908 14140
rect 3964 14084 4012 14140
rect 3804 14074 4068 14084
rect 4956 13860 5012 13870
rect 4284 13746 4340 13758
rect 4284 13694 4286 13746
rect 4338 13694 4340 13746
rect 4284 13300 4340 13694
rect 4464 13356 4728 13366
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4464 13290 4728 13300
rect 4284 13234 4340 13244
rect 3724 13076 3780 13086
rect 3724 13074 4340 13076
rect 3724 13022 3726 13074
rect 3778 13022 4340 13074
rect 3724 13020 4340 13022
rect 3724 13010 3780 13020
rect 4284 12964 4340 13020
rect 4508 12964 4564 12974
rect 4284 12962 4564 12964
rect 4284 12910 4510 12962
rect 4562 12910 4564 12962
rect 4284 12908 4564 12910
rect 4508 12898 4564 12908
rect 4956 12962 5012 13804
rect 5068 13636 5124 23324
rect 5180 20804 5236 23660
rect 5404 23604 5460 23884
rect 5292 23548 5460 23604
rect 5292 22596 5348 23548
rect 5516 23156 5572 27244
rect 5628 26908 5684 27468
rect 5852 27300 5908 29932
rect 5964 28642 6020 28654
rect 5964 28590 5966 28642
rect 6018 28590 6020 28642
rect 5964 27746 6020 28590
rect 5964 27694 5966 27746
rect 6018 27694 6020 27746
rect 5964 27682 6020 27694
rect 5852 27234 5908 27244
rect 5628 26852 5796 26908
rect 5628 24498 5684 24510
rect 5628 24446 5630 24498
rect 5682 24446 5684 24498
rect 5628 24162 5684 24446
rect 5628 24110 5630 24162
rect 5682 24110 5684 24162
rect 5628 24098 5684 24110
rect 5628 23604 5684 23614
rect 5628 23492 5684 23548
rect 5628 23426 5684 23436
rect 5292 22530 5348 22540
rect 5404 23100 5572 23156
rect 5740 23156 5796 26852
rect 5852 26628 5908 26638
rect 5852 23604 5908 26572
rect 6076 24050 6132 30156
rect 6300 26516 6356 26526
rect 6188 26292 6244 26302
rect 6188 24834 6244 26236
rect 6300 25506 6356 26460
rect 6300 25454 6302 25506
rect 6354 25454 6356 25506
rect 6300 25442 6356 25454
rect 6188 24782 6190 24834
rect 6242 24782 6244 24834
rect 6188 24770 6244 24782
rect 6076 23998 6078 24050
rect 6130 23998 6132 24050
rect 6076 23986 6132 23998
rect 6188 24164 6244 24174
rect 5852 23538 5908 23548
rect 6076 23604 6132 23614
rect 5852 23156 5908 23166
rect 5740 23100 5852 23156
rect 5292 22372 5348 22382
rect 5292 22278 5348 22316
rect 5292 20804 5348 20814
rect 5180 20802 5348 20804
rect 5180 20750 5294 20802
rect 5346 20750 5348 20802
rect 5180 20748 5348 20750
rect 5292 20738 5348 20748
rect 5292 20132 5348 20142
rect 5292 16996 5348 20076
rect 5404 17220 5460 23100
rect 5852 23090 5908 23100
rect 5628 23044 5684 23054
rect 5628 23042 5796 23044
rect 5628 22990 5630 23042
rect 5682 22990 5796 23042
rect 5628 22988 5796 22990
rect 5628 22978 5684 22988
rect 5740 22820 5796 22988
rect 5740 22764 6020 22820
rect 5852 22596 5908 22606
rect 5852 22370 5908 22540
rect 5964 22594 6020 22764
rect 5964 22542 5966 22594
rect 6018 22542 6020 22594
rect 5964 22530 6020 22542
rect 5852 22318 5854 22370
rect 5906 22318 5908 22370
rect 5516 22036 5572 22046
rect 5516 21698 5572 21980
rect 5516 21646 5518 21698
rect 5570 21646 5572 21698
rect 5516 21634 5572 21646
rect 5740 21700 5796 21710
rect 5740 21028 5796 21644
rect 5740 20962 5796 20972
rect 5628 20916 5684 20926
rect 5628 19794 5684 20860
rect 5628 19742 5630 19794
rect 5682 19742 5684 19794
rect 5628 19236 5684 19742
rect 5740 20804 5796 20814
rect 5740 19458 5796 20748
rect 5852 20468 5908 22318
rect 5964 21364 6020 21374
rect 5964 21270 6020 21308
rect 6076 21140 6132 23548
rect 6188 23266 6244 24108
rect 6412 23380 6468 39900
rect 6636 39844 6692 41020
rect 6524 39788 6692 39844
rect 6972 40290 7028 40302
rect 6972 40238 6974 40290
rect 7026 40238 7028 40290
rect 6972 39844 7028 40238
rect 6524 28196 6580 39788
rect 6972 39778 7028 39788
rect 6636 39620 6692 39630
rect 6636 36372 6692 39564
rect 6748 39618 6804 39630
rect 6748 39566 6750 39618
rect 6802 39566 6804 39618
rect 6748 39060 6804 39566
rect 6748 38994 6804 39004
rect 7084 39618 7140 39630
rect 7084 39566 7086 39618
rect 7138 39566 7140 39618
rect 6748 38050 6804 38062
rect 6748 37998 6750 38050
rect 6802 37998 6804 38050
rect 6748 37940 6804 37998
rect 6748 37874 6804 37884
rect 6748 37492 6804 37502
rect 6748 37398 6804 37436
rect 6636 36306 6692 36316
rect 6748 36370 6804 36382
rect 6748 36318 6750 36370
rect 6802 36318 6804 36370
rect 6748 35924 6804 36318
rect 6748 35858 6804 35868
rect 6860 36036 6916 36046
rect 6748 34914 6804 34926
rect 6748 34862 6750 34914
rect 6802 34862 6804 34914
rect 6748 34354 6804 34862
rect 6748 34302 6750 34354
rect 6802 34302 6804 34354
rect 6748 34290 6804 34302
rect 6748 32564 6804 32574
rect 6748 32470 6804 32508
rect 6636 31106 6692 31118
rect 6636 31054 6638 31106
rect 6690 31054 6692 31106
rect 6636 30884 6692 31054
rect 6636 30818 6692 30828
rect 6748 30210 6804 30222
rect 6748 30158 6750 30210
rect 6802 30158 6804 30210
rect 6748 29650 6804 30158
rect 6748 29598 6750 29650
rect 6802 29598 6804 29650
rect 6748 29586 6804 29598
rect 6748 28980 6804 28990
rect 6636 28532 6692 28542
rect 6636 28438 6692 28476
rect 6524 28140 6692 28196
rect 6524 27858 6580 27870
rect 6524 27806 6526 27858
rect 6578 27806 6580 27858
rect 6524 27298 6580 27806
rect 6524 27246 6526 27298
rect 6578 27246 6580 27298
rect 6524 27234 6580 27246
rect 6636 26908 6692 28140
rect 6412 23314 6468 23324
rect 6524 26852 6692 26908
rect 6748 26964 6804 28924
rect 6748 26898 6804 26908
rect 6188 23214 6190 23266
rect 6242 23214 6244 23266
rect 6188 23202 6244 23214
rect 6524 23156 6580 26852
rect 6636 25620 6692 25630
rect 6636 25526 6692 25564
rect 6748 25060 6804 25070
rect 6636 24276 6692 24286
rect 6636 23938 6692 24220
rect 6636 23886 6638 23938
rect 6690 23886 6692 23938
rect 6636 23380 6692 23886
rect 6636 23314 6692 23324
rect 6524 23090 6580 23100
rect 6748 23266 6804 25004
rect 6748 23214 6750 23266
rect 6802 23214 6804 23266
rect 6524 22932 6580 22942
rect 6412 22370 6468 22382
rect 6412 22318 6414 22370
rect 6466 22318 6468 22370
rect 6300 21474 6356 21486
rect 6300 21422 6302 21474
rect 6354 21422 6356 21474
rect 6076 21084 6244 21140
rect 6188 20692 6244 21084
rect 6300 21028 6356 21422
rect 6300 20962 6356 20972
rect 6412 20804 6468 22318
rect 6524 20916 6580 22876
rect 6748 21812 6804 23214
rect 6524 20850 6580 20860
rect 6636 21756 6804 21812
rect 6860 21812 6916 35980
rect 7084 35588 7140 39566
rect 7196 39284 7252 48972
rect 7308 40290 7364 40302
rect 7308 40238 7310 40290
rect 7362 40238 7364 40290
rect 7308 39618 7364 40238
rect 7308 39566 7310 39618
rect 7362 39566 7364 39618
rect 7308 39554 7364 39566
rect 7196 39228 7364 39284
rect 7196 39060 7252 39070
rect 7196 38966 7252 39004
rect 7308 38668 7364 39228
rect 7084 35522 7140 35532
rect 7196 38612 7364 38668
rect 7196 35140 7252 38612
rect 7308 38164 7364 38174
rect 7420 38164 7476 49532
rect 7308 38162 7476 38164
rect 7308 38110 7310 38162
rect 7362 38110 7476 38162
rect 7308 38108 7476 38110
rect 7308 38098 7364 38108
rect 7532 37828 7588 55246
rect 9996 54628 10052 55918
rect 11452 55188 11508 57344
rect 12796 56644 12852 57344
rect 14140 56756 14196 57344
rect 14140 56700 14644 56756
rect 12796 56588 13076 56644
rect 13020 56306 13076 56588
rect 13020 56254 13022 56306
rect 13074 56254 13076 56306
rect 13020 56242 13076 56254
rect 14588 56306 14644 56700
rect 14588 56254 14590 56306
rect 14642 56254 14644 56306
rect 14588 56242 14644 56254
rect 15484 56308 15540 57344
rect 16828 57204 16884 57344
rect 16828 57148 16996 57204
rect 15484 56242 15540 56252
rect 16492 56308 16548 56318
rect 16492 56214 16548 56252
rect 11564 55970 11620 55982
rect 11564 55918 11566 55970
rect 11618 55918 11620 55970
rect 11564 55412 11620 55918
rect 11564 55346 11620 55356
rect 14028 55970 14084 55982
rect 14028 55918 14030 55970
rect 14082 55918 14084 55970
rect 12908 55298 12964 55310
rect 12908 55246 12910 55298
rect 12962 55246 12964 55298
rect 11900 55188 11956 55198
rect 11452 55186 11956 55188
rect 11452 55134 11902 55186
rect 11954 55134 11956 55186
rect 11452 55132 11956 55134
rect 11900 55122 11956 55132
rect 12908 55076 12964 55246
rect 12908 55010 12964 55020
rect 9996 54562 10052 54572
rect 8652 54292 8708 54302
rect 8652 50428 8708 54236
rect 14028 53956 14084 55918
rect 15596 55970 15652 55982
rect 15596 55918 15598 55970
rect 15650 55918 15652 55970
rect 15596 55524 15652 55918
rect 15596 55458 15652 55468
rect 16940 55468 16996 57148
rect 18172 56308 18228 57344
rect 18508 56308 18564 56318
rect 18172 56306 18564 56308
rect 18172 56254 18510 56306
rect 18562 56254 18564 56306
rect 18172 56252 18564 56254
rect 18508 56242 18564 56252
rect 19516 56308 19572 57344
rect 19516 56242 19572 56252
rect 20636 56308 20692 56318
rect 20636 56214 20692 56252
rect 20860 56308 20916 57344
rect 22204 57204 22260 57344
rect 22204 57148 22708 57204
rect 20860 56242 20916 56252
rect 21868 56308 21924 56318
rect 21868 56214 21924 56252
rect 22540 56196 22596 56206
rect 20188 56082 20244 56094
rect 20188 56030 20190 56082
rect 20242 56030 20244 56082
rect 17500 55970 17556 55982
rect 17500 55918 17502 55970
rect 17554 55918 17556 55970
rect 16940 55412 17332 55468
rect 17276 55186 17332 55412
rect 17276 55134 17278 55186
rect 17330 55134 17332 55186
rect 17276 55122 17332 55134
rect 14028 53890 14084 53900
rect 14700 54404 14756 54414
rect 14252 53508 14308 53518
rect 12684 52500 12740 52510
rect 10108 52388 10164 52398
rect 8652 50372 9044 50428
rect 7980 44100 8036 44110
rect 7756 43428 7812 43438
rect 7644 40402 7700 40414
rect 7644 40350 7646 40402
rect 7698 40350 7700 40402
rect 7644 38948 7700 40350
rect 7644 38882 7700 38892
rect 7532 37762 7588 37772
rect 7644 38612 7700 38622
rect 7532 37156 7588 37166
rect 6972 35084 7252 35140
rect 7308 37100 7532 37156
rect 7644 37156 7700 38556
rect 7756 38162 7812 43372
rect 7756 38110 7758 38162
rect 7810 38110 7812 38162
rect 7756 38098 7812 38110
rect 7868 40516 7924 40526
rect 7756 37492 7812 37502
rect 7868 37492 7924 40460
rect 7980 37604 8036 44044
rect 8876 41186 8932 41198
rect 8876 41134 8878 41186
rect 8930 41134 8932 41186
rect 8876 40740 8932 41134
rect 8428 40684 8932 40740
rect 8092 40402 8148 40414
rect 8092 40350 8094 40402
rect 8146 40350 8148 40402
rect 8092 40180 8148 40350
rect 8092 37716 8148 40124
rect 8204 40292 8260 40302
rect 8204 39618 8260 40236
rect 8316 40292 8372 40302
rect 8428 40292 8484 40684
rect 8764 40404 8820 40414
rect 8764 40310 8820 40348
rect 8316 40290 8484 40292
rect 8316 40238 8318 40290
rect 8370 40238 8484 40290
rect 8316 40236 8484 40238
rect 8316 40226 8372 40236
rect 8988 40180 9044 50372
rect 8204 39566 8206 39618
rect 8258 39566 8260 39618
rect 8204 39554 8260 39566
rect 8652 40124 9044 40180
rect 9100 48804 9156 48814
rect 8652 38668 8708 40124
rect 8988 38836 9044 38846
rect 8652 38612 8820 38668
rect 8316 38052 8372 38062
rect 8316 38050 8596 38052
rect 8316 37998 8318 38050
rect 8370 37998 8596 38050
rect 8316 37996 8596 37998
rect 8316 37986 8372 37996
rect 8092 37660 8372 37716
rect 7980 37548 8148 37604
rect 7868 37436 8036 37492
rect 7756 37268 7812 37436
rect 7868 37268 7924 37278
rect 7756 37266 7924 37268
rect 7756 37214 7870 37266
rect 7922 37214 7924 37266
rect 7756 37212 7924 37214
rect 7868 37202 7924 37212
rect 7644 37100 7812 37156
rect 6972 28980 7028 35084
rect 7196 34914 7252 34926
rect 7196 34862 7198 34914
rect 7250 34862 7252 34914
rect 7084 34468 7140 34478
rect 7084 32562 7140 34412
rect 7196 33460 7252 34862
rect 7308 33796 7364 37100
rect 7532 37062 7588 37100
rect 7420 35812 7476 35822
rect 7420 35810 7700 35812
rect 7420 35758 7422 35810
rect 7474 35758 7700 35810
rect 7420 35756 7700 35758
rect 7420 35746 7476 35756
rect 7644 35700 7700 35756
rect 7644 35634 7700 35644
rect 7756 35476 7812 37100
rect 7868 36370 7924 36382
rect 7868 36318 7870 36370
rect 7922 36318 7924 36370
rect 7868 36148 7924 36318
rect 7868 36082 7924 36092
rect 7868 35588 7924 35598
rect 7868 35494 7924 35532
rect 7420 35420 7812 35476
rect 7420 33908 7476 35420
rect 7420 33842 7476 33852
rect 7532 33908 7588 33918
rect 7532 33906 7812 33908
rect 7532 33854 7534 33906
rect 7586 33854 7812 33906
rect 7532 33852 7812 33854
rect 7532 33842 7588 33852
rect 7308 33730 7364 33740
rect 7196 33394 7252 33404
rect 7644 33348 7700 33358
rect 7308 33346 7700 33348
rect 7308 33294 7646 33346
rect 7698 33294 7700 33346
rect 7308 33292 7700 33294
rect 7084 32510 7086 32562
rect 7138 32510 7140 32562
rect 7084 31556 7140 32510
rect 7196 33122 7252 33134
rect 7196 33070 7198 33122
rect 7250 33070 7252 33122
rect 7196 32564 7252 33070
rect 7196 32498 7252 32508
rect 7308 32450 7364 33292
rect 7644 33282 7700 33292
rect 7308 32398 7310 32450
rect 7362 32398 7364 32450
rect 7308 32386 7364 32398
rect 7420 32788 7476 32798
rect 7308 31780 7364 31790
rect 7308 31686 7364 31724
rect 7084 31500 7364 31556
rect 7196 31106 7252 31118
rect 7196 31054 7198 31106
rect 7250 31054 7252 31106
rect 7084 30548 7140 30558
rect 7084 30210 7140 30492
rect 7084 30158 7086 30210
rect 7138 30158 7140 30210
rect 7084 30146 7140 30158
rect 6972 28914 7028 28924
rect 6972 28754 7028 28766
rect 6972 28702 6974 28754
rect 7026 28702 7028 28754
rect 6972 28644 7028 28702
rect 6972 28578 7028 28588
rect 7196 28420 7252 31054
rect 6972 28364 7252 28420
rect 6972 23604 7028 28364
rect 6972 23538 7028 23548
rect 7084 27860 7140 27870
rect 6972 23380 7028 23390
rect 6972 22370 7028 23324
rect 6972 22318 6974 22370
rect 7026 22318 7028 22370
rect 6972 22306 7028 22318
rect 6412 20738 6468 20748
rect 6300 20692 6356 20702
rect 6188 20690 6356 20692
rect 6188 20638 6302 20690
rect 6354 20638 6356 20690
rect 6188 20636 6356 20638
rect 5852 20402 5908 20412
rect 6188 19906 6244 19918
rect 6188 19854 6190 19906
rect 6242 19854 6244 19906
rect 6188 19684 6244 19854
rect 6188 19618 6244 19628
rect 5740 19406 5742 19458
rect 5794 19406 5796 19458
rect 5740 19394 5796 19406
rect 5628 19180 5908 19236
rect 5404 17154 5460 17164
rect 5628 18900 5684 18910
rect 5628 18450 5684 18844
rect 5628 18398 5630 18450
rect 5682 18398 5684 18450
rect 5292 16940 5460 16996
rect 5404 16660 5460 16940
rect 5516 16660 5572 16670
rect 5404 16658 5572 16660
rect 5404 16606 5518 16658
rect 5570 16606 5572 16658
rect 5404 16604 5572 16606
rect 5516 16594 5572 16604
rect 5628 16660 5684 18398
rect 5628 16594 5684 16604
rect 5740 16884 5796 16894
rect 5292 15876 5348 15886
rect 5292 14530 5348 15820
rect 5740 15426 5796 16828
rect 5852 16660 5908 19180
rect 6300 18900 6356 20636
rect 6636 19236 6692 21756
rect 6860 21746 6916 21756
rect 6748 21588 6804 21598
rect 7084 21588 7140 27804
rect 7196 27858 7252 27870
rect 7196 27806 7198 27858
rect 7250 27806 7252 27858
rect 7196 24836 7252 27806
rect 7196 24770 7252 24780
rect 7196 22932 7252 22942
rect 7196 22838 7252 22876
rect 6748 21586 6916 21588
rect 6748 21534 6750 21586
rect 6802 21534 6916 21586
rect 6748 21532 6916 21534
rect 6748 21522 6804 21532
rect 6748 20916 6804 20926
rect 6748 20822 6804 20860
rect 6748 20132 6804 20142
rect 6748 20038 6804 20076
rect 6860 19572 6916 21532
rect 7084 21494 7140 21532
rect 7196 21812 7252 21822
rect 7196 20020 7252 21756
rect 7308 21588 7364 31500
rect 7420 21700 7476 32732
rect 7756 32562 7812 33852
rect 7756 32510 7758 32562
rect 7810 32510 7812 32562
rect 7756 32498 7812 32510
rect 7868 33796 7924 33806
rect 7868 32004 7924 33740
rect 7980 32788 8036 37436
rect 8092 36036 8148 37548
rect 8092 35970 8148 35980
rect 8204 37492 8260 37502
rect 8316 37492 8372 37660
rect 8316 37436 8484 37492
rect 8092 35364 8148 35374
rect 8092 34914 8148 35308
rect 8092 34862 8094 34914
rect 8146 34862 8148 34914
rect 8092 34850 8148 34862
rect 8204 33458 8260 37436
rect 8316 37268 8372 37278
rect 8316 37174 8372 37212
rect 8316 36482 8372 36494
rect 8316 36430 8318 36482
rect 8370 36430 8372 36482
rect 8316 36036 8372 36430
rect 8316 35970 8372 35980
rect 8316 35700 8372 35710
rect 8428 35700 8484 37436
rect 8540 37154 8596 37996
rect 8540 37102 8542 37154
rect 8594 37102 8596 37154
rect 8540 37090 8596 37102
rect 8652 35700 8708 35710
rect 8428 35698 8708 35700
rect 8428 35646 8654 35698
rect 8706 35646 8708 35698
rect 8428 35644 8708 35646
rect 8316 35606 8372 35644
rect 8652 35364 8708 35644
rect 8652 35298 8708 35308
rect 8652 33906 8708 33918
rect 8652 33854 8654 33906
rect 8706 33854 8708 33906
rect 8540 33684 8596 33694
rect 8204 33406 8206 33458
rect 8258 33406 8260 33458
rect 8204 33394 8260 33406
rect 8316 33460 8372 33470
rect 7980 32722 8036 32732
rect 8316 32564 8372 33404
rect 8428 32564 8484 32574
rect 8316 32562 8484 32564
rect 8316 32510 8430 32562
rect 8482 32510 8484 32562
rect 8316 32508 8484 32510
rect 7868 31948 8260 32004
rect 7644 31780 7700 31790
rect 7644 30770 7700 31724
rect 7644 30718 7646 30770
rect 7698 30718 7700 30770
rect 7644 30324 7700 30718
rect 7980 31666 8036 31678
rect 7980 31614 7982 31666
rect 8034 31614 8036 31666
rect 7980 30996 8036 31614
rect 7980 30324 8036 30940
rect 8092 31668 8148 31678
rect 8092 30994 8148 31612
rect 8092 30942 8094 30994
rect 8146 30942 8148 30994
rect 8092 30930 8148 30942
rect 7644 30268 7924 30324
rect 7756 30100 7812 30110
rect 7644 26516 7700 26526
rect 7644 26402 7700 26460
rect 7644 26350 7646 26402
rect 7698 26350 7700 26402
rect 7644 26338 7700 26350
rect 7532 24836 7588 24846
rect 7532 24388 7588 24780
rect 7532 24322 7588 24332
rect 7756 24164 7812 30044
rect 7868 26908 7924 30268
rect 7980 30258 8036 30268
rect 8204 30212 8260 31948
rect 8204 30118 8260 30156
rect 8316 30100 8372 32508
rect 8428 32498 8484 32508
rect 8540 31668 8596 33628
rect 8540 31602 8596 31612
rect 8652 33348 8708 33854
rect 8652 32340 8708 33292
rect 8652 30882 8708 32284
rect 8652 30830 8654 30882
rect 8706 30830 8708 30882
rect 8652 30818 8708 30830
rect 8316 30034 8372 30044
rect 8540 29428 8596 29438
rect 8540 29426 8708 29428
rect 8540 29374 8542 29426
rect 8594 29374 8708 29426
rect 8540 29372 8708 29374
rect 8540 29362 8596 29372
rect 8652 28532 8708 29372
rect 8204 28418 8260 28430
rect 8204 28366 8206 28418
rect 8258 28366 8260 28418
rect 8092 27858 8148 27870
rect 8092 27806 8094 27858
rect 8146 27806 8148 27858
rect 8092 27412 8148 27806
rect 8204 27860 8260 28366
rect 8204 27794 8260 27804
rect 8092 27356 8596 27412
rect 8316 27076 8372 27086
rect 7868 26852 8036 26908
rect 7868 25282 7924 25294
rect 7868 25230 7870 25282
rect 7922 25230 7924 25282
rect 7868 24722 7924 25230
rect 7868 24670 7870 24722
rect 7922 24670 7924 24722
rect 7868 24658 7924 24670
rect 7644 24108 7812 24164
rect 7644 21924 7700 24108
rect 7644 21858 7700 21868
rect 7756 23938 7812 23950
rect 7756 23886 7758 23938
rect 7810 23886 7812 23938
rect 7420 21644 7700 21700
rect 7308 21522 7364 21532
rect 7308 21364 7364 21374
rect 7308 21270 7364 21308
rect 7196 19954 7252 19964
rect 7196 19796 7252 19806
rect 7252 19740 7364 19796
rect 7196 19702 7252 19740
rect 6860 19516 7252 19572
rect 6636 19142 6692 19180
rect 6972 19346 7028 19358
rect 6972 19294 6974 19346
rect 7026 19294 7028 19346
rect 6300 18834 6356 18844
rect 5964 18340 6020 18350
rect 5964 18246 6020 18284
rect 6972 18340 7028 19294
rect 7196 18674 7252 19516
rect 7196 18622 7198 18674
rect 7250 18622 7252 18674
rect 7196 18610 7252 18622
rect 6972 17778 7028 18284
rect 7308 18228 7364 19740
rect 7644 19460 7700 21644
rect 7644 19394 7700 19404
rect 6972 17726 6974 17778
rect 7026 17726 7028 17778
rect 6972 17714 7028 17726
rect 7196 18172 7364 18228
rect 7420 19236 7476 19246
rect 6636 17668 6692 17678
rect 5852 16100 5908 16604
rect 5852 16034 5908 16044
rect 5964 17442 6020 17454
rect 5964 17390 5966 17442
rect 6018 17390 6020 17442
rect 5740 15374 5742 15426
rect 5794 15374 5796 15426
rect 5740 15362 5796 15374
rect 5852 15874 5908 15886
rect 5852 15822 5854 15874
rect 5906 15822 5908 15874
rect 5628 14756 5684 14766
rect 5292 14478 5294 14530
rect 5346 14478 5348 14530
rect 5292 13860 5348 14478
rect 5292 13794 5348 13804
rect 5516 14642 5572 14654
rect 5516 14590 5518 14642
rect 5570 14590 5572 14642
rect 5068 13570 5124 13580
rect 5180 13746 5236 13758
rect 5180 13694 5182 13746
rect 5234 13694 5236 13746
rect 5180 13412 5236 13694
rect 4956 12910 4958 12962
rect 5010 12910 5012 12962
rect 4956 12898 5012 12910
rect 5068 13356 5180 13412
rect 5068 12964 5124 13356
rect 5180 13346 5236 13356
rect 5292 13636 5348 13646
rect 5068 12898 5124 12908
rect 5180 13074 5236 13086
rect 5180 13022 5182 13074
rect 5234 13022 5236 13074
rect 4172 12852 4228 12862
rect 4172 12758 4228 12796
rect 3804 12572 4068 12582
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 3804 12506 4068 12516
rect 4464 11788 4728 11798
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4464 11722 4728 11732
rect 4844 11506 4900 11518
rect 4844 11454 4846 11506
rect 4898 11454 4900 11506
rect 4284 11396 4340 11406
rect 3804 11004 4068 11014
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 3804 10938 4068 10948
rect 4284 10500 4340 11340
rect 4844 11396 4900 11454
rect 4844 11330 4900 11340
rect 4284 10434 4340 10444
rect 4464 10220 4728 10230
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4464 10154 4728 10164
rect 4732 9940 4788 9950
rect 4732 9846 4788 9884
rect 5180 9826 5236 13022
rect 5292 12292 5348 13580
rect 5292 12226 5348 12236
rect 5516 12178 5572 14590
rect 5628 13634 5684 14700
rect 5852 13748 5908 15822
rect 5964 14642 6020 17390
rect 6188 17220 6244 17230
rect 6076 15204 6132 15242
rect 6076 15138 6132 15148
rect 6188 14980 6244 17164
rect 6636 17108 6692 17612
rect 6636 17042 6692 17052
rect 6972 17444 7028 17454
rect 6636 16884 6692 16894
rect 6524 16100 6580 16110
rect 6636 16100 6692 16828
rect 6860 16212 6916 16222
rect 6860 16118 6916 16156
rect 6524 16098 6692 16100
rect 6524 16046 6526 16098
rect 6578 16046 6692 16098
rect 6524 16044 6692 16046
rect 6524 16034 6580 16044
rect 5964 14590 5966 14642
rect 6018 14590 6020 14642
rect 5964 14578 6020 14590
rect 6076 14924 6244 14980
rect 5852 13682 5908 13692
rect 5628 13582 5630 13634
rect 5682 13582 5684 13634
rect 5628 13570 5684 13582
rect 5852 13524 5908 13534
rect 5852 12962 5908 13468
rect 5852 12910 5854 12962
rect 5906 12910 5908 12962
rect 5852 12898 5908 12910
rect 5964 12516 6020 12526
rect 5964 12290 6020 12460
rect 5964 12238 5966 12290
rect 6018 12238 6020 12290
rect 5964 12226 6020 12238
rect 5516 12126 5518 12178
rect 5570 12126 5572 12178
rect 5516 12114 5572 12126
rect 5404 11396 5460 11406
rect 5404 10610 5460 11340
rect 6076 11396 6132 14924
rect 6524 14532 6580 14542
rect 6412 14530 6580 14532
rect 6412 14478 6526 14530
rect 6578 14478 6580 14530
rect 6412 14476 6580 14478
rect 6412 13188 6468 14476
rect 6524 14466 6580 14476
rect 6748 13524 6804 13534
rect 6748 13430 6804 13468
rect 6412 12962 6468 13132
rect 6412 12910 6414 12962
rect 6466 12910 6468 12962
rect 6412 12292 6468 12910
rect 6412 12226 6468 12236
rect 6860 12852 6916 12862
rect 6860 12178 6916 12796
rect 6860 12126 6862 12178
rect 6914 12126 6916 12178
rect 6860 12068 6916 12126
rect 6636 12012 6916 12068
rect 6076 11330 6132 11340
rect 6188 11844 6244 11854
rect 5964 11170 6020 11182
rect 5964 11118 5966 11170
rect 6018 11118 6020 11170
rect 5852 10724 5908 10734
rect 5852 10630 5908 10668
rect 5404 10558 5406 10610
rect 5458 10558 5460 10610
rect 5404 10546 5460 10558
rect 5964 10612 6020 11118
rect 5964 10546 6020 10556
rect 5180 9774 5182 9826
rect 5234 9774 5236 9826
rect 5180 9762 5236 9774
rect 3804 9436 4068 9446
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 3804 9370 4068 9380
rect 4464 8652 4728 8662
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4464 8586 4728 8596
rect 3804 7868 4068 7878
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 3804 7802 4068 7812
rect 4464 7084 4728 7094
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4464 7018 4728 7028
rect 3804 6300 4068 6310
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 3804 6234 4068 6244
rect 4464 5516 4728 5526
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4464 5450 4728 5460
rect 3804 4732 4068 4742
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 3804 4666 4068 4676
rect 4464 3948 4728 3958
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4464 3882 4728 3892
rect 6188 3388 6244 11788
rect 6636 11394 6692 12012
rect 6636 11342 6638 11394
rect 6690 11342 6692 11394
rect 6636 11330 6692 11342
rect 6972 11506 7028 17388
rect 7084 17220 7140 17230
rect 7084 16770 7140 17164
rect 7084 16718 7086 16770
rect 7138 16718 7140 16770
rect 7084 16706 7140 16718
rect 7196 13188 7252 18172
rect 7308 15090 7364 15102
rect 7308 15038 7310 15090
rect 7362 15038 7364 15090
rect 7308 14868 7364 15038
rect 7308 14802 7364 14812
rect 7420 13970 7476 19180
rect 7756 19236 7812 23886
rect 7980 22596 8036 26852
rect 8092 26068 8148 26078
rect 8092 25974 8148 26012
rect 8316 25060 8372 27020
rect 8540 25620 8596 27356
rect 8652 27076 8708 28476
rect 8652 27010 8708 27020
rect 8316 24994 8372 25004
rect 8428 25564 8596 25620
rect 8316 24724 8372 24734
rect 8204 24722 8372 24724
rect 8204 24670 8318 24722
rect 8370 24670 8372 24722
rect 8204 24668 8372 24670
rect 8204 22708 8260 24668
rect 8316 24658 8372 24668
rect 8316 22932 8372 22942
rect 8316 22838 8372 22876
rect 8204 22652 8372 22708
rect 7868 22540 8036 22596
rect 7868 21812 7924 22540
rect 8092 22370 8148 22382
rect 8092 22318 8094 22370
rect 8146 22318 8148 22370
rect 8092 22260 8148 22318
rect 8092 22194 8148 22204
rect 8204 22372 8260 22382
rect 8092 21812 8148 21822
rect 7868 21756 8036 21812
rect 7868 21586 7924 21598
rect 7868 21534 7870 21586
rect 7922 21534 7924 21586
rect 7868 21026 7924 21534
rect 7868 20974 7870 21026
rect 7922 20974 7924 21026
rect 7868 20962 7924 20974
rect 7756 19170 7812 19180
rect 7868 20804 7924 20814
rect 7868 17108 7924 20748
rect 7756 17052 7924 17108
rect 7756 15428 7812 17052
rect 7756 15362 7812 15372
rect 7868 16884 7924 16894
rect 7868 15314 7924 16828
rect 7980 15652 8036 21756
rect 8092 20804 8148 21756
rect 8092 20738 8148 20748
rect 8204 19458 8260 22316
rect 8316 21028 8372 22652
rect 8428 21588 8484 25564
rect 8764 25172 8820 38612
rect 8988 37266 9044 38780
rect 8988 37214 8990 37266
rect 9042 37214 9044 37266
rect 8988 37202 9044 37214
rect 9100 36484 9156 48748
rect 9772 42756 9828 42766
rect 9436 41074 9492 41086
rect 9436 41022 9438 41074
rect 9490 41022 9492 41074
rect 9324 40402 9380 40414
rect 9324 40350 9326 40402
rect 9378 40350 9380 40402
rect 9324 40292 9380 40350
rect 9324 40226 9380 40236
rect 9436 39844 9492 41022
rect 9324 39788 9492 39844
rect 9548 41076 9604 41086
rect 8876 36428 9156 36484
rect 9212 38052 9268 38062
rect 9212 37716 9268 37996
rect 8876 35700 8932 36428
rect 8988 36260 9044 36270
rect 8988 36166 9044 36204
rect 9100 36036 9156 36046
rect 8876 35644 9044 35700
rect 8876 35476 8932 35486
rect 8876 35382 8932 35420
rect 8988 32788 9044 35644
rect 9100 35476 9156 35980
rect 9100 35410 9156 35420
rect 9212 34130 9268 37660
rect 9324 37604 9380 39788
rect 9436 39620 9492 39630
rect 9548 39620 9604 41020
rect 9436 39618 9604 39620
rect 9436 39566 9438 39618
rect 9490 39566 9604 39618
rect 9436 39564 9604 39566
rect 9436 39554 9492 39564
rect 9548 38668 9604 39564
rect 9772 38668 9828 42700
rect 9996 40292 10052 40302
rect 9884 39956 9940 39966
rect 9884 39842 9940 39900
rect 9884 39790 9886 39842
rect 9938 39790 9940 39842
rect 9884 39778 9940 39790
rect 9996 38668 10052 40236
rect 9324 37538 9380 37548
rect 9436 38612 9604 38668
rect 9660 38612 9828 38668
rect 9884 38612 10052 38668
rect 10108 38668 10164 52332
rect 10892 50820 10948 50830
rect 10892 42084 10948 50764
rect 12684 50428 12740 52444
rect 12684 50372 13076 50428
rect 11788 48916 11844 48926
rect 10892 42018 10948 42028
rect 11340 43652 11396 43662
rect 10556 41298 10612 41310
rect 10556 41246 10558 41298
rect 10610 41246 10612 41298
rect 10556 41188 10612 41246
rect 10556 41122 10612 41132
rect 10220 41076 10276 41086
rect 10220 40982 10276 41020
rect 10444 40402 10500 40414
rect 10444 40350 10446 40402
rect 10498 40350 10500 40402
rect 10108 38612 10388 38668
rect 9436 37380 9492 38612
rect 9548 38052 9604 38062
rect 9548 37958 9604 37996
rect 9324 37324 9492 37380
rect 9324 36484 9380 37324
rect 9548 37268 9604 37278
rect 9324 36418 9380 36428
rect 9436 37266 9604 37268
rect 9436 37214 9550 37266
rect 9602 37214 9604 37266
rect 9436 37212 9604 37214
rect 9324 36260 9380 36270
rect 9324 35698 9380 36204
rect 9324 35646 9326 35698
rect 9378 35646 9380 35698
rect 9324 35634 9380 35646
rect 9212 34078 9214 34130
rect 9266 34078 9268 34130
rect 9212 33236 9268 34078
rect 9212 33170 9268 33180
rect 9324 35364 9380 35374
rect 8988 32732 9156 32788
rect 8876 31780 8932 31790
rect 8876 31686 8932 31724
rect 8988 29204 9044 29214
rect 8988 29110 9044 29148
rect 8988 27972 9044 27982
rect 8764 25106 8820 25116
rect 8876 25506 8932 25518
rect 8876 25454 8878 25506
rect 8930 25454 8932 25506
rect 8876 24724 8932 25454
rect 8540 24668 8932 24724
rect 8540 24610 8596 24668
rect 8540 24558 8542 24610
rect 8594 24558 8596 24610
rect 8540 24546 8596 24558
rect 8764 24500 8820 24510
rect 8652 23380 8708 23390
rect 8428 21522 8484 21532
rect 8540 22484 8596 22494
rect 8540 21586 8596 22428
rect 8540 21534 8542 21586
rect 8594 21534 8596 21586
rect 8540 21522 8596 21534
rect 8316 20962 8372 20972
rect 8316 20132 8372 20142
rect 8316 20038 8372 20076
rect 8204 19406 8206 19458
rect 8258 19406 8260 19458
rect 8204 19394 8260 19406
rect 8092 18450 8148 18462
rect 8092 18398 8094 18450
rect 8146 18398 8148 18450
rect 8092 17668 8148 18398
rect 8092 17602 8148 17612
rect 8428 18338 8484 18350
rect 8428 18286 8430 18338
rect 8482 18286 8484 18338
rect 8204 17442 8260 17454
rect 8204 17390 8206 17442
rect 8258 17390 8260 17442
rect 8204 16324 8260 17390
rect 8316 16996 8372 17006
rect 8316 16902 8372 16940
rect 8428 16660 8484 18286
rect 8428 16594 8484 16604
rect 8204 16258 8260 16268
rect 8316 16212 8372 16222
rect 8092 15988 8148 15998
rect 8092 15894 8148 15932
rect 7980 15596 8148 15652
rect 7868 15262 7870 15314
rect 7922 15262 7924 15314
rect 7868 15250 7924 15262
rect 7980 15428 8036 15438
rect 7644 14756 7700 14766
rect 7420 13918 7422 13970
rect 7474 13918 7476 13970
rect 7420 13906 7476 13918
rect 7532 14532 7588 14542
rect 7196 13132 7364 13188
rect 7196 12962 7252 12974
rect 7196 12910 7198 12962
rect 7250 12910 7252 12962
rect 7196 12628 7252 12910
rect 7196 12562 7252 12572
rect 6972 11454 6974 11506
rect 7026 11454 7028 11506
rect 6748 10836 6804 10846
rect 6748 10722 6804 10780
rect 6748 10670 6750 10722
rect 6802 10670 6804 10722
rect 6748 10658 6804 10670
rect 6972 9940 7028 11454
rect 7308 12066 7364 13132
rect 7308 12014 7310 12066
rect 7362 12014 7364 12066
rect 7308 11508 7364 12014
rect 7308 11442 7364 11452
rect 7532 10836 7588 14476
rect 7644 14530 7700 14700
rect 7644 14478 7646 14530
rect 7698 14478 7700 14530
rect 7644 14466 7700 14478
rect 7308 10780 7588 10836
rect 7644 14308 7700 14318
rect 7084 10612 7140 10622
rect 7084 10518 7140 10556
rect 6972 9884 7140 9940
rect 6972 9716 7028 9726
rect 6972 9622 7028 9660
rect 7084 8932 7140 9884
rect 7308 9156 7364 10780
rect 7532 10612 7588 10622
rect 7644 10612 7700 14252
rect 7756 13412 7812 13422
rect 7756 13186 7812 13356
rect 7756 13134 7758 13186
rect 7810 13134 7812 13186
rect 7756 13122 7812 13134
rect 7980 10836 8036 15372
rect 7980 10770 8036 10780
rect 7308 9062 7364 9100
rect 7420 10610 7700 10612
rect 7420 10558 7534 10610
rect 7586 10558 7700 10610
rect 7420 10556 7700 10558
rect 7420 10052 7476 10556
rect 7532 10546 7588 10556
rect 7756 10386 7812 10398
rect 7756 10334 7758 10386
rect 7810 10334 7812 10386
rect 7084 8866 7140 8876
rect 7420 8036 7476 9996
rect 7532 10052 7588 10062
rect 7756 10052 7812 10334
rect 7532 10050 7812 10052
rect 7532 9998 7534 10050
rect 7586 9998 7812 10050
rect 7532 9996 7812 9998
rect 7532 9986 7588 9996
rect 7644 8932 7700 8942
rect 7644 8484 7700 8876
rect 7756 8484 7812 8494
rect 7644 8482 7812 8484
rect 7644 8430 7758 8482
rect 7810 8430 7812 8482
rect 7644 8428 7812 8430
rect 7756 8418 7812 8428
rect 7420 7970 7476 7980
rect 8092 3388 8148 15596
rect 8316 15202 8372 16156
rect 8316 15150 8318 15202
rect 8370 15150 8372 15202
rect 8316 15138 8372 15150
rect 8652 13860 8708 23324
rect 8652 13794 8708 13804
rect 8204 13746 8260 13758
rect 8204 13694 8206 13746
rect 8258 13694 8260 13746
rect 8204 12852 8260 13694
rect 8204 12758 8260 12796
rect 8316 13748 8372 13758
rect 8204 11396 8260 11406
rect 8204 11302 8260 11340
rect 8316 10610 8372 13692
rect 8540 12180 8596 12190
rect 8540 12086 8596 12124
rect 8764 10836 8820 24444
rect 8876 24388 8932 24398
rect 8876 22258 8932 24332
rect 8988 23380 9044 27916
rect 8988 23314 9044 23324
rect 8876 22206 8878 22258
rect 8930 22206 8932 22258
rect 8876 21140 8932 22206
rect 8876 21074 8932 21084
rect 8988 23154 9044 23166
rect 8988 23102 8990 23154
rect 9042 23102 9044 23154
rect 8988 20130 9044 23102
rect 8988 20078 8990 20130
rect 9042 20078 9044 20130
rect 8988 20066 9044 20078
rect 8876 20020 8932 20030
rect 8876 18564 8932 19964
rect 9100 19796 9156 32732
rect 9212 32564 9268 32574
rect 9212 31668 9268 32508
rect 9324 32562 9380 35308
rect 9324 32510 9326 32562
rect 9378 32510 9380 32562
rect 9324 32228 9380 32510
rect 9324 32162 9380 32172
rect 9436 31892 9492 37212
rect 9548 37202 9604 37212
rect 9548 36484 9604 36494
rect 9548 33684 9604 36428
rect 9548 33346 9604 33628
rect 9548 33294 9550 33346
rect 9602 33294 9604 33346
rect 9548 33282 9604 33294
rect 9436 31836 9604 31892
rect 9324 31668 9380 31678
rect 9212 31666 9380 31668
rect 9212 31614 9326 31666
rect 9378 31614 9380 31666
rect 9212 31612 9380 31614
rect 9324 31602 9380 31612
rect 9436 30212 9492 30222
rect 9548 30212 9604 31836
rect 9436 30210 9604 30212
rect 9436 30158 9438 30210
rect 9490 30158 9604 30210
rect 9436 30156 9604 30158
rect 9436 27972 9492 30156
rect 9436 27906 9492 27916
rect 9548 29316 9604 29326
rect 9324 27860 9380 27870
rect 9324 27766 9380 27804
rect 9212 26066 9268 26078
rect 9212 26014 9214 26066
rect 9266 26014 9268 26066
rect 9212 24722 9268 26014
rect 9324 26068 9380 26078
rect 9324 25060 9380 26012
rect 9436 25620 9492 25630
rect 9548 25620 9604 29260
rect 9436 25618 9604 25620
rect 9436 25566 9438 25618
rect 9490 25566 9604 25618
rect 9436 25564 9604 25566
rect 9436 25554 9492 25564
rect 9324 25004 9492 25060
rect 9212 24670 9214 24722
rect 9266 24670 9268 24722
rect 9212 24658 9268 24670
rect 9324 24724 9380 24734
rect 9324 24050 9380 24668
rect 9324 23998 9326 24050
rect 9378 23998 9380 24050
rect 9324 23986 9380 23998
rect 9436 23042 9492 25004
rect 9660 24948 9716 38612
rect 9772 37604 9828 37614
rect 9772 35476 9828 37548
rect 9884 35700 9940 38612
rect 9996 38162 10052 38174
rect 9996 38110 9998 38162
rect 10050 38110 10052 38162
rect 9996 36596 10052 38110
rect 10108 36708 10164 36718
rect 10108 36614 10164 36652
rect 9996 36530 10052 36540
rect 9996 35700 10052 35710
rect 9884 35698 10052 35700
rect 9884 35646 9998 35698
rect 10050 35646 10052 35698
rect 9884 35644 10052 35646
rect 9772 35420 9940 35476
rect 9772 30770 9828 30782
rect 9772 30718 9774 30770
rect 9826 30718 9828 30770
rect 9772 30210 9828 30718
rect 9772 30158 9774 30210
rect 9826 30158 9828 30210
rect 9772 30146 9828 30158
rect 9772 29428 9828 29438
rect 9772 27858 9828 29372
rect 9772 27806 9774 27858
rect 9826 27806 9828 27858
rect 9772 27794 9828 27806
rect 9884 26964 9940 35420
rect 9996 35140 10052 35644
rect 9996 35074 10052 35084
rect 9996 33572 10052 33582
rect 9996 33478 10052 33516
rect 10332 32340 10388 38612
rect 10444 32788 10500 40350
rect 11004 39508 11060 39518
rect 11004 39414 11060 39452
rect 10556 38834 10612 38846
rect 10556 38782 10558 38834
rect 10610 38782 10612 38834
rect 10556 38052 10612 38782
rect 10556 37986 10612 37996
rect 11004 38722 11060 38734
rect 11004 38670 11006 38722
rect 11058 38670 11060 38722
rect 11004 37940 11060 38670
rect 11116 38052 11172 38062
rect 11116 37958 11172 37996
rect 10668 37266 10724 37278
rect 10668 37214 10670 37266
rect 10722 37214 10724 37266
rect 10556 36372 10612 36382
rect 10556 35812 10612 36316
rect 10556 35746 10612 35756
rect 10556 34802 10612 34814
rect 10556 34750 10558 34802
rect 10610 34750 10612 34802
rect 10556 33012 10612 34750
rect 10668 33124 10724 37214
rect 10668 33058 10724 33068
rect 10892 35698 10948 35710
rect 10892 35646 10894 35698
rect 10946 35646 10948 35698
rect 10556 32946 10612 32956
rect 10444 32732 10836 32788
rect 10444 32564 10500 32574
rect 10444 32470 10500 32508
rect 10332 32284 10612 32340
rect 9996 32228 10052 32238
rect 9996 30100 10052 32172
rect 10444 30994 10500 31006
rect 10444 30942 10446 30994
rect 10498 30942 10500 30994
rect 10444 30434 10500 30942
rect 10444 30382 10446 30434
rect 10498 30382 10500 30434
rect 10444 30370 10500 30382
rect 9996 29876 10052 30044
rect 9996 29810 10052 29820
rect 10220 30212 10276 30222
rect 10220 29428 10276 30156
rect 10220 29362 10276 29372
rect 10108 29204 10164 29214
rect 10108 29202 10500 29204
rect 10108 29150 10110 29202
rect 10162 29150 10500 29202
rect 10108 29148 10500 29150
rect 10108 29138 10164 29148
rect 10444 27858 10500 29148
rect 10444 27806 10446 27858
rect 10498 27806 10500 27858
rect 10444 27794 10500 27806
rect 9996 27636 10052 27646
rect 10556 27636 10612 32284
rect 9996 27634 10164 27636
rect 9996 27582 9998 27634
rect 10050 27582 10164 27634
rect 9996 27580 10164 27582
rect 9996 27570 10052 27580
rect 10108 27300 10164 27580
rect 10444 27580 10612 27636
rect 10668 31332 10724 31342
rect 10220 27300 10276 27310
rect 10108 27298 10276 27300
rect 10108 27246 10222 27298
rect 10274 27246 10276 27298
rect 10108 27244 10276 27246
rect 10220 27234 10276 27244
rect 10444 26908 10500 27580
rect 9884 26898 9940 26908
rect 9660 24882 9716 24892
rect 10220 26852 10500 26908
rect 10556 27300 10612 27310
rect 9436 22990 9438 23042
rect 9490 22990 9492 23042
rect 9436 22978 9492 22990
rect 9772 24722 9828 24734
rect 9772 24670 9774 24722
rect 9826 24670 9828 24722
rect 9772 22484 9828 24670
rect 9884 23938 9940 23950
rect 9884 23886 9886 23938
rect 9938 23886 9940 23938
rect 9884 22594 9940 23886
rect 9884 22542 9886 22594
rect 9938 22542 9940 22594
rect 9884 22530 9940 22542
rect 10220 22596 10276 26852
rect 10332 25620 10388 25630
rect 10332 24724 10388 25564
rect 10444 25394 10500 25406
rect 10444 25342 10446 25394
rect 10498 25342 10500 25394
rect 10444 25172 10500 25342
rect 10444 25106 10500 25116
rect 10332 24668 10500 24724
rect 10220 22530 10276 22540
rect 10332 22932 10388 22942
rect 9772 22418 9828 22428
rect 10332 22482 10388 22876
rect 10332 22430 10334 22482
rect 10386 22430 10388 22482
rect 10332 22418 10388 22430
rect 9212 22372 9268 22382
rect 9212 22278 9268 22316
rect 9660 22370 9716 22382
rect 9660 22318 9662 22370
rect 9714 22318 9716 22370
rect 9436 21588 9492 21598
rect 9436 20692 9492 21532
rect 9660 21028 9716 22318
rect 10108 21588 10164 21598
rect 10108 21586 10276 21588
rect 10108 21534 10110 21586
rect 10162 21534 10276 21586
rect 10108 21532 10276 21534
rect 10108 21522 10164 21532
rect 9436 20626 9492 20636
rect 9548 20914 9604 20926
rect 9548 20862 9550 20914
rect 9602 20862 9604 20914
rect 9324 20580 9380 20590
rect 9324 19908 9380 20524
rect 9548 20356 9604 20862
rect 9660 20580 9716 20972
rect 9772 21364 9828 21374
rect 9772 21026 9828 21308
rect 9772 20974 9774 21026
rect 9826 20974 9828 21026
rect 9772 20962 9828 20974
rect 9884 20804 9940 20814
rect 9884 20710 9940 20748
rect 9996 20802 10052 20814
rect 9996 20750 9998 20802
rect 10050 20750 10052 20802
rect 9660 20524 9940 20580
rect 9548 20290 9604 20300
rect 8876 18498 8932 18508
rect 8988 19740 9156 19796
rect 9212 19906 9380 19908
rect 9212 19854 9326 19906
rect 9378 19854 9380 19906
rect 9212 19852 9380 19854
rect 8988 14420 9044 19740
rect 9100 16098 9156 16110
rect 9100 16046 9102 16098
rect 9154 16046 9156 16098
rect 9100 15540 9156 16046
rect 9100 15474 9156 15484
rect 8988 14354 9044 14364
rect 9212 13076 9268 19852
rect 9324 19842 9380 19852
rect 9548 19796 9604 19806
rect 9548 19234 9604 19740
rect 9548 19182 9550 19234
rect 9602 19182 9604 19234
rect 9548 19170 9604 19182
rect 9436 18676 9492 18686
rect 9324 16100 9380 16110
rect 9324 16006 9380 16044
rect 9436 15148 9492 18620
rect 9548 18564 9604 18574
rect 9548 17666 9604 18508
rect 9660 18228 9716 18238
rect 9660 18226 9828 18228
rect 9660 18174 9662 18226
rect 9714 18174 9828 18226
rect 9660 18172 9828 18174
rect 9660 18162 9716 18172
rect 9548 17614 9550 17666
rect 9602 17614 9604 17666
rect 9548 17602 9604 17614
rect 9660 17554 9716 17566
rect 9660 17502 9662 17554
rect 9714 17502 9716 17554
rect 9660 16884 9716 17502
rect 9660 16818 9716 16828
rect 9548 16210 9604 16222
rect 9548 16158 9550 16210
rect 9602 16158 9604 16210
rect 9548 15428 9604 16158
rect 9772 16212 9828 18172
rect 9884 17444 9940 20524
rect 9996 19460 10052 20750
rect 9996 19394 10052 19404
rect 10220 18564 10276 21532
rect 10444 21474 10500 24668
rect 10556 23268 10612 27244
rect 10668 25060 10724 31276
rect 10780 27412 10836 32732
rect 10892 31444 10948 35646
rect 11004 35138 11060 37884
rect 11340 35812 11396 43596
rect 11788 42980 11844 48860
rect 11788 42914 11844 42924
rect 12012 44548 12068 44558
rect 11788 40964 11844 40974
rect 11788 40962 11956 40964
rect 11788 40910 11790 40962
rect 11842 40910 11956 40962
rect 11788 40908 11956 40910
rect 11788 40898 11844 40908
rect 11900 39732 11956 40908
rect 11900 39666 11956 39676
rect 11788 39618 11844 39630
rect 11788 39566 11790 39618
rect 11842 39566 11844 39618
rect 11452 39506 11508 39518
rect 11452 39454 11454 39506
rect 11506 39454 11508 39506
rect 11452 38668 11508 39454
rect 11788 39508 11844 39566
rect 11788 39442 11844 39452
rect 11452 38612 11620 38668
rect 11564 37938 11620 38612
rect 11900 38052 11956 38062
rect 11900 37958 11956 37996
rect 11564 37886 11566 37938
rect 11618 37886 11620 37938
rect 11452 35812 11508 35822
rect 11340 35810 11508 35812
rect 11340 35758 11454 35810
rect 11506 35758 11508 35810
rect 11340 35756 11508 35758
rect 11452 35746 11508 35756
rect 11004 35086 11006 35138
rect 11058 35086 11060 35138
rect 11004 35074 11060 35086
rect 11116 33122 11172 33134
rect 11116 33070 11118 33122
rect 11170 33070 11172 33122
rect 10892 31378 10948 31388
rect 11004 32338 11060 32350
rect 11004 32286 11006 32338
rect 11058 32286 11060 32338
rect 11004 31108 11060 32286
rect 11004 31042 11060 31052
rect 10892 30882 10948 30894
rect 10892 30830 10894 30882
rect 10946 30830 10948 30882
rect 10892 30436 10948 30830
rect 10892 30370 10948 30380
rect 11116 30210 11172 33070
rect 11452 33124 11508 33134
rect 11340 31108 11396 31118
rect 11340 30994 11396 31052
rect 11340 30942 11342 30994
rect 11394 30942 11396 30994
rect 11340 30930 11396 30942
rect 11116 30158 11118 30210
rect 11170 30158 11172 30210
rect 11116 30146 11172 30158
rect 11452 30210 11508 33068
rect 11452 30158 11454 30210
rect 11506 30158 11508 30210
rect 11452 30100 11508 30158
rect 11228 30044 11508 30100
rect 11004 28868 11060 28878
rect 10892 28532 10948 28542
rect 10892 28438 10948 28476
rect 10780 27346 10836 27356
rect 10892 27972 10948 27982
rect 10780 27188 10836 27198
rect 10892 27188 10948 27916
rect 10780 27186 10948 27188
rect 10780 27134 10782 27186
rect 10834 27134 10948 27186
rect 10780 27132 10948 27134
rect 10780 27122 10836 27132
rect 11004 26908 11060 28812
rect 10892 26852 11060 26908
rect 11228 27858 11284 30044
rect 11340 28868 11396 28878
rect 11340 28774 11396 28812
rect 11228 27806 11230 27858
rect 11282 27806 11284 27858
rect 10892 25618 10948 26852
rect 10892 25566 10894 25618
rect 10946 25566 10948 25618
rect 10668 24994 10724 25004
rect 10780 25172 10836 25182
rect 10668 24722 10724 24734
rect 10668 24670 10670 24722
rect 10722 24670 10724 24722
rect 10668 23492 10724 24670
rect 10780 23826 10836 25116
rect 10780 23774 10782 23826
rect 10834 23774 10836 23826
rect 10780 23716 10836 23774
rect 10780 23650 10836 23660
rect 10668 23426 10724 23436
rect 10556 23212 10836 23268
rect 10556 23044 10612 23054
rect 10556 22950 10612 22988
rect 10444 21422 10446 21474
rect 10498 21422 10500 21474
rect 10444 21410 10500 21422
rect 10444 20804 10500 20814
rect 10780 20804 10836 23212
rect 10892 21476 10948 25566
rect 10892 21410 10948 21420
rect 11004 24388 11060 24398
rect 11004 21028 11060 24332
rect 11228 24276 11284 27806
rect 11340 28532 11396 28542
rect 11340 27076 11396 28476
rect 11340 26982 11396 27020
rect 11564 24388 11620 37886
rect 11788 36370 11844 36382
rect 11788 36318 11790 36370
rect 11842 36318 11844 36370
rect 11788 35700 11844 36318
rect 11900 35700 11956 35710
rect 11788 35698 11956 35700
rect 11788 35646 11902 35698
rect 11954 35646 11956 35698
rect 11788 35644 11956 35646
rect 12012 35700 12068 44492
rect 12236 41860 12292 41870
rect 12124 41300 12180 41310
rect 12124 39396 12180 41244
rect 12124 39330 12180 39340
rect 12124 38610 12180 38622
rect 12124 38558 12126 38610
rect 12178 38558 12180 38610
rect 12124 38052 12180 38558
rect 12124 37986 12180 37996
rect 12124 36596 12180 36606
rect 12124 36502 12180 36540
rect 12012 35644 12180 35700
rect 11788 33346 11844 35644
rect 11900 35634 11956 35644
rect 12124 35252 12180 35644
rect 12124 35186 12180 35196
rect 12124 34916 12180 34926
rect 12124 34822 12180 34860
rect 12236 34244 12292 41804
rect 12908 40180 12964 40190
rect 12460 40178 12964 40180
rect 12460 40126 12910 40178
rect 12962 40126 12964 40178
rect 12460 40124 12964 40126
rect 12460 39842 12516 40124
rect 12908 40114 12964 40124
rect 13020 39956 13076 50372
rect 13916 42868 13972 42878
rect 12460 39790 12462 39842
rect 12514 39790 12516 39842
rect 12460 39778 12516 39790
rect 12796 39900 13076 39956
rect 13132 42644 13188 42654
rect 12348 39620 12404 39630
rect 12348 39618 12516 39620
rect 12348 39566 12350 39618
rect 12402 39566 12516 39618
rect 12348 39564 12516 39566
rect 12348 39554 12404 39564
rect 12236 34178 12292 34188
rect 12348 39396 12404 39406
rect 12348 33684 12404 39340
rect 12460 38612 12516 39564
rect 12796 38668 12852 39900
rect 13132 39844 13188 42588
rect 13356 40516 13412 40526
rect 13020 39788 13188 39844
rect 13244 40514 13412 40516
rect 13244 40462 13358 40514
rect 13410 40462 13412 40514
rect 13244 40460 13412 40462
rect 12908 39732 12964 39742
rect 12908 39638 12964 39676
rect 12460 38056 12516 38556
rect 12684 38612 12852 38668
rect 12572 38276 12628 38286
rect 12572 38182 12628 38220
rect 12460 38004 12462 38056
rect 12514 38004 12516 38056
rect 12460 37940 12516 38004
rect 12460 37874 12516 37884
rect 12572 34802 12628 34814
rect 12572 34750 12574 34802
rect 12626 34750 12628 34802
rect 12572 34692 12628 34750
rect 12572 34132 12628 34636
rect 12684 34244 12740 38612
rect 12908 38610 12964 38622
rect 12908 38558 12910 38610
rect 12962 38558 12964 38610
rect 12908 38276 12964 38558
rect 12908 38210 12964 38220
rect 12796 36708 12852 36718
rect 12796 35588 12852 36652
rect 12908 35812 12964 35822
rect 13020 35812 13076 39788
rect 13132 38052 13188 38062
rect 13132 37958 13188 37996
rect 13244 36708 13300 40460
rect 13356 40450 13412 40460
rect 13580 39618 13636 39630
rect 13580 39566 13582 39618
rect 13634 39566 13636 39618
rect 13356 38946 13412 38958
rect 13356 38894 13358 38946
rect 13410 38894 13412 38946
rect 13356 38276 13412 38894
rect 13356 38210 13412 38220
rect 13580 38050 13636 39566
rect 13916 38668 13972 42812
rect 13916 38612 14196 38668
rect 13580 37998 13582 38050
rect 13634 37998 13636 38050
rect 13580 37156 13636 37998
rect 13580 37090 13636 37100
rect 13244 36642 13300 36652
rect 13916 36370 13972 36382
rect 13916 36318 13918 36370
rect 13970 36318 13972 36370
rect 13356 36260 13412 36270
rect 12908 35810 13076 35812
rect 12908 35758 12910 35810
rect 12962 35758 13076 35810
rect 12908 35756 13076 35758
rect 13244 36258 13412 36260
rect 13244 36206 13358 36258
rect 13410 36206 13412 36258
rect 13244 36204 13412 36206
rect 12908 35746 12964 35756
rect 12796 35532 13076 35588
rect 12908 34916 12964 34926
rect 12908 34822 12964 34860
rect 13020 34804 13076 35532
rect 13020 34738 13076 34748
rect 13132 35364 13188 35374
rect 13132 34468 13188 35308
rect 13244 35028 13300 36204
rect 13356 36194 13412 36204
rect 13356 35474 13412 35486
rect 13356 35422 13358 35474
rect 13410 35422 13412 35474
rect 13356 35140 13412 35422
rect 13580 35140 13636 35150
rect 13356 35138 13636 35140
rect 13356 35086 13582 35138
rect 13634 35086 13636 35138
rect 13356 35084 13636 35086
rect 13580 35074 13636 35084
rect 13244 34962 13300 34972
rect 13356 34914 13412 34926
rect 13356 34862 13358 34914
rect 13410 34862 13412 34914
rect 13356 34468 13412 34862
rect 13132 34412 13412 34468
rect 13692 34692 13748 34702
rect 12684 34188 12964 34244
rect 12572 34066 12628 34076
rect 12348 33628 12740 33684
rect 12348 33460 12404 33470
rect 12348 33458 12516 33460
rect 12348 33406 12350 33458
rect 12402 33406 12516 33458
rect 12348 33404 12516 33406
rect 12348 33394 12404 33404
rect 11788 33294 11790 33346
rect 11842 33294 11844 33346
rect 11788 32564 11844 33294
rect 11788 32498 11844 32508
rect 12124 32338 12180 32350
rect 12124 32286 12126 32338
rect 12178 32286 12180 32338
rect 12124 32228 12180 32286
rect 12124 32172 12404 32228
rect 12348 31778 12404 32172
rect 12348 31726 12350 31778
rect 12402 31726 12404 31778
rect 12348 31714 12404 31726
rect 12012 31666 12068 31678
rect 12012 31614 12014 31666
rect 12066 31614 12068 31666
rect 12012 31556 12068 31614
rect 12012 31490 12068 31500
rect 11564 24322 11620 24332
rect 11676 31108 11732 31118
rect 11676 27186 11732 31052
rect 11900 31108 11956 31118
rect 11900 31014 11956 31052
rect 12124 29652 12180 29662
rect 12124 29538 12180 29596
rect 12124 29486 12126 29538
rect 12178 29486 12180 29538
rect 12124 29474 12180 29486
rect 11788 29428 11844 29438
rect 11788 28868 11844 29372
rect 12460 29428 12516 33404
rect 12460 29362 12516 29372
rect 12572 30210 12628 30222
rect 12572 30158 12574 30210
rect 12626 30158 12628 30210
rect 11788 28802 11844 28812
rect 11676 27134 11678 27186
rect 11730 27134 11732 27186
rect 11116 24220 11284 24276
rect 11116 22820 11172 24220
rect 11676 24164 11732 27134
rect 11116 22754 11172 22764
rect 11228 24108 11732 24164
rect 11900 28644 11956 28654
rect 11228 24050 11284 24108
rect 11228 23998 11230 24050
rect 11282 23998 11284 24050
rect 11116 22484 11172 22494
rect 11116 22370 11172 22428
rect 11116 22318 11118 22370
rect 11170 22318 11172 22370
rect 11116 22306 11172 22318
rect 11004 20972 11172 21028
rect 10780 20748 10948 20804
rect 10444 20710 10500 20748
rect 10780 20578 10836 20590
rect 10780 20526 10782 20578
rect 10834 20526 10836 20578
rect 10556 20356 10612 20366
rect 10556 20130 10612 20300
rect 10556 20078 10558 20130
rect 10610 20078 10612 20130
rect 10556 20066 10612 20078
rect 10332 19236 10388 19246
rect 10332 19142 10388 19180
rect 10780 19012 10836 20526
rect 10892 19572 10948 20748
rect 10892 19506 10948 19516
rect 11004 20802 11060 20814
rect 11004 20750 11006 20802
rect 11058 20750 11060 20802
rect 10780 18946 10836 18956
rect 11004 18788 11060 20750
rect 11116 19572 11172 20972
rect 11228 19908 11284 23998
rect 11676 23380 11732 23390
rect 11564 23378 11732 23380
rect 11564 23326 11678 23378
rect 11730 23326 11732 23378
rect 11564 23324 11732 23326
rect 11452 23154 11508 23166
rect 11452 23102 11454 23154
rect 11506 23102 11508 23154
rect 11228 19842 11284 19852
rect 11340 22820 11396 22830
rect 11116 19516 11284 19572
rect 11116 19348 11172 19358
rect 11116 19254 11172 19292
rect 11004 18722 11060 18732
rect 10332 18564 10388 18574
rect 10220 18508 10332 18564
rect 10332 18470 10388 18508
rect 10108 18452 10164 18462
rect 9996 17778 10052 17790
rect 9996 17726 9998 17778
rect 10050 17726 10052 17778
rect 9996 17668 10052 17726
rect 9996 17602 10052 17612
rect 9884 17378 9940 17388
rect 9772 16146 9828 16156
rect 9884 16770 9940 16782
rect 9884 16718 9886 16770
rect 9938 16718 9940 16770
rect 9884 16098 9940 16718
rect 10108 16770 10164 18396
rect 11228 18340 11284 19516
rect 11340 19236 11396 22764
rect 11452 21812 11508 23102
rect 11452 21746 11508 21756
rect 11452 21588 11508 21598
rect 11452 20804 11508 21532
rect 11564 21140 11620 23324
rect 11676 23314 11732 23324
rect 11788 22930 11844 22942
rect 11788 22878 11790 22930
rect 11842 22878 11844 22930
rect 11676 21812 11732 21822
rect 11676 21718 11732 21756
rect 11564 21084 11732 21140
rect 11564 20804 11620 20814
rect 11452 20802 11620 20804
rect 11452 20750 11566 20802
rect 11618 20750 11620 20802
rect 11452 20748 11620 20750
rect 11564 20738 11620 20748
rect 11676 20468 11732 21084
rect 11788 20690 11844 22878
rect 11900 22596 11956 28588
rect 12460 28644 12516 28654
rect 12460 28550 12516 28588
rect 12012 27858 12068 27870
rect 12012 27806 12014 27858
rect 12066 27806 12068 27858
rect 12012 25732 12068 27806
rect 12012 25666 12068 25676
rect 12012 25284 12068 25294
rect 12012 25282 12404 25284
rect 12012 25230 12014 25282
rect 12066 25230 12404 25282
rect 12012 25228 12404 25230
rect 12012 25218 12068 25228
rect 12236 24610 12292 24622
rect 12236 24558 12238 24610
rect 12290 24558 12292 24610
rect 12012 24500 12068 24510
rect 12012 24406 12068 24444
rect 12124 24498 12180 24510
rect 12124 24446 12126 24498
rect 12178 24446 12180 24498
rect 12012 23044 12068 23054
rect 12012 22950 12068 22988
rect 11900 22540 12068 22596
rect 11900 22372 11956 22382
rect 11900 22278 11956 22316
rect 11788 20638 11790 20690
rect 11842 20638 11844 20690
rect 11788 20626 11844 20638
rect 11900 20802 11956 20814
rect 11900 20750 11902 20802
rect 11954 20750 11956 20802
rect 11676 20412 11844 20468
rect 11452 20020 11508 20030
rect 11452 19926 11508 19964
rect 11676 19908 11732 19918
rect 11676 19814 11732 19852
rect 11788 19794 11844 20412
rect 11900 20356 11956 20750
rect 11900 20290 11956 20300
rect 11788 19742 11790 19794
rect 11842 19742 11844 19794
rect 11788 19730 11844 19742
rect 11900 20018 11956 20030
rect 11900 19966 11902 20018
rect 11954 19966 11956 20018
rect 11676 19572 11732 19582
rect 11564 19460 11620 19470
rect 11564 19366 11620 19404
rect 11340 19180 11620 19236
rect 11228 18284 11396 18340
rect 10780 18226 10836 18238
rect 10780 18174 10782 18226
rect 10834 18174 10836 18226
rect 10780 17668 10836 18174
rect 11228 18116 11284 18126
rect 11228 17890 11284 18060
rect 11228 17838 11230 17890
rect 11282 17838 11284 17890
rect 11228 17826 11284 17838
rect 10780 17602 10836 17612
rect 11340 17444 11396 18284
rect 11340 17378 11396 17388
rect 10220 16994 10276 17006
rect 10220 16942 10222 16994
rect 10274 16942 10276 16994
rect 10220 16884 10276 16942
rect 10556 16884 10612 16894
rect 10220 16882 10612 16884
rect 10220 16830 10558 16882
rect 10610 16830 10612 16882
rect 10220 16828 10612 16830
rect 10556 16818 10612 16828
rect 10892 16882 10948 16894
rect 10892 16830 10894 16882
rect 10946 16830 10948 16882
rect 10108 16718 10110 16770
rect 10162 16718 10164 16770
rect 10108 16706 10164 16718
rect 10332 16660 10388 16670
rect 10108 16436 10164 16446
rect 10108 16322 10164 16380
rect 10108 16270 10110 16322
rect 10162 16270 10164 16322
rect 10108 16258 10164 16270
rect 10332 16212 10388 16604
rect 10892 16660 10948 16830
rect 10892 16594 10948 16604
rect 11004 16882 11060 16894
rect 11004 16830 11006 16882
rect 11058 16830 11060 16882
rect 10220 16210 10388 16212
rect 10220 16158 10334 16210
rect 10386 16158 10388 16210
rect 10220 16156 10388 16158
rect 9884 16046 9886 16098
rect 9938 16046 9940 16098
rect 9884 15988 9940 16046
rect 9996 16100 10052 16110
rect 9996 16006 10052 16044
rect 9660 15874 9716 15886
rect 9660 15822 9662 15874
rect 9714 15822 9716 15874
rect 9660 15652 9716 15822
rect 9660 15586 9716 15596
rect 9548 15334 9604 15372
rect 9884 15316 9940 15932
rect 10108 15316 10164 15326
rect 9884 15260 10108 15316
rect 10108 15222 10164 15260
rect 9436 15092 9828 15148
rect 9436 14756 9492 14766
rect 9436 14662 9492 14700
rect 9548 14644 9604 14654
rect 9548 14550 9604 14588
rect 9436 14308 9492 14318
rect 9436 14214 9492 14252
rect 9212 13010 9268 13020
rect 9324 13746 9380 13758
rect 9324 13694 9326 13746
rect 9378 13694 9380 13746
rect 9100 12852 9156 12862
rect 9324 12852 9380 13694
rect 9772 13636 9828 15092
rect 9996 15092 10052 15102
rect 9996 15090 10164 15092
rect 9996 15038 9998 15090
rect 10050 15038 10164 15090
rect 9996 15036 10164 15038
rect 9996 15026 10052 15036
rect 10108 14644 10164 15036
rect 10108 14550 10164 14588
rect 10220 14868 10276 16156
rect 10332 16146 10388 16156
rect 10780 15986 10836 15998
rect 10780 15934 10782 15986
rect 10834 15934 10836 15986
rect 10780 15876 10836 15934
rect 11004 15988 11060 16830
rect 11340 16770 11396 16782
rect 11340 16718 11342 16770
rect 11394 16718 11396 16770
rect 11228 16658 11284 16670
rect 11228 16606 11230 16658
rect 11282 16606 11284 16658
rect 11116 16324 11172 16334
rect 11116 16098 11172 16268
rect 11116 16046 11118 16098
rect 11170 16046 11172 16098
rect 11116 16034 11172 16046
rect 11004 15922 11060 15932
rect 10780 15810 10836 15820
rect 10556 15652 10612 15662
rect 10556 15314 10612 15596
rect 11228 15538 11284 16606
rect 11228 15486 11230 15538
rect 11282 15486 11284 15538
rect 11228 15474 11284 15486
rect 11004 15428 11060 15438
rect 11004 15334 11060 15372
rect 10556 15262 10558 15314
rect 10610 15262 10612 15314
rect 10556 15250 10612 15262
rect 11340 15316 11396 16718
rect 11340 15250 11396 15260
rect 11452 15314 11508 15326
rect 11452 15262 11454 15314
rect 11506 15262 11508 15314
rect 10780 15204 10836 15214
rect 10780 15202 11172 15204
rect 10780 15150 10782 15202
rect 10834 15150 11172 15202
rect 10780 15148 11172 15150
rect 11452 15148 11508 15262
rect 10780 15138 10836 15148
rect 10668 15092 10724 15102
rect 10220 14642 10276 14812
rect 10220 14590 10222 14642
rect 10274 14590 10276 14642
rect 10220 14578 10276 14590
rect 10444 15090 10724 15092
rect 10444 15038 10670 15090
rect 10722 15038 10724 15090
rect 10444 15036 10724 15038
rect 9996 14532 10052 14542
rect 9996 14438 10052 14476
rect 9772 13542 9828 13580
rect 9884 13748 9940 13758
rect 9436 13076 9492 13086
rect 9436 12982 9492 13020
rect 9156 12796 9380 12852
rect 9100 12758 9156 12796
rect 9884 12404 9940 13692
rect 9772 12348 9940 12404
rect 10108 12964 10164 12974
rect 9324 12180 9380 12190
rect 9324 12086 9380 12124
rect 8316 10558 8318 10610
rect 8370 10558 8372 10610
rect 8316 10546 8372 10558
rect 8652 10780 8820 10836
rect 8988 12066 9044 12078
rect 8988 12014 8990 12066
rect 9042 12014 9044 12066
rect 8988 11956 9044 12014
rect 9772 11956 9828 12348
rect 9884 12178 9940 12190
rect 9884 12126 9886 12178
rect 9938 12126 9940 12178
rect 9884 12068 9940 12126
rect 9884 12002 9940 12012
rect 9996 12068 10052 12078
rect 10108 12068 10164 12908
rect 9996 12066 10164 12068
rect 9996 12014 9998 12066
rect 10050 12014 10164 12066
rect 9996 12012 10164 12014
rect 10220 12068 10276 12078
rect 9996 12002 10052 12012
rect 8988 11900 9828 11956
rect 8316 8148 8372 8158
rect 8316 8054 8372 8092
rect 6076 3332 6244 3388
rect 7980 3332 8148 3388
rect 8652 3388 8708 10780
rect 8988 10610 9044 11900
rect 9772 11508 9828 11900
rect 10220 11788 10276 12012
rect 10108 11732 10276 11788
rect 9884 11508 9940 11518
rect 9772 11506 9940 11508
rect 9772 11454 9886 11506
rect 9938 11454 9940 11506
rect 9772 11452 9940 11454
rect 9884 11442 9940 11452
rect 8988 10558 8990 10610
rect 9042 10558 9044 10610
rect 8988 10546 9044 10558
rect 9884 10610 9940 10622
rect 9884 10558 9886 10610
rect 9938 10558 9940 10610
rect 9548 10500 9604 10510
rect 8876 9268 8932 9278
rect 8876 9174 8932 9212
rect 9548 9154 9604 10444
rect 9884 9828 9940 10558
rect 10108 9938 10164 11732
rect 10444 11620 10500 15036
rect 10668 15026 10724 15036
rect 11116 14754 11172 15148
rect 11340 15092 11508 15148
rect 11116 14702 11118 14754
rect 11170 14702 11172 14754
rect 11116 14690 11172 14702
rect 11228 14868 11284 14878
rect 11228 14754 11284 14812
rect 11228 14702 11230 14754
rect 11282 14702 11284 14754
rect 11228 14690 11284 14702
rect 10668 14532 10724 14542
rect 11340 14532 11396 15092
rect 10668 14530 11396 14532
rect 10668 14478 10670 14530
rect 10722 14478 11396 14530
rect 10668 14476 11396 14478
rect 10668 14466 10724 14476
rect 11004 14308 11060 14318
rect 11004 14214 11060 14252
rect 10444 11554 10500 11564
rect 10556 13636 10612 13646
rect 10220 11396 10276 11406
rect 10220 11302 10276 11340
rect 10556 10948 10612 13580
rect 10780 13636 10836 13646
rect 10668 12738 10724 12750
rect 10668 12686 10670 12738
rect 10722 12686 10724 12738
rect 10668 12178 10724 12686
rect 10668 12126 10670 12178
rect 10722 12126 10724 12178
rect 10668 12114 10724 12126
rect 10780 12068 10836 13580
rect 11004 13524 11060 13534
rect 11004 13522 11508 13524
rect 11004 13470 11006 13522
rect 11058 13470 11508 13522
rect 11004 13468 11508 13470
rect 11004 13458 11060 13468
rect 11340 12964 11396 12974
rect 10780 11394 10836 12012
rect 10892 12962 11396 12964
rect 10892 12910 11342 12962
rect 11394 12910 11396 12962
rect 10892 12908 11396 12910
rect 10892 11618 10948 12908
rect 11340 12898 11396 12908
rect 10892 11566 10894 11618
rect 10946 11566 10948 11618
rect 10892 11554 10948 11566
rect 11228 12178 11284 12190
rect 11228 12126 11230 12178
rect 11282 12126 11284 12178
rect 10780 11342 10782 11394
rect 10834 11342 10836 11394
rect 10780 11330 10836 11342
rect 11228 11396 11284 12126
rect 11228 11330 11284 11340
rect 11452 11394 11508 13468
rect 11452 11342 11454 11394
rect 11506 11342 11508 11394
rect 11452 11330 11508 11342
rect 11564 11172 11620 19180
rect 11676 16436 11732 19516
rect 11900 19460 11956 19966
rect 11900 19394 11956 19404
rect 11788 19236 11844 19246
rect 11788 19142 11844 19180
rect 11900 18228 11956 18238
rect 11900 18134 11956 18172
rect 12012 16996 12068 22540
rect 12124 21588 12180 24446
rect 12236 23380 12292 24558
rect 12348 24388 12404 25228
rect 12572 24836 12628 30158
rect 12684 26908 12740 33628
rect 12796 31780 12852 31790
rect 12796 27076 12852 31724
rect 12908 29988 12964 34188
rect 13020 32562 13076 32574
rect 13020 32510 13022 32562
rect 13074 32510 13076 32562
rect 13020 32002 13076 32510
rect 13020 31950 13022 32002
rect 13074 31950 13076 32002
rect 13020 31938 13076 31950
rect 13244 31780 13300 34412
rect 13356 34244 13412 34254
rect 13356 32674 13412 34188
rect 13468 33124 13524 33134
rect 13468 33122 13636 33124
rect 13468 33070 13470 33122
rect 13522 33070 13636 33122
rect 13468 33068 13636 33070
rect 13468 33058 13524 33068
rect 13356 32622 13358 32674
rect 13410 32622 13412 32674
rect 13356 32610 13412 32622
rect 13244 31714 13300 31724
rect 13580 31778 13636 33068
rect 13580 31726 13582 31778
rect 13634 31726 13636 31778
rect 13580 31714 13636 31726
rect 12908 29922 12964 29932
rect 13580 29428 13636 29438
rect 13468 29426 13636 29428
rect 13468 29374 13582 29426
rect 13634 29374 13636 29426
rect 13468 29372 13636 29374
rect 12908 28868 12964 28878
rect 12908 28754 12964 28812
rect 12908 28702 12910 28754
rect 12962 28702 12964 28754
rect 12908 28690 12964 28702
rect 13244 28644 13300 28654
rect 13020 28642 13300 28644
rect 13020 28590 13246 28642
rect 13298 28590 13300 28642
rect 13020 28588 13300 28590
rect 12908 27300 12964 27310
rect 13020 27300 13076 28588
rect 13244 28578 13300 28588
rect 12908 27298 13076 27300
rect 12908 27246 12910 27298
rect 12962 27246 13076 27298
rect 12908 27244 13076 27246
rect 12908 27234 12964 27244
rect 12796 27020 13076 27076
rect 13020 26908 13076 27020
rect 13468 27074 13524 29372
rect 13580 29362 13636 29372
rect 13468 27022 13470 27074
rect 13522 27022 13524 27074
rect 12684 26852 12964 26908
rect 13020 26852 13300 26908
rect 12908 26290 12964 26796
rect 12908 26238 12910 26290
rect 12962 26238 12964 26290
rect 12908 25620 12964 26238
rect 13244 26180 13300 26852
rect 13468 26516 13524 27022
rect 13468 26450 13524 26460
rect 13580 28868 13636 28878
rect 13580 27970 13636 28812
rect 13580 27918 13582 27970
rect 13634 27918 13636 27970
rect 13356 26404 13412 26414
rect 13356 26310 13412 26348
rect 13244 26114 13300 26124
rect 13132 25620 13188 25630
rect 12908 25618 13188 25620
rect 12908 25566 13134 25618
rect 13186 25566 13188 25618
rect 12908 25564 13188 25566
rect 12684 25394 12740 25406
rect 12684 25342 12686 25394
rect 12738 25342 12740 25394
rect 12684 25172 12740 25342
rect 13132 25284 13188 25564
rect 13132 25228 13524 25284
rect 12684 25106 12740 25116
rect 12572 24780 13300 24836
rect 12908 24612 12964 24622
rect 12796 24610 12964 24612
rect 12796 24558 12910 24610
rect 12962 24558 12964 24610
rect 12796 24556 12964 24558
rect 12348 24322 12404 24332
rect 12460 24500 12516 24510
rect 12348 23940 12404 23950
rect 12348 23846 12404 23884
rect 12236 23314 12292 23324
rect 12236 23042 12292 23054
rect 12236 22990 12238 23042
rect 12290 22990 12292 23042
rect 12236 22596 12292 22990
rect 12236 22530 12292 22540
rect 12124 21522 12180 21532
rect 12236 22036 12292 22046
rect 12236 21474 12292 21980
rect 12460 22036 12516 24444
rect 12796 23826 12852 24556
rect 12908 24546 12964 24556
rect 13132 24388 13188 24398
rect 13132 23938 13188 24332
rect 13132 23886 13134 23938
rect 13186 23886 13188 23938
rect 13132 23874 13188 23886
rect 12796 23774 12798 23826
rect 12850 23774 12852 23826
rect 12796 23044 12852 23774
rect 13132 23154 13188 23166
rect 13132 23102 13134 23154
rect 13186 23102 13188 23154
rect 12796 23042 12964 23044
rect 12796 22990 12798 23042
rect 12850 22990 12964 23042
rect 12796 22988 12964 22990
rect 12796 22978 12852 22988
rect 12460 21970 12516 21980
rect 12796 21812 12852 21822
rect 12236 21422 12238 21474
rect 12290 21422 12292 21474
rect 12124 21364 12180 21374
rect 12124 21270 12180 21308
rect 12236 20244 12292 21422
rect 12236 20178 12292 20188
rect 12460 21810 12852 21812
rect 12460 21758 12798 21810
rect 12850 21758 12852 21810
rect 12460 21756 12852 21758
rect 12124 20020 12180 20030
rect 12124 19234 12180 19964
rect 12236 20020 12292 20030
rect 12460 20020 12516 21756
rect 12796 21746 12852 21756
rect 12908 21588 12964 22988
rect 13020 22370 13076 22382
rect 13020 22318 13022 22370
rect 13074 22318 13076 22370
rect 13020 22148 13076 22318
rect 13020 22082 13076 22092
rect 12796 21532 12964 21588
rect 13132 21812 13188 23102
rect 12236 20018 12516 20020
rect 12236 19966 12238 20018
rect 12290 19966 12516 20018
rect 12236 19964 12516 19966
rect 12572 21252 12628 21262
rect 12236 19954 12292 19964
rect 12572 19908 12628 21196
rect 12796 20692 12852 21532
rect 12908 21364 12964 21374
rect 12908 21270 12964 21308
rect 12908 20692 12964 20702
rect 12460 19852 12628 19908
rect 12684 20690 12964 20692
rect 12684 20638 12910 20690
rect 12962 20638 12964 20690
rect 12684 20636 12964 20638
rect 12124 19182 12126 19234
rect 12178 19182 12180 19234
rect 12124 19170 12180 19182
rect 12348 19796 12404 19806
rect 12348 17666 12404 19740
rect 12348 17614 12350 17666
rect 12402 17614 12404 17666
rect 12124 16996 12180 17006
rect 12012 16994 12180 16996
rect 12012 16942 12126 16994
rect 12178 16942 12180 16994
rect 12012 16940 12180 16942
rect 12124 16930 12180 16940
rect 11676 16098 11732 16380
rect 11788 16882 11844 16894
rect 11788 16830 11790 16882
rect 11842 16830 11844 16882
rect 11788 16322 11844 16830
rect 11788 16270 11790 16322
rect 11842 16270 11844 16322
rect 11788 16258 11844 16270
rect 12236 16212 12292 16222
rect 12236 16118 12292 16156
rect 11676 16046 11678 16098
rect 11730 16046 11732 16098
rect 11676 16034 11732 16046
rect 12012 15876 12068 15886
rect 11900 15540 11956 15550
rect 11900 15446 11956 15484
rect 11788 15316 11844 15326
rect 11788 15222 11844 15260
rect 11900 15204 11956 15214
rect 12012 15204 12068 15820
rect 12348 15876 12404 17614
rect 12348 15810 12404 15820
rect 11900 15202 12068 15204
rect 11900 15150 11902 15202
rect 11954 15150 12068 15202
rect 11900 15148 12068 15150
rect 11900 15138 11956 15148
rect 12460 15092 12516 19852
rect 12572 19572 12628 19582
rect 12572 19346 12628 19516
rect 12572 19294 12574 19346
rect 12626 19294 12628 19346
rect 12572 19282 12628 19294
rect 12460 15026 12516 15036
rect 11900 13188 11956 13198
rect 11900 13074 11956 13132
rect 11900 13022 11902 13074
rect 11954 13022 11956 13074
rect 11900 13010 11956 13022
rect 12236 12964 12292 12974
rect 12236 12870 12292 12908
rect 12124 12180 12180 12190
rect 12124 12086 12180 12124
rect 12124 11844 12180 11854
rect 11564 11106 11620 11116
rect 12012 11396 12068 11406
rect 10108 9886 10110 9938
rect 10162 9886 10164 9938
rect 10108 9874 10164 9886
rect 10220 10892 10948 10948
rect 9884 9762 9940 9772
rect 9548 9102 9550 9154
rect 9602 9102 9604 9154
rect 9548 9090 9604 9102
rect 9660 9156 9716 9166
rect 9660 8258 9716 9100
rect 9884 8932 9940 8942
rect 9884 8838 9940 8876
rect 9660 8206 9662 8258
rect 9714 8206 9716 8258
rect 9660 8194 9716 8206
rect 10220 8370 10276 10892
rect 10444 10610 10500 10622
rect 10444 10558 10446 10610
rect 10498 10558 10500 10610
rect 10444 10500 10500 10558
rect 10444 10434 10500 10444
rect 10892 10498 10948 10892
rect 10892 10446 10894 10498
rect 10946 10446 10948 10498
rect 10892 10434 10948 10446
rect 11228 10500 11284 10510
rect 10892 10052 10948 10062
rect 10444 9826 10500 9838
rect 10444 9774 10446 9826
rect 10498 9774 10500 9826
rect 10444 9268 10500 9774
rect 10892 9826 10948 9996
rect 11116 9940 11172 9950
rect 10892 9774 10894 9826
rect 10946 9774 10948 9826
rect 10892 9762 10948 9774
rect 11004 9938 11172 9940
rect 11004 9886 11118 9938
rect 11170 9886 11172 9938
rect 11004 9884 11172 9886
rect 10444 9202 10500 9212
rect 10220 8318 10222 8370
rect 10274 8318 10276 8370
rect 10220 7474 10276 8318
rect 10220 7422 10222 7474
rect 10274 7422 10276 7474
rect 10220 7410 10276 7422
rect 11004 7474 11060 9884
rect 11116 9874 11172 9884
rect 11116 9268 11172 9278
rect 11228 9268 11284 10444
rect 11116 9266 11284 9268
rect 11116 9214 11118 9266
rect 11170 9214 11284 9266
rect 11116 9212 11284 9214
rect 11564 9826 11620 9838
rect 11564 9774 11566 9826
rect 11618 9774 11620 9826
rect 11116 9202 11172 9212
rect 11340 8484 11396 8494
rect 11564 8484 11620 9774
rect 12012 9828 12068 11340
rect 12124 10834 12180 11788
rect 12684 11396 12740 20636
rect 12908 20626 12964 20636
rect 12908 20468 12964 20478
rect 12796 20244 12852 20254
rect 12796 19012 12852 20188
rect 12908 20242 12964 20412
rect 12908 20190 12910 20242
rect 12962 20190 12964 20242
rect 12908 20178 12964 20190
rect 13132 20020 13188 21756
rect 13244 20356 13300 24780
rect 13356 24722 13412 24734
rect 13356 24670 13358 24722
rect 13410 24670 13412 24722
rect 13356 24500 13412 24670
rect 13356 24434 13412 24444
rect 13356 20804 13412 20814
rect 13356 20710 13412 20748
rect 13244 20300 13412 20356
rect 13244 20132 13300 20142
rect 13244 20038 13300 20076
rect 13132 19954 13188 19964
rect 13356 19796 13412 20300
rect 13468 20244 13524 25228
rect 13580 24052 13636 27918
rect 13692 28642 13748 34636
rect 13804 32340 13860 32350
rect 13804 30772 13860 32284
rect 13916 31444 13972 36318
rect 14028 35028 14084 35038
rect 14028 34934 14084 34972
rect 13916 31378 13972 31388
rect 13804 30706 13860 30716
rect 14140 30436 14196 38612
rect 14252 36932 14308 53452
rect 14252 36866 14308 36876
rect 14364 48244 14420 48254
rect 14364 36708 14420 48188
rect 14700 47068 14756 54348
rect 17500 53620 17556 55918
rect 19516 55970 19572 55982
rect 19516 55918 19518 55970
rect 19570 55918 19572 55970
rect 18844 55412 18900 55422
rect 18844 55318 18900 55356
rect 18284 55298 18340 55310
rect 19292 55300 19348 55310
rect 18284 55246 18286 55298
rect 18338 55246 18340 55298
rect 17500 53554 17556 53564
rect 18060 55188 18116 55198
rect 15148 52948 15204 52958
rect 14252 36652 14420 36708
rect 14476 47012 14756 47068
rect 14924 47908 14980 47918
rect 14252 35588 14308 36652
rect 14364 36484 14420 36494
rect 14364 36390 14420 36428
rect 14252 35532 14420 35588
rect 14364 32674 14420 35532
rect 14476 35308 14532 47012
rect 14588 39620 14644 39630
rect 14588 39618 14756 39620
rect 14588 39566 14590 39618
rect 14642 39566 14756 39618
rect 14588 39564 14756 39566
rect 14588 39554 14644 39564
rect 14700 38050 14756 39564
rect 14700 37998 14702 38050
rect 14754 37998 14756 38050
rect 14700 36820 14756 37998
rect 14700 36754 14756 36764
rect 14700 36596 14756 36606
rect 14700 35308 14756 36540
rect 14812 36484 14868 36494
rect 14812 36390 14868 36428
rect 14476 35252 14644 35308
rect 14700 35252 14868 35308
rect 14588 35140 14644 35252
rect 14588 35084 14756 35140
rect 14588 34916 14644 34926
rect 14364 32622 14366 32674
rect 14418 32622 14420 32674
rect 14364 32610 14420 32622
rect 14476 34914 14644 34916
rect 14476 34862 14590 34914
rect 14642 34862 14644 34914
rect 14476 34860 14644 34862
rect 14476 32340 14532 34860
rect 14588 34850 14644 34860
rect 14588 33460 14644 33470
rect 14588 33366 14644 33404
rect 14476 32284 14644 32340
rect 14252 31780 14308 31790
rect 14252 31778 14420 31780
rect 14252 31726 14254 31778
rect 14306 31726 14420 31778
rect 14252 31724 14420 31726
rect 14252 31714 14308 31724
rect 14252 31444 14308 31454
rect 14252 30996 14308 31388
rect 14252 30902 14308 30940
rect 14140 30380 14308 30436
rect 14140 30212 14196 30222
rect 13916 30210 14196 30212
rect 13916 30158 14142 30210
rect 14194 30158 14196 30210
rect 13916 30156 14196 30158
rect 13916 28866 13972 30156
rect 14140 30146 14196 30156
rect 13916 28814 13918 28866
rect 13970 28814 13972 28866
rect 13916 28802 13972 28814
rect 14140 29316 14196 29326
rect 14252 29316 14308 30380
rect 14140 29314 14308 29316
rect 14140 29262 14142 29314
rect 14194 29262 14308 29314
rect 14140 29260 14308 29262
rect 13692 28590 13694 28642
rect 13746 28590 13748 28642
rect 13692 27412 13748 28590
rect 14028 27860 14084 27870
rect 14028 27766 14084 27804
rect 13692 27346 13748 27356
rect 13916 27186 13972 27198
rect 13916 27134 13918 27186
rect 13970 27134 13972 27186
rect 13916 26852 13972 27134
rect 13916 26786 13972 26796
rect 14028 26066 14084 26078
rect 14028 26014 14030 26066
rect 14082 26014 14084 26066
rect 13804 25060 13860 25070
rect 13804 24724 13860 25004
rect 13580 23986 13636 23996
rect 13692 24722 13860 24724
rect 13692 24670 13806 24722
rect 13858 24670 13860 24722
rect 13692 24668 13860 24670
rect 13692 23940 13748 24668
rect 13804 24658 13860 24668
rect 13916 24612 13972 24622
rect 13916 24518 13972 24556
rect 13804 24164 13860 24174
rect 14028 24164 14084 26014
rect 14140 24388 14196 29260
rect 14364 28868 14420 31724
rect 14364 28802 14420 28812
rect 14364 28644 14420 28654
rect 14364 28550 14420 28588
rect 14588 28644 14644 32284
rect 14700 30996 14756 35084
rect 14812 31668 14868 35252
rect 14924 33236 14980 47852
rect 15036 38836 15092 38846
rect 15036 33460 15092 38780
rect 15148 38274 15204 52892
rect 17612 52164 17668 52174
rect 16380 48132 16436 48142
rect 16380 47068 16436 48076
rect 17612 47908 17668 52108
rect 17612 47842 17668 47852
rect 16156 47012 16436 47068
rect 16044 41188 16100 41198
rect 15484 40514 15540 40526
rect 15484 40462 15486 40514
rect 15538 40462 15540 40514
rect 15148 38222 15150 38274
rect 15202 38222 15204 38274
rect 15148 38210 15204 38222
rect 15372 40404 15428 40414
rect 15148 36260 15204 36270
rect 15372 36260 15428 40348
rect 15484 38668 15540 40462
rect 15820 39620 15876 39630
rect 15820 38834 15876 39564
rect 15820 38782 15822 38834
rect 15874 38782 15876 38834
rect 15820 38770 15876 38782
rect 15484 38612 15652 38668
rect 15148 36258 15428 36260
rect 15148 36206 15150 36258
rect 15202 36206 15428 36258
rect 15148 36204 15428 36206
rect 15484 38050 15540 38062
rect 15484 37998 15486 38050
rect 15538 37998 15540 38050
rect 15148 34468 15204 36204
rect 15484 35810 15540 37998
rect 15596 37268 15652 38612
rect 15596 37202 15652 37212
rect 15484 35758 15486 35810
rect 15538 35758 15540 35810
rect 15484 35746 15540 35758
rect 15708 36594 15764 36606
rect 15708 36542 15710 36594
rect 15762 36542 15764 36594
rect 15148 34402 15204 34412
rect 15708 34914 15764 36542
rect 15932 36482 15988 36494
rect 15932 36430 15934 36482
rect 15986 36430 15988 36482
rect 15932 35252 15988 36430
rect 15932 35186 15988 35196
rect 15708 34862 15710 34914
rect 15762 34862 15764 34914
rect 15596 33572 15652 33582
rect 15036 33404 15204 33460
rect 15036 33236 15092 33246
rect 14924 33234 15092 33236
rect 14924 33182 15038 33234
rect 15090 33182 15092 33234
rect 14924 33180 15092 33182
rect 15036 33170 15092 33180
rect 15148 33012 15204 33404
rect 14812 31602 14868 31612
rect 14924 32956 15204 33012
rect 14700 30940 14868 30996
rect 14700 30772 14756 30782
rect 14700 30678 14756 30716
rect 14588 28578 14644 28588
rect 14700 30098 14756 30110
rect 14700 30046 14702 30098
rect 14754 30046 14756 30098
rect 14476 27858 14532 27870
rect 14476 27806 14478 27858
rect 14530 27806 14532 27858
rect 14476 27412 14532 27806
rect 14588 27636 14644 27646
rect 14588 27542 14644 27580
rect 14476 27346 14532 27356
rect 14700 27300 14756 30046
rect 14700 27234 14756 27244
rect 14812 26908 14868 30940
rect 14924 29988 14980 32956
rect 15148 32562 15204 32574
rect 15148 32510 15150 32562
rect 15202 32510 15204 32562
rect 15036 31780 15092 31790
rect 15036 31686 15092 31724
rect 15148 31444 15204 32510
rect 15596 32450 15652 33516
rect 15596 32398 15598 32450
rect 15650 32398 15652 32450
rect 15596 32386 15652 32398
rect 15148 31378 15204 31388
rect 15372 32004 15428 32014
rect 14924 29932 15092 29988
rect 14924 28644 14980 28654
rect 14924 28550 14980 28588
rect 14700 26852 14868 26908
rect 14588 26516 14644 26526
rect 14588 26402 14644 26460
rect 14588 26350 14590 26402
rect 14642 26350 14644 26402
rect 14588 26338 14644 26350
rect 14700 26404 14756 26852
rect 14700 26338 14756 26348
rect 14924 25732 14980 25742
rect 14700 25506 14756 25518
rect 14700 25454 14702 25506
rect 14754 25454 14756 25506
rect 14252 25282 14308 25294
rect 14252 25230 14254 25282
rect 14306 25230 14308 25282
rect 14252 24724 14308 25230
rect 14364 24724 14420 24734
rect 14252 24722 14420 24724
rect 14252 24670 14366 24722
rect 14418 24670 14420 24722
rect 14252 24668 14420 24670
rect 14364 24658 14420 24668
rect 14700 24612 14756 25454
rect 14700 24546 14756 24556
rect 14924 24722 14980 25676
rect 14924 24670 14926 24722
rect 14978 24670 14980 24722
rect 14140 24322 14196 24332
rect 13804 24162 14084 24164
rect 13804 24110 13806 24162
rect 13858 24110 14084 24162
rect 13804 24108 14084 24110
rect 13804 24098 13860 24108
rect 14140 24052 14196 24062
rect 14028 23996 14140 24052
rect 13692 23938 13972 23940
rect 13692 23886 13694 23938
rect 13746 23886 13972 23938
rect 13692 23884 13972 23886
rect 13692 23874 13748 23884
rect 13804 23380 13860 23390
rect 13692 23154 13748 23166
rect 13692 23102 13694 23154
rect 13746 23102 13748 23154
rect 13692 22372 13748 23102
rect 13804 23042 13860 23324
rect 13804 22990 13806 23042
rect 13858 22990 13860 23042
rect 13804 22978 13860 22990
rect 13916 22596 13972 23884
rect 13580 21924 13636 21934
rect 13580 21586 13636 21868
rect 13580 21534 13582 21586
rect 13634 21534 13636 21586
rect 13580 21522 13636 21534
rect 13692 21364 13748 22316
rect 13804 22540 13972 22596
rect 13804 21476 13860 22540
rect 13916 22370 13972 22382
rect 13916 22318 13918 22370
rect 13970 22318 13972 22370
rect 13916 22260 13972 22318
rect 13916 22194 13972 22204
rect 13804 21420 13972 21476
rect 13692 21298 13748 21308
rect 13916 21140 13972 21420
rect 13692 21084 13972 21140
rect 13468 20188 13636 20244
rect 13356 19730 13412 19740
rect 13468 20020 13524 20030
rect 13468 19906 13524 19964
rect 13468 19854 13470 19906
rect 13522 19854 13524 19906
rect 12908 19236 12964 19246
rect 13356 19236 13412 19246
rect 13468 19236 13524 19854
rect 12908 19234 13076 19236
rect 12908 19182 12910 19234
rect 12962 19182 13076 19234
rect 12908 19180 13076 19182
rect 12908 19170 12964 19180
rect 12796 18956 12964 19012
rect 12796 18788 12852 18798
rect 12796 17106 12852 18732
rect 12796 17054 12798 17106
rect 12850 17054 12852 17106
rect 12796 17042 12852 17054
rect 12908 16770 12964 18956
rect 12908 16718 12910 16770
rect 12962 16718 12964 16770
rect 12908 16706 12964 16718
rect 13020 17220 13076 19180
rect 13356 19234 13524 19236
rect 13356 19182 13358 19234
rect 13410 19182 13524 19234
rect 13356 19180 13524 19182
rect 13356 19170 13412 19180
rect 13020 16098 13076 17164
rect 13244 19124 13300 19134
rect 13244 17666 13300 19068
rect 13244 17614 13246 17666
rect 13298 17614 13300 17666
rect 13132 17108 13188 17118
rect 13132 17014 13188 17052
rect 13020 16046 13022 16098
rect 13074 16046 13076 16098
rect 13020 16034 13076 16046
rect 13132 16884 13188 16894
rect 13132 13746 13188 16828
rect 13132 13694 13134 13746
rect 13186 13694 13188 13746
rect 13132 13682 13188 13694
rect 13244 14532 13300 17614
rect 13356 18900 13412 18910
rect 13356 17332 13412 18844
rect 13468 18226 13524 18238
rect 13468 18174 13470 18226
rect 13522 18174 13524 18226
rect 13468 17668 13524 18174
rect 13468 17602 13524 17612
rect 13356 16884 13412 17276
rect 13356 16818 13412 16828
rect 13580 16436 13636 20188
rect 13692 19908 13748 21084
rect 13804 20916 13860 20926
rect 13804 20802 13860 20860
rect 13804 20750 13806 20802
rect 13858 20750 13860 20802
rect 13804 20738 13860 20750
rect 13916 20914 13972 20926
rect 13916 20862 13918 20914
rect 13970 20862 13972 20914
rect 13804 19908 13860 19918
rect 13692 19906 13860 19908
rect 13692 19854 13806 19906
rect 13858 19854 13860 19906
rect 13692 19852 13860 19854
rect 13692 18452 13748 19852
rect 13804 19842 13860 19852
rect 13916 19572 13972 20862
rect 13916 19506 13972 19516
rect 13804 19348 13860 19358
rect 13804 19234 13860 19292
rect 13804 19182 13806 19234
rect 13858 19182 13860 19234
rect 13804 19170 13860 19182
rect 13916 19346 13972 19358
rect 13916 19294 13918 19346
rect 13970 19294 13972 19346
rect 13804 18676 13860 18686
rect 13804 18582 13860 18620
rect 13692 18386 13748 18396
rect 13804 18228 13860 18238
rect 13692 17668 13748 17678
rect 13692 16884 13748 17612
rect 13804 17666 13860 18172
rect 13804 17614 13806 17666
rect 13858 17614 13860 17666
rect 13804 17602 13860 17614
rect 13916 17108 13972 19294
rect 14028 18228 14084 23996
rect 14140 23986 14196 23996
rect 14252 23940 14308 23950
rect 14252 23846 14308 23884
rect 14924 23938 14980 24670
rect 14924 23886 14926 23938
rect 14978 23886 14980 23938
rect 14700 23716 14756 23726
rect 14140 23492 14196 23502
rect 14140 19348 14196 23436
rect 14364 23154 14420 23166
rect 14364 23102 14366 23154
rect 14418 23102 14420 23154
rect 14364 23044 14420 23102
rect 14252 21252 14308 21262
rect 14252 20916 14308 21196
rect 14252 20850 14308 20860
rect 14140 19124 14196 19292
rect 14140 19058 14196 19068
rect 14252 19796 14308 19806
rect 14028 18162 14084 18172
rect 14140 18564 14196 18574
rect 13916 17042 13972 17052
rect 14028 17666 14084 17678
rect 14028 17614 14030 17666
rect 14082 17614 14084 17666
rect 13804 16884 13860 16894
rect 13692 16882 13860 16884
rect 13692 16830 13806 16882
rect 13858 16830 13860 16882
rect 13692 16828 13860 16830
rect 13804 16818 13860 16828
rect 14028 16884 14084 17614
rect 14028 16790 14084 16828
rect 14140 16660 14196 18508
rect 14252 17106 14308 19740
rect 14364 19460 14420 22988
rect 14700 22482 14756 23660
rect 14700 22430 14702 22482
rect 14754 22430 14756 22482
rect 14700 22418 14756 22430
rect 14812 23156 14868 23166
rect 14476 22260 14532 22270
rect 14476 21586 14532 22204
rect 14476 21534 14478 21586
rect 14530 21534 14532 21586
rect 14476 21522 14532 21534
rect 14812 21924 14868 23100
rect 14700 21364 14756 21374
rect 14476 20804 14532 20814
rect 14476 19572 14532 20748
rect 14588 20802 14644 20814
rect 14588 20750 14590 20802
rect 14642 20750 14644 20802
rect 14588 20468 14644 20750
rect 14588 20402 14644 20412
rect 14700 20018 14756 21308
rect 14700 19966 14702 20018
rect 14754 19966 14756 20018
rect 14700 19954 14756 19966
rect 14812 20804 14868 21868
rect 14924 21476 14980 23886
rect 14924 21028 14980 21420
rect 14924 20962 14980 20972
rect 14924 20804 14980 20814
rect 14812 20802 14980 20804
rect 14812 20750 14926 20802
rect 14978 20750 14980 20802
rect 14812 20748 14980 20750
rect 14476 19516 14644 19572
rect 14364 19346 14420 19404
rect 14364 19294 14366 19346
rect 14418 19294 14420 19346
rect 14364 19282 14420 19294
rect 14364 18452 14420 18462
rect 14364 18338 14420 18396
rect 14588 18452 14644 19516
rect 14588 18386 14644 18396
rect 14700 19236 14756 19246
rect 14364 18286 14366 18338
rect 14418 18286 14420 18338
rect 14364 18274 14420 18286
rect 14588 18228 14644 18238
rect 14252 17054 14254 17106
rect 14306 17054 14308 17106
rect 14252 17042 14308 17054
rect 14364 18004 14420 18014
rect 14364 16882 14420 17948
rect 14476 17892 14532 17902
rect 14476 17798 14532 17836
rect 14588 17668 14644 18172
rect 14364 16830 14366 16882
rect 14418 16830 14420 16882
rect 14364 16818 14420 16830
rect 14476 17612 14644 17668
rect 14700 17666 14756 19180
rect 14700 17614 14702 17666
rect 14754 17614 14756 17666
rect 13580 16370 13636 16380
rect 13692 16604 14196 16660
rect 14364 16660 14420 16670
rect 13580 15876 13636 15886
rect 13580 15148 13636 15820
rect 13692 15314 13748 16604
rect 13692 15262 13694 15314
rect 13746 15262 13748 15314
rect 13692 15250 13748 15262
rect 13804 16436 13860 16446
rect 12796 12964 12852 12974
rect 12796 12870 12852 12908
rect 13244 12404 13300 14476
rect 12796 12348 13300 12404
rect 12796 12290 12852 12348
rect 12796 12238 12798 12290
rect 12850 12238 12852 12290
rect 12796 12226 12852 12238
rect 13132 12178 13188 12190
rect 13132 12126 13134 12178
rect 13186 12126 13188 12178
rect 13020 11396 13076 11406
rect 12684 11394 13076 11396
rect 12684 11342 13022 11394
rect 13074 11342 13076 11394
rect 12684 11340 13076 11342
rect 12124 10782 12126 10834
rect 12178 10782 12180 10834
rect 12124 10770 12180 10782
rect 12124 9828 12180 9838
rect 12012 9826 12180 9828
rect 12012 9774 12126 9826
rect 12178 9774 12180 9826
rect 12012 9772 12180 9774
rect 12124 9762 12180 9772
rect 11340 8482 11620 8484
rect 11340 8430 11342 8482
rect 11394 8430 11620 8482
rect 11340 8428 11620 8430
rect 11676 9380 11732 9390
rect 11340 8418 11396 8428
rect 11564 7588 11620 7598
rect 11676 7588 11732 9324
rect 11564 7586 11732 7588
rect 11564 7534 11566 7586
rect 11618 7534 11732 7586
rect 11564 7532 11732 7534
rect 12124 8932 12180 8942
rect 11564 7522 11620 7532
rect 11004 7422 11006 7474
rect 11058 7422 11060 7474
rect 11004 7410 11060 7422
rect 10668 7364 10724 7374
rect 10668 7270 10724 7308
rect 11452 6020 11508 6030
rect 10108 5124 10164 5134
rect 8652 3332 8820 3388
rect 3804 3164 4068 3174
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 3804 3098 4068 3108
rect 4464 2380 4728 2390
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4464 2314 4728 2324
rect 3804 1596 4068 1606
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 3804 1530 4068 1540
rect 4464 812 4728 822
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4464 746 4728 756
rect 3612 130 3668 140
rect 4732 196 4788 206
rect 4732 112 4788 140
rect 6076 112 6132 3332
rect 7420 3108 7476 3118
rect 7420 112 7476 3052
rect 7980 1428 8036 3332
rect 8764 3108 8820 3332
rect 8764 3042 8820 3052
rect 7980 1362 8036 1372
rect 8764 1652 8820 1662
rect 8764 112 8820 1596
rect 10108 112 10164 5068
rect 11452 112 11508 5964
rect 12124 1652 12180 8876
rect 13020 2996 13076 11340
rect 13132 10500 13188 12126
rect 13132 10434 13188 10444
rect 13132 9828 13188 9838
rect 13132 9734 13188 9772
rect 13244 8036 13300 12348
rect 13356 15090 13412 15102
rect 13356 15038 13358 15090
rect 13410 15038 13412 15090
rect 13356 12404 13412 15038
rect 13356 12338 13412 12348
rect 13468 15092 13636 15148
rect 13244 7970 13300 7980
rect 13468 3388 13524 15092
rect 13804 14756 13860 16380
rect 14364 16324 14420 16604
rect 14476 16436 14532 17612
rect 14588 17108 14644 17118
rect 14588 16658 14644 17052
rect 14588 16606 14590 16658
rect 14642 16606 14644 16658
rect 14588 16594 14644 16606
rect 14476 16380 14644 16436
rect 14364 16268 14532 16324
rect 13916 16212 13972 16222
rect 13916 16098 13972 16156
rect 13916 16046 13918 16098
rect 13970 16046 13972 16098
rect 13916 16034 13972 16046
rect 14364 14756 14420 14766
rect 13804 14754 14420 14756
rect 13804 14702 14366 14754
rect 14418 14702 14420 14754
rect 13804 14700 14420 14702
rect 13580 14084 13636 14094
rect 13580 12628 13636 14028
rect 13692 13636 13748 13646
rect 13804 13636 13860 14700
rect 14364 14690 14420 14700
rect 13916 14418 13972 14430
rect 13916 14366 13918 14418
rect 13970 14366 13972 14418
rect 13916 14308 13972 14366
rect 13916 14242 13972 14252
rect 13692 13634 13860 13636
rect 13692 13582 13694 13634
rect 13746 13582 13860 13634
rect 13692 13580 13860 13582
rect 13692 13570 13748 13580
rect 13580 12180 13636 12572
rect 14140 13300 14196 13310
rect 14476 13300 14532 16268
rect 13580 12178 13972 12180
rect 13580 12126 13582 12178
rect 13634 12126 13972 12178
rect 13580 12124 13972 12126
rect 13580 12114 13636 12124
rect 13804 11956 13860 11966
rect 13580 11954 13860 11956
rect 13580 11902 13806 11954
rect 13858 11902 13860 11954
rect 13580 11900 13860 11902
rect 13580 10610 13636 11900
rect 13804 11890 13860 11900
rect 13580 10558 13582 10610
rect 13634 10558 13636 10610
rect 13580 10546 13636 10558
rect 13916 8820 13972 12124
rect 14140 11620 14196 13244
rect 14364 13244 14532 13300
rect 14588 13300 14644 16380
rect 14700 14084 14756 17614
rect 14812 15876 14868 20748
rect 14924 20738 14980 20748
rect 15036 20130 15092 29932
rect 15260 29202 15316 29214
rect 15260 29150 15262 29202
rect 15314 29150 15316 29202
rect 15148 27860 15204 27870
rect 15148 27298 15204 27804
rect 15260 27858 15316 29150
rect 15260 27806 15262 27858
rect 15314 27806 15316 27858
rect 15260 27794 15316 27806
rect 15148 27246 15150 27298
rect 15202 27246 15204 27298
rect 15148 27234 15204 27246
rect 15372 26908 15428 31948
rect 15708 31780 15764 34862
rect 15708 31714 15764 31724
rect 15932 31444 15988 31454
rect 15820 31220 15876 31230
rect 15820 31126 15876 31164
rect 15708 30212 15764 30222
rect 15932 30212 15988 31388
rect 15708 30210 15876 30212
rect 15708 30158 15710 30210
rect 15762 30158 15876 30210
rect 15708 30156 15876 30158
rect 15708 30146 15764 30156
rect 15596 28644 15652 28654
rect 15596 27860 15652 28588
rect 15820 28532 15876 30156
rect 15932 29538 15988 30156
rect 15932 29486 15934 29538
rect 15986 29486 15988 29538
rect 15932 29474 15988 29486
rect 15820 28466 15876 28476
rect 15932 28642 15988 28654
rect 15932 28590 15934 28642
rect 15986 28590 15988 28642
rect 15260 26852 15428 26908
rect 15484 27858 15652 27860
rect 15484 27806 15598 27858
rect 15650 27806 15652 27858
rect 15484 27804 15652 27806
rect 15260 25618 15316 26852
rect 15484 26740 15540 27804
rect 15596 27794 15652 27804
rect 15596 27636 15652 27646
rect 15596 27298 15652 27580
rect 15596 27246 15598 27298
rect 15650 27246 15652 27298
rect 15596 27234 15652 27246
rect 15932 26908 15988 28590
rect 15260 25566 15262 25618
rect 15314 25566 15316 25618
rect 15260 25554 15316 25566
rect 15372 26684 15540 26740
rect 15708 26852 15988 26908
rect 15148 22596 15204 22606
rect 15148 22502 15204 22540
rect 15260 22372 15316 22382
rect 15036 20078 15038 20130
rect 15090 20078 15092 20130
rect 15036 20066 15092 20078
rect 15148 22370 15316 22372
rect 15148 22318 15262 22370
rect 15314 22318 15316 22370
rect 15148 22316 15316 22318
rect 15148 21588 15204 22316
rect 15260 22306 15316 22316
rect 15148 20132 15204 21532
rect 15260 21476 15316 21486
rect 15260 21382 15316 21420
rect 14924 19348 14980 19358
rect 14924 19234 14980 19292
rect 14924 19182 14926 19234
rect 14978 19182 14980 19234
rect 14924 17668 14980 19182
rect 15148 18676 15204 20076
rect 15372 19460 15428 26684
rect 15484 23492 15540 23502
rect 15484 20916 15540 23436
rect 15708 23156 15764 26852
rect 16044 26628 16100 41132
rect 16156 30322 16212 47012
rect 17836 45668 17892 45678
rect 17052 44324 17108 44334
rect 16268 41972 16324 41982
rect 16268 41970 16548 41972
rect 16268 41918 16270 41970
rect 16322 41918 16548 41970
rect 16268 41916 16548 41918
rect 16268 41906 16324 41916
rect 16492 37378 16548 41916
rect 16716 39620 16772 39630
rect 16716 39526 16772 39564
rect 16492 37326 16494 37378
rect 16546 37326 16548 37378
rect 16492 37314 16548 37326
rect 16716 38050 16772 38062
rect 16716 37998 16718 38050
rect 16770 37998 16772 38050
rect 16604 37154 16660 37166
rect 16604 37102 16606 37154
rect 16658 37102 16660 37154
rect 16604 34132 16660 37102
rect 16716 34242 16772 37998
rect 16828 35252 16884 35262
rect 16828 35138 16884 35196
rect 16828 35086 16830 35138
rect 16882 35086 16884 35138
rect 16828 35074 16884 35086
rect 16716 34190 16718 34242
rect 16770 34190 16772 34242
rect 16716 34178 16772 34190
rect 16604 34066 16660 34076
rect 16940 33236 16996 33246
rect 17052 33236 17108 44268
rect 17724 40404 17780 40414
rect 17724 40310 17780 40348
rect 17276 40180 17332 40190
rect 16940 33234 17108 33236
rect 16940 33182 16942 33234
rect 16994 33182 17108 33234
rect 16940 33180 17108 33182
rect 17164 37268 17220 37278
rect 16940 33170 16996 33180
rect 17164 32676 17220 37212
rect 16828 32338 16884 32350
rect 16828 32286 16830 32338
rect 16882 32286 16884 32338
rect 16828 31892 16884 32286
rect 16828 31826 16884 31836
rect 16156 30270 16158 30322
rect 16210 30270 16212 30322
rect 16156 30258 16212 30270
rect 16268 31780 16324 31790
rect 16156 28420 16212 28430
rect 16156 27186 16212 28364
rect 16156 27134 16158 27186
rect 16210 27134 16212 27186
rect 16156 27122 16212 27134
rect 16044 26562 16100 26572
rect 15708 23090 15764 23100
rect 15932 24722 15988 24734
rect 15932 24670 15934 24722
rect 15986 24670 15988 24722
rect 15932 23938 15988 24670
rect 15932 23886 15934 23938
rect 15986 23886 15988 23938
rect 15932 23154 15988 23886
rect 15932 23102 15934 23154
rect 15986 23102 15988 23154
rect 15820 22372 15876 22382
rect 15820 22278 15876 22316
rect 15820 21588 15876 21598
rect 15820 21494 15876 21532
rect 15708 21364 15764 21374
rect 15708 21270 15764 21308
rect 15484 20860 15652 20916
rect 15596 20132 15652 20860
rect 15596 20066 15652 20076
rect 15820 20804 15876 20814
rect 15484 20020 15540 20030
rect 15484 19926 15540 19964
rect 15820 20018 15876 20748
rect 15932 20802 15988 23102
rect 16156 22258 16212 22270
rect 16156 22206 16158 22258
rect 16210 22206 16212 22258
rect 16156 21364 16212 22206
rect 16268 21924 16324 31724
rect 17052 31778 17108 31790
rect 17052 31726 17054 31778
rect 17106 31726 17108 31778
rect 16716 31668 16772 31678
rect 16716 31574 16772 31612
rect 17052 31220 17108 31726
rect 17164 31780 17220 32620
rect 17276 32674 17332 40124
rect 17836 38668 17892 45612
rect 17724 38612 17892 38668
rect 17948 44212 18004 44222
rect 17500 37940 17556 37950
rect 17500 37846 17556 37884
rect 17388 36260 17444 36270
rect 17388 36166 17444 36204
rect 17724 33572 17780 38612
rect 17724 33506 17780 33516
rect 17836 36482 17892 36494
rect 17836 36430 17838 36482
rect 17890 36430 17892 36482
rect 17388 33348 17444 33358
rect 17388 33346 17780 33348
rect 17388 33294 17390 33346
rect 17442 33294 17780 33346
rect 17388 33292 17780 33294
rect 17388 33282 17444 33292
rect 17276 32622 17278 32674
rect 17330 32622 17332 32674
rect 17276 32610 17332 32622
rect 17612 32340 17668 32350
rect 17500 31780 17556 31790
rect 17164 31778 17556 31780
rect 17164 31726 17502 31778
rect 17554 31726 17556 31778
rect 17164 31724 17556 31726
rect 17052 31154 17108 31164
rect 17164 30996 17220 31006
rect 17164 30994 17444 30996
rect 17164 30942 17166 30994
rect 17218 30942 17444 30994
rect 17164 30940 17444 30942
rect 17164 30930 17220 30940
rect 16716 30882 16772 30894
rect 16716 30830 16718 30882
rect 16770 30830 16772 30882
rect 16716 30660 16772 30830
rect 16380 29202 16436 29214
rect 16380 29150 16382 29202
rect 16434 29150 16436 29202
rect 16380 28532 16436 29150
rect 16380 28466 16436 28476
rect 16716 28308 16772 30604
rect 17276 30324 17332 30334
rect 17164 30322 17332 30324
rect 17164 30270 17278 30322
rect 17330 30270 17332 30322
rect 17164 30268 17332 30270
rect 16828 30212 16884 30222
rect 16828 30118 16884 30156
rect 16380 28252 16772 28308
rect 16940 28532 16996 28542
rect 16380 23492 16436 28252
rect 16604 27858 16660 27870
rect 16604 27806 16606 27858
rect 16658 27806 16660 27858
rect 16492 27076 16548 27086
rect 16492 26402 16548 27020
rect 16492 26350 16494 26402
rect 16546 26350 16548 26402
rect 16492 26338 16548 26350
rect 16604 24724 16660 27806
rect 16940 26068 16996 28476
rect 17164 26852 17220 30268
rect 17276 30258 17332 30268
rect 17388 29652 17444 30940
rect 17500 30994 17556 31724
rect 17500 30942 17502 30994
rect 17554 30942 17556 30994
rect 17500 30930 17556 30942
rect 17500 29652 17556 29662
rect 17388 29650 17556 29652
rect 17388 29598 17502 29650
rect 17554 29598 17556 29650
rect 17388 29596 17556 29598
rect 17500 29586 17556 29596
rect 17612 29428 17668 32284
rect 17724 32002 17780 33292
rect 17836 33346 17892 36430
rect 17948 35028 18004 44156
rect 18060 40292 18116 55132
rect 18284 53172 18340 55246
rect 18284 53106 18340 53116
rect 18956 55298 19348 55300
rect 18956 55246 19294 55298
rect 19346 55246 19348 55298
rect 18956 55244 19348 55246
rect 18508 52724 18564 52734
rect 18508 47124 18564 52668
rect 18060 40226 18116 40236
rect 18172 47068 18564 47124
rect 18172 38668 18228 47068
rect 18060 38612 18228 38668
rect 18284 46900 18340 46910
rect 18060 35308 18116 38612
rect 18284 36708 18340 46844
rect 18396 41858 18452 41870
rect 18396 41806 18398 41858
rect 18450 41806 18452 41858
rect 18396 40402 18452 41806
rect 18396 40350 18398 40402
rect 18450 40350 18452 40402
rect 18396 40338 18452 40350
rect 18732 39508 18788 39518
rect 18508 39506 18788 39508
rect 18508 39454 18734 39506
rect 18786 39454 18788 39506
rect 18508 39452 18788 39454
rect 18508 38668 18564 39452
rect 18732 39442 18788 39452
rect 18284 36642 18340 36652
rect 18396 38612 18564 38668
rect 18620 38722 18676 38734
rect 18620 38670 18622 38722
rect 18674 38670 18676 38722
rect 18284 36482 18340 36494
rect 18284 36430 18286 36482
rect 18338 36430 18340 36482
rect 18284 36260 18340 36430
rect 18060 35252 18228 35308
rect 17948 34934 18004 34972
rect 17836 33294 17838 33346
rect 17890 33294 17892 33346
rect 17836 33282 17892 33294
rect 17948 33236 18004 33246
rect 17948 33142 18004 33180
rect 17724 31950 17726 32002
rect 17778 31950 17780 32002
rect 17724 31938 17780 31950
rect 17836 32338 17892 32350
rect 17836 32286 17838 32338
rect 17890 32286 17892 32338
rect 17724 30884 17780 30894
rect 17836 30884 17892 32286
rect 18172 32116 18228 35252
rect 18284 34804 18340 36204
rect 18396 35698 18452 38612
rect 18620 37266 18676 38670
rect 18620 37214 18622 37266
rect 18674 37214 18676 37266
rect 18620 37202 18676 37214
rect 18844 37828 18900 37838
rect 18844 36594 18900 37772
rect 18844 36542 18846 36594
rect 18898 36542 18900 36594
rect 18844 36530 18900 36542
rect 18396 35646 18398 35698
rect 18450 35646 18452 35698
rect 18396 35634 18452 35646
rect 18956 35140 19012 55244
rect 19292 55234 19348 55244
rect 19404 54628 19460 54638
rect 19404 54534 19460 54572
rect 19068 54514 19124 54526
rect 19068 54462 19070 54514
rect 19122 54462 19124 54514
rect 19068 38668 19124 54462
rect 19516 53284 19572 55918
rect 20188 55412 20244 56030
rect 20188 55346 20244 55356
rect 21084 55972 21140 55982
rect 20076 55298 20132 55310
rect 20076 55246 20078 55298
rect 20130 55246 20132 55298
rect 19516 53218 19572 53228
rect 19964 53618 20020 53630
rect 19964 53566 19966 53618
rect 20018 53566 20020 53618
rect 19964 52276 20020 53566
rect 19964 52210 20020 52220
rect 20076 50428 20132 55246
rect 20524 55300 20580 55310
rect 20860 55300 20916 55310
rect 20524 55206 20580 55244
rect 20748 55298 20916 55300
rect 20748 55246 20862 55298
rect 20914 55246 20916 55298
rect 20748 55244 20916 55246
rect 20636 54292 20692 54302
rect 20636 54198 20692 54236
rect 20524 53732 20580 53742
rect 20524 53638 20580 53676
rect 20748 50428 20804 55244
rect 20860 55234 20916 55244
rect 21084 54626 21140 55916
rect 21980 55972 22036 55982
rect 21644 55860 21700 55870
rect 21644 55410 21700 55804
rect 21644 55358 21646 55410
rect 21698 55358 21700 55410
rect 21644 55346 21700 55358
rect 21084 54574 21086 54626
rect 21138 54574 21140 54626
rect 21084 54562 21140 54574
rect 21532 54402 21588 54414
rect 21532 54350 21534 54402
rect 21586 54350 21588 54402
rect 19964 50372 20132 50428
rect 20300 50372 20804 50428
rect 20860 53730 20916 53742
rect 20860 53678 20862 53730
rect 20914 53678 20916 53730
rect 20860 50484 20916 53678
rect 21308 53620 21364 53630
rect 21308 53526 21364 53564
rect 21420 52948 21476 52958
rect 21420 52854 21476 52892
rect 20860 50418 20916 50428
rect 21084 51156 21140 51166
rect 19628 40292 19684 40302
rect 19068 38612 19348 38668
rect 18844 35084 19012 35140
rect 18396 34804 18452 34814
rect 18284 34802 18452 34804
rect 18284 34750 18398 34802
rect 18450 34750 18452 34802
rect 18284 34748 18452 34750
rect 18284 33012 18340 34748
rect 18396 34738 18452 34748
rect 18508 34132 18564 34142
rect 18508 34038 18564 34076
rect 18396 33572 18452 33582
rect 18452 33516 18564 33572
rect 18396 33478 18452 33516
rect 18284 32956 18452 33012
rect 18284 32788 18340 32798
rect 18284 32694 18340 32732
rect 18396 32564 18452 32956
rect 17724 30882 17892 30884
rect 17724 30830 17726 30882
rect 17778 30830 17892 30882
rect 17724 30828 17892 30830
rect 18060 32060 18228 32116
rect 18284 32508 18452 32564
rect 17724 30818 17780 30828
rect 16940 26066 17108 26068
rect 16940 26014 16942 26066
rect 16994 26014 17108 26066
rect 16940 26012 17108 26014
rect 16940 26002 16996 26012
rect 16380 23426 16436 23436
rect 16492 24668 16660 24724
rect 16940 25284 16996 25294
rect 16380 22930 16436 22942
rect 16380 22878 16382 22930
rect 16434 22878 16436 22930
rect 16380 22596 16436 22878
rect 16380 22530 16436 22540
rect 16268 21858 16324 21868
rect 16380 21588 16436 21598
rect 16380 21494 16436 21532
rect 16156 21298 16212 21308
rect 16492 21140 16548 24668
rect 16604 24500 16660 24510
rect 16604 24406 16660 24444
rect 16828 23716 16884 23726
rect 16828 23622 16884 23660
rect 16940 23266 16996 25228
rect 16940 23214 16942 23266
rect 16994 23214 16996 23266
rect 16940 23202 16996 23214
rect 17052 22708 17108 26012
rect 17164 23828 17220 26796
rect 17164 23762 17220 23772
rect 17276 29372 17668 29428
rect 17836 30660 17892 30670
rect 17052 22642 17108 22652
rect 16828 22370 16884 22382
rect 16828 22318 16830 22370
rect 16882 22318 16884 22370
rect 16716 22148 16772 22158
rect 15932 20750 15934 20802
rect 15986 20750 15988 20802
rect 15932 20356 15988 20750
rect 16156 21084 16548 21140
rect 16604 22146 16772 22148
rect 16604 22094 16718 22146
rect 16770 22094 16772 22146
rect 16604 22092 16772 22094
rect 15932 20290 15988 20300
rect 16044 20580 16100 20590
rect 16044 20242 16100 20524
rect 16044 20190 16046 20242
rect 16098 20190 16100 20242
rect 16044 20178 16100 20190
rect 15820 19966 15822 20018
rect 15874 19966 15876 20018
rect 15820 19954 15876 19966
rect 15596 19796 15652 19806
rect 15596 19702 15652 19740
rect 15372 19394 15428 19404
rect 16156 19348 16212 21084
rect 16268 20468 16324 20478
rect 16268 20020 16324 20412
rect 16604 20020 16660 22092
rect 16716 22082 16772 22092
rect 16828 22148 16884 22318
rect 16716 21474 16772 21486
rect 16716 21422 16718 21474
rect 16770 21422 16772 21474
rect 16716 21364 16772 21422
rect 16716 21298 16772 21308
rect 16716 20804 16772 20842
rect 16716 20738 16772 20748
rect 16716 20580 16772 20590
rect 16716 20486 16772 20524
rect 16268 20018 16436 20020
rect 16268 19966 16270 20018
rect 16322 19966 16436 20018
rect 16268 19964 16436 19966
rect 16268 19954 16324 19964
rect 16156 19282 16212 19292
rect 15148 18610 15204 18620
rect 15708 19236 15764 19246
rect 14924 17602 14980 17612
rect 15036 18452 15092 18462
rect 15036 17668 15092 18396
rect 15596 18450 15652 18462
rect 15596 18398 15598 18450
rect 15650 18398 15652 18450
rect 15260 18338 15316 18350
rect 15260 18286 15262 18338
rect 15314 18286 15316 18338
rect 15148 18226 15204 18238
rect 15148 18174 15150 18226
rect 15202 18174 15204 18226
rect 15148 18004 15204 18174
rect 15260 18116 15316 18286
rect 15260 18050 15316 18060
rect 15148 17938 15204 17948
rect 15036 17666 15316 17668
rect 15036 17614 15038 17666
rect 15090 17614 15316 17666
rect 15036 17612 15316 17614
rect 15036 17602 15092 17612
rect 14924 17220 14980 17230
rect 14924 16996 14980 17164
rect 14924 16994 15092 16996
rect 14924 16942 14926 16994
rect 14978 16942 15092 16994
rect 14924 16940 15092 16942
rect 14924 16930 14980 16940
rect 14812 15810 14868 15820
rect 14924 15204 14980 15242
rect 14924 15138 14980 15148
rect 15036 15092 15092 16940
rect 15260 16882 15316 17612
rect 15484 17556 15540 17566
rect 15260 16830 15262 16882
rect 15314 16830 15316 16882
rect 15260 16818 15316 16830
rect 15372 17554 15540 17556
rect 15372 17502 15486 17554
rect 15538 17502 15540 17554
rect 15372 17500 15540 17502
rect 15372 16660 15428 17500
rect 15484 17490 15540 17500
rect 15596 17108 15652 18398
rect 15596 17042 15652 17052
rect 15708 16884 15764 19180
rect 16044 19234 16100 19246
rect 16044 19182 16046 19234
rect 16098 19182 16100 19234
rect 16044 19124 16100 19182
rect 16044 19058 16100 19068
rect 15820 18676 15876 18686
rect 15820 18582 15876 18620
rect 16044 18564 16100 18574
rect 15932 18562 16100 18564
rect 15932 18510 16046 18562
rect 16098 18510 16100 18562
rect 15932 18508 16100 18510
rect 15932 18116 15988 18508
rect 16044 18498 16100 18508
rect 16268 18564 16324 18574
rect 16268 18470 16324 18508
rect 15932 17668 15988 18060
rect 16044 18228 16100 18238
rect 16044 17890 16100 18172
rect 16044 17838 16046 17890
rect 16098 17838 16100 17890
rect 16044 17826 16100 17838
rect 16268 18226 16324 18238
rect 16268 18174 16270 18226
rect 16322 18174 16324 18226
rect 15932 17612 16100 17668
rect 15820 17444 15876 17454
rect 15820 17442 15988 17444
rect 15820 17390 15822 17442
rect 15874 17390 15988 17442
rect 15820 17388 15988 17390
rect 15820 17378 15876 17388
rect 15708 16882 15876 16884
rect 15708 16830 15710 16882
rect 15762 16830 15876 16882
rect 15708 16828 15876 16830
rect 15708 16818 15764 16828
rect 15372 16594 15428 16604
rect 15260 16548 15316 16558
rect 15260 16212 15316 16492
rect 15260 16118 15316 16156
rect 15708 16212 15764 16222
rect 15708 16118 15764 16156
rect 15372 15988 15428 15998
rect 15372 15874 15428 15932
rect 15372 15822 15374 15874
rect 15426 15822 15428 15874
rect 15372 15764 15428 15822
rect 15372 15698 15428 15708
rect 15708 15988 15764 15998
rect 15148 15652 15204 15662
rect 15148 15314 15204 15596
rect 15260 15428 15316 15438
rect 15260 15334 15316 15372
rect 15148 15262 15150 15314
rect 15202 15262 15204 15314
rect 15148 15250 15204 15262
rect 15484 15204 15540 15214
rect 15372 15148 15484 15204
rect 15036 15036 15204 15092
rect 14700 14018 14756 14028
rect 15036 14756 15092 14766
rect 14812 13524 14868 13534
rect 14252 12066 14308 12078
rect 14252 12014 14254 12066
rect 14306 12014 14308 12066
rect 14252 11844 14308 12014
rect 14252 11778 14308 11788
rect 14140 11564 14308 11620
rect 14252 11284 14308 11564
rect 14364 11396 14420 13244
rect 14588 13234 14644 13244
rect 14700 13522 14868 13524
rect 14700 13470 14814 13522
rect 14866 13470 14868 13522
rect 14700 13468 14868 13470
rect 14476 13074 14532 13086
rect 14476 13022 14478 13074
rect 14530 13022 14532 13074
rect 14476 11956 14532 13022
rect 14476 11890 14532 11900
rect 14700 11506 14756 13468
rect 14812 13458 14868 13468
rect 14924 13524 14980 13534
rect 14812 13076 14868 13086
rect 14924 13076 14980 13468
rect 14812 13074 14980 13076
rect 14812 13022 14814 13074
rect 14866 13022 14980 13074
rect 14812 13020 14980 13022
rect 14812 13010 14868 13020
rect 15036 12628 15092 14700
rect 14700 11454 14702 11506
rect 14754 11454 14756 11506
rect 14700 11442 14756 11454
rect 14924 12572 15092 12628
rect 15148 14532 15204 15036
rect 15372 15090 15428 15148
rect 15484 15138 15540 15148
rect 15372 15038 15374 15090
rect 15426 15038 15428 15090
rect 15372 15026 15428 15038
rect 15484 14980 15540 14990
rect 14364 11340 14644 11396
rect 14252 11228 14532 11284
rect 14140 11172 14196 11182
rect 14140 11170 14420 11172
rect 14140 11118 14142 11170
rect 14194 11118 14420 11170
rect 14140 11116 14420 11118
rect 14140 11106 14196 11116
rect 14028 10836 14084 10846
rect 14028 10722 14084 10780
rect 14028 10670 14030 10722
rect 14082 10670 14084 10722
rect 14028 10658 14084 10670
rect 14364 10610 14420 11116
rect 14476 11170 14532 11228
rect 14476 11118 14478 11170
rect 14530 11118 14532 11170
rect 14476 11106 14532 11118
rect 14364 10558 14366 10610
rect 14418 10558 14420 10610
rect 14364 10546 14420 10558
rect 13916 8754 13972 8764
rect 14588 4900 14644 11340
rect 14924 10722 14980 12572
rect 15036 12178 15092 12190
rect 15036 12126 15038 12178
rect 15090 12126 15092 12178
rect 15036 12068 15092 12126
rect 15148 12180 15204 14476
rect 15260 14868 15316 14878
rect 15260 13634 15316 14812
rect 15484 14754 15540 14924
rect 15708 14868 15764 15932
rect 15820 15314 15876 16828
rect 15932 16770 15988 17388
rect 16044 16996 16100 17612
rect 16156 17556 16212 17566
rect 16268 17556 16324 18174
rect 16156 17554 16324 17556
rect 16156 17502 16158 17554
rect 16210 17502 16324 17554
rect 16156 17500 16324 17502
rect 16156 17490 16212 17500
rect 16044 16930 16100 16940
rect 16156 17108 16212 17118
rect 15932 16718 15934 16770
rect 15986 16718 15988 16770
rect 15932 16706 15988 16718
rect 15932 16098 15988 16110
rect 15932 16046 15934 16098
rect 15986 16046 15988 16098
rect 15932 15428 15988 16046
rect 16156 15988 16212 17052
rect 16380 16884 16436 19964
rect 16604 19954 16660 19964
rect 16828 19908 16884 22092
rect 17164 21476 17220 21486
rect 17164 21382 17220 21420
rect 17052 20916 17108 20926
rect 17052 20580 17108 20860
rect 17052 20486 17108 20524
rect 16828 19852 17108 19908
rect 16716 19572 16772 19582
rect 16604 19460 16660 19470
rect 16492 18228 16548 18238
rect 16492 18134 16548 18172
rect 16380 16790 16436 16828
rect 16156 15922 16212 15932
rect 16268 16098 16324 16110
rect 16268 16046 16270 16098
rect 16322 16046 16324 16098
rect 16044 15876 16100 15886
rect 16044 15782 16100 15820
rect 15932 15362 15988 15372
rect 15820 15262 15822 15314
rect 15874 15262 15876 15314
rect 15820 14980 15876 15262
rect 16044 15316 16100 15326
rect 16044 15222 16100 15260
rect 15932 15202 15988 15214
rect 15932 15150 15934 15202
rect 15986 15150 15988 15202
rect 15932 15148 15988 15150
rect 15932 15092 16212 15148
rect 15820 14924 16100 14980
rect 15708 14802 15764 14812
rect 16044 14868 16100 14924
rect 16044 14802 16100 14812
rect 15484 14702 15486 14754
rect 15538 14702 15540 14754
rect 15484 14690 15540 14702
rect 15932 14644 15988 14654
rect 15932 14550 15988 14588
rect 16044 14642 16100 14654
rect 16044 14590 16046 14642
rect 16098 14590 16100 14642
rect 16044 14532 16100 14590
rect 16044 14466 16100 14476
rect 16156 14308 16212 15092
rect 16268 14754 16324 16046
rect 16604 16100 16660 19404
rect 16716 19346 16772 19516
rect 16716 19294 16718 19346
rect 16770 19294 16772 19346
rect 16716 19282 16772 19294
rect 16940 19346 16996 19358
rect 16940 19294 16942 19346
rect 16994 19294 16996 19346
rect 16716 19124 16772 19134
rect 16716 16884 16772 19068
rect 16828 19122 16884 19134
rect 16828 19070 16830 19122
rect 16882 19070 16884 19122
rect 16828 18676 16884 19070
rect 16828 18610 16884 18620
rect 16940 18452 16996 19294
rect 17052 18676 17108 19852
rect 17052 18610 17108 18620
rect 16940 18386 16996 18396
rect 16940 18226 16996 18238
rect 16940 18174 16942 18226
rect 16994 18174 16996 18226
rect 16940 17892 16996 18174
rect 17052 18228 17108 18238
rect 17052 18134 17108 18172
rect 17164 18226 17220 18238
rect 17164 18174 17166 18226
rect 17218 18174 17220 18226
rect 17164 18004 17220 18174
rect 17276 18004 17332 29372
rect 17500 27972 17556 27982
rect 17500 27878 17556 27916
rect 17724 27972 17780 27982
rect 17388 27748 17444 27758
rect 17388 23156 17444 27692
rect 17724 27076 17780 27916
rect 17724 26982 17780 27020
rect 17836 27746 17892 30604
rect 17836 27694 17838 27746
rect 17890 27694 17892 27746
rect 17500 25732 17556 25742
rect 17500 25618 17556 25676
rect 17500 25566 17502 25618
rect 17554 25566 17556 25618
rect 17500 23268 17556 25566
rect 17724 24498 17780 24510
rect 17724 24446 17726 24498
rect 17778 24446 17780 24498
rect 17724 24388 17780 24446
rect 17724 24322 17780 24332
rect 17500 23212 17780 23268
rect 17388 23100 17556 23156
rect 17388 22930 17444 22942
rect 17388 22878 17390 22930
rect 17442 22878 17444 22930
rect 17388 22372 17444 22878
rect 17388 22306 17444 22316
rect 17388 22146 17444 22158
rect 17388 22094 17390 22146
rect 17442 22094 17444 22146
rect 17388 20804 17444 22094
rect 17388 20738 17444 20748
rect 17388 18228 17444 18238
rect 17388 18134 17444 18172
rect 17276 17948 17444 18004
rect 17164 17938 17220 17948
rect 16940 17826 16996 17836
rect 16716 16548 16772 16828
rect 16940 17668 16996 17678
rect 16940 17108 16996 17612
rect 16940 16882 16996 17052
rect 16940 16830 16942 16882
rect 16994 16830 16996 16882
rect 16940 16818 16996 16830
rect 16716 16482 16772 16492
rect 16604 16034 16660 16044
rect 16828 15876 16884 15886
rect 16716 15874 16884 15876
rect 16716 15822 16830 15874
rect 16882 15822 16884 15874
rect 16716 15820 16884 15822
rect 16492 15428 16548 15438
rect 16492 15334 16548 15372
rect 16716 15204 16772 15820
rect 16828 15810 16884 15820
rect 17276 15764 17332 15774
rect 16716 15138 16772 15148
rect 16828 15316 16884 15326
rect 16828 15204 16884 15260
rect 16940 15204 16996 15214
rect 16828 15202 16996 15204
rect 16828 15150 16942 15202
rect 16994 15150 16996 15202
rect 16828 15148 16996 15150
rect 16268 14702 16270 14754
rect 16322 14702 16324 14754
rect 16268 14690 16324 14702
rect 16492 14644 16548 14654
rect 15932 14252 16212 14308
rect 16268 14420 16324 14430
rect 15708 13748 15764 13758
rect 15484 13746 15764 13748
rect 15484 13694 15710 13746
rect 15762 13694 15764 13746
rect 15484 13692 15764 13694
rect 15260 13582 15262 13634
rect 15314 13582 15316 13634
rect 15260 13412 15316 13582
rect 15372 13636 15428 13646
rect 15372 13542 15428 13580
rect 15260 13346 15316 13356
rect 15484 13300 15540 13692
rect 15708 13682 15764 13692
rect 15372 13244 15540 13300
rect 15820 13412 15876 13422
rect 15372 13186 15428 13244
rect 15372 13134 15374 13186
rect 15426 13134 15428 13186
rect 15372 13122 15428 13134
rect 15148 12114 15204 12124
rect 15260 13076 15316 13086
rect 15036 12002 15092 12012
rect 14924 10670 14926 10722
rect 14978 10670 14980 10722
rect 14924 10658 14980 10670
rect 15148 11506 15204 11518
rect 15148 11454 15150 11506
rect 15202 11454 15204 11506
rect 14588 4834 14644 4844
rect 15148 9828 15204 11454
rect 14140 3668 14196 3678
rect 13468 3332 13636 3388
rect 13020 2930 13076 2940
rect 13580 2548 13636 3332
rect 13580 2482 13636 2492
rect 12124 1586 12180 1596
rect 12796 1652 12852 1662
rect 12796 112 12852 1596
rect 14140 112 14196 3612
rect 15148 1428 15204 9772
rect 15260 5236 15316 13020
rect 15484 12852 15540 12862
rect 15484 12758 15540 12796
rect 15820 12180 15876 13356
rect 15932 13188 15988 14252
rect 16268 14196 16324 14364
rect 16044 14140 16324 14196
rect 16044 13746 16100 14140
rect 16380 14084 16436 14094
rect 16380 13858 16436 14028
rect 16380 13806 16382 13858
rect 16434 13806 16436 13858
rect 16380 13794 16436 13806
rect 16044 13694 16046 13746
rect 16098 13694 16100 13746
rect 16044 13682 16100 13694
rect 16156 13746 16212 13758
rect 16156 13694 16158 13746
rect 16210 13694 16212 13746
rect 16156 13636 16212 13694
rect 16156 13570 16212 13580
rect 16492 13748 16548 14588
rect 16716 14532 16772 14542
rect 16716 14438 16772 14476
rect 16828 14420 16884 15148
rect 16940 15138 16996 15148
rect 16828 13972 16884 14364
rect 17052 14980 17108 14990
rect 16940 14306 16996 14318
rect 16940 14254 16942 14306
rect 16994 14254 16996 14306
rect 16940 14196 16996 14254
rect 16940 14130 16996 14140
rect 16940 13972 16996 13982
rect 16828 13970 16996 13972
rect 16828 13918 16942 13970
rect 16994 13918 16996 13970
rect 16828 13916 16996 13918
rect 17052 13972 17108 14924
rect 17164 14868 17220 14878
rect 17164 14530 17220 14812
rect 17164 14478 17166 14530
rect 17218 14478 17220 14530
rect 17164 14466 17220 14478
rect 17052 13916 17220 13972
rect 16940 13906 16996 13916
rect 17052 13748 17108 13758
rect 16492 13746 17108 13748
rect 16492 13694 16494 13746
rect 16546 13694 17054 13746
rect 17106 13694 17108 13746
rect 16492 13692 17108 13694
rect 16492 13412 16548 13692
rect 17052 13682 17108 13692
rect 16156 13356 16548 13412
rect 16716 13412 16772 13422
rect 16044 13188 16100 13198
rect 15932 13186 16100 13188
rect 15932 13134 16046 13186
rect 16098 13134 16100 13186
rect 15932 13132 16100 13134
rect 16044 13122 16100 13132
rect 16156 13074 16212 13356
rect 16156 13022 16158 13074
rect 16210 13022 16212 13074
rect 16156 12964 16212 13022
rect 16044 12908 16212 12964
rect 16044 12852 16100 12908
rect 16044 12786 16100 12796
rect 16156 12740 16212 12750
rect 15932 12180 15988 12190
rect 15820 12178 15988 12180
rect 15820 12126 15934 12178
rect 15986 12126 15988 12178
rect 15820 12124 15988 12126
rect 15932 6132 15988 12124
rect 16156 10724 16212 12684
rect 16604 12180 16660 12190
rect 16156 10658 16212 10668
rect 16492 12068 16548 12078
rect 16492 7252 16548 12012
rect 16492 7186 16548 7196
rect 16604 6580 16660 12124
rect 16716 9716 16772 13356
rect 17164 9940 17220 13916
rect 17276 13970 17332 15708
rect 17388 14868 17444 17948
rect 17500 14980 17556 23100
rect 17612 21588 17668 21598
rect 17612 21026 17668 21532
rect 17612 20974 17614 21026
rect 17666 20974 17668 21026
rect 17612 20962 17668 20974
rect 17500 14914 17556 14924
rect 17612 15876 17668 15886
rect 17388 14802 17444 14812
rect 17612 14754 17668 15820
rect 17612 14702 17614 14754
rect 17666 14702 17668 14754
rect 17612 14690 17668 14702
rect 17276 13918 17278 13970
rect 17330 13918 17332 13970
rect 17276 13906 17332 13918
rect 17388 14530 17444 14542
rect 17388 14478 17390 14530
rect 17442 14478 17444 14530
rect 17388 13970 17444 14478
rect 17388 13918 17390 13970
rect 17442 13918 17444 13970
rect 17388 13906 17444 13918
rect 17500 14418 17556 14430
rect 17500 14366 17502 14418
rect 17554 14366 17556 14418
rect 17500 13524 17556 14366
rect 17500 13458 17556 13468
rect 17724 12852 17780 23212
rect 17836 21476 17892 27694
rect 18060 26292 18116 32060
rect 18172 31892 18228 31902
rect 18172 31798 18228 31836
rect 18172 29426 18228 29438
rect 18172 29374 18174 29426
rect 18226 29374 18228 29426
rect 18172 27972 18228 29374
rect 18172 27906 18228 27916
rect 18172 27186 18228 27198
rect 18172 27134 18174 27186
rect 18226 27134 18228 27186
rect 18172 26852 18228 27134
rect 18172 26786 18228 26796
rect 18060 26236 18228 26292
rect 18060 26066 18116 26078
rect 18060 26014 18062 26066
rect 18114 26014 18116 26066
rect 17948 25508 18004 25518
rect 18060 25508 18116 26014
rect 17948 25506 18116 25508
rect 17948 25454 17950 25506
rect 18002 25454 18116 25506
rect 17948 25452 18116 25454
rect 17948 25442 18004 25452
rect 18172 25396 18228 26236
rect 18060 25340 18228 25396
rect 17948 24050 18004 24062
rect 17948 23998 17950 24050
rect 18002 23998 18004 24050
rect 17948 22708 18004 23998
rect 17948 22642 18004 22652
rect 18060 21588 18116 25340
rect 18172 25060 18228 25070
rect 18172 24834 18228 25004
rect 18172 24782 18174 24834
rect 18226 24782 18228 24834
rect 18172 24770 18228 24782
rect 18172 24388 18228 24398
rect 18172 22820 18228 24332
rect 18172 22754 18228 22764
rect 18284 21700 18340 32508
rect 18396 30994 18452 31006
rect 18396 30942 18398 30994
rect 18450 30942 18452 30994
rect 18396 30100 18452 30942
rect 18508 30324 18564 33516
rect 18620 32676 18676 32686
rect 18620 32582 18676 32620
rect 18732 30994 18788 31006
rect 18732 30942 18734 30994
rect 18786 30942 18788 30994
rect 18508 30268 18676 30324
rect 18508 30100 18564 30110
rect 18396 30098 18564 30100
rect 18396 30046 18510 30098
rect 18562 30046 18564 30098
rect 18396 30044 18564 30046
rect 18508 30034 18564 30044
rect 18620 29314 18676 30268
rect 18620 29262 18622 29314
rect 18674 29262 18676 29314
rect 18396 29092 18452 29102
rect 18396 28754 18452 29036
rect 18396 28702 18398 28754
rect 18450 28702 18452 28754
rect 18396 25732 18452 28702
rect 18396 25666 18452 25676
rect 18620 26068 18676 29262
rect 18732 29092 18788 30942
rect 18732 29026 18788 29036
rect 18844 28868 18900 35084
rect 18956 34914 19012 34926
rect 18956 34862 18958 34914
rect 19010 34862 19012 34914
rect 18956 32788 19012 34862
rect 18956 32722 19012 32732
rect 19068 32564 19124 32574
rect 19068 32470 19124 32508
rect 19180 32450 19236 32462
rect 19180 32398 19182 32450
rect 19234 32398 19236 32450
rect 18732 28812 18900 28868
rect 18956 31778 19012 31790
rect 18956 31726 18958 31778
rect 19010 31726 19012 31778
rect 18956 28868 19012 31726
rect 19180 31780 19236 32398
rect 19180 31714 19236 31724
rect 19068 31668 19124 31678
rect 19068 29764 19124 31612
rect 19068 29708 19236 29764
rect 18732 26908 18788 28812
rect 18956 28802 19012 28812
rect 18844 28644 18900 28654
rect 18844 28642 19124 28644
rect 18844 28590 18846 28642
rect 18898 28590 19124 28642
rect 18844 28588 19124 28590
rect 18844 28578 18900 28588
rect 19068 28082 19124 28588
rect 19068 28030 19070 28082
rect 19122 28030 19124 28082
rect 19068 28018 19124 28030
rect 19180 28642 19236 29708
rect 19180 28590 19182 28642
rect 19234 28590 19236 28642
rect 19068 27636 19124 27646
rect 18732 26852 18900 26908
rect 18508 25620 18564 25630
rect 18508 25526 18564 25564
rect 18396 25506 18452 25518
rect 18396 25454 18398 25506
rect 18450 25454 18452 25506
rect 18396 25396 18452 25454
rect 18396 25330 18452 25340
rect 18396 25060 18452 25070
rect 18396 23938 18452 25004
rect 18396 23886 18398 23938
rect 18450 23886 18452 23938
rect 18396 23604 18452 23886
rect 18396 23538 18452 23548
rect 18508 23828 18564 23838
rect 18508 23042 18564 23772
rect 18508 22990 18510 23042
rect 18562 22990 18564 23042
rect 18508 22978 18564 22990
rect 18508 22820 18564 22830
rect 18284 21644 18452 21700
rect 18060 21532 18228 21588
rect 17892 21420 18004 21476
rect 17836 21410 17892 21420
rect 17724 12786 17780 12796
rect 17836 20580 17892 20590
rect 17164 9874 17220 9884
rect 16716 9650 16772 9660
rect 16604 6514 16660 6524
rect 15932 6066 15988 6076
rect 15260 5170 15316 5180
rect 16828 4564 16884 4574
rect 15148 1362 15204 1372
rect 15484 1652 15540 1662
rect 15484 112 15540 1596
rect 16828 112 16884 4508
rect 17836 4116 17892 20524
rect 17948 19796 18004 21420
rect 18172 21364 18228 21532
rect 18284 21476 18340 21486
rect 18284 21382 18340 21420
rect 18060 21308 18228 21364
rect 18060 19908 18116 21308
rect 18396 21252 18452 21644
rect 18172 21196 18452 21252
rect 18172 20132 18228 21196
rect 18172 20130 18340 20132
rect 18172 20078 18174 20130
rect 18226 20078 18340 20130
rect 18172 20076 18340 20078
rect 18172 20066 18228 20076
rect 18060 19852 18228 19908
rect 17948 19740 18116 19796
rect 17948 16884 18004 16894
rect 17948 16790 18004 16828
rect 17948 16548 18004 16558
rect 17948 16322 18004 16492
rect 17948 16270 17950 16322
rect 18002 16270 18004 16322
rect 17948 16258 18004 16270
rect 18060 15202 18116 19740
rect 18060 15150 18062 15202
rect 18114 15150 18116 15202
rect 18060 15138 18116 15150
rect 17948 14868 18004 14878
rect 17948 10836 18004 14812
rect 17948 10770 18004 10780
rect 17836 4050 17892 4060
rect 18172 112 18228 19852
rect 18284 18900 18340 20076
rect 18284 18834 18340 18844
rect 18508 19906 18564 22764
rect 18620 22482 18676 26012
rect 18620 22430 18622 22482
rect 18674 22430 18676 22482
rect 18620 21028 18676 22430
rect 18732 23604 18788 23614
rect 18732 21700 18788 23548
rect 18732 21606 18788 21644
rect 18732 21028 18788 21038
rect 18620 21026 18788 21028
rect 18620 20974 18734 21026
rect 18786 20974 18788 21026
rect 18620 20972 18788 20974
rect 18732 20962 18788 20972
rect 18508 19854 18510 19906
rect 18562 19854 18564 19906
rect 18284 18676 18340 18686
rect 18284 4340 18340 18620
rect 18396 18452 18452 18462
rect 18396 16098 18452 18396
rect 18508 18228 18564 19854
rect 18844 18564 18900 26852
rect 18956 25620 19012 25630
rect 18956 24722 19012 25564
rect 18956 24670 18958 24722
rect 19010 24670 19012 24722
rect 18956 24658 19012 24670
rect 18956 23604 19012 23614
rect 18956 23266 19012 23548
rect 18956 23214 18958 23266
rect 19010 23214 19012 23266
rect 18956 23202 19012 23214
rect 18508 16548 18564 18172
rect 18508 16482 18564 16492
rect 18620 18508 18900 18564
rect 18956 22258 19012 22270
rect 18956 22206 18958 22258
rect 19010 22206 19012 22258
rect 18396 16046 18398 16098
rect 18450 16046 18452 16098
rect 18396 15428 18452 16046
rect 18508 15428 18564 15438
rect 18396 15426 18564 15428
rect 18396 15374 18510 15426
rect 18562 15374 18564 15426
rect 18396 15372 18564 15374
rect 18396 14308 18452 15372
rect 18508 15362 18564 15372
rect 18620 15148 18676 18508
rect 18956 18452 19012 22206
rect 18956 18386 19012 18396
rect 18956 18228 19012 18238
rect 18956 18134 19012 18172
rect 18620 15092 18900 15148
rect 18396 14242 18452 14252
rect 18284 4274 18340 4284
rect 672 0 784 112
rect 2016 0 2128 112
rect 3360 0 3472 112
rect 4704 0 4816 112
rect 6048 0 6160 112
rect 7392 0 7504 112
rect 8736 0 8848 112
rect 10080 0 10192 112
rect 11424 0 11536 112
rect 12768 0 12880 112
rect 14112 0 14224 112
rect 15456 0 15568 112
rect 16800 0 16912 112
rect 18144 0 18256 112
rect 18844 84 18900 15092
rect 19068 8932 19124 27580
rect 19180 26908 19236 28590
rect 19292 27636 19348 38612
rect 19404 34802 19460 34814
rect 19404 34750 19406 34802
rect 19458 34750 19460 34802
rect 19404 30884 19460 34750
rect 19516 33122 19572 33134
rect 19516 33070 19518 33122
rect 19570 33070 19572 33122
rect 19516 32564 19572 33070
rect 19516 32498 19572 32508
rect 19404 30828 19572 30884
rect 19404 28754 19460 28766
rect 19404 28702 19406 28754
rect 19458 28702 19460 28754
rect 19404 27748 19460 28702
rect 19516 28196 19572 30828
rect 19628 28196 19684 40236
rect 19740 37938 19796 37950
rect 19740 37886 19742 37938
rect 19794 37886 19796 37938
rect 19740 35364 19796 37886
rect 19740 35298 19796 35308
rect 19852 35028 19908 35038
rect 19852 34934 19908 34972
rect 19852 31780 19908 31790
rect 19852 30996 19908 31724
rect 19852 30902 19908 30940
rect 19740 29428 19796 29438
rect 19740 29334 19796 29372
rect 19964 29428 20020 50372
rect 19964 29362 20020 29372
rect 20076 46452 20132 46462
rect 19740 28980 19796 28990
rect 19740 28644 19796 28924
rect 20076 28980 20132 46396
rect 20076 28914 20132 28924
rect 20188 29428 20244 29438
rect 20076 28644 20132 28654
rect 19740 28588 19908 28644
rect 19628 28140 19796 28196
rect 19516 28130 19572 28140
rect 19516 27748 19572 27758
rect 19404 27746 19572 27748
rect 19404 27694 19518 27746
rect 19570 27694 19572 27746
rect 19404 27692 19572 27694
rect 19516 27682 19572 27692
rect 19292 27570 19348 27580
rect 19516 27524 19572 27534
rect 19180 26852 19348 26908
rect 19180 26068 19236 26078
rect 19180 25974 19236 26012
rect 19292 25732 19348 26852
rect 19292 25666 19348 25676
rect 19404 26850 19460 26862
rect 19404 26798 19406 26850
rect 19458 26798 19460 26850
rect 19180 25508 19236 25518
rect 19404 25508 19460 26798
rect 19180 25506 19460 25508
rect 19180 25454 19182 25506
rect 19234 25454 19460 25506
rect 19180 25452 19460 25454
rect 19180 25442 19236 25452
rect 19516 25396 19572 27468
rect 19740 26908 19796 28140
rect 19628 26852 19796 26908
rect 19628 26402 19684 26852
rect 19628 26350 19630 26402
rect 19682 26350 19684 26402
rect 19628 26338 19684 26350
rect 19404 25340 19572 25396
rect 19628 26180 19684 26190
rect 19404 24164 19460 25340
rect 19516 24836 19572 24846
rect 19628 24836 19684 26124
rect 19740 25508 19796 25518
rect 19740 25414 19796 25452
rect 19516 24834 19684 24836
rect 19516 24782 19518 24834
rect 19570 24782 19684 24834
rect 19516 24780 19684 24782
rect 19516 24770 19572 24780
rect 19404 24098 19460 24108
rect 19404 23938 19460 23950
rect 19404 23886 19406 23938
rect 19458 23886 19460 23938
rect 19404 23828 19460 23886
rect 19404 23762 19460 23772
rect 19852 23826 19908 28588
rect 20076 28550 20132 28588
rect 20076 28084 20132 28094
rect 20076 27970 20132 28028
rect 20076 27918 20078 27970
rect 20130 27918 20132 27970
rect 20076 27906 20132 27918
rect 20188 27748 20244 29372
rect 20076 27692 20244 27748
rect 19852 23774 19854 23826
rect 19906 23774 19908 23826
rect 19852 23762 19908 23774
rect 19964 25396 20020 25406
rect 19404 21924 19460 21934
rect 19180 21700 19236 21710
rect 19180 20802 19236 21644
rect 19292 21476 19348 21486
rect 19292 21382 19348 21420
rect 19180 20750 19182 20802
rect 19234 20750 19236 20802
rect 19180 20738 19236 20750
rect 19068 8866 19124 8876
rect 19404 980 19460 21868
rect 19852 21362 19908 21374
rect 19852 21310 19854 21362
rect 19906 21310 19908 21362
rect 19852 21026 19908 21310
rect 19852 20974 19854 21026
rect 19906 20974 19908 21026
rect 19852 20962 19908 20974
rect 19740 20916 19796 20926
rect 19740 20130 19796 20860
rect 19740 20078 19742 20130
rect 19794 20078 19796 20130
rect 19740 20066 19796 20078
rect 19516 18452 19572 18462
rect 19516 18358 19572 18396
rect 19964 16660 20020 25340
rect 19964 16594 20020 16604
rect 20076 5124 20132 27692
rect 20188 25956 20244 25966
rect 20188 20802 20244 25900
rect 20188 20750 20190 20802
rect 20242 20750 20244 20802
rect 20188 20738 20244 20750
rect 20300 12740 20356 50372
rect 20972 45892 21028 45902
rect 20412 44436 20468 44446
rect 20412 35026 20468 44380
rect 20412 34974 20414 35026
rect 20466 34974 20468 35026
rect 20412 34962 20468 34974
rect 20412 28868 20468 28878
rect 20412 28642 20468 28812
rect 20412 28590 20414 28642
rect 20466 28590 20468 28642
rect 20412 28578 20468 28590
rect 20636 28642 20692 28654
rect 20636 28590 20638 28642
rect 20690 28590 20692 28642
rect 20524 25506 20580 25518
rect 20524 25454 20526 25506
rect 20578 25454 20580 25506
rect 20412 20916 20468 20926
rect 20412 20822 20468 20860
rect 20524 20356 20580 25454
rect 20636 25508 20692 28590
rect 20636 25442 20692 25452
rect 20524 20290 20580 20300
rect 20748 21140 20804 21150
rect 20748 20914 20804 21084
rect 20748 20862 20750 20914
rect 20802 20862 20804 20914
rect 20300 12674 20356 12684
rect 20076 5058 20132 5068
rect 20748 1204 20804 20862
rect 20972 7364 21028 45836
rect 20972 7298 21028 7308
rect 21084 6020 21140 51100
rect 21532 37380 21588 54350
rect 21532 37314 21588 37324
rect 21644 53732 21700 53742
rect 21532 35476 21588 35486
rect 21420 28642 21476 28654
rect 21420 28590 21422 28642
rect 21474 28590 21476 28642
rect 21308 25508 21364 25518
rect 21084 5954 21140 5964
rect 21196 20356 21252 20366
rect 20748 1138 20804 1148
rect 20860 3332 20916 3342
rect 19404 914 19460 924
rect 19180 196 19236 206
rect 19180 84 19236 140
rect 19516 196 19572 206
rect 19516 112 19572 140
rect 20860 112 20916 3276
rect 21196 2100 21252 20300
rect 21308 9268 21364 25452
rect 21308 9202 21364 9212
rect 21420 16884 21476 28590
rect 21532 21588 21588 35420
rect 21532 21522 21588 21532
rect 21420 5684 21476 16828
rect 21644 16772 21700 53676
rect 21868 53730 21924 53742
rect 21868 53678 21870 53730
rect 21922 53678 21924 53730
rect 21868 53508 21924 53678
rect 21868 53442 21924 53452
rect 21756 53172 21812 53182
rect 21756 53058 21812 53116
rect 21756 53006 21758 53058
rect 21810 53006 21812 53058
rect 21756 52994 21812 53006
rect 21868 52276 21924 52286
rect 21980 52276 22036 55916
rect 22540 54738 22596 56140
rect 22652 55186 22708 57148
rect 23548 56308 23604 57344
rect 23804 56476 24068 56486
rect 23860 56420 23908 56476
rect 23964 56420 24012 56476
rect 23804 56410 24068 56420
rect 23548 56242 23604 56252
rect 24444 56308 24500 56318
rect 24444 56214 24500 56252
rect 24892 56308 24948 57344
rect 25452 57316 25508 57326
rect 24892 56242 24948 56252
rect 25116 57204 25172 57214
rect 23548 56084 23604 56094
rect 22876 55970 22932 55982
rect 22876 55918 22878 55970
rect 22930 55918 22932 55970
rect 22876 55468 22932 55918
rect 23436 55524 23492 55534
rect 22876 55412 23044 55468
rect 22652 55134 22654 55186
rect 22706 55134 22708 55186
rect 22652 55122 22708 55134
rect 22540 54686 22542 54738
rect 22594 54686 22596 54738
rect 22540 54674 22596 54686
rect 22316 53956 22372 53966
rect 22316 53730 22372 53900
rect 22316 53678 22318 53730
rect 22370 53678 22372 53730
rect 22316 53666 22372 53678
rect 22876 53730 22932 53742
rect 22876 53678 22878 53730
rect 22930 53678 22932 53730
rect 22652 53284 22708 53294
rect 22652 53058 22708 53228
rect 22652 53006 22654 53058
rect 22706 53006 22708 53058
rect 22652 52994 22708 53006
rect 22204 52724 22260 52734
rect 22204 52630 22260 52668
rect 21868 52274 22036 52276
rect 21868 52222 21870 52274
rect 21922 52222 22036 52274
rect 21868 52220 22036 52222
rect 22764 52276 22820 52286
rect 21868 52210 21924 52220
rect 22764 52182 22820 52220
rect 22428 52162 22484 52174
rect 22428 52110 22430 52162
rect 22482 52110 22484 52162
rect 22204 36708 22260 36718
rect 21868 27412 21924 27422
rect 21868 21700 21924 27356
rect 21868 21634 21924 21644
rect 21644 16706 21700 16716
rect 21420 5618 21476 5628
rect 21196 2034 21252 2044
rect 22204 112 22260 36652
rect 22428 1316 22484 52110
rect 22876 51492 22932 53678
rect 22876 51426 22932 51436
rect 22764 51154 22820 51166
rect 22764 51102 22766 51154
rect 22818 51102 22820 51154
rect 22652 40404 22708 40414
rect 22652 9380 22708 40348
rect 22652 9314 22708 9324
rect 22764 3668 22820 51102
rect 22988 49924 23044 55412
rect 23100 54402 23156 54414
rect 23100 54350 23102 54402
rect 23154 54350 23156 54402
rect 23100 51380 23156 54350
rect 23100 51314 23156 51324
rect 23212 52946 23268 52958
rect 23212 52894 23214 52946
rect 23266 52894 23268 52946
rect 22988 49858 23044 49868
rect 23212 39396 23268 52894
rect 23324 51492 23380 51502
rect 23436 51492 23492 55468
rect 23548 52274 23604 56028
rect 23884 55972 23940 55982
rect 23884 55878 23940 55916
rect 24464 55692 24728 55702
rect 24520 55636 24568 55692
rect 24624 55636 24672 55692
rect 24464 55626 24728 55636
rect 24780 55412 24836 55422
rect 23660 55300 23716 55310
rect 23660 55206 23716 55244
rect 24668 55298 24724 55310
rect 24668 55246 24670 55298
rect 24722 55246 24724 55298
rect 24668 55188 24724 55246
rect 24668 55122 24724 55132
rect 24332 55076 24388 55086
rect 24220 54964 24276 54974
rect 23804 54908 24068 54918
rect 23860 54852 23908 54908
rect 23964 54852 24012 54908
rect 23804 54842 24068 54852
rect 24108 54740 24164 54750
rect 24220 54740 24276 54908
rect 24108 54738 24276 54740
rect 24108 54686 24110 54738
rect 24162 54686 24276 54738
rect 24108 54684 24276 54686
rect 24108 54674 24164 54684
rect 23548 52222 23550 52274
rect 23602 52222 23604 52274
rect 23548 52210 23604 52222
rect 23660 54516 23716 54526
rect 23324 51490 23492 51492
rect 23324 51438 23326 51490
rect 23378 51438 23492 51490
rect 23324 51436 23492 51438
rect 23324 51426 23380 51436
rect 23436 50708 23492 50718
rect 23660 50708 23716 54460
rect 23772 54180 23828 54190
rect 23772 53618 23828 54124
rect 23772 53566 23774 53618
rect 23826 53566 23828 53618
rect 23772 53554 23828 53566
rect 23804 53340 24068 53350
rect 23860 53284 23908 53340
rect 23964 53284 24012 53340
rect 23804 53274 24068 53284
rect 24108 53172 24164 53182
rect 24108 53078 24164 53116
rect 23804 51772 24068 51782
rect 23860 51716 23908 51772
rect 23964 51716 24012 51772
rect 23804 51706 24068 51716
rect 24332 51490 24388 55020
rect 24668 54516 24724 54526
rect 24668 54422 24724 54460
rect 24780 54292 24836 55356
rect 24780 54226 24836 54236
rect 25004 55300 25060 55310
rect 24464 54124 24728 54134
rect 24520 54068 24568 54124
rect 24624 54068 24672 54124
rect 24464 54058 24728 54068
rect 24892 53732 24948 53742
rect 24892 53638 24948 53676
rect 24668 53060 24724 53070
rect 24668 52946 24724 53004
rect 24668 52894 24670 52946
rect 24722 52894 24724 52946
rect 24668 52882 24724 52894
rect 24464 52556 24728 52566
rect 24520 52500 24568 52556
rect 24624 52500 24672 52556
rect 24464 52490 24728 52500
rect 24668 52388 24724 52398
rect 24668 52274 24724 52332
rect 24668 52222 24670 52274
rect 24722 52222 24724 52274
rect 24668 52210 24724 52222
rect 24332 51438 24334 51490
rect 24386 51438 24388 51490
rect 24332 51426 24388 51438
rect 24668 51268 24724 51278
rect 24668 51174 24724 51212
rect 23772 51156 23828 51166
rect 23772 51062 23828 51100
rect 24464 50988 24728 50998
rect 24520 50932 24568 50988
rect 24624 50932 24672 50988
rect 24464 50922 24728 50932
rect 23436 50706 23716 50708
rect 23436 50654 23438 50706
rect 23490 50654 23716 50706
rect 23436 50652 23716 50654
rect 23436 50642 23492 50652
rect 23884 50596 23940 50606
rect 23548 50594 23940 50596
rect 23548 50542 23886 50594
rect 23938 50542 23940 50594
rect 23548 50540 23940 50542
rect 23548 50428 23604 50540
rect 23884 50530 23940 50540
rect 24892 50594 24948 50606
rect 24892 50542 24894 50594
rect 24946 50542 24948 50594
rect 23212 39330 23268 39340
rect 23436 50372 23604 50428
rect 22764 3602 22820 3612
rect 22876 30996 22932 31006
rect 22428 1250 22484 1260
rect 22876 308 22932 30940
rect 23100 29988 23156 29998
rect 22988 21364 23044 21374
rect 22988 3444 23044 21308
rect 23100 19124 23156 29932
rect 23100 19058 23156 19068
rect 23436 11284 23492 50372
rect 23804 50204 24068 50214
rect 23860 50148 23908 50204
rect 23964 50148 24012 50204
rect 23804 50138 24068 50148
rect 24220 49924 24276 49934
rect 24220 49830 24276 49868
rect 24668 49698 24724 49710
rect 24668 49646 24670 49698
rect 24722 49646 24724 49698
rect 23772 49586 23828 49598
rect 23772 49534 23774 49586
rect 23826 49534 23828 49586
rect 23772 49252 23828 49534
rect 24668 49588 24724 49646
rect 24668 49522 24724 49532
rect 24464 49420 24728 49430
rect 24520 49364 24568 49420
rect 24624 49364 24672 49420
rect 24464 49354 24728 49364
rect 23772 49186 23828 49196
rect 24668 49026 24724 49038
rect 24668 48974 24670 49026
rect 24722 48974 24724 49026
rect 24668 48916 24724 48974
rect 24668 48850 24724 48860
rect 23804 48636 24068 48646
rect 23860 48580 23908 48636
rect 23964 48580 24012 48636
rect 23804 48570 24068 48580
rect 24892 48244 24948 50542
rect 25004 48354 25060 55244
rect 25116 53172 25172 57148
rect 25116 53106 25172 53116
rect 25340 56756 25396 56766
rect 25340 51490 25396 56700
rect 25452 54626 25508 57260
rect 26236 57316 26292 57344
rect 26236 57250 26292 57260
rect 26012 56308 26068 56318
rect 26012 56214 26068 56252
rect 25676 56082 25732 56094
rect 25676 56030 25678 56082
rect 25730 56030 25732 56082
rect 25452 54574 25454 54626
rect 25506 54574 25508 54626
rect 25452 54562 25508 54574
rect 25564 55186 25620 55198
rect 25564 55134 25566 55186
rect 25618 55134 25620 55186
rect 25564 54516 25620 55134
rect 25564 54450 25620 54460
rect 25564 53620 25620 53630
rect 25564 53526 25620 53564
rect 25452 52834 25508 52846
rect 25452 52782 25454 52834
rect 25506 52782 25508 52834
rect 25452 52724 25508 52782
rect 25452 52658 25508 52668
rect 25564 52050 25620 52062
rect 25564 51998 25566 52050
rect 25618 51998 25620 52050
rect 25564 51828 25620 51998
rect 25564 51762 25620 51772
rect 25340 51438 25342 51490
rect 25394 51438 25396 51490
rect 25340 51426 25396 51438
rect 25564 50484 25620 50494
rect 25564 50390 25620 50428
rect 25676 50428 25732 56030
rect 27580 56084 27636 57344
rect 27580 56018 27636 56028
rect 26236 55300 26292 55310
rect 25900 55298 26292 55300
rect 25900 55246 26238 55298
rect 26290 55246 26292 55298
rect 25900 55244 26292 55246
rect 25676 50372 25844 50428
rect 25676 49922 25732 49934
rect 25676 49870 25678 49922
rect 25730 49870 25732 49922
rect 25676 49588 25732 49870
rect 25676 49522 25732 49532
rect 25676 48802 25732 48814
rect 25676 48750 25678 48802
rect 25730 48750 25732 48802
rect 25676 48692 25732 48750
rect 25676 48626 25732 48636
rect 25004 48302 25006 48354
rect 25058 48302 25060 48354
rect 25004 48290 25060 48302
rect 25788 48354 25844 50372
rect 25788 48302 25790 48354
rect 25842 48302 25844 48354
rect 25788 48290 25844 48302
rect 24892 48178 24948 48188
rect 24444 48020 24500 48030
rect 24332 48018 24500 48020
rect 24332 47966 24446 48018
rect 24498 47966 24500 48018
rect 24332 47964 24500 47966
rect 24332 47236 24388 47964
rect 24444 47954 24500 47964
rect 25340 48020 25396 48030
rect 25340 47926 25396 47964
rect 24464 47852 24728 47862
rect 24520 47796 24568 47852
rect 24624 47796 24672 47852
rect 24464 47786 24728 47796
rect 24332 47170 24388 47180
rect 24668 47458 24724 47470
rect 24668 47406 24670 47458
rect 24722 47406 24724 47458
rect 23804 47068 24068 47078
rect 23860 47012 23908 47068
rect 23964 47012 24012 47068
rect 23804 47002 24068 47012
rect 24668 46452 24724 47406
rect 25676 47348 25732 47358
rect 25676 47254 25732 47292
rect 25676 46786 25732 46798
rect 25676 46734 25678 46786
rect 25730 46734 25732 46786
rect 24668 46386 24724 46396
rect 24892 46674 24948 46686
rect 24892 46622 24894 46674
rect 24946 46622 24948 46674
rect 24464 46284 24728 46294
rect 24520 46228 24568 46284
rect 24624 46228 24672 46284
rect 24464 46218 24728 46228
rect 24668 45892 24724 45902
rect 24668 45798 24724 45836
rect 23804 45500 24068 45510
rect 23860 45444 23908 45500
rect 23964 45444 24012 45500
rect 23804 45434 24068 45444
rect 24464 44716 24728 44726
rect 24520 44660 24568 44716
rect 24624 44660 24672 44716
rect 24464 44650 24728 44660
rect 24892 44548 24948 46622
rect 25676 46452 25732 46734
rect 25676 46386 25732 46396
rect 25676 45666 25732 45678
rect 25676 45614 25678 45666
rect 25730 45614 25732 45666
rect 25676 45556 25732 45614
rect 25676 45490 25732 45500
rect 24892 44482 24948 44492
rect 25900 44436 25956 55244
rect 26236 55234 26292 55244
rect 27244 55074 27300 55086
rect 27244 55022 27246 55074
rect 27298 55022 27300 55074
rect 26236 54404 26292 54414
rect 26236 54310 26292 54348
rect 27020 54402 27076 54414
rect 27020 54350 27022 54402
rect 27074 54350 27076 54402
rect 26236 53732 26292 53742
rect 26124 53730 26292 53732
rect 26124 53678 26238 53730
rect 26290 53678 26292 53730
rect 26124 53676 26292 53678
rect 26124 46116 26180 53676
rect 26236 53666 26292 53676
rect 26796 53732 26852 53742
rect 26236 52836 26292 52846
rect 26236 52742 26292 52780
rect 26236 52164 26292 52174
rect 26236 52070 26292 52108
rect 26348 51940 26404 51950
rect 26236 51266 26292 51278
rect 26236 51214 26238 51266
rect 26290 51214 26292 51266
rect 26236 50820 26292 51214
rect 26236 50754 26292 50764
rect 26348 50594 26404 51884
rect 26348 50542 26350 50594
rect 26402 50542 26404 50594
rect 26348 50530 26404 50542
rect 26348 49810 26404 49822
rect 26348 49758 26350 49810
rect 26402 49758 26404 49810
rect 26236 49028 26292 49038
rect 26236 48934 26292 48972
rect 26348 48804 26404 49758
rect 26348 48738 26404 48748
rect 26236 48132 26292 48142
rect 26236 48038 26292 48076
rect 26460 47460 26516 47470
rect 26460 47458 26628 47460
rect 26460 47406 26462 47458
rect 26514 47406 26628 47458
rect 26460 47404 26628 47406
rect 26460 47394 26516 47404
rect 26124 46050 26180 46060
rect 26348 46674 26404 46686
rect 26348 46622 26350 46674
rect 26402 46622 26404 46674
rect 26236 45892 26292 45902
rect 25900 44370 25956 44380
rect 26012 45890 26292 45892
rect 26012 45838 26238 45890
rect 26290 45838 26292 45890
rect 26012 45836 26292 45838
rect 24668 44322 24724 44334
rect 24668 44270 24670 44322
rect 24722 44270 24724 44322
rect 24668 44100 24724 44270
rect 25676 44212 25732 44222
rect 25676 44118 25732 44156
rect 24668 44034 24724 44044
rect 23804 43932 24068 43942
rect 23860 43876 23908 43932
rect 23964 43876 24012 43932
rect 23804 43866 24068 43876
rect 25676 43650 25732 43662
rect 25676 43598 25678 43650
rect 25730 43598 25732 43650
rect 24892 43538 24948 43550
rect 24892 43486 24894 43538
rect 24946 43486 24948 43538
rect 24464 43148 24728 43158
rect 24520 43092 24568 43148
rect 24624 43092 24672 43148
rect 24464 43082 24728 43092
rect 24668 42754 24724 42766
rect 24668 42702 24670 42754
rect 24722 42702 24724 42754
rect 24668 42644 24724 42702
rect 24668 42578 24724 42588
rect 23804 42364 24068 42374
rect 23860 42308 23908 42364
rect 23964 42308 24012 42364
rect 23804 42298 24068 42308
rect 24464 41580 24728 41590
rect 24520 41524 24568 41580
rect 24624 41524 24672 41580
rect 24464 41514 24728 41524
rect 24780 41186 24836 41198
rect 24780 41134 24782 41186
rect 24834 41134 24836 41186
rect 23804 40796 24068 40806
rect 23860 40740 23908 40796
rect 23964 40740 24012 40796
rect 23804 40730 24068 40740
rect 24668 40404 24724 40414
rect 24668 40310 24724 40348
rect 24780 40180 24836 41134
rect 24892 40628 24948 43486
rect 25676 43316 25732 43598
rect 25676 43250 25732 43260
rect 25676 42530 25732 42542
rect 25676 42478 25678 42530
rect 25730 42478 25732 42530
rect 25676 42420 25732 42478
rect 25676 42354 25732 42364
rect 25676 41076 25732 41086
rect 25676 40982 25732 41020
rect 24892 40562 24948 40572
rect 24780 40114 24836 40124
rect 25676 40514 25732 40526
rect 25676 40462 25678 40514
rect 25730 40462 25732 40514
rect 25676 40180 25732 40462
rect 25676 40114 25732 40124
rect 24464 40012 24728 40022
rect 24520 39956 24568 40012
rect 24624 39956 24672 40012
rect 24464 39946 24728 39956
rect 24668 39732 24724 39742
rect 24668 39638 24724 39676
rect 25676 39394 25732 39406
rect 25676 39342 25678 39394
rect 25730 39342 25732 39394
rect 25676 39284 25732 39342
rect 23804 39228 24068 39238
rect 23860 39172 23908 39228
rect 23964 39172 24012 39228
rect 25676 39218 25732 39228
rect 23804 39162 24068 39172
rect 24464 38444 24728 38454
rect 24520 38388 24568 38444
rect 24624 38388 24672 38444
rect 24464 38378 24728 38388
rect 24892 38052 24948 38062
rect 25564 38052 25620 38062
rect 24892 38050 25172 38052
rect 24892 37998 24894 38050
rect 24946 37998 25172 38050
rect 24892 37996 25172 37998
rect 24892 37986 24948 37996
rect 23804 37660 24068 37670
rect 23860 37604 23908 37660
rect 23964 37604 24012 37660
rect 23804 37594 24068 37604
rect 24668 37156 24724 37166
rect 24332 37154 24724 37156
rect 24332 37102 24670 37154
rect 24722 37102 24724 37154
rect 24332 37100 24724 37102
rect 23660 36148 23716 36158
rect 23548 33908 23604 33918
rect 23548 25284 23604 33852
rect 23660 30772 23716 36092
rect 23804 36092 24068 36102
rect 23860 36036 23908 36092
rect 23964 36036 24012 36092
rect 23804 36026 24068 36036
rect 23804 34524 24068 34534
rect 23860 34468 23908 34524
rect 23964 34468 24012 34524
rect 23804 34458 24068 34468
rect 23804 32956 24068 32966
rect 23860 32900 23908 32956
rect 23964 32900 24012 32956
rect 23804 32890 24068 32900
rect 24332 32004 24388 37100
rect 24668 37090 24724 37100
rect 24464 36876 24728 36886
rect 24520 36820 24568 36876
rect 24624 36820 24672 36876
rect 24464 36810 24728 36820
rect 24892 36484 24948 36494
rect 24892 36482 25060 36484
rect 24892 36430 24894 36482
rect 24946 36430 25060 36482
rect 24892 36428 25060 36430
rect 24892 36418 24948 36428
rect 24464 35308 24728 35318
rect 24520 35252 24568 35308
rect 24624 35252 24672 35308
rect 24464 35242 24728 35252
rect 24668 34914 24724 34926
rect 24668 34862 24670 34914
rect 24722 34862 24724 34914
rect 24668 34356 24724 34862
rect 24668 34290 24724 34300
rect 24892 34804 24948 34814
rect 24668 34018 24724 34030
rect 24668 33966 24670 34018
rect 24722 33966 24724 34018
rect 24668 33908 24724 33966
rect 24668 33842 24724 33852
rect 24464 33740 24728 33750
rect 24520 33684 24568 33740
rect 24624 33684 24672 33740
rect 24464 33674 24728 33684
rect 24668 33346 24724 33358
rect 24668 33294 24670 33346
rect 24722 33294 24724 33346
rect 24668 32340 24724 33294
rect 24668 32274 24724 32284
rect 24464 32172 24728 32182
rect 24520 32116 24568 32172
rect 24624 32116 24672 32172
rect 24464 32106 24728 32116
rect 24332 31938 24388 31948
rect 24668 31780 24724 31790
rect 24220 31778 24724 31780
rect 24220 31726 24670 31778
rect 24722 31726 24724 31778
rect 24220 31724 24724 31726
rect 23804 31388 24068 31398
rect 23860 31332 23908 31388
rect 23964 31332 24012 31388
rect 23804 31322 24068 31332
rect 23660 30706 23716 30716
rect 23804 29820 24068 29830
rect 23860 29764 23908 29820
rect 23964 29764 24012 29820
rect 23804 29754 24068 29764
rect 23804 28252 24068 28262
rect 23860 28196 23908 28252
rect 23964 28196 24012 28252
rect 23804 28186 24068 28196
rect 23804 26684 24068 26694
rect 23860 26628 23908 26684
rect 23964 26628 24012 26684
rect 23804 26618 24068 26628
rect 23548 25218 23604 25228
rect 23804 25116 24068 25126
rect 23860 25060 23908 25116
rect 23964 25060 24012 25116
rect 23804 25050 24068 25060
rect 23804 23548 24068 23558
rect 23860 23492 23908 23548
rect 23964 23492 24012 23548
rect 23804 23482 24068 23492
rect 24220 23268 24276 31724
rect 24668 31714 24724 31724
rect 24892 30994 24948 34748
rect 24892 30942 24894 30994
rect 24946 30942 24948 30994
rect 24892 30930 24948 30942
rect 24892 30772 24948 30782
rect 24464 30604 24728 30614
rect 24520 30548 24568 30604
rect 24624 30548 24672 30604
rect 24464 30538 24728 30548
rect 24464 29036 24728 29046
rect 24520 28980 24568 29036
rect 24624 28980 24672 29036
rect 24464 28970 24728 28980
rect 24332 27860 24388 27870
rect 24332 25620 24388 27804
rect 24668 27748 24724 27758
rect 24668 27654 24724 27692
rect 24464 27468 24728 27478
rect 24520 27412 24568 27468
rect 24624 27412 24672 27468
rect 24464 27402 24728 27412
rect 24668 27300 24724 27310
rect 24668 27186 24724 27244
rect 24668 27134 24670 27186
rect 24722 27134 24724 27186
rect 24668 27122 24724 27134
rect 24464 25900 24728 25910
rect 24520 25844 24568 25900
rect 24624 25844 24672 25900
rect 24464 25834 24728 25844
rect 24668 25620 24724 25630
rect 24332 25618 24724 25620
rect 24332 25566 24670 25618
rect 24722 25566 24724 25618
rect 24332 25564 24724 25566
rect 24668 25554 24724 25564
rect 24892 24722 24948 30716
rect 25004 29540 25060 36428
rect 25004 29474 25060 29484
rect 25116 29204 25172 37996
rect 25452 37154 25508 37166
rect 25452 37102 25454 37154
rect 25506 37102 25508 37154
rect 25452 37044 25508 37102
rect 25452 36978 25508 36988
rect 25452 30882 25508 30894
rect 25452 30830 25454 30882
rect 25506 30830 25508 30882
rect 25452 30772 25508 30830
rect 25452 30706 25508 30716
rect 25116 29138 25172 29148
rect 25564 28756 25620 37996
rect 25676 37940 25732 37950
rect 25676 37846 25732 37884
rect 25676 36258 25732 36270
rect 25676 36206 25678 36258
rect 25730 36206 25732 36258
rect 25676 36148 25732 36206
rect 25676 36082 25732 36092
rect 25900 35588 25956 35598
rect 25676 34804 25732 34814
rect 25676 34710 25732 34748
rect 25676 34242 25732 34254
rect 25676 34190 25678 34242
rect 25730 34190 25732 34242
rect 25676 33908 25732 34190
rect 25676 33842 25732 33852
rect 25676 33122 25732 33134
rect 25676 33070 25678 33122
rect 25730 33070 25732 33122
rect 25676 33012 25732 33070
rect 25676 32946 25732 32956
rect 25676 31668 25732 31678
rect 25676 31574 25732 31612
rect 25900 30996 25956 35532
rect 25900 30930 25956 30940
rect 25564 28690 25620 28700
rect 25676 30884 25732 30894
rect 25676 28420 25732 30828
rect 25788 30436 25844 30446
rect 25788 28756 25844 30380
rect 25788 28690 25844 28700
rect 25900 30212 25956 30222
rect 25676 28354 25732 28364
rect 25676 27970 25732 27982
rect 25676 27918 25678 27970
rect 25730 27918 25732 27970
rect 25676 27188 25732 27918
rect 25676 27122 25732 27132
rect 25676 26850 25732 26862
rect 25676 26798 25678 26850
rect 25730 26798 25732 26850
rect 25676 26292 25732 26798
rect 25676 26226 25732 26236
rect 24892 24670 24894 24722
rect 24946 24670 24948 24722
rect 24892 24658 24948 24670
rect 25564 25508 25620 25518
rect 25452 24610 25508 24622
rect 25452 24558 25454 24610
rect 25506 24558 25508 24610
rect 24464 24332 24728 24342
rect 24520 24276 24568 24332
rect 24624 24276 24672 24332
rect 24464 24266 24728 24276
rect 24668 24052 24724 24062
rect 24668 23958 24724 23996
rect 25452 24052 25508 24558
rect 25452 23986 25508 23996
rect 24220 23202 24276 23212
rect 24464 22764 24728 22774
rect 24520 22708 24568 22764
rect 24624 22708 24672 22764
rect 24464 22698 24728 22708
rect 24892 22370 24948 22382
rect 24892 22318 24894 22370
rect 24946 22318 24948 22370
rect 23804 21980 24068 21990
rect 23860 21924 23908 21980
rect 23964 21924 24012 21980
rect 23804 21914 24068 21924
rect 24464 21196 24728 21206
rect 24520 21140 24568 21196
rect 24624 21140 24672 21196
rect 24464 21130 24728 21140
rect 23804 20412 24068 20422
rect 23860 20356 23908 20412
rect 23964 20356 24012 20412
rect 23804 20346 24068 20356
rect 24464 19628 24728 19638
rect 24520 19572 24568 19628
rect 24624 19572 24672 19628
rect 24464 19562 24728 19572
rect 23804 18844 24068 18854
rect 23860 18788 23908 18844
rect 23964 18788 24012 18844
rect 23804 18778 24068 18788
rect 24464 18060 24728 18070
rect 24520 18004 24568 18060
rect 24624 18004 24672 18060
rect 24464 17994 24728 18004
rect 23804 17276 24068 17286
rect 23860 17220 23908 17276
rect 23964 17220 24012 17276
rect 23804 17210 24068 17220
rect 24464 16492 24728 16502
rect 24520 16436 24568 16492
rect 24624 16436 24672 16492
rect 24464 16426 24728 16436
rect 23804 15708 24068 15718
rect 23860 15652 23908 15708
rect 23964 15652 24012 15708
rect 23804 15642 24068 15652
rect 24464 14924 24728 14934
rect 24520 14868 24568 14924
rect 24624 14868 24672 14924
rect 24464 14858 24728 14868
rect 24892 14756 24948 22318
rect 24892 14690 24948 14700
rect 25004 22260 25060 22270
rect 23804 14140 24068 14150
rect 23860 14084 23908 14140
rect 23964 14084 24012 14140
rect 23804 14074 24068 14084
rect 24464 13356 24728 13366
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24464 13290 24728 13300
rect 23804 12572 24068 12582
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 23804 12506 24068 12516
rect 24464 11788 24728 11798
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24464 11722 24728 11732
rect 23436 11218 23492 11228
rect 23804 11004 24068 11014
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 23804 10938 24068 10948
rect 25004 10612 25060 22204
rect 25564 13076 25620 25452
rect 25676 25282 25732 25294
rect 25676 25230 25678 25282
rect 25730 25230 25732 25282
rect 25676 24948 25732 25230
rect 25676 24882 25732 24892
rect 25676 23714 25732 23726
rect 25676 23662 25678 23714
rect 25730 23662 25732 23714
rect 25676 23156 25732 23662
rect 25676 23090 25732 23100
rect 25676 22146 25732 22158
rect 25676 22094 25678 22146
rect 25730 22094 25732 22146
rect 25676 21812 25732 22094
rect 25676 21746 25732 21756
rect 25564 13010 25620 13020
rect 25900 12964 25956 30156
rect 26012 19796 26068 45836
rect 26236 45826 26292 45836
rect 26236 44996 26292 45006
rect 26236 44902 26292 44940
rect 26236 44324 26292 44334
rect 26236 44230 26292 44268
rect 26236 43428 26292 43438
rect 26236 43334 26292 43372
rect 26348 43092 26404 46622
rect 26572 44884 26628 47404
rect 26572 44818 26628 44828
rect 26796 44660 26852 53676
rect 27020 53172 27076 54350
rect 27244 54068 27300 55022
rect 27244 54002 27300 54012
rect 27020 53106 27076 53116
rect 27244 53506 27300 53518
rect 27244 53454 27246 53506
rect 27298 53454 27300 53506
rect 27132 53058 27188 53070
rect 27132 53006 27134 53058
rect 27186 53006 27188 53058
rect 26012 19730 26068 19740
rect 26124 43036 26404 43092
rect 26572 44604 26852 44660
rect 26908 52948 26964 52958
rect 25900 12898 25956 12908
rect 26012 16772 26068 16782
rect 25004 10546 25060 10556
rect 24464 10220 24728 10230
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24464 10154 24728 10164
rect 23804 9436 24068 9446
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 23804 9370 24068 9380
rect 24464 8652 24728 8662
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24464 8586 24728 8596
rect 23804 7868 24068 7878
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 23804 7802 24068 7812
rect 24464 7084 24728 7094
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 24464 7018 24728 7028
rect 23804 6300 24068 6310
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 23804 6234 24068 6244
rect 24464 5516 24728 5526
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24464 5450 24728 5460
rect 23804 4732 24068 4742
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 23804 4666 24068 4676
rect 24464 3948 24728 3958
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24464 3882 24728 3892
rect 22988 3378 23044 3388
rect 23804 3164 24068 3174
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 23804 3098 24068 3108
rect 24464 2380 24728 2390
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24464 2314 24728 2324
rect 24892 1652 24948 1662
rect 23804 1596 24068 1606
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 23804 1530 24068 1540
rect 22876 242 22932 252
rect 23548 1316 23604 1326
rect 23548 112 23604 1260
rect 24464 812 24728 822
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24464 746 24728 756
rect 24892 112 24948 1596
rect 26012 1540 26068 16716
rect 26124 8148 26180 43036
rect 26236 42756 26292 42766
rect 26236 42662 26292 42700
rect 26460 42644 26516 42654
rect 26236 41860 26292 41870
rect 26236 41766 26292 41804
rect 26236 41188 26292 41198
rect 26236 41094 26292 41132
rect 26236 40516 26292 40526
rect 26236 40402 26292 40460
rect 26236 40350 26238 40402
rect 26290 40350 26292 40402
rect 26236 40338 26292 40350
rect 26236 39618 26292 39630
rect 26236 39566 26238 39618
rect 26290 39566 26292 39618
rect 26236 39060 26292 39566
rect 26236 38994 26292 39004
rect 26236 38836 26292 38846
rect 26236 38742 26292 38780
rect 26348 38276 26404 38286
rect 26236 38052 26292 38062
rect 26236 37958 26292 37996
rect 26236 37492 26292 37502
rect 26236 37266 26292 37436
rect 26236 37214 26238 37266
rect 26290 37214 26292 37266
rect 26236 37202 26292 37214
rect 26348 36482 26404 38220
rect 26348 36430 26350 36482
rect 26402 36430 26404 36482
rect 26348 36418 26404 36430
rect 26348 35924 26404 35934
rect 26236 35588 26292 35598
rect 26236 35494 26292 35532
rect 26236 34916 26292 34926
rect 26236 34822 26292 34860
rect 26236 34020 26292 34030
rect 26236 33926 26292 33964
rect 26348 33796 26404 35868
rect 26236 33740 26404 33796
rect 26236 32562 26292 33740
rect 26236 32510 26238 32562
rect 26290 32510 26292 32562
rect 26236 32498 26292 32510
rect 26348 33346 26404 33358
rect 26348 33294 26350 33346
rect 26402 33294 26404 33346
rect 26348 32452 26404 33294
rect 26348 32386 26404 32396
rect 26348 31778 26404 31790
rect 26348 31726 26350 31778
rect 26402 31726 26404 31778
rect 26236 30884 26292 30894
rect 26236 30790 26292 30828
rect 26236 30212 26292 30222
rect 26236 30118 26292 30156
rect 26236 29316 26292 29326
rect 26236 29222 26292 29260
rect 26236 28756 26292 28766
rect 26236 28662 26292 28700
rect 26348 28084 26404 31726
rect 26348 28018 26404 28028
rect 26348 27858 26404 27870
rect 26348 27806 26350 27858
rect 26402 27806 26404 27858
rect 26236 27074 26292 27086
rect 26236 27022 26238 27074
rect 26290 27022 26292 27074
rect 26236 26964 26292 27022
rect 26236 26898 26292 26908
rect 26348 26404 26404 27806
rect 26348 26338 26404 26348
rect 26236 26180 26292 26190
rect 26236 26086 26292 26124
rect 26236 25508 26292 25518
rect 26236 25414 26292 25452
rect 26348 24836 26404 24846
rect 26236 24724 26292 24734
rect 26236 24630 26292 24668
rect 26236 23940 26292 23950
rect 26236 23846 26292 23884
rect 26348 23716 26404 24780
rect 26236 23660 26404 23716
rect 26236 22482 26292 23660
rect 26236 22430 26238 22482
rect 26290 22430 26292 22482
rect 26236 22418 26292 22430
rect 26348 23154 26404 23166
rect 26348 23102 26350 23154
rect 26402 23102 26404 23154
rect 26236 21476 26292 21486
rect 26236 21382 26292 21420
rect 26348 12292 26404 23102
rect 26460 21028 26516 42588
rect 26572 26908 26628 44604
rect 26684 44436 26740 44446
rect 26684 31108 26740 44380
rect 26908 43708 26964 52892
rect 27132 51380 27188 53006
rect 27244 52276 27300 53454
rect 27244 52210 27300 52220
rect 27132 51314 27188 51324
rect 27244 51938 27300 51950
rect 27244 51886 27246 51938
rect 27298 51886 27300 51938
rect 27020 51266 27076 51278
rect 27020 51214 27022 51266
rect 27074 51214 27076 51266
rect 27020 50036 27076 51214
rect 27244 50932 27300 51886
rect 27244 50866 27300 50876
rect 27020 49970 27076 49980
rect 27244 50370 27300 50382
rect 27244 50318 27246 50370
rect 27298 50318 27300 50370
rect 27132 49922 27188 49934
rect 27132 49870 27134 49922
rect 27186 49870 27188 49922
rect 27132 48244 27188 49870
rect 27244 49140 27300 50318
rect 27244 49074 27300 49084
rect 27468 49252 27524 49262
rect 27132 48178 27188 48188
rect 27244 48802 27300 48814
rect 27244 48750 27246 48802
rect 27298 48750 27300 48802
rect 27020 48130 27076 48142
rect 27020 48078 27022 48130
rect 27074 48078 27076 48130
rect 27020 46900 27076 48078
rect 27244 47796 27300 48750
rect 27244 47730 27300 47740
rect 27356 48020 27412 48030
rect 27020 46834 27076 46844
rect 27244 47234 27300 47246
rect 27244 47182 27246 47234
rect 27298 47182 27300 47234
rect 27132 46786 27188 46798
rect 27132 46734 27134 46786
rect 27186 46734 27188 46786
rect 27132 45108 27188 46734
rect 27244 46004 27300 47182
rect 27244 45938 27300 45948
rect 27132 45042 27188 45052
rect 27244 45666 27300 45678
rect 27244 45614 27246 45666
rect 27298 45614 27300 45666
rect 27020 44994 27076 45006
rect 27020 44942 27022 44994
rect 27074 44942 27076 44994
rect 27020 43876 27076 44942
rect 27244 44660 27300 45614
rect 27244 44594 27300 44604
rect 27356 44436 27412 47964
rect 27020 43810 27076 43820
rect 27132 44380 27412 44436
rect 26908 43652 27076 43708
rect 26796 43316 26852 43326
rect 26796 43314 26964 43316
rect 26796 43262 26798 43314
rect 26850 43262 26964 43314
rect 26796 43260 26964 43262
rect 26796 43250 26852 43260
rect 26908 41972 26964 43260
rect 26908 41906 26964 41916
rect 26796 41748 26852 41758
rect 26796 41746 26964 41748
rect 26796 41694 26798 41746
rect 26850 41694 26964 41746
rect 26796 41692 26964 41694
rect 26796 41682 26852 41692
rect 26908 40628 26964 41692
rect 26908 40562 26964 40572
rect 26796 40180 26852 40190
rect 26796 40178 26964 40180
rect 26796 40126 26798 40178
rect 26850 40126 26964 40178
rect 26796 40124 26964 40126
rect 26796 40114 26852 40124
rect 26908 39172 26964 40124
rect 26908 39106 26964 39116
rect 26908 38946 26964 38958
rect 26908 38894 26910 38946
rect 26962 38894 26964 38946
rect 26908 37492 26964 38894
rect 26908 37426 26964 37436
rect 26796 37044 26852 37054
rect 26796 37042 26964 37044
rect 26796 36990 26798 37042
rect 26850 36990 26964 37042
rect 26796 36988 26964 36990
rect 26796 36978 26852 36988
rect 26908 36036 26964 36988
rect 26908 35970 26964 35980
rect 26908 35810 26964 35822
rect 26908 35758 26910 35810
rect 26962 35758 26964 35810
rect 26908 34356 26964 35758
rect 26908 34290 26964 34300
rect 26796 33908 26852 33918
rect 26796 33906 26964 33908
rect 26796 33854 26798 33906
rect 26850 33854 26964 33906
rect 26796 33852 26964 33854
rect 26796 33842 26852 33852
rect 26908 32900 26964 33852
rect 26908 32834 26964 32844
rect 26908 32674 26964 32686
rect 26908 32622 26910 32674
rect 26962 32622 26964 32674
rect 26908 31892 26964 32622
rect 26908 31826 26964 31836
rect 26684 31042 26740 31052
rect 26908 31666 26964 31678
rect 26908 31614 26910 31666
rect 26962 31614 26964 31666
rect 26908 30324 26964 31614
rect 26908 30258 26964 30268
rect 26908 30098 26964 30110
rect 26908 30046 26910 30098
rect 26962 30046 26964 30098
rect 26908 29428 26964 30046
rect 26908 29362 26964 29372
rect 26572 26852 26740 26908
rect 26460 20972 26628 21028
rect 26572 12740 26628 20972
rect 26684 18452 26740 26852
rect 26684 18386 26740 18396
rect 26572 12674 26628 12684
rect 26348 12226 26404 12236
rect 26124 8082 26180 8092
rect 26236 11284 26292 11294
rect 26012 1474 26068 1484
rect 26236 112 26292 11228
rect 27020 4564 27076 43652
rect 27020 4498 27076 4508
rect 27132 1652 27188 44380
rect 27244 44098 27300 44110
rect 27244 44046 27246 44098
rect 27298 44046 27300 44098
rect 27244 42868 27300 44046
rect 27244 42802 27300 42812
rect 27244 42530 27300 42542
rect 27244 42478 27246 42530
rect 27298 42478 27300 42530
rect 27244 41524 27300 42478
rect 27244 41458 27300 41468
rect 27244 40962 27300 40974
rect 27244 40910 27246 40962
rect 27298 40910 27300 40962
rect 27244 39732 27300 40910
rect 27244 39666 27300 39676
rect 27244 39394 27300 39406
rect 27244 39342 27246 39394
rect 27298 39342 27300 39394
rect 27244 38388 27300 39342
rect 27244 38322 27300 38332
rect 27356 39396 27412 39406
rect 27244 37826 27300 37838
rect 27244 37774 27246 37826
rect 27298 37774 27300 37826
rect 27244 36596 27300 37774
rect 27244 36530 27300 36540
rect 27244 36258 27300 36270
rect 27244 36206 27246 36258
rect 27298 36206 27300 36258
rect 27244 35252 27300 36206
rect 27244 35186 27300 35196
rect 27244 34690 27300 34702
rect 27244 34638 27246 34690
rect 27298 34638 27300 34690
rect 27244 33460 27300 34638
rect 27244 33394 27300 33404
rect 27244 33122 27300 33134
rect 27244 33070 27246 33122
rect 27298 33070 27300 33122
rect 27244 32340 27300 33070
rect 27244 32274 27300 32284
rect 27356 32116 27412 39340
rect 27244 32060 27412 32116
rect 27244 31332 27300 32060
rect 27468 31948 27524 49196
rect 27356 31892 27524 31948
rect 28140 35140 28196 35150
rect 28028 31892 28084 31902
rect 27356 31444 27412 31892
rect 27804 31556 27860 31566
rect 27356 31388 27748 31444
rect 27244 31266 27300 31276
rect 27468 31220 27524 31230
rect 27244 31106 27300 31118
rect 27244 31054 27246 31106
rect 27298 31054 27300 31106
rect 27244 29876 27300 31054
rect 27244 29810 27300 29820
rect 27244 29538 27300 29550
rect 27244 29486 27246 29538
rect 27298 29486 27300 29538
rect 27244 28980 27300 29486
rect 27244 28914 27300 28924
rect 27244 28532 27300 28542
rect 27244 28438 27300 28476
rect 27244 28084 27300 28094
rect 27244 27990 27300 28028
rect 27244 27636 27300 27646
rect 27244 26962 27300 27580
rect 27244 26910 27246 26962
rect 27298 26910 27300 26962
rect 27244 26898 27300 26910
rect 27468 26908 27524 31164
rect 27468 26852 27636 26908
rect 27244 26740 27300 26750
rect 27244 26514 27300 26684
rect 27244 26462 27246 26514
rect 27298 26462 27300 26514
rect 27244 26450 27300 26462
rect 27244 25844 27300 25854
rect 27244 25394 27300 25788
rect 27244 25342 27246 25394
rect 27298 25342 27300 25394
rect 27244 25330 27300 25342
rect 27356 25396 27412 25406
rect 27244 24948 27300 24958
rect 27356 24948 27412 25340
rect 27244 24946 27412 24948
rect 27244 24894 27246 24946
rect 27298 24894 27412 24946
rect 27244 24892 27412 24894
rect 27244 24882 27300 24892
rect 27244 24500 27300 24510
rect 27244 23826 27300 24444
rect 27244 23774 27246 23826
rect 27298 23774 27300 23826
rect 27244 23762 27300 23774
rect 27356 23604 27412 23614
rect 27244 23380 27300 23390
rect 27356 23380 27412 23548
rect 27244 23378 27412 23380
rect 27244 23326 27246 23378
rect 27298 23326 27412 23378
rect 27244 23324 27412 23326
rect 27244 23314 27300 23324
rect 27244 22708 27300 22718
rect 27244 22258 27300 22652
rect 27244 22206 27246 22258
rect 27298 22206 27300 22258
rect 27244 22194 27300 22206
rect 27356 22260 27412 22270
rect 27244 21812 27300 21822
rect 27356 21812 27412 22204
rect 27244 21810 27412 21812
rect 27244 21758 27246 21810
rect 27298 21758 27412 21810
rect 27244 21756 27412 21758
rect 27244 21746 27300 21756
rect 27468 21700 27524 21710
rect 27356 21140 27412 21150
rect 27356 3332 27412 21084
rect 27468 16884 27524 21644
rect 27468 16818 27524 16828
rect 27580 13972 27636 26852
rect 27692 21140 27748 31388
rect 27692 21074 27748 21084
rect 27804 20468 27860 31500
rect 28028 31220 28084 31836
rect 28028 31154 28084 31164
rect 27804 20402 27860 20412
rect 27916 21588 27972 21598
rect 27916 15540 27972 21532
rect 27916 15474 27972 15484
rect 27580 13906 27636 13916
rect 28140 11956 28196 35084
rect 28252 24164 28308 24174
rect 28308 24108 28420 24164
rect 28252 24098 28308 24108
rect 28140 11890 28196 11900
rect 28252 16324 28308 16334
rect 28252 8428 28308 16268
rect 28364 11508 28420 24108
rect 28364 11442 28420 11452
rect 28252 8372 28532 8428
rect 28420 8316 28532 8372
rect 28364 8306 28420 8316
rect 27356 3266 27412 3276
rect 27132 1586 27188 1596
rect 27580 1540 27636 1550
rect 27580 112 27636 1484
rect 18844 28 19236 84
rect 19488 0 19600 112
rect 20832 0 20944 112
rect 22176 0 22288 112
rect 23520 0 23632 112
rect 24864 0 24976 112
rect 26208 0 26320 112
rect 27552 0 27664 112
<< via2 >>
rect 364 53564 420 53620
rect 252 36092 308 36148
rect 140 29148 196 29204
rect 252 26124 308 26180
rect 4732 57260 4788 57316
rect 5516 57260 5572 57316
rect 3804 56474 3860 56476
rect 3804 56422 3806 56474
rect 3806 56422 3858 56474
rect 3858 56422 3860 56474
rect 3804 56420 3860 56422
rect 3908 56474 3964 56476
rect 3908 56422 3910 56474
rect 3910 56422 3962 56474
rect 3962 56422 3964 56474
rect 3908 56420 3964 56422
rect 4012 56474 4068 56476
rect 4012 56422 4014 56474
rect 4014 56422 4066 56474
rect 4066 56422 4068 56474
rect 4012 56420 4068 56422
rect 3052 55970 3108 55972
rect 3052 55918 3054 55970
rect 3054 55918 3106 55970
rect 3106 55918 3108 55970
rect 3052 55916 3108 55918
rect 4464 55690 4520 55692
rect 4464 55638 4466 55690
rect 4466 55638 4518 55690
rect 4518 55638 4520 55690
rect 4464 55636 4520 55638
rect 4568 55690 4624 55692
rect 4568 55638 4570 55690
rect 4570 55638 4622 55690
rect 4622 55638 4624 55690
rect 4568 55636 4624 55638
rect 4672 55690 4728 55692
rect 4672 55638 4674 55690
rect 4674 55638 4726 55690
rect 4726 55638 4728 55690
rect 4672 55636 4728 55638
rect 1372 52892 1428 52948
rect 1820 52220 1876 52276
rect 1484 42924 1540 42980
rect 812 40124 868 40180
rect 588 38780 644 38836
rect 476 36988 532 37044
rect 476 28028 532 28084
rect 588 28700 644 28756
rect 588 19740 644 19796
rect 700 30940 756 30996
rect 364 19292 420 19348
rect 1260 37548 1316 37604
rect 812 29260 868 29316
rect 924 37436 980 37492
rect 1036 37042 1092 37044
rect 1036 36990 1038 37042
rect 1038 36990 1090 37042
rect 1090 36990 1092 37042
rect 1036 36988 1092 36990
rect 1708 41244 1764 41300
rect 1708 40402 1764 40404
rect 1708 40350 1710 40402
rect 1710 40350 1762 40402
rect 1762 40350 1764 40402
rect 1708 40348 1764 40350
rect 1708 38668 1764 38724
rect 1708 38556 1764 38612
rect 1596 37996 1652 38052
rect 1596 36876 1652 36932
rect 1708 36540 1764 36596
rect 924 27692 980 27748
rect 1708 34300 1764 34356
rect 1708 33180 1764 33236
rect 1260 32508 1316 32564
rect 1260 31612 1316 31668
rect 1260 30994 1316 30996
rect 1260 30942 1262 30994
rect 1262 30942 1314 30994
rect 1314 30942 1316 30994
rect 1260 30940 1316 30942
rect 1148 30156 1204 30212
rect 812 20524 868 20580
rect 924 26908 980 26964
rect 700 13804 756 13860
rect 140 13244 196 13300
rect 1596 32562 1652 32564
rect 1596 32510 1598 32562
rect 1598 32510 1650 32562
rect 1650 32510 1652 32562
rect 1596 32508 1652 32510
rect 1932 50876 1988 50932
rect 3276 46844 3332 46900
rect 2268 44940 2324 44996
rect 1932 40572 1988 40628
rect 2044 42028 2100 42084
rect 1932 40348 1988 40404
rect 2156 40572 2212 40628
rect 2156 40236 2212 40292
rect 3804 54906 3860 54908
rect 3804 54854 3806 54906
rect 3806 54854 3858 54906
rect 3858 54854 3860 54906
rect 3804 54852 3860 54854
rect 3908 54906 3964 54908
rect 3908 54854 3910 54906
rect 3910 54854 3962 54906
rect 3962 54854 3964 54906
rect 3908 54852 3964 54854
rect 4012 54906 4068 54908
rect 4012 54854 4014 54906
rect 4014 54854 4066 54906
rect 4066 54854 4068 54906
rect 4012 54852 4068 54854
rect 4464 54122 4520 54124
rect 4464 54070 4466 54122
rect 4466 54070 4518 54122
rect 4518 54070 4520 54122
rect 4464 54068 4520 54070
rect 4568 54122 4624 54124
rect 4568 54070 4570 54122
rect 4570 54070 4622 54122
rect 4622 54070 4624 54122
rect 4568 54068 4624 54070
rect 4672 54122 4728 54124
rect 4672 54070 4674 54122
rect 4674 54070 4726 54122
rect 4726 54070 4728 54122
rect 4672 54068 4728 54070
rect 3804 53338 3860 53340
rect 3804 53286 3806 53338
rect 3806 53286 3858 53338
rect 3858 53286 3860 53338
rect 3804 53284 3860 53286
rect 3908 53338 3964 53340
rect 3908 53286 3910 53338
rect 3910 53286 3962 53338
rect 3962 53286 3964 53338
rect 3908 53284 3964 53286
rect 4012 53338 4068 53340
rect 4012 53286 4014 53338
rect 4014 53286 4066 53338
rect 4066 53286 4068 53338
rect 4012 53284 4068 53286
rect 6300 53004 6356 53060
rect 4464 52554 4520 52556
rect 4464 52502 4466 52554
rect 4466 52502 4518 52554
rect 4518 52502 4520 52554
rect 4464 52500 4520 52502
rect 4568 52554 4624 52556
rect 4568 52502 4570 52554
rect 4570 52502 4622 52554
rect 4622 52502 4624 52554
rect 4568 52500 4624 52502
rect 4672 52554 4728 52556
rect 4672 52502 4674 52554
rect 4674 52502 4726 52554
rect 4726 52502 4728 52554
rect 4672 52500 4728 52502
rect 5964 51884 6020 51940
rect 3804 51770 3860 51772
rect 3804 51718 3806 51770
rect 3806 51718 3858 51770
rect 3858 51718 3860 51770
rect 3804 51716 3860 51718
rect 3908 51770 3964 51772
rect 3908 51718 3910 51770
rect 3910 51718 3962 51770
rect 3962 51718 3964 51770
rect 3908 51716 3964 51718
rect 4012 51770 4068 51772
rect 4012 51718 4014 51770
rect 4014 51718 4066 51770
rect 4066 51718 4068 51770
rect 4012 51716 4068 51718
rect 4172 51324 4228 51380
rect 3804 50202 3860 50204
rect 3804 50150 3806 50202
rect 3806 50150 3858 50202
rect 3858 50150 3860 50202
rect 3804 50148 3860 50150
rect 3908 50202 3964 50204
rect 3908 50150 3910 50202
rect 3910 50150 3962 50202
rect 3962 50150 3964 50202
rect 3908 50148 3964 50150
rect 4012 50202 4068 50204
rect 4012 50150 4014 50202
rect 4014 50150 4066 50202
rect 4066 50150 4068 50202
rect 4012 50148 4068 50150
rect 3804 48634 3860 48636
rect 3804 48582 3806 48634
rect 3806 48582 3858 48634
rect 3858 48582 3860 48634
rect 3804 48580 3860 48582
rect 3908 48634 3964 48636
rect 3908 48582 3910 48634
rect 3910 48582 3962 48634
rect 3962 48582 3964 48634
rect 3908 48580 3964 48582
rect 4012 48634 4068 48636
rect 4012 48582 4014 48634
rect 4014 48582 4066 48634
rect 4066 48582 4068 48634
rect 4012 48580 4068 48582
rect 3804 47066 3860 47068
rect 3804 47014 3806 47066
rect 3806 47014 3858 47066
rect 3858 47014 3860 47066
rect 3804 47012 3860 47014
rect 3908 47066 3964 47068
rect 3908 47014 3910 47066
rect 3910 47014 3962 47066
rect 3962 47014 3964 47066
rect 3908 47012 3964 47014
rect 4012 47066 4068 47068
rect 4012 47014 4014 47066
rect 4014 47014 4066 47066
rect 4066 47014 4068 47066
rect 4012 47012 4068 47014
rect 3804 45498 3860 45500
rect 3804 45446 3806 45498
rect 3806 45446 3858 45498
rect 3858 45446 3860 45498
rect 3804 45444 3860 45446
rect 3908 45498 3964 45500
rect 3908 45446 3910 45498
rect 3910 45446 3962 45498
rect 3962 45446 3964 45498
rect 3908 45444 3964 45446
rect 4012 45498 4068 45500
rect 4012 45446 4014 45498
rect 4014 45446 4066 45498
rect 4066 45446 4068 45498
rect 4012 45444 4068 45446
rect 3804 43930 3860 43932
rect 3804 43878 3806 43930
rect 3806 43878 3858 43930
rect 3858 43878 3860 43930
rect 3804 43876 3860 43878
rect 3908 43930 3964 43932
rect 3908 43878 3910 43930
rect 3910 43878 3962 43930
rect 3962 43878 3964 43930
rect 3908 43876 3964 43878
rect 4012 43930 4068 43932
rect 4012 43878 4014 43930
rect 4014 43878 4066 43930
rect 4066 43878 4068 43930
rect 4012 43876 4068 43878
rect 3500 43596 3556 43652
rect 3804 42362 3860 42364
rect 3804 42310 3806 42362
rect 3806 42310 3858 42362
rect 3858 42310 3860 42362
rect 3804 42308 3860 42310
rect 3908 42362 3964 42364
rect 3908 42310 3910 42362
rect 3910 42310 3962 42362
rect 3962 42310 3964 42362
rect 3908 42308 3964 42310
rect 4012 42362 4068 42364
rect 4012 42310 4014 42362
rect 4014 42310 4066 42362
rect 4066 42310 4068 42362
rect 4012 42308 4068 42310
rect 4464 50986 4520 50988
rect 4464 50934 4466 50986
rect 4466 50934 4518 50986
rect 4518 50934 4520 50986
rect 4464 50932 4520 50934
rect 4568 50986 4624 50988
rect 4568 50934 4570 50986
rect 4570 50934 4622 50986
rect 4622 50934 4624 50986
rect 4568 50932 4624 50934
rect 4672 50986 4728 50988
rect 4672 50934 4674 50986
rect 4674 50934 4726 50986
rect 4726 50934 4728 50986
rect 4672 50932 4728 50934
rect 5740 49532 5796 49588
rect 4464 49418 4520 49420
rect 4464 49366 4466 49418
rect 4466 49366 4518 49418
rect 4518 49366 4520 49418
rect 4464 49364 4520 49366
rect 4568 49418 4624 49420
rect 4568 49366 4570 49418
rect 4570 49366 4622 49418
rect 4622 49366 4624 49418
rect 4568 49364 4624 49366
rect 4672 49418 4728 49420
rect 4672 49366 4674 49418
rect 4674 49366 4726 49418
rect 4726 49366 4728 49418
rect 4672 49364 4728 49366
rect 4464 47850 4520 47852
rect 4464 47798 4466 47850
rect 4466 47798 4518 47850
rect 4518 47798 4520 47850
rect 4464 47796 4520 47798
rect 4568 47850 4624 47852
rect 4568 47798 4570 47850
rect 4570 47798 4622 47850
rect 4622 47798 4624 47850
rect 4568 47796 4624 47798
rect 4672 47850 4728 47852
rect 4672 47798 4674 47850
rect 4674 47798 4726 47850
rect 4726 47798 4728 47850
rect 4672 47796 4728 47798
rect 4464 46282 4520 46284
rect 4464 46230 4466 46282
rect 4466 46230 4518 46282
rect 4518 46230 4520 46282
rect 4464 46228 4520 46230
rect 4568 46282 4624 46284
rect 4568 46230 4570 46282
rect 4570 46230 4622 46282
rect 4622 46230 4624 46282
rect 4568 46228 4624 46230
rect 4672 46282 4728 46284
rect 4672 46230 4674 46282
rect 4674 46230 4726 46282
rect 4726 46230 4728 46282
rect 4672 46228 4728 46230
rect 4464 44714 4520 44716
rect 4464 44662 4466 44714
rect 4466 44662 4518 44714
rect 4518 44662 4520 44714
rect 4464 44660 4520 44662
rect 4568 44714 4624 44716
rect 4568 44662 4570 44714
rect 4570 44662 4622 44714
rect 4622 44662 4624 44714
rect 4568 44660 4624 44662
rect 4672 44714 4728 44716
rect 4672 44662 4674 44714
rect 4674 44662 4726 44714
rect 4726 44662 4728 44714
rect 4672 44660 4728 44662
rect 4464 43146 4520 43148
rect 4464 43094 4466 43146
rect 4466 43094 4518 43146
rect 4518 43094 4520 43146
rect 4464 43092 4520 43094
rect 4568 43146 4624 43148
rect 4568 43094 4570 43146
rect 4570 43094 4622 43146
rect 4622 43094 4624 43146
rect 4568 43092 4624 43094
rect 4672 43146 4728 43148
rect 4672 43094 4674 43146
rect 4674 43094 4726 43146
rect 4726 43094 4728 43146
rect 4672 43092 4728 43094
rect 4464 41578 4520 41580
rect 4464 41526 4466 41578
rect 4466 41526 4518 41578
rect 4518 41526 4520 41578
rect 4464 41524 4520 41526
rect 4568 41578 4624 41580
rect 4568 41526 4570 41578
rect 4570 41526 4622 41578
rect 4622 41526 4624 41578
rect 4568 41524 4624 41526
rect 4672 41578 4728 41580
rect 4672 41526 4674 41578
rect 4674 41526 4726 41578
rect 4726 41526 4728 41578
rect 4672 41524 4728 41526
rect 5292 41356 5348 41412
rect 4284 41298 4340 41300
rect 4284 41246 4286 41298
rect 4286 41246 4338 41298
rect 4338 41246 4340 41298
rect 4284 41244 4340 41246
rect 3276 41132 3332 41188
rect 1932 37212 1988 37268
rect 2380 38162 2436 38164
rect 2380 38110 2382 38162
rect 2382 38110 2434 38162
rect 2434 38110 2436 38162
rect 2380 38108 2436 38110
rect 2268 37212 2324 37268
rect 1932 36652 1988 36708
rect 2044 36540 2100 36596
rect 1932 33180 1988 33236
rect 1708 31612 1764 31668
rect 1820 31164 1876 31220
rect 1596 29314 1652 29316
rect 1596 29262 1598 29314
rect 1598 29262 1650 29314
rect 1650 29262 1652 29314
rect 1596 29260 1652 29262
rect 1484 29148 1540 29204
rect 1596 28754 1652 28756
rect 1596 28702 1598 28754
rect 1598 28702 1650 28754
rect 1650 28702 1652 28754
rect 1596 28700 1652 28702
rect 1820 28588 1876 28644
rect 1260 27074 1316 27076
rect 1260 27022 1262 27074
rect 1262 27022 1314 27074
rect 1314 27022 1316 27074
rect 1260 27020 1316 27022
rect 1484 27692 1540 27748
rect 1036 26124 1092 26180
rect 1708 27020 1764 27076
rect 1484 26012 1540 26068
rect 1148 24892 1204 24948
rect 1260 24722 1316 24724
rect 1260 24670 1262 24722
rect 1262 24670 1314 24722
rect 1314 24670 1316 24722
rect 1260 24668 1316 24670
rect 1708 25452 1764 25508
rect 1708 23212 1764 23268
rect 1596 23154 1652 23156
rect 1596 23102 1598 23154
rect 1598 23102 1650 23154
rect 1650 23102 1652 23154
rect 1596 23100 1652 23102
rect 1596 22428 1652 22484
rect 2268 32396 2324 32452
rect 2044 32060 2100 32116
rect 2268 32060 2324 32116
rect 2716 38946 2772 38948
rect 2716 38894 2718 38946
rect 2718 38894 2770 38946
rect 2770 38894 2772 38946
rect 2716 38892 2772 38894
rect 3164 39730 3220 39732
rect 3164 39678 3166 39730
rect 3166 39678 3218 39730
rect 3218 39678 3220 39730
rect 3164 39676 3220 39678
rect 2604 38108 2660 38164
rect 2716 37772 2772 37828
rect 2492 37378 2548 37380
rect 2492 37326 2494 37378
rect 2494 37326 2546 37378
rect 2546 37326 2548 37378
rect 2492 37324 2548 37326
rect 2716 37548 2772 37604
rect 3164 37884 3220 37940
rect 2604 36428 2660 36484
rect 3052 36652 3108 36708
rect 2492 34188 2548 34244
rect 2156 30156 2212 30212
rect 2044 29484 2100 29540
rect 2044 26178 2100 26180
rect 2044 26126 2046 26178
rect 2046 26126 2098 26178
rect 2098 26126 2100 26178
rect 2044 26124 2100 26126
rect 2044 25564 2100 25620
rect 2380 30716 2436 30772
rect 2268 29820 2324 29876
rect 2604 32396 2660 32452
rect 2268 29596 2324 29652
rect 2044 24108 2100 24164
rect 2268 23772 2324 23828
rect 2156 23660 2212 23716
rect 1932 22540 1988 22596
rect 2044 23548 2100 23604
rect 1932 20914 1988 20916
rect 1932 20862 1934 20914
rect 1934 20862 1986 20914
rect 1986 20862 1988 20914
rect 1932 20860 1988 20862
rect 2828 32060 2884 32116
rect 2828 31890 2884 31892
rect 2828 31838 2830 31890
rect 2830 31838 2882 31890
rect 2882 31838 2884 31890
rect 2828 31836 2884 31838
rect 2716 31778 2772 31780
rect 2716 31726 2718 31778
rect 2718 31726 2770 31778
rect 2770 31726 2772 31778
rect 2716 31724 2772 31726
rect 3804 40794 3860 40796
rect 3804 40742 3806 40794
rect 3806 40742 3858 40794
rect 3858 40742 3860 40794
rect 3804 40740 3860 40742
rect 3908 40794 3964 40796
rect 3908 40742 3910 40794
rect 3910 40742 3962 40794
rect 3962 40742 3964 40794
rect 3908 40740 3964 40742
rect 4012 40794 4068 40796
rect 4012 40742 4014 40794
rect 4014 40742 4066 40794
rect 4066 40742 4068 40794
rect 4012 40740 4068 40742
rect 4284 40402 4340 40404
rect 4284 40350 4286 40402
rect 4286 40350 4338 40402
rect 4338 40350 4340 40402
rect 4284 40348 4340 40350
rect 5068 40124 5124 40180
rect 4464 40010 4520 40012
rect 4464 39958 4466 40010
rect 4466 39958 4518 40010
rect 4518 39958 4520 40010
rect 4464 39956 4520 39958
rect 4568 40010 4624 40012
rect 4568 39958 4570 40010
rect 4570 39958 4622 40010
rect 4622 39958 4624 40010
rect 4568 39956 4624 39958
rect 4672 40010 4728 40012
rect 4672 39958 4674 40010
rect 4674 39958 4726 40010
rect 4726 39958 4728 40010
rect 4672 39956 4728 39958
rect 5292 39900 5348 39956
rect 3804 39226 3860 39228
rect 3804 39174 3806 39226
rect 3806 39174 3858 39226
rect 3858 39174 3860 39226
rect 3804 39172 3860 39174
rect 3908 39226 3964 39228
rect 3908 39174 3910 39226
rect 3910 39174 3962 39226
rect 3962 39174 3964 39226
rect 3908 39172 3964 39174
rect 4012 39226 4068 39228
rect 4012 39174 4014 39226
rect 4014 39174 4066 39226
rect 4066 39174 4068 39226
rect 4012 39172 4068 39174
rect 3612 38892 3668 38948
rect 5180 38892 5236 38948
rect 4284 38834 4340 38836
rect 4284 38782 4286 38834
rect 4286 38782 4338 38834
rect 4338 38782 4340 38834
rect 4284 38780 4340 38782
rect 4464 38442 4520 38444
rect 4464 38390 4466 38442
rect 4466 38390 4518 38442
rect 4518 38390 4520 38442
rect 4464 38388 4520 38390
rect 4568 38442 4624 38444
rect 4568 38390 4570 38442
rect 4570 38390 4622 38442
rect 4622 38390 4624 38442
rect 4568 38388 4624 38390
rect 4672 38442 4728 38444
rect 4672 38390 4674 38442
rect 4674 38390 4726 38442
rect 4726 38390 4728 38442
rect 4672 38388 4728 38390
rect 3500 37212 3556 37268
rect 3388 36482 3444 36484
rect 3388 36430 3390 36482
rect 3390 36430 3442 36482
rect 3442 36430 3444 36482
rect 3388 36428 3444 36430
rect 2828 30828 2884 30884
rect 2492 28588 2548 28644
rect 2604 29484 2660 29540
rect 2828 30044 2884 30100
rect 2716 28700 2772 28756
rect 2604 27916 2660 27972
rect 3276 33516 3332 33572
rect 3500 31724 3556 31780
rect 3804 37658 3860 37660
rect 3804 37606 3806 37658
rect 3806 37606 3858 37658
rect 3858 37606 3860 37658
rect 3804 37604 3860 37606
rect 3908 37658 3964 37660
rect 3908 37606 3910 37658
rect 3910 37606 3962 37658
rect 3962 37606 3964 37658
rect 3908 37604 3964 37606
rect 4012 37658 4068 37660
rect 4012 37606 4014 37658
rect 4014 37606 4066 37658
rect 4066 37606 4068 37658
rect 4012 37604 4068 37606
rect 5068 36988 5124 37044
rect 5628 38946 5684 38948
rect 5628 38894 5630 38946
rect 5630 38894 5682 38946
rect 5682 38894 5684 38946
rect 5628 38892 5684 38894
rect 4464 36874 4520 36876
rect 4464 36822 4466 36874
rect 4466 36822 4518 36874
rect 4518 36822 4520 36874
rect 4464 36820 4520 36822
rect 4568 36874 4624 36876
rect 4568 36822 4570 36874
rect 4570 36822 4622 36874
rect 4622 36822 4624 36874
rect 4568 36820 4624 36822
rect 4672 36874 4728 36876
rect 4672 36822 4674 36874
rect 4674 36822 4726 36874
rect 4726 36822 4728 36874
rect 4672 36820 4728 36822
rect 3948 36594 4004 36596
rect 3948 36542 3950 36594
rect 3950 36542 4002 36594
rect 4002 36542 4004 36594
rect 3948 36540 4004 36542
rect 3804 36090 3860 36092
rect 3804 36038 3806 36090
rect 3806 36038 3858 36090
rect 3858 36038 3860 36090
rect 3804 36036 3860 36038
rect 3908 36090 3964 36092
rect 3908 36038 3910 36090
rect 3910 36038 3962 36090
rect 3962 36038 3964 36090
rect 3908 36036 3964 36038
rect 4012 36090 4068 36092
rect 4012 36038 4014 36090
rect 4014 36038 4066 36090
rect 4066 36038 4068 36090
rect 4012 36036 4068 36038
rect 4464 35306 4520 35308
rect 4464 35254 4466 35306
rect 4466 35254 4518 35306
rect 4518 35254 4520 35306
rect 4464 35252 4520 35254
rect 4568 35306 4624 35308
rect 4568 35254 4570 35306
rect 4570 35254 4622 35306
rect 4622 35254 4624 35306
rect 4568 35252 4624 35254
rect 4672 35306 4728 35308
rect 4672 35254 4674 35306
rect 4674 35254 4726 35306
rect 4726 35254 4728 35306
rect 4672 35252 4728 35254
rect 4284 34914 4340 34916
rect 4284 34862 4286 34914
rect 4286 34862 4338 34914
rect 4338 34862 4340 34914
rect 4284 34860 4340 34862
rect 3804 34522 3860 34524
rect 3804 34470 3806 34522
rect 3806 34470 3858 34522
rect 3858 34470 3860 34522
rect 3804 34468 3860 34470
rect 3908 34522 3964 34524
rect 3908 34470 3910 34522
rect 3910 34470 3962 34522
rect 3962 34470 3964 34522
rect 3908 34468 3964 34470
rect 4012 34522 4068 34524
rect 4012 34470 4014 34522
rect 4014 34470 4066 34522
rect 4066 34470 4068 34522
rect 4012 34468 4068 34470
rect 4284 34130 4340 34132
rect 4284 34078 4286 34130
rect 4286 34078 4338 34130
rect 4338 34078 4340 34130
rect 4284 34076 4340 34078
rect 4464 33738 4520 33740
rect 4464 33686 4466 33738
rect 4466 33686 4518 33738
rect 4518 33686 4520 33738
rect 4464 33684 4520 33686
rect 4568 33738 4624 33740
rect 4568 33686 4570 33738
rect 4570 33686 4622 33738
rect 4622 33686 4624 33738
rect 4568 33684 4624 33686
rect 4672 33738 4728 33740
rect 4672 33686 4674 33738
rect 4674 33686 4726 33738
rect 4726 33686 4728 33738
rect 4672 33684 4728 33686
rect 4172 33516 4228 33572
rect 3804 32954 3860 32956
rect 3804 32902 3806 32954
rect 3806 32902 3858 32954
rect 3858 32902 3860 32954
rect 3804 32900 3860 32902
rect 3908 32954 3964 32956
rect 3908 32902 3910 32954
rect 3910 32902 3962 32954
rect 3962 32902 3964 32954
rect 3908 32900 3964 32902
rect 4012 32954 4068 32956
rect 4012 32902 4014 32954
rect 4014 32902 4066 32954
rect 4066 32902 4068 32954
rect 4012 32900 4068 32902
rect 3724 31836 3780 31892
rect 4060 31778 4116 31780
rect 4060 31726 4062 31778
rect 4062 31726 4114 31778
rect 4114 31726 4116 31778
rect 4060 31724 4116 31726
rect 3804 31386 3860 31388
rect 3804 31334 3806 31386
rect 3806 31334 3858 31386
rect 3858 31334 3860 31386
rect 3804 31332 3860 31334
rect 3908 31386 3964 31388
rect 3908 31334 3910 31386
rect 3910 31334 3962 31386
rect 3962 31334 3964 31386
rect 3908 31332 3964 31334
rect 4012 31386 4068 31388
rect 4012 31334 4014 31386
rect 4014 31334 4066 31386
rect 4066 31334 4068 31386
rect 4012 31332 4068 31334
rect 3948 30044 4004 30100
rect 3804 29818 3860 29820
rect 3804 29766 3806 29818
rect 3806 29766 3858 29818
rect 3858 29766 3860 29818
rect 3804 29764 3860 29766
rect 3908 29818 3964 29820
rect 3908 29766 3910 29818
rect 3910 29766 3962 29818
rect 3962 29766 3964 29818
rect 3908 29764 3964 29766
rect 4012 29818 4068 29820
rect 4012 29766 4014 29818
rect 4014 29766 4066 29818
rect 4066 29766 4068 29818
rect 4012 29764 4068 29766
rect 4060 29484 4116 29540
rect 3500 28530 3556 28532
rect 3500 28478 3502 28530
rect 3502 28478 3554 28530
rect 3554 28478 3556 28530
rect 3500 28476 3556 28478
rect 2492 26796 2548 26852
rect 2828 26850 2884 26852
rect 2828 26798 2830 26850
rect 2830 26798 2882 26850
rect 2882 26798 2884 26850
rect 2828 26796 2884 26798
rect 3388 28028 3444 28084
rect 2828 26124 2884 26180
rect 2716 25340 2772 25396
rect 2828 25228 2884 25284
rect 2268 21644 2324 21700
rect 2156 20972 2212 21028
rect 2156 20748 2212 20804
rect 1708 19852 1764 19908
rect 1596 19458 1652 19460
rect 1596 19406 1598 19458
rect 1598 19406 1650 19458
rect 1650 19406 1652 19458
rect 1596 19404 1652 19406
rect 1596 17052 1652 17108
rect 1148 13858 1204 13860
rect 1148 13806 1150 13858
rect 1150 13806 1202 13858
rect 1202 13806 1204 13858
rect 1148 13804 1204 13806
rect 924 12236 980 12292
rect 1148 13132 1204 13188
rect 1260 10556 1316 10612
rect 1260 9212 1316 9268
rect 1596 15036 1652 15092
rect 2044 17836 2100 17892
rect 2380 20188 2436 20244
rect 2268 18732 2324 18788
rect 2716 22594 2772 22596
rect 2716 22542 2718 22594
rect 2718 22542 2770 22594
rect 2770 22542 2772 22594
rect 2716 22540 2772 22542
rect 3276 25788 3332 25844
rect 3052 25730 3108 25732
rect 3052 25678 3054 25730
rect 3054 25678 3106 25730
rect 3106 25678 3108 25730
rect 3052 25676 3108 25678
rect 3500 26460 3556 26516
rect 4284 32450 4340 32452
rect 4284 32398 4286 32450
rect 4286 32398 4338 32450
rect 4338 32398 4340 32450
rect 4284 32396 4340 32398
rect 4464 32170 4520 32172
rect 4464 32118 4466 32170
rect 4466 32118 4518 32170
rect 4518 32118 4520 32170
rect 4464 32116 4520 32118
rect 4568 32170 4624 32172
rect 4568 32118 4570 32170
rect 4570 32118 4622 32170
rect 4622 32118 4624 32170
rect 4568 32116 4624 32118
rect 4672 32170 4728 32172
rect 4672 32118 4674 32170
rect 4674 32118 4726 32170
rect 4726 32118 4728 32170
rect 4672 32116 4728 32118
rect 4284 31724 4340 31780
rect 4844 31612 4900 31668
rect 4396 31500 4452 31556
rect 4396 31164 4452 31220
rect 4284 30716 4340 30772
rect 4844 30716 4900 30772
rect 4464 30602 4520 30604
rect 4464 30550 4466 30602
rect 4466 30550 4518 30602
rect 4518 30550 4520 30602
rect 4464 30548 4520 30550
rect 4568 30602 4624 30604
rect 4568 30550 4570 30602
rect 4570 30550 4622 30602
rect 4622 30550 4624 30602
rect 4568 30548 4624 30550
rect 4672 30602 4728 30604
rect 4672 30550 4674 30602
rect 4674 30550 4726 30602
rect 4726 30550 4728 30602
rect 4672 30548 4728 30550
rect 4464 29034 4520 29036
rect 4464 28982 4466 29034
rect 4466 28982 4518 29034
rect 4518 28982 4520 29034
rect 4464 28980 4520 28982
rect 4568 29034 4624 29036
rect 4568 28982 4570 29034
rect 4570 28982 4622 29034
rect 4622 28982 4624 29034
rect 4568 28980 4624 28982
rect 4672 29034 4728 29036
rect 4672 28982 4674 29034
rect 4674 28982 4726 29034
rect 4726 28982 4728 29034
rect 4672 28980 4728 28982
rect 3804 28250 3860 28252
rect 3804 28198 3806 28250
rect 3806 28198 3858 28250
rect 3858 28198 3860 28250
rect 3804 28196 3860 28198
rect 3908 28250 3964 28252
rect 3908 28198 3910 28250
rect 3910 28198 3962 28250
rect 3962 28198 3964 28250
rect 3908 28196 3964 28198
rect 4012 28250 4068 28252
rect 4012 28198 4014 28250
rect 4014 28198 4066 28250
rect 4066 28198 4068 28250
rect 4012 28196 4068 28198
rect 3612 26684 3668 26740
rect 3500 25788 3556 25844
rect 3500 25228 3556 25284
rect 3052 23660 3108 23716
rect 3052 22540 3108 22596
rect 3804 26682 3860 26684
rect 3804 26630 3806 26682
rect 3806 26630 3858 26682
rect 3858 26630 3860 26682
rect 3804 26628 3860 26630
rect 3908 26682 3964 26684
rect 3908 26630 3910 26682
rect 3910 26630 3962 26682
rect 3962 26630 3964 26682
rect 3908 26628 3964 26630
rect 4012 26682 4068 26684
rect 4012 26630 4014 26682
rect 4014 26630 4066 26682
rect 4066 26630 4068 26682
rect 4012 26628 4068 26630
rect 3836 26460 3892 26516
rect 3724 25676 3780 25732
rect 4284 27858 4340 27860
rect 4284 27806 4286 27858
rect 4286 27806 4338 27858
rect 4338 27806 4340 27858
rect 4284 27804 4340 27806
rect 5180 34188 5236 34244
rect 5180 33628 5236 33684
rect 5068 31836 5124 31892
rect 5180 33180 5236 33236
rect 5068 29820 5124 29876
rect 5404 35532 5460 35588
rect 5404 34914 5460 34916
rect 5404 34862 5406 34914
rect 5406 34862 5458 34914
rect 5458 34862 5460 34914
rect 5404 34860 5460 34862
rect 5292 31612 5348 31668
rect 5404 34076 5460 34132
rect 5404 30380 5460 30436
rect 5180 29596 5236 29652
rect 5628 37042 5684 37044
rect 5628 36990 5630 37042
rect 5630 36990 5682 37042
rect 5682 36990 5684 37042
rect 5628 36988 5684 36990
rect 6076 48188 6132 48244
rect 6076 41410 6132 41412
rect 6076 41358 6078 41410
rect 6078 41358 6130 41410
rect 6130 41358 6132 41410
rect 6076 41356 6132 41358
rect 8092 55970 8148 55972
rect 8092 55918 8094 55970
rect 8094 55918 8146 55970
rect 8146 55918 8148 55970
rect 8092 55916 8148 55918
rect 6636 51436 6692 51492
rect 7420 49532 7476 49588
rect 7196 48972 7252 49028
rect 5964 39676 6020 39732
rect 6188 38892 6244 38948
rect 5964 38722 6020 38724
rect 5964 38670 5966 38722
rect 5966 38670 6018 38722
rect 6018 38670 6020 38722
rect 5964 38668 6020 38670
rect 5852 35810 5908 35812
rect 5852 35758 5854 35810
rect 5854 35758 5906 35810
rect 5906 35758 5908 35810
rect 5852 35756 5908 35758
rect 5740 35420 5796 35476
rect 5628 33234 5684 33236
rect 5628 33182 5630 33234
rect 5630 33182 5682 33234
rect 5682 33182 5684 33234
rect 5628 33180 5684 33182
rect 5628 30380 5684 30436
rect 5852 35532 5908 35588
rect 6300 35474 6356 35476
rect 6300 35422 6302 35474
rect 6302 35422 6354 35474
rect 6354 35422 6356 35474
rect 6300 35420 6356 35422
rect 5964 34412 6020 34468
rect 6076 34748 6132 34804
rect 6076 33570 6132 33572
rect 6076 33518 6078 33570
rect 6078 33518 6130 33570
rect 6130 33518 6132 33570
rect 6076 33516 6132 33518
rect 6300 31836 6356 31892
rect 5852 30380 5908 30436
rect 5964 31612 6020 31668
rect 5852 30210 5908 30212
rect 5852 30158 5854 30210
rect 5854 30158 5906 30210
rect 5906 30158 5908 30210
rect 5852 30156 5908 30158
rect 6300 30604 6356 30660
rect 4956 28028 5012 28084
rect 4844 27916 4900 27972
rect 3836 25452 3892 25508
rect 4464 27466 4520 27468
rect 4464 27414 4466 27466
rect 4466 27414 4518 27466
rect 4518 27414 4520 27466
rect 4464 27412 4520 27414
rect 4568 27466 4624 27468
rect 4568 27414 4570 27466
rect 4570 27414 4622 27466
rect 4622 27414 4624 27466
rect 4568 27412 4624 27414
rect 4672 27466 4728 27468
rect 4672 27414 4674 27466
rect 4674 27414 4726 27466
rect 4726 27414 4728 27466
rect 4672 27412 4728 27414
rect 5068 28364 5124 28420
rect 4464 25898 4520 25900
rect 4464 25846 4466 25898
rect 4466 25846 4518 25898
rect 4518 25846 4520 25898
rect 4464 25844 4520 25846
rect 4568 25898 4624 25900
rect 4568 25846 4570 25898
rect 4570 25846 4622 25898
rect 4622 25846 4624 25898
rect 4568 25844 4624 25846
rect 4672 25898 4728 25900
rect 4672 25846 4674 25898
rect 4674 25846 4726 25898
rect 4726 25846 4728 25898
rect 4672 25844 4728 25846
rect 3804 25114 3860 25116
rect 3804 25062 3806 25114
rect 3806 25062 3858 25114
rect 3858 25062 3860 25114
rect 3804 25060 3860 25062
rect 3908 25114 3964 25116
rect 3908 25062 3910 25114
rect 3910 25062 3962 25114
rect 3962 25062 3964 25114
rect 3908 25060 3964 25062
rect 4012 25114 4068 25116
rect 4012 25062 4014 25114
rect 4014 25062 4066 25114
rect 4066 25062 4068 25114
rect 4012 25060 4068 25062
rect 3276 23100 3332 23156
rect 2940 20748 2996 20804
rect 3052 21196 3108 21252
rect 2828 20242 2884 20244
rect 2828 20190 2830 20242
rect 2830 20190 2882 20242
rect 2882 20190 2884 20242
rect 2828 20188 2884 20190
rect 3276 21196 3332 21252
rect 3276 21026 3332 21028
rect 3276 20974 3278 21026
rect 3278 20974 3330 21026
rect 3330 20974 3332 21026
rect 3276 20972 3332 20974
rect 2604 19404 2660 19460
rect 2716 19346 2772 19348
rect 2716 19294 2718 19346
rect 2718 19294 2770 19346
rect 2770 19294 2772 19346
rect 2716 19292 2772 19294
rect 2716 18732 2772 18788
rect 2492 18396 2548 18452
rect 2156 17724 2212 17780
rect 2604 17778 2660 17780
rect 2604 17726 2606 17778
rect 2606 17726 2658 17778
rect 2658 17726 2660 17778
rect 2604 17724 2660 17726
rect 2604 17500 2660 17556
rect 1932 16156 1988 16212
rect 1932 15090 1988 15092
rect 1932 15038 1934 15090
rect 1934 15038 1986 15090
rect 1986 15038 1988 15090
rect 1932 15036 1988 15038
rect 1932 14812 1988 14868
rect 1932 13468 1988 13524
rect 2492 13916 2548 13972
rect 1708 12908 1764 12964
rect 1596 12290 1652 12292
rect 1596 12238 1598 12290
rect 1598 12238 1650 12290
rect 1650 12238 1652 12290
rect 1596 12236 1652 12238
rect 2044 13020 2100 13076
rect 2156 12962 2212 12964
rect 2156 12910 2158 12962
rect 2158 12910 2210 12962
rect 2210 12910 2212 12962
rect 2156 12908 2212 12910
rect 2828 17836 2884 17892
rect 2940 19404 2996 19460
rect 2828 14754 2884 14756
rect 2828 14702 2830 14754
rect 2830 14702 2882 14754
rect 2882 14702 2884 14754
rect 2828 14700 2884 14702
rect 3052 19292 3108 19348
rect 3164 18732 3220 18788
rect 3164 18562 3220 18564
rect 3164 18510 3166 18562
rect 3166 18510 3218 18562
rect 3218 18510 3220 18562
rect 3164 18508 3220 18510
rect 3052 15148 3108 15204
rect 3164 16156 3220 16212
rect 3052 14812 3108 14868
rect 4060 23660 4116 23716
rect 3804 23546 3860 23548
rect 3804 23494 3806 23546
rect 3806 23494 3858 23546
rect 3858 23494 3860 23546
rect 3804 23492 3860 23494
rect 3908 23546 3964 23548
rect 3908 23494 3910 23546
rect 3910 23494 3962 23546
rect 3962 23494 3964 23546
rect 3908 23492 3964 23494
rect 4012 23546 4068 23548
rect 4012 23494 4014 23546
rect 4014 23494 4066 23546
rect 4066 23494 4068 23546
rect 4012 23492 4068 23494
rect 4464 24330 4520 24332
rect 4464 24278 4466 24330
rect 4466 24278 4518 24330
rect 4518 24278 4520 24330
rect 4464 24276 4520 24278
rect 4568 24330 4624 24332
rect 4568 24278 4570 24330
rect 4570 24278 4622 24330
rect 4622 24278 4624 24330
rect 4568 24276 4624 24278
rect 4672 24330 4728 24332
rect 4672 24278 4674 24330
rect 4674 24278 4726 24330
rect 4726 24278 4728 24330
rect 4672 24276 4728 24278
rect 4844 23884 4900 23940
rect 4620 23826 4676 23828
rect 4620 23774 4622 23826
rect 4622 23774 4674 23826
rect 4674 23774 4676 23826
rect 4620 23772 4676 23774
rect 4284 23660 4340 23716
rect 3804 21978 3860 21980
rect 3804 21926 3806 21978
rect 3806 21926 3858 21978
rect 3858 21926 3860 21978
rect 3804 21924 3860 21926
rect 3908 21978 3964 21980
rect 3908 21926 3910 21978
rect 3910 21926 3962 21978
rect 3962 21926 3964 21978
rect 3908 21924 3964 21926
rect 4012 21978 4068 21980
rect 4012 21926 4014 21978
rect 4014 21926 4066 21978
rect 4066 21926 4068 21978
rect 4012 21924 4068 21926
rect 3804 20410 3860 20412
rect 3804 20358 3806 20410
rect 3806 20358 3858 20410
rect 3858 20358 3860 20410
rect 3804 20356 3860 20358
rect 3908 20410 3964 20412
rect 3908 20358 3910 20410
rect 3910 20358 3962 20410
rect 3962 20358 3964 20410
rect 3908 20356 3964 20358
rect 4012 20410 4068 20412
rect 4012 20358 4014 20410
rect 4014 20358 4066 20410
rect 4066 20358 4068 20410
rect 4012 20356 4068 20358
rect 3500 19852 3556 19908
rect 5292 27858 5348 27860
rect 5292 27806 5294 27858
rect 5294 27806 5346 27858
rect 5346 27806 5348 27858
rect 5292 27804 5348 27806
rect 5516 29036 5572 29092
rect 5740 28364 5796 28420
rect 5740 27858 5796 27860
rect 5740 27806 5742 27858
rect 5742 27806 5794 27858
rect 5794 27806 5796 27858
rect 5740 27804 5796 27806
rect 5516 27244 5572 27300
rect 5292 25340 5348 25396
rect 5404 23938 5460 23940
rect 5404 23886 5406 23938
rect 5406 23886 5458 23938
rect 5458 23886 5460 23938
rect 5404 23884 5460 23886
rect 5068 23324 5124 23380
rect 4464 22762 4520 22764
rect 4464 22710 4466 22762
rect 4466 22710 4518 22762
rect 4518 22710 4520 22762
rect 4464 22708 4520 22710
rect 4568 22762 4624 22764
rect 4568 22710 4570 22762
rect 4570 22710 4622 22762
rect 4622 22710 4624 22762
rect 4568 22708 4624 22710
rect 4672 22762 4728 22764
rect 4672 22710 4674 22762
rect 4674 22710 4726 22762
rect 4726 22710 4728 22762
rect 4672 22708 4728 22710
rect 4284 22316 4340 22372
rect 4464 21194 4520 21196
rect 4464 21142 4466 21194
rect 4466 21142 4518 21194
rect 4518 21142 4520 21194
rect 4464 21140 4520 21142
rect 4568 21194 4624 21196
rect 4568 21142 4570 21194
rect 4570 21142 4622 21194
rect 4622 21142 4624 21194
rect 4568 21140 4624 21142
rect 4672 21194 4728 21196
rect 4672 21142 4674 21194
rect 4674 21142 4726 21194
rect 4726 21142 4728 21194
rect 4956 21196 5012 21252
rect 4672 21140 4728 21142
rect 4508 20412 4564 20468
rect 4172 19852 4228 19908
rect 4956 19964 5012 20020
rect 4464 19626 4520 19628
rect 4464 19574 4466 19626
rect 4466 19574 4518 19626
rect 4518 19574 4520 19626
rect 4464 19572 4520 19574
rect 4568 19626 4624 19628
rect 4568 19574 4570 19626
rect 4570 19574 4622 19626
rect 4622 19574 4624 19626
rect 4568 19572 4624 19574
rect 4672 19626 4728 19628
rect 4672 19574 4674 19626
rect 4674 19574 4726 19626
rect 4726 19574 4728 19626
rect 4672 19572 4728 19574
rect 4508 19346 4564 19348
rect 4508 19294 4510 19346
rect 4510 19294 4562 19346
rect 4562 19294 4564 19346
rect 4508 19292 4564 19294
rect 3612 18732 3668 18788
rect 3804 18842 3860 18844
rect 3804 18790 3806 18842
rect 3806 18790 3858 18842
rect 3858 18790 3860 18842
rect 3804 18788 3860 18790
rect 3908 18842 3964 18844
rect 3908 18790 3910 18842
rect 3910 18790 3962 18842
rect 3962 18790 3964 18842
rect 3908 18788 3964 18790
rect 4012 18842 4068 18844
rect 4012 18790 4014 18842
rect 4014 18790 4066 18842
rect 4066 18790 4068 18842
rect 4012 18788 4068 18790
rect 4284 18732 4340 18788
rect 4956 18732 5012 18788
rect 3948 18284 4004 18340
rect 4464 18058 4520 18060
rect 4464 18006 4466 18058
rect 4466 18006 4518 18058
rect 4518 18006 4520 18058
rect 4464 18004 4520 18006
rect 4568 18058 4624 18060
rect 4568 18006 4570 18058
rect 4570 18006 4622 18058
rect 4622 18006 4624 18058
rect 4568 18004 4624 18006
rect 4672 18058 4728 18060
rect 4672 18006 4674 18058
rect 4674 18006 4726 18058
rect 4726 18006 4728 18058
rect 4672 18004 4728 18006
rect 4284 17836 4340 17892
rect 3724 17666 3780 17668
rect 3724 17614 3726 17666
rect 3726 17614 3778 17666
rect 3778 17614 3780 17666
rect 3724 17612 3780 17614
rect 3612 17276 3668 17332
rect 3804 17274 3860 17276
rect 3804 17222 3806 17274
rect 3806 17222 3858 17274
rect 3858 17222 3860 17274
rect 3804 17220 3860 17222
rect 3908 17274 3964 17276
rect 3908 17222 3910 17274
rect 3910 17222 3962 17274
rect 3962 17222 3964 17274
rect 3908 17220 3964 17222
rect 4012 17274 4068 17276
rect 4012 17222 4014 17274
rect 4014 17222 4066 17274
rect 4066 17222 4068 17274
rect 4012 17220 4068 17222
rect 3836 16882 3892 16884
rect 3836 16830 3838 16882
rect 3838 16830 3890 16882
rect 3890 16830 3892 16882
rect 3836 16828 3892 16830
rect 4844 17890 4900 17892
rect 4844 17838 4846 17890
rect 4846 17838 4898 17890
rect 4898 17838 4900 17890
rect 4844 17836 4900 17838
rect 4844 17612 4900 17668
rect 4508 17276 4564 17332
rect 4396 16658 4452 16660
rect 4396 16606 4398 16658
rect 4398 16606 4450 16658
rect 4450 16606 4452 16658
rect 4396 16604 4452 16606
rect 4464 16490 4520 16492
rect 4464 16438 4466 16490
rect 4466 16438 4518 16490
rect 4518 16438 4520 16490
rect 4464 16436 4520 16438
rect 4568 16490 4624 16492
rect 4568 16438 4570 16490
rect 4570 16438 4622 16490
rect 4622 16438 4624 16490
rect 4568 16436 4624 16438
rect 4672 16490 4728 16492
rect 4672 16438 4674 16490
rect 4674 16438 4726 16490
rect 4726 16438 4728 16490
rect 4672 16436 4728 16438
rect 3388 14812 3444 14868
rect 3500 15708 3556 15764
rect 3804 15706 3860 15708
rect 3388 14588 3444 14644
rect 2604 13186 2660 13188
rect 2604 13134 2606 13186
rect 2606 13134 2658 13186
rect 2658 13134 2660 13186
rect 2604 13132 2660 13134
rect 2940 14252 2996 14308
rect 2156 12348 2212 12404
rect 1932 11900 1988 11956
rect 2492 12290 2548 12292
rect 2492 12238 2494 12290
rect 2494 12238 2546 12290
rect 2546 12238 2548 12290
rect 2492 12236 2548 12238
rect 2380 11900 2436 11956
rect 2268 11564 2324 11620
rect 2604 11506 2660 11508
rect 2604 11454 2606 11506
rect 2606 11454 2658 11506
rect 2658 11454 2660 11506
rect 2604 11452 2660 11454
rect 3276 14418 3332 14420
rect 3276 14366 3278 14418
rect 3278 14366 3330 14418
rect 3330 14366 3332 14418
rect 3276 14364 3332 14366
rect 3052 13468 3108 13524
rect 1260 6578 1316 6580
rect 1260 6526 1262 6578
rect 1262 6526 1314 6578
rect 1314 6526 1316 6578
rect 1260 6524 1316 6526
rect 1260 5180 1316 5236
rect 3164 12684 3220 12740
rect 3388 12796 3444 12852
rect 3500 11340 3556 11396
rect 3612 15596 3668 15652
rect 3804 15654 3806 15706
rect 3806 15654 3858 15706
rect 3858 15654 3860 15706
rect 3804 15652 3860 15654
rect 3908 15706 3964 15708
rect 3908 15654 3910 15706
rect 3910 15654 3962 15706
rect 3962 15654 3964 15706
rect 3908 15652 3964 15654
rect 4012 15706 4068 15708
rect 4012 15654 4014 15706
rect 4014 15654 4066 15706
rect 4066 15654 4068 15706
rect 4012 15652 4068 15654
rect 3052 3836 3108 3892
rect 1372 2380 1428 2436
rect 3388 2380 3444 2436
rect 700 1596 756 1652
rect 2044 1372 2100 1428
rect 4732 16322 4788 16324
rect 4732 16270 4734 16322
rect 4734 16270 4786 16322
rect 4786 16270 4788 16322
rect 4732 16268 4788 16270
rect 4396 15036 4452 15092
rect 4464 14922 4520 14924
rect 4464 14870 4466 14922
rect 4466 14870 4518 14922
rect 4518 14870 4520 14922
rect 4464 14868 4520 14870
rect 4568 14922 4624 14924
rect 4568 14870 4570 14922
rect 4570 14870 4622 14922
rect 4622 14870 4624 14922
rect 4568 14868 4624 14870
rect 4672 14922 4728 14924
rect 4672 14870 4674 14922
rect 4674 14870 4726 14922
rect 4726 14870 4728 14922
rect 4672 14868 4728 14870
rect 4508 14642 4564 14644
rect 4508 14590 4510 14642
rect 4510 14590 4562 14642
rect 4562 14590 4564 14642
rect 4508 14588 4564 14590
rect 4956 16882 5012 16884
rect 4956 16830 4958 16882
rect 4958 16830 5010 16882
rect 5010 16830 5012 16882
rect 4956 16828 5012 16830
rect 4956 15708 5012 15764
rect 4956 14588 5012 14644
rect 3804 14138 3860 14140
rect 3804 14086 3806 14138
rect 3806 14086 3858 14138
rect 3858 14086 3860 14138
rect 3804 14084 3860 14086
rect 3908 14138 3964 14140
rect 3908 14086 3910 14138
rect 3910 14086 3962 14138
rect 3962 14086 3964 14138
rect 3908 14084 3964 14086
rect 4012 14138 4068 14140
rect 4012 14086 4014 14138
rect 4014 14086 4066 14138
rect 4066 14086 4068 14138
rect 4012 14084 4068 14086
rect 4956 13804 5012 13860
rect 4284 13244 4340 13300
rect 4464 13354 4520 13356
rect 4464 13302 4466 13354
rect 4466 13302 4518 13354
rect 4518 13302 4520 13354
rect 4464 13300 4520 13302
rect 4568 13354 4624 13356
rect 4568 13302 4570 13354
rect 4570 13302 4622 13354
rect 4622 13302 4624 13354
rect 4568 13300 4624 13302
rect 4672 13354 4728 13356
rect 4672 13302 4674 13354
rect 4674 13302 4726 13354
rect 4726 13302 4728 13354
rect 4672 13300 4728 13302
rect 5852 27244 5908 27300
rect 5628 23548 5684 23604
rect 5628 23436 5684 23492
rect 5292 22540 5348 22596
rect 5852 26572 5908 26628
rect 6300 26460 6356 26516
rect 6188 26236 6244 26292
rect 6188 24108 6244 24164
rect 5852 23548 5908 23604
rect 6076 23548 6132 23604
rect 5852 23100 5908 23156
rect 5292 22370 5348 22372
rect 5292 22318 5294 22370
rect 5294 22318 5346 22370
rect 5346 22318 5348 22370
rect 5292 22316 5348 22318
rect 5292 20076 5348 20132
rect 5852 22540 5908 22596
rect 5516 21980 5572 22036
rect 5740 21644 5796 21700
rect 5740 20972 5796 21028
rect 5628 20860 5684 20916
rect 5740 20748 5796 20804
rect 5964 21362 6020 21364
rect 5964 21310 5966 21362
rect 5966 21310 6018 21362
rect 6018 21310 6020 21362
rect 5964 21308 6020 21310
rect 6972 39788 7028 39844
rect 6636 39564 6692 39620
rect 6748 39004 6804 39060
rect 6748 37884 6804 37940
rect 6748 37490 6804 37492
rect 6748 37438 6750 37490
rect 6750 37438 6802 37490
rect 6802 37438 6804 37490
rect 6748 37436 6804 37438
rect 6636 36316 6692 36372
rect 6748 35868 6804 35924
rect 6860 35980 6916 36036
rect 6748 32562 6804 32564
rect 6748 32510 6750 32562
rect 6750 32510 6802 32562
rect 6802 32510 6804 32562
rect 6748 32508 6804 32510
rect 6636 30828 6692 30884
rect 6748 28924 6804 28980
rect 6636 28530 6692 28532
rect 6636 28478 6638 28530
rect 6638 28478 6690 28530
rect 6690 28478 6692 28530
rect 6636 28476 6692 28478
rect 6412 23324 6468 23380
rect 6748 26908 6804 26964
rect 6636 25618 6692 25620
rect 6636 25566 6638 25618
rect 6638 25566 6690 25618
rect 6690 25566 6692 25618
rect 6636 25564 6692 25566
rect 6748 25004 6804 25060
rect 6636 24220 6692 24276
rect 6636 23324 6692 23380
rect 6524 23100 6580 23156
rect 6524 22876 6580 22932
rect 6300 20972 6356 21028
rect 6524 20860 6580 20916
rect 7196 39058 7252 39060
rect 7196 39006 7198 39058
rect 7198 39006 7250 39058
rect 7250 39006 7252 39058
rect 7196 39004 7252 39006
rect 7084 35532 7140 35588
rect 15484 56252 15540 56308
rect 16492 56306 16548 56308
rect 16492 56254 16494 56306
rect 16494 56254 16546 56306
rect 16546 56254 16548 56306
rect 16492 56252 16548 56254
rect 11564 55356 11620 55412
rect 12908 55020 12964 55076
rect 9996 54572 10052 54628
rect 8652 54236 8708 54292
rect 15596 55468 15652 55524
rect 19516 56252 19572 56308
rect 20636 56306 20692 56308
rect 20636 56254 20638 56306
rect 20638 56254 20690 56306
rect 20690 56254 20692 56306
rect 20636 56252 20692 56254
rect 20860 56252 20916 56308
rect 21868 56306 21924 56308
rect 21868 56254 21870 56306
rect 21870 56254 21922 56306
rect 21922 56254 21924 56306
rect 21868 56252 21924 56254
rect 22540 56140 22596 56196
rect 14028 53900 14084 53956
rect 14700 54348 14756 54404
rect 14252 53452 14308 53508
rect 12684 52444 12740 52500
rect 10108 52332 10164 52388
rect 7980 44044 8036 44100
rect 7756 43372 7812 43428
rect 7644 38892 7700 38948
rect 7532 37772 7588 37828
rect 7644 38556 7700 38612
rect 7532 37154 7588 37156
rect 7532 37102 7534 37154
rect 7534 37102 7586 37154
rect 7586 37102 7588 37154
rect 7532 37100 7588 37102
rect 7868 40460 7924 40516
rect 7756 37436 7812 37492
rect 8092 40124 8148 40180
rect 8204 40236 8260 40292
rect 8764 40402 8820 40404
rect 8764 40350 8766 40402
rect 8766 40350 8818 40402
rect 8818 40350 8820 40402
rect 8764 40348 8820 40350
rect 9100 48748 9156 48804
rect 8988 38780 9044 38836
rect 7084 34412 7140 34468
rect 7644 35644 7700 35700
rect 7868 36092 7924 36148
rect 7868 35586 7924 35588
rect 7868 35534 7870 35586
rect 7870 35534 7922 35586
rect 7922 35534 7924 35586
rect 7868 35532 7924 35534
rect 7420 33852 7476 33908
rect 7308 33740 7364 33796
rect 7196 33404 7252 33460
rect 7196 32508 7252 32564
rect 7420 32732 7476 32788
rect 7308 31778 7364 31780
rect 7308 31726 7310 31778
rect 7310 31726 7362 31778
rect 7362 31726 7364 31778
rect 7308 31724 7364 31726
rect 7084 30492 7140 30548
rect 6972 28924 7028 28980
rect 6972 28588 7028 28644
rect 6972 23548 7028 23604
rect 7084 27804 7140 27860
rect 6972 23324 7028 23380
rect 6860 21756 6916 21812
rect 6412 20748 6468 20804
rect 5852 20412 5908 20468
rect 6188 19628 6244 19684
rect 5404 17164 5460 17220
rect 5628 18844 5684 18900
rect 5628 16604 5684 16660
rect 5740 16828 5796 16884
rect 5292 15820 5348 15876
rect 7196 24780 7252 24836
rect 7196 22930 7252 22932
rect 7196 22878 7198 22930
rect 7198 22878 7250 22930
rect 7250 22878 7252 22930
rect 7196 22876 7252 22878
rect 6748 20914 6804 20916
rect 6748 20862 6750 20914
rect 6750 20862 6802 20914
rect 6802 20862 6804 20914
rect 6748 20860 6804 20862
rect 6748 20130 6804 20132
rect 6748 20078 6750 20130
rect 6750 20078 6802 20130
rect 6802 20078 6804 20130
rect 6748 20076 6804 20078
rect 7084 21586 7140 21588
rect 7084 21534 7086 21586
rect 7086 21534 7138 21586
rect 7138 21534 7140 21586
rect 7084 21532 7140 21534
rect 7196 21756 7252 21812
rect 7868 33740 7924 33796
rect 8092 35980 8148 36036
rect 8204 37436 8260 37492
rect 8092 35308 8148 35364
rect 8316 37266 8372 37268
rect 8316 37214 8318 37266
rect 8318 37214 8370 37266
rect 8370 37214 8372 37266
rect 8316 37212 8372 37214
rect 8316 35980 8372 36036
rect 8316 35698 8372 35700
rect 8316 35646 8318 35698
rect 8318 35646 8370 35698
rect 8370 35646 8372 35698
rect 8316 35644 8372 35646
rect 8652 35308 8708 35364
rect 8540 33628 8596 33684
rect 8316 33404 8372 33460
rect 7980 32732 8036 32788
rect 7644 31724 7700 31780
rect 7980 30940 8036 30996
rect 8092 31612 8148 31668
rect 7756 30044 7812 30100
rect 7644 26460 7700 26516
rect 7532 24834 7588 24836
rect 7532 24782 7534 24834
rect 7534 24782 7586 24834
rect 7586 24782 7588 24834
rect 7532 24780 7588 24782
rect 7532 24332 7588 24388
rect 7980 30268 8036 30324
rect 8204 30210 8260 30212
rect 8204 30158 8206 30210
rect 8206 30158 8258 30210
rect 8258 30158 8260 30210
rect 8204 30156 8260 30158
rect 8540 31612 8596 31668
rect 8652 33292 8708 33348
rect 8652 32284 8708 32340
rect 8316 30044 8372 30100
rect 8652 28476 8708 28532
rect 8204 27804 8260 27860
rect 8316 27020 8372 27076
rect 7644 21868 7700 21924
rect 7308 21532 7364 21588
rect 7308 21362 7364 21364
rect 7308 21310 7310 21362
rect 7310 21310 7362 21362
rect 7362 21310 7364 21362
rect 7308 21308 7364 21310
rect 7196 19964 7252 20020
rect 7196 19794 7252 19796
rect 7196 19742 7198 19794
rect 7198 19742 7250 19794
rect 7250 19742 7252 19794
rect 7196 19740 7252 19742
rect 6636 19234 6692 19236
rect 6636 19182 6638 19234
rect 6638 19182 6690 19234
rect 6690 19182 6692 19234
rect 6636 19180 6692 19182
rect 6300 18844 6356 18900
rect 5964 18338 6020 18340
rect 5964 18286 5966 18338
rect 5966 18286 6018 18338
rect 6018 18286 6020 18338
rect 5964 18284 6020 18286
rect 6972 18284 7028 18340
rect 7644 19404 7700 19460
rect 7420 19180 7476 19236
rect 6636 17666 6692 17668
rect 6636 17614 6638 17666
rect 6638 17614 6690 17666
rect 6690 17614 6692 17666
rect 6636 17612 6692 17614
rect 5852 16604 5908 16660
rect 5852 16044 5908 16100
rect 5628 14700 5684 14756
rect 5292 13804 5348 13860
rect 5068 13580 5124 13636
rect 5180 13356 5236 13412
rect 5292 13580 5348 13636
rect 5068 12908 5124 12964
rect 4172 12850 4228 12852
rect 4172 12798 4174 12850
rect 4174 12798 4226 12850
rect 4226 12798 4228 12850
rect 4172 12796 4228 12798
rect 3804 12570 3860 12572
rect 3804 12518 3806 12570
rect 3806 12518 3858 12570
rect 3858 12518 3860 12570
rect 3804 12516 3860 12518
rect 3908 12570 3964 12572
rect 3908 12518 3910 12570
rect 3910 12518 3962 12570
rect 3962 12518 3964 12570
rect 3908 12516 3964 12518
rect 4012 12570 4068 12572
rect 4012 12518 4014 12570
rect 4014 12518 4066 12570
rect 4066 12518 4068 12570
rect 4012 12516 4068 12518
rect 4464 11786 4520 11788
rect 4464 11734 4466 11786
rect 4466 11734 4518 11786
rect 4518 11734 4520 11786
rect 4464 11732 4520 11734
rect 4568 11786 4624 11788
rect 4568 11734 4570 11786
rect 4570 11734 4622 11786
rect 4622 11734 4624 11786
rect 4568 11732 4624 11734
rect 4672 11786 4728 11788
rect 4672 11734 4674 11786
rect 4674 11734 4726 11786
rect 4726 11734 4728 11786
rect 4672 11732 4728 11734
rect 4284 11394 4340 11396
rect 4284 11342 4286 11394
rect 4286 11342 4338 11394
rect 4338 11342 4340 11394
rect 4284 11340 4340 11342
rect 3804 11002 3860 11004
rect 3804 10950 3806 11002
rect 3806 10950 3858 11002
rect 3858 10950 3860 11002
rect 3804 10948 3860 10950
rect 3908 11002 3964 11004
rect 3908 10950 3910 11002
rect 3910 10950 3962 11002
rect 3962 10950 3964 11002
rect 3908 10948 3964 10950
rect 4012 11002 4068 11004
rect 4012 10950 4014 11002
rect 4014 10950 4066 11002
rect 4066 10950 4068 11002
rect 4012 10948 4068 10950
rect 4844 11340 4900 11396
rect 4284 10444 4340 10500
rect 4464 10218 4520 10220
rect 4464 10166 4466 10218
rect 4466 10166 4518 10218
rect 4518 10166 4520 10218
rect 4464 10164 4520 10166
rect 4568 10218 4624 10220
rect 4568 10166 4570 10218
rect 4570 10166 4622 10218
rect 4622 10166 4624 10218
rect 4568 10164 4624 10166
rect 4672 10218 4728 10220
rect 4672 10166 4674 10218
rect 4674 10166 4726 10218
rect 4726 10166 4728 10218
rect 4672 10164 4728 10166
rect 4732 9938 4788 9940
rect 4732 9886 4734 9938
rect 4734 9886 4786 9938
rect 4786 9886 4788 9938
rect 4732 9884 4788 9886
rect 5292 12236 5348 12292
rect 6188 17164 6244 17220
rect 6076 15202 6132 15204
rect 6076 15150 6078 15202
rect 6078 15150 6130 15202
rect 6130 15150 6132 15202
rect 6076 15148 6132 15150
rect 6636 17052 6692 17108
rect 6972 17388 7028 17444
rect 6636 16882 6692 16884
rect 6636 16830 6638 16882
rect 6638 16830 6690 16882
rect 6690 16830 6692 16882
rect 6636 16828 6692 16830
rect 6860 16210 6916 16212
rect 6860 16158 6862 16210
rect 6862 16158 6914 16210
rect 6914 16158 6916 16210
rect 6860 16156 6916 16158
rect 5852 13692 5908 13748
rect 5852 13468 5908 13524
rect 5964 12460 6020 12516
rect 5404 11340 5460 11396
rect 6748 13522 6804 13524
rect 6748 13470 6750 13522
rect 6750 13470 6802 13522
rect 6802 13470 6804 13522
rect 6748 13468 6804 13470
rect 6412 13132 6468 13188
rect 6412 12236 6468 12292
rect 6860 12796 6916 12852
rect 6076 11340 6132 11396
rect 6188 11788 6244 11844
rect 5852 10722 5908 10724
rect 5852 10670 5854 10722
rect 5854 10670 5906 10722
rect 5906 10670 5908 10722
rect 5852 10668 5908 10670
rect 5964 10556 6020 10612
rect 3804 9434 3860 9436
rect 3804 9382 3806 9434
rect 3806 9382 3858 9434
rect 3858 9382 3860 9434
rect 3804 9380 3860 9382
rect 3908 9434 3964 9436
rect 3908 9382 3910 9434
rect 3910 9382 3962 9434
rect 3962 9382 3964 9434
rect 3908 9380 3964 9382
rect 4012 9434 4068 9436
rect 4012 9382 4014 9434
rect 4014 9382 4066 9434
rect 4066 9382 4068 9434
rect 4012 9380 4068 9382
rect 4464 8650 4520 8652
rect 4464 8598 4466 8650
rect 4466 8598 4518 8650
rect 4518 8598 4520 8650
rect 4464 8596 4520 8598
rect 4568 8650 4624 8652
rect 4568 8598 4570 8650
rect 4570 8598 4622 8650
rect 4622 8598 4624 8650
rect 4568 8596 4624 8598
rect 4672 8650 4728 8652
rect 4672 8598 4674 8650
rect 4674 8598 4726 8650
rect 4726 8598 4728 8650
rect 4672 8596 4728 8598
rect 3804 7866 3860 7868
rect 3804 7814 3806 7866
rect 3806 7814 3858 7866
rect 3858 7814 3860 7866
rect 3804 7812 3860 7814
rect 3908 7866 3964 7868
rect 3908 7814 3910 7866
rect 3910 7814 3962 7866
rect 3962 7814 3964 7866
rect 3908 7812 3964 7814
rect 4012 7866 4068 7868
rect 4012 7814 4014 7866
rect 4014 7814 4066 7866
rect 4066 7814 4068 7866
rect 4012 7812 4068 7814
rect 4464 7082 4520 7084
rect 4464 7030 4466 7082
rect 4466 7030 4518 7082
rect 4518 7030 4520 7082
rect 4464 7028 4520 7030
rect 4568 7082 4624 7084
rect 4568 7030 4570 7082
rect 4570 7030 4622 7082
rect 4622 7030 4624 7082
rect 4568 7028 4624 7030
rect 4672 7082 4728 7084
rect 4672 7030 4674 7082
rect 4674 7030 4726 7082
rect 4726 7030 4728 7082
rect 4672 7028 4728 7030
rect 3804 6298 3860 6300
rect 3804 6246 3806 6298
rect 3806 6246 3858 6298
rect 3858 6246 3860 6298
rect 3804 6244 3860 6246
rect 3908 6298 3964 6300
rect 3908 6246 3910 6298
rect 3910 6246 3962 6298
rect 3962 6246 3964 6298
rect 3908 6244 3964 6246
rect 4012 6298 4068 6300
rect 4012 6246 4014 6298
rect 4014 6246 4066 6298
rect 4066 6246 4068 6298
rect 4012 6244 4068 6246
rect 4464 5514 4520 5516
rect 4464 5462 4466 5514
rect 4466 5462 4518 5514
rect 4518 5462 4520 5514
rect 4464 5460 4520 5462
rect 4568 5514 4624 5516
rect 4568 5462 4570 5514
rect 4570 5462 4622 5514
rect 4622 5462 4624 5514
rect 4568 5460 4624 5462
rect 4672 5514 4728 5516
rect 4672 5462 4674 5514
rect 4674 5462 4726 5514
rect 4726 5462 4728 5514
rect 4672 5460 4728 5462
rect 3804 4730 3860 4732
rect 3804 4678 3806 4730
rect 3806 4678 3858 4730
rect 3858 4678 3860 4730
rect 3804 4676 3860 4678
rect 3908 4730 3964 4732
rect 3908 4678 3910 4730
rect 3910 4678 3962 4730
rect 3962 4678 3964 4730
rect 3908 4676 3964 4678
rect 4012 4730 4068 4732
rect 4012 4678 4014 4730
rect 4014 4678 4066 4730
rect 4066 4678 4068 4730
rect 4012 4676 4068 4678
rect 4464 3946 4520 3948
rect 4464 3894 4466 3946
rect 4466 3894 4518 3946
rect 4518 3894 4520 3946
rect 4464 3892 4520 3894
rect 4568 3946 4624 3948
rect 4568 3894 4570 3946
rect 4570 3894 4622 3946
rect 4622 3894 4624 3946
rect 4568 3892 4624 3894
rect 4672 3946 4728 3948
rect 4672 3894 4674 3946
rect 4674 3894 4726 3946
rect 4726 3894 4728 3946
rect 4672 3892 4728 3894
rect 7084 17164 7140 17220
rect 7308 14812 7364 14868
rect 8092 26066 8148 26068
rect 8092 26014 8094 26066
rect 8094 26014 8146 26066
rect 8146 26014 8148 26066
rect 8092 26012 8148 26014
rect 8652 27020 8708 27076
rect 8316 25004 8372 25060
rect 8316 22930 8372 22932
rect 8316 22878 8318 22930
rect 8318 22878 8370 22930
rect 8370 22878 8372 22930
rect 8316 22876 8372 22878
rect 8092 22204 8148 22260
rect 8204 22316 8260 22372
rect 7756 19180 7812 19236
rect 7868 20748 7924 20804
rect 7756 15372 7812 15428
rect 7868 16828 7924 16884
rect 8092 21756 8148 21812
rect 8092 20748 8148 20804
rect 9772 42700 9828 42756
rect 9324 40236 9380 40292
rect 9548 41020 9604 41076
rect 9212 37996 9268 38052
rect 9212 37660 9268 37716
rect 8988 36258 9044 36260
rect 8988 36206 8990 36258
rect 8990 36206 9042 36258
rect 9042 36206 9044 36258
rect 8988 36204 9044 36206
rect 9100 35980 9156 36036
rect 8876 35474 8932 35476
rect 8876 35422 8878 35474
rect 8878 35422 8930 35474
rect 8930 35422 8932 35474
rect 8876 35420 8932 35422
rect 9100 35420 9156 35476
rect 9996 40236 10052 40292
rect 9884 39900 9940 39956
rect 9324 37548 9380 37604
rect 10892 50764 10948 50820
rect 11788 48860 11844 48916
rect 10892 42028 10948 42084
rect 11340 43596 11396 43652
rect 10556 41132 10612 41188
rect 10220 41074 10276 41076
rect 10220 41022 10222 41074
rect 10222 41022 10274 41074
rect 10274 41022 10276 41074
rect 10220 41020 10276 41022
rect 9548 38050 9604 38052
rect 9548 37998 9550 38050
rect 9550 37998 9602 38050
rect 9602 37998 9604 38050
rect 9548 37996 9604 37998
rect 9324 36428 9380 36484
rect 9324 36204 9380 36260
rect 9212 33180 9268 33236
rect 9324 35308 9380 35364
rect 8876 31778 8932 31780
rect 8876 31726 8878 31778
rect 8878 31726 8930 31778
rect 8930 31726 8932 31778
rect 8876 31724 8932 31726
rect 8988 29202 9044 29204
rect 8988 29150 8990 29202
rect 8990 29150 9042 29202
rect 9042 29150 9044 29202
rect 8988 29148 9044 29150
rect 8988 27970 9044 27972
rect 8988 27918 8990 27970
rect 8990 27918 9042 27970
rect 9042 27918 9044 27970
rect 8988 27916 9044 27918
rect 8764 25116 8820 25172
rect 8764 24444 8820 24500
rect 8652 23324 8708 23380
rect 8428 21532 8484 21588
rect 8540 22428 8596 22484
rect 8316 20972 8372 21028
rect 8316 20130 8372 20132
rect 8316 20078 8318 20130
rect 8318 20078 8370 20130
rect 8370 20078 8372 20130
rect 8316 20076 8372 20078
rect 8092 17612 8148 17668
rect 8316 16994 8372 16996
rect 8316 16942 8318 16994
rect 8318 16942 8370 16994
rect 8370 16942 8372 16994
rect 8316 16940 8372 16942
rect 8428 16604 8484 16660
rect 8204 16268 8260 16324
rect 8316 16156 8372 16212
rect 8092 15986 8148 15988
rect 8092 15934 8094 15986
rect 8094 15934 8146 15986
rect 8146 15934 8148 15986
rect 8092 15932 8148 15934
rect 7980 15372 8036 15428
rect 7644 14700 7700 14756
rect 7532 14476 7588 14532
rect 7196 12572 7252 12628
rect 6748 10780 6804 10836
rect 7308 11452 7364 11508
rect 7644 14252 7700 14308
rect 7084 10610 7140 10612
rect 7084 10558 7086 10610
rect 7086 10558 7138 10610
rect 7138 10558 7140 10610
rect 7084 10556 7140 10558
rect 6972 9714 7028 9716
rect 6972 9662 6974 9714
rect 6974 9662 7026 9714
rect 7026 9662 7028 9714
rect 6972 9660 7028 9662
rect 7756 13356 7812 13412
rect 7980 10780 8036 10836
rect 7308 9154 7364 9156
rect 7308 9102 7310 9154
rect 7310 9102 7362 9154
rect 7362 9102 7364 9154
rect 7308 9100 7364 9102
rect 7420 9996 7476 10052
rect 7084 8876 7140 8932
rect 7644 8930 7700 8932
rect 7644 8878 7646 8930
rect 7646 8878 7698 8930
rect 7698 8878 7700 8930
rect 7644 8876 7700 8878
rect 7420 7980 7476 8036
rect 8652 13804 8708 13860
rect 8204 12850 8260 12852
rect 8204 12798 8206 12850
rect 8206 12798 8258 12850
rect 8258 12798 8260 12850
rect 8204 12796 8260 12798
rect 8316 13692 8372 13748
rect 8204 11394 8260 11396
rect 8204 11342 8206 11394
rect 8206 11342 8258 11394
rect 8258 11342 8260 11394
rect 8204 11340 8260 11342
rect 8540 12178 8596 12180
rect 8540 12126 8542 12178
rect 8542 12126 8594 12178
rect 8594 12126 8596 12178
rect 8540 12124 8596 12126
rect 8876 24332 8932 24388
rect 8988 23324 9044 23380
rect 8876 21084 8932 21140
rect 8876 20018 8932 20020
rect 8876 19966 8878 20018
rect 8878 19966 8930 20018
rect 8930 19966 8932 20018
rect 8876 19964 8932 19966
rect 9212 32508 9268 32564
rect 9324 32172 9380 32228
rect 9548 36428 9604 36484
rect 9548 33628 9604 33684
rect 9436 27916 9492 27972
rect 9548 29260 9604 29316
rect 9324 27858 9380 27860
rect 9324 27806 9326 27858
rect 9326 27806 9378 27858
rect 9378 27806 9380 27858
rect 9324 27804 9380 27806
rect 9324 26012 9380 26068
rect 9324 24668 9380 24724
rect 9772 37548 9828 37604
rect 10108 36706 10164 36708
rect 10108 36654 10110 36706
rect 10110 36654 10162 36706
rect 10162 36654 10164 36706
rect 10108 36652 10164 36654
rect 9996 36540 10052 36596
rect 9772 29372 9828 29428
rect 9996 35084 10052 35140
rect 9996 33570 10052 33572
rect 9996 33518 9998 33570
rect 9998 33518 10050 33570
rect 10050 33518 10052 33570
rect 9996 33516 10052 33518
rect 11004 39506 11060 39508
rect 11004 39454 11006 39506
rect 11006 39454 11058 39506
rect 11058 39454 11060 39506
rect 11004 39452 11060 39454
rect 10556 37996 10612 38052
rect 11116 38050 11172 38052
rect 11116 37998 11118 38050
rect 11118 37998 11170 38050
rect 11170 37998 11172 38050
rect 11116 37996 11172 37998
rect 11004 37884 11060 37940
rect 10556 36370 10612 36372
rect 10556 36318 10558 36370
rect 10558 36318 10610 36370
rect 10610 36318 10612 36370
rect 10556 36316 10612 36318
rect 10556 35756 10612 35812
rect 10668 33068 10724 33124
rect 10556 32956 10612 33012
rect 10444 32562 10500 32564
rect 10444 32510 10446 32562
rect 10446 32510 10498 32562
rect 10498 32510 10500 32562
rect 10444 32508 10500 32510
rect 9996 32172 10052 32228
rect 9996 30044 10052 30100
rect 9996 29820 10052 29876
rect 10220 30210 10276 30212
rect 10220 30158 10222 30210
rect 10222 30158 10274 30210
rect 10274 30158 10276 30210
rect 10220 30156 10276 30158
rect 10220 29372 10276 29428
rect 10668 31276 10724 31332
rect 9884 26908 9940 26964
rect 9660 24892 9716 24948
rect 10556 27244 10612 27300
rect 10332 25564 10388 25620
rect 10444 25116 10500 25172
rect 10220 22540 10276 22596
rect 10332 22876 10388 22932
rect 9772 22428 9828 22484
rect 9212 22370 9268 22372
rect 9212 22318 9214 22370
rect 9214 22318 9266 22370
rect 9266 22318 9268 22370
rect 9212 22316 9268 22318
rect 9436 21586 9492 21588
rect 9436 21534 9438 21586
rect 9438 21534 9490 21586
rect 9490 21534 9492 21586
rect 9436 21532 9492 21534
rect 9660 20972 9716 21028
rect 9436 20636 9492 20692
rect 9324 20524 9380 20580
rect 9772 21308 9828 21364
rect 9884 20802 9940 20804
rect 9884 20750 9886 20802
rect 9886 20750 9938 20802
rect 9938 20750 9940 20802
rect 9884 20748 9940 20750
rect 9548 20300 9604 20356
rect 8876 18508 8932 18564
rect 9100 15484 9156 15540
rect 8988 14364 9044 14420
rect 9548 19740 9604 19796
rect 9436 18620 9492 18676
rect 9324 16098 9380 16100
rect 9324 16046 9326 16098
rect 9326 16046 9378 16098
rect 9378 16046 9380 16098
rect 9324 16044 9380 16046
rect 9548 18508 9604 18564
rect 9660 16828 9716 16884
rect 9996 19404 10052 19460
rect 11788 42924 11844 42980
rect 12012 44492 12068 44548
rect 11900 39676 11956 39732
rect 11788 39452 11844 39508
rect 11900 38050 11956 38052
rect 11900 37998 11902 38050
rect 11902 37998 11954 38050
rect 11954 37998 11956 38050
rect 11900 37996 11956 37998
rect 10892 31388 10948 31444
rect 11004 31052 11060 31108
rect 10892 30380 10948 30436
rect 11452 33068 11508 33124
rect 11340 31052 11396 31108
rect 11004 28812 11060 28868
rect 10892 28530 10948 28532
rect 10892 28478 10894 28530
rect 10894 28478 10946 28530
rect 10946 28478 10948 28530
rect 10892 28476 10948 28478
rect 10780 27356 10836 27412
rect 10892 27916 10948 27972
rect 11340 28866 11396 28868
rect 11340 28814 11342 28866
rect 11342 28814 11394 28866
rect 11394 28814 11396 28866
rect 11340 28812 11396 28814
rect 10668 25004 10724 25060
rect 10780 25116 10836 25172
rect 10780 23660 10836 23716
rect 10668 23436 10724 23492
rect 10556 23042 10612 23044
rect 10556 22990 10558 23042
rect 10558 22990 10610 23042
rect 10610 22990 10612 23042
rect 10556 22988 10612 22990
rect 10444 20802 10500 20804
rect 10444 20750 10446 20802
rect 10446 20750 10498 20802
rect 10498 20750 10500 20802
rect 10444 20748 10500 20750
rect 10892 21420 10948 21476
rect 11004 24332 11060 24388
rect 11340 28476 11396 28532
rect 11340 27074 11396 27076
rect 11340 27022 11342 27074
rect 11342 27022 11394 27074
rect 11394 27022 11396 27074
rect 11340 27020 11396 27022
rect 12236 41804 12292 41860
rect 12124 41244 12180 41300
rect 12124 39340 12180 39396
rect 12124 37996 12180 38052
rect 12124 36594 12180 36596
rect 12124 36542 12126 36594
rect 12126 36542 12178 36594
rect 12178 36542 12180 36594
rect 12124 36540 12180 36542
rect 12124 35196 12180 35252
rect 12124 34914 12180 34916
rect 12124 34862 12126 34914
rect 12126 34862 12178 34914
rect 12178 34862 12180 34914
rect 12124 34860 12180 34862
rect 13916 42812 13972 42868
rect 13132 42588 13188 42644
rect 12236 34188 12292 34244
rect 12348 39340 12404 39396
rect 12908 39730 12964 39732
rect 12908 39678 12910 39730
rect 12910 39678 12962 39730
rect 12962 39678 12964 39730
rect 12908 39676 12964 39678
rect 12460 38556 12516 38612
rect 12572 38274 12628 38276
rect 12572 38222 12574 38274
rect 12574 38222 12626 38274
rect 12626 38222 12628 38274
rect 12572 38220 12628 38222
rect 12460 37884 12516 37940
rect 12572 34636 12628 34692
rect 12908 38220 12964 38276
rect 12796 36652 12852 36708
rect 13132 38050 13188 38052
rect 13132 37998 13134 38050
rect 13134 37998 13186 38050
rect 13186 37998 13188 38050
rect 13132 37996 13188 37998
rect 13356 38220 13412 38276
rect 13580 37100 13636 37156
rect 13244 36652 13300 36708
rect 12908 34914 12964 34916
rect 12908 34862 12910 34914
rect 12910 34862 12962 34914
rect 12962 34862 12964 34914
rect 12908 34860 12964 34862
rect 13020 34748 13076 34804
rect 13132 35308 13188 35364
rect 13244 34972 13300 35028
rect 13692 34636 13748 34692
rect 12572 34076 12628 34132
rect 11788 32508 11844 32564
rect 12012 31500 12068 31556
rect 11564 24332 11620 24388
rect 11676 31052 11732 31108
rect 11900 31106 11956 31108
rect 11900 31054 11902 31106
rect 11902 31054 11954 31106
rect 11954 31054 11956 31106
rect 11900 31052 11956 31054
rect 12124 29596 12180 29652
rect 11788 29426 11844 29428
rect 11788 29374 11790 29426
rect 11790 29374 11842 29426
rect 11842 29374 11844 29426
rect 11788 29372 11844 29374
rect 12460 29372 12516 29428
rect 11788 28812 11844 28868
rect 11116 22764 11172 22820
rect 11900 28588 11956 28644
rect 11116 22428 11172 22484
rect 10556 20300 10612 20356
rect 10332 19234 10388 19236
rect 10332 19182 10334 19234
rect 10334 19182 10386 19234
rect 10386 19182 10388 19234
rect 10332 19180 10388 19182
rect 10892 19516 10948 19572
rect 10780 18956 10836 19012
rect 11228 19852 11284 19908
rect 11340 22764 11396 22820
rect 11116 19346 11172 19348
rect 11116 19294 11118 19346
rect 11118 19294 11170 19346
rect 11170 19294 11172 19346
rect 11116 19292 11172 19294
rect 11004 18732 11060 18788
rect 10332 18562 10388 18564
rect 10332 18510 10334 18562
rect 10334 18510 10386 18562
rect 10386 18510 10388 18562
rect 10332 18508 10388 18510
rect 10108 18396 10164 18452
rect 9996 17612 10052 17668
rect 9884 17388 9940 17444
rect 9772 16156 9828 16212
rect 11452 21756 11508 21812
rect 11452 21532 11508 21588
rect 11676 21810 11732 21812
rect 11676 21758 11678 21810
rect 11678 21758 11730 21810
rect 11730 21758 11732 21810
rect 11676 21756 11732 21758
rect 12460 28642 12516 28644
rect 12460 28590 12462 28642
rect 12462 28590 12514 28642
rect 12514 28590 12516 28642
rect 12460 28588 12516 28590
rect 12012 25676 12068 25732
rect 12012 24498 12068 24500
rect 12012 24446 12014 24498
rect 12014 24446 12066 24498
rect 12066 24446 12068 24498
rect 12012 24444 12068 24446
rect 12012 23042 12068 23044
rect 12012 22990 12014 23042
rect 12014 22990 12066 23042
rect 12066 22990 12068 23042
rect 12012 22988 12068 22990
rect 11900 22370 11956 22372
rect 11900 22318 11902 22370
rect 11902 22318 11954 22370
rect 11954 22318 11956 22370
rect 11900 22316 11956 22318
rect 11452 20018 11508 20020
rect 11452 19966 11454 20018
rect 11454 19966 11506 20018
rect 11506 19966 11508 20018
rect 11452 19964 11508 19966
rect 11676 19906 11732 19908
rect 11676 19854 11678 19906
rect 11678 19854 11730 19906
rect 11730 19854 11732 19906
rect 11676 19852 11732 19854
rect 11900 20300 11956 20356
rect 11676 19516 11732 19572
rect 11564 19458 11620 19460
rect 11564 19406 11566 19458
rect 11566 19406 11618 19458
rect 11618 19406 11620 19458
rect 11564 19404 11620 19406
rect 11228 18060 11284 18116
rect 10780 17612 10836 17668
rect 11340 17388 11396 17444
rect 10332 16604 10388 16660
rect 10108 16380 10164 16436
rect 10892 16604 10948 16660
rect 9996 16098 10052 16100
rect 9996 16046 9998 16098
rect 9998 16046 10050 16098
rect 10050 16046 10052 16098
rect 9996 16044 10052 16046
rect 9884 15932 9940 15988
rect 9660 15596 9716 15652
rect 9548 15426 9604 15428
rect 9548 15374 9550 15426
rect 9550 15374 9602 15426
rect 9602 15374 9604 15426
rect 9548 15372 9604 15374
rect 10108 15314 10164 15316
rect 10108 15262 10110 15314
rect 10110 15262 10162 15314
rect 10162 15262 10164 15314
rect 10108 15260 10164 15262
rect 9436 14754 9492 14756
rect 9436 14702 9438 14754
rect 9438 14702 9490 14754
rect 9490 14702 9492 14754
rect 9436 14700 9492 14702
rect 9548 14642 9604 14644
rect 9548 14590 9550 14642
rect 9550 14590 9602 14642
rect 9602 14590 9604 14642
rect 9548 14588 9604 14590
rect 9436 14306 9492 14308
rect 9436 14254 9438 14306
rect 9438 14254 9490 14306
rect 9490 14254 9492 14306
rect 9436 14252 9492 14254
rect 9212 13020 9268 13076
rect 10108 14642 10164 14644
rect 10108 14590 10110 14642
rect 10110 14590 10162 14642
rect 10162 14590 10164 14642
rect 10108 14588 10164 14590
rect 11116 16268 11172 16324
rect 11004 15932 11060 15988
rect 10780 15820 10836 15876
rect 10556 15596 10612 15652
rect 11004 15426 11060 15428
rect 11004 15374 11006 15426
rect 11006 15374 11058 15426
rect 11058 15374 11060 15426
rect 11004 15372 11060 15374
rect 11340 15260 11396 15316
rect 10220 14812 10276 14868
rect 9996 14530 10052 14532
rect 9996 14478 9998 14530
rect 9998 14478 10050 14530
rect 10050 14478 10052 14530
rect 9996 14476 10052 14478
rect 9772 13634 9828 13636
rect 9772 13582 9774 13634
rect 9774 13582 9826 13634
rect 9826 13582 9828 13634
rect 9772 13580 9828 13582
rect 9884 13692 9940 13748
rect 9436 13074 9492 13076
rect 9436 13022 9438 13074
rect 9438 13022 9490 13074
rect 9490 13022 9492 13074
rect 9436 13020 9492 13022
rect 9100 12850 9156 12852
rect 9100 12798 9102 12850
rect 9102 12798 9154 12850
rect 9154 12798 9156 12850
rect 9100 12796 9156 12798
rect 10108 12908 10164 12964
rect 9324 12178 9380 12180
rect 9324 12126 9326 12178
rect 9326 12126 9378 12178
rect 9378 12126 9380 12178
rect 9324 12124 9380 12126
rect 9884 12012 9940 12068
rect 10220 12012 10276 12068
rect 8316 8146 8372 8148
rect 8316 8094 8318 8146
rect 8318 8094 8370 8146
rect 8370 8094 8372 8146
rect 8316 8092 8372 8094
rect 9548 10444 9604 10500
rect 8876 9266 8932 9268
rect 8876 9214 8878 9266
rect 8878 9214 8930 9266
rect 8930 9214 8932 9266
rect 8876 9212 8932 9214
rect 11228 14812 11284 14868
rect 11004 14306 11060 14308
rect 11004 14254 11006 14306
rect 11006 14254 11058 14306
rect 11058 14254 11060 14306
rect 11004 14252 11060 14254
rect 10444 11564 10500 11620
rect 10556 13580 10612 13636
rect 10220 11394 10276 11396
rect 10220 11342 10222 11394
rect 10222 11342 10274 11394
rect 10274 11342 10276 11394
rect 10220 11340 10276 11342
rect 10780 13580 10836 13636
rect 10780 12012 10836 12068
rect 11228 11340 11284 11396
rect 11900 19404 11956 19460
rect 11788 19234 11844 19236
rect 11788 19182 11790 19234
rect 11790 19182 11842 19234
rect 11842 19182 11844 19234
rect 11788 19180 11844 19182
rect 11900 18226 11956 18228
rect 11900 18174 11902 18226
rect 11902 18174 11954 18226
rect 11954 18174 11956 18226
rect 11900 18172 11956 18174
rect 12796 31778 12852 31780
rect 12796 31726 12798 31778
rect 12798 31726 12850 31778
rect 12850 31726 12852 31778
rect 12796 31724 12852 31726
rect 13356 34188 13412 34244
rect 13244 31724 13300 31780
rect 12908 29932 12964 29988
rect 12908 28812 12964 28868
rect 12908 26796 12964 26852
rect 13468 26460 13524 26516
rect 13580 28812 13636 28868
rect 13356 26402 13412 26404
rect 13356 26350 13358 26402
rect 13358 26350 13410 26402
rect 13410 26350 13412 26402
rect 13356 26348 13412 26350
rect 13244 26124 13300 26180
rect 12684 25116 12740 25172
rect 12348 24332 12404 24388
rect 12460 24444 12516 24500
rect 12348 23938 12404 23940
rect 12348 23886 12350 23938
rect 12350 23886 12402 23938
rect 12402 23886 12404 23938
rect 12348 23884 12404 23886
rect 12236 23324 12292 23380
rect 12236 22540 12292 22596
rect 12124 21532 12180 21588
rect 12236 21980 12292 22036
rect 13132 24332 13188 24388
rect 12460 21980 12516 22036
rect 12124 21362 12180 21364
rect 12124 21310 12126 21362
rect 12126 21310 12178 21362
rect 12178 21310 12180 21362
rect 12124 21308 12180 21310
rect 12236 20188 12292 20244
rect 12124 19964 12180 20020
rect 13020 22092 13076 22148
rect 13132 21810 13188 21812
rect 13132 21758 13134 21810
rect 13134 21758 13186 21810
rect 13186 21758 13188 21810
rect 13132 21756 13188 21758
rect 12572 21196 12628 21252
rect 12908 21362 12964 21364
rect 12908 21310 12910 21362
rect 12910 21310 12962 21362
rect 12962 21310 12964 21362
rect 12908 21308 12964 21310
rect 12348 19740 12404 19796
rect 11676 16380 11732 16436
rect 12236 16210 12292 16212
rect 12236 16158 12238 16210
rect 12238 16158 12290 16210
rect 12290 16158 12292 16210
rect 12236 16156 12292 16158
rect 12012 15820 12068 15876
rect 11900 15538 11956 15540
rect 11900 15486 11902 15538
rect 11902 15486 11954 15538
rect 11954 15486 11956 15538
rect 11900 15484 11956 15486
rect 11788 15314 11844 15316
rect 11788 15262 11790 15314
rect 11790 15262 11842 15314
rect 11842 15262 11844 15314
rect 11788 15260 11844 15262
rect 12348 15820 12404 15876
rect 12572 19516 12628 19572
rect 12460 15036 12516 15092
rect 11900 13132 11956 13188
rect 12236 12962 12292 12964
rect 12236 12910 12238 12962
rect 12238 12910 12290 12962
rect 12290 12910 12292 12962
rect 12236 12908 12292 12910
rect 12124 12178 12180 12180
rect 12124 12126 12126 12178
rect 12126 12126 12178 12178
rect 12178 12126 12180 12178
rect 12124 12124 12180 12126
rect 12124 11788 12180 11844
rect 11564 11116 11620 11172
rect 12012 11394 12068 11396
rect 12012 11342 12014 11394
rect 12014 11342 12066 11394
rect 12066 11342 12068 11394
rect 12012 11340 12068 11342
rect 9884 9772 9940 9828
rect 9660 9100 9716 9156
rect 9884 8930 9940 8932
rect 9884 8878 9886 8930
rect 9886 8878 9938 8930
rect 9938 8878 9940 8930
rect 9884 8876 9940 8878
rect 10444 10444 10500 10500
rect 11228 10444 11284 10500
rect 10892 9996 10948 10052
rect 10444 9212 10500 9268
rect 12908 20412 12964 20468
rect 12796 20188 12852 20244
rect 13356 24444 13412 24500
rect 13356 20802 13412 20804
rect 13356 20750 13358 20802
rect 13358 20750 13410 20802
rect 13410 20750 13412 20802
rect 13356 20748 13412 20750
rect 13244 20130 13300 20132
rect 13244 20078 13246 20130
rect 13246 20078 13298 20130
rect 13298 20078 13300 20130
rect 13244 20076 13300 20078
rect 13132 19964 13188 20020
rect 13804 32338 13860 32340
rect 13804 32286 13806 32338
rect 13806 32286 13858 32338
rect 13858 32286 13860 32338
rect 13804 32284 13860 32286
rect 14028 35026 14084 35028
rect 14028 34974 14030 35026
rect 14030 34974 14082 35026
rect 14082 34974 14084 35026
rect 14028 34972 14084 34974
rect 13916 31388 13972 31444
rect 13804 30716 13860 30772
rect 14252 36876 14308 36932
rect 14364 48188 14420 48244
rect 18844 55410 18900 55412
rect 18844 55358 18846 55410
rect 18846 55358 18898 55410
rect 18898 55358 18900 55410
rect 18844 55356 18900 55358
rect 17500 53564 17556 53620
rect 18060 55132 18116 55188
rect 15148 52892 15204 52948
rect 14924 47852 14980 47908
rect 14364 36482 14420 36484
rect 14364 36430 14366 36482
rect 14366 36430 14418 36482
rect 14418 36430 14420 36482
rect 14364 36428 14420 36430
rect 14700 36764 14756 36820
rect 14700 36540 14756 36596
rect 14812 36482 14868 36484
rect 14812 36430 14814 36482
rect 14814 36430 14866 36482
rect 14866 36430 14868 36482
rect 14812 36428 14868 36430
rect 14588 33458 14644 33460
rect 14588 33406 14590 33458
rect 14590 33406 14642 33458
rect 14642 33406 14644 33458
rect 14588 33404 14644 33406
rect 14252 31388 14308 31444
rect 14252 30994 14308 30996
rect 14252 30942 14254 30994
rect 14254 30942 14306 30994
rect 14306 30942 14308 30994
rect 14252 30940 14308 30942
rect 14028 27858 14084 27860
rect 14028 27806 14030 27858
rect 14030 27806 14082 27858
rect 14082 27806 14084 27858
rect 14028 27804 14084 27806
rect 13692 27356 13748 27412
rect 13916 26796 13972 26852
rect 13804 25004 13860 25060
rect 13580 23996 13636 24052
rect 13916 24610 13972 24612
rect 13916 24558 13918 24610
rect 13918 24558 13970 24610
rect 13970 24558 13972 24610
rect 13916 24556 13972 24558
rect 14364 28812 14420 28868
rect 14364 28642 14420 28644
rect 14364 28590 14366 28642
rect 14366 28590 14418 28642
rect 14418 28590 14420 28642
rect 14364 28588 14420 28590
rect 15036 38780 15092 38836
rect 17612 52108 17668 52164
rect 16380 48076 16436 48132
rect 17612 47852 17668 47908
rect 16044 41132 16100 41188
rect 15372 40348 15428 40404
rect 15820 39564 15876 39620
rect 15596 37212 15652 37268
rect 15148 34412 15204 34468
rect 15932 35196 15988 35252
rect 15596 33516 15652 33572
rect 14812 31612 14868 31668
rect 14700 30770 14756 30772
rect 14700 30718 14702 30770
rect 14702 30718 14754 30770
rect 14754 30718 14756 30770
rect 14700 30716 14756 30718
rect 14588 28588 14644 28644
rect 14588 27634 14644 27636
rect 14588 27582 14590 27634
rect 14590 27582 14642 27634
rect 14642 27582 14644 27634
rect 14588 27580 14644 27582
rect 14476 27356 14532 27412
rect 14700 27244 14756 27300
rect 15036 31778 15092 31780
rect 15036 31726 15038 31778
rect 15038 31726 15090 31778
rect 15090 31726 15092 31778
rect 15036 31724 15092 31726
rect 15148 31388 15204 31444
rect 15372 31948 15428 32004
rect 14924 28642 14980 28644
rect 14924 28590 14926 28642
rect 14926 28590 14978 28642
rect 14978 28590 14980 28642
rect 14924 28588 14980 28590
rect 14588 26460 14644 26516
rect 14700 26348 14756 26404
rect 14924 25676 14980 25732
rect 14700 24556 14756 24612
rect 14140 24332 14196 24388
rect 14140 23996 14196 24052
rect 13804 23324 13860 23380
rect 13692 22316 13748 22372
rect 13580 21868 13636 21924
rect 13916 22204 13972 22260
rect 13692 21308 13748 21364
rect 13356 19740 13412 19796
rect 13468 19964 13524 20020
rect 12796 18732 12852 18788
rect 13020 17164 13076 17220
rect 13244 19068 13300 19124
rect 13132 17106 13188 17108
rect 13132 17054 13134 17106
rect 13134 17054 13186 17106
rect 13186 17054 13188 17106
rect 13132 17052 13188 17054
rect 13132 16828 13188 16884
rect 13356 18844 13412 18900
rect 13468 17612 13524 17668
rect 13356 17276 13412 17332
rect 13356 16828 13412 16884
rect 13804 20860 13860 20916
rect 13916 19516 13972 19572
rect 13804 19292 13860 19348
rect 13804 18674 13860 18676
rect 13804 18622 13806 18674
rect 13806 18622 13858 18674
rect 13858 18622 13860 18674
rect 13804 18620 13860 18622
rect 13692 18396 13748 18452
rect 13804 18172 13860 18228
rect 13692 17612 13748 17668
rect 14252 23938 14308 23940
rect 14252 23886 14254 23938
rect 14254 23886 14306 23938
rect 14306 23886 14308 23938
rect 14252 23884 14308 23886
rect 14700 23660 14756 23716
rect 14140 23436 14196 23492
rect 14364 22988 14420 23044
rect 14252 21196 14308 21252
rect 14252 20860 14308 20916
rect 14140 19292 14196 19348
rect 14140 19068 14196 19124
rect 14252 19740 14308 19796
rect 14028 18172 14084 18228
rect 14140 18508 14196 18564
rect 13916 17052 13972 17108
rect 14028 16882 14084 16884
rect 14028 16830 14030 16882
rect 14030 16830 14082 16882
rect 14082 16830 14084 16882
rect 14028 16828 14084 16830
rect 14812 23154 14868 23156
rect 14812 23102 14814 23154
rect 14814 23102 14866 23154
rect 14866 23102 14868 23154
rect 14812 23100 14868 23102
rect 14476 22204 14532 22260
rect 14812 21868 14868 21924
rect 14700 21308 14756 21364
rect 14476 20748 14532 20804
rect 14588 20412 14644 20468
rect 14924 21420 14980 21476
rect 14924 20972 14980 21028
rect 14364 19404 14420 19460
rect 14364 18396 14420 18452
rect 14588 18450 14644 18452
rect 14588 18398 14590 18450
rect 14590 18398 14642 18450
rect 14642 18398 14644 18450
rect 14588 18396 14644 18398
rect 14700 19180 14756 19236
rect 14588 18172 14644 18228
rect 14364 17948 14420 18004
rect 14476 17890 14532 17892
rect 14476 17838 14478 17890
rect 14478 17838 14530 17890
rect 14530 17838 14532 17890
rect 14476 17836 14532 17838
rect 13580 16380 13636 16436
rect 14364 16604 14420 16660
rect 13580 15820 13636 15876
rect 13804 16380 13860 16436
rect 13244 14476 13300 14532
rect 12796 12962 12852 12964
rect 12796 12910 12798 12962
rect 12798 12910 12850 12962
rect 12850 12910 12852 12962
rect 12796 12908 12852 12910
rect 11676 9324 11732 9380
rect 12124 8876 12180 8932
rect 10668 7362 10724 7364
rect 10668 7310 10670 7362
rect 10670 7310 10722 7362
rect 10722 7310 10724 7362
rect 10668 7308 10724 7310
rect 11452 5964 11508 6020
rect 10108 5068 10164 5124
rect 3804 3162 3860 3164
rect 3804 3110 3806 3162
rect 3806 3110 3858 3162
rect 3858 3110 3860 3162
rect 3804 3108 3860 3110
rect 3908 3162 3964 3164
rect 3908 3110 3910 3162
rect 3910 3110 3962 3162
rect 3962 3110 3964 3162
rect 3908 3108 3964 3110
rect 4012 3162 4068 3164
rect 4012 3110 4014 3162
rect 4014 3110 4066 3162
rect 4066 3110 4068 3162
rect 4012 3108 4068 3110
rect 4464 2378 4520 2380
rect 4464 2326 4466 2378
rect 4466 2326 4518 2378
rect 4518 2326 4520 2378
rect 4464 2324 4520 2326
rect 4568 2378 4624 2380
rect 4568 2326 4570 2378
rect 4570 2326 4622 2378
rect 4622 2326 4624 2378
rect 4568 2324 4624 2326
rect 4672 2378 4728 2380
rect 4672 2326 4674 2378
rect 4674 2326 4726 2378
rect 4726 2326 4728 2378
rect 4672 2324 4728 2326
rect 3804 1594 3860 1596
rect 3804 1542 3806 1594
rect 3806 1542 3858 1594
rect 3858 1542 3860 1594
rect 3804 1540 3860 1542
rect 3908 1594 3964 1596
rect 3908 1542 3910 1594
rect 3910 1542 3962 1594
rect 3962 1542 3964 1594
rect 3908 1540 3964 1542
rect 4012 1594 4068 1596
rect 4012 1542 4014 1594
rect 4014 1542 4066 1594
rect 4066 1542 4068 1594
rect 4012 1540 4068 1542
rect 4464 810 4520 812
rect 4464 758 4466 810
rect 4466 758 4518 810
rect 4518 758 4520 810
rect 4464 756 4520 758
rect 4568 810 4624 812
rect 4568 758 4570 810
rect 4570 758 4622 810
rect 4622 758 4624 810
rect 4568 756 4624 758
rect 4672 810 4728 812
rect 4672 758 4674 810
rect 4674 758 4726 810
rect 4726 758 4728 810
rect 4672 756 4728 758
rect 3612 140 3668 196
rect 4732 140 4788 196
rect 7420 3052 7476 3108
rect 8764 3052 8820 3108
rect 7980 1372 8036 1428
rect 8764 1596 8820 1652
rect 13132 10444 13188 10500
rect 13132 9826 13188 9828
rect 13132 9774 13134 9826
rect 13134 9774 13186 9826
rect 13186 9774 13188 9826
rect 13132 9772 13188 9774
rect 13356 12348 13412 12404
rect 13244 7980 13300 8036
rect 14588 17052 14644 17108
rect 13916 16156 13972 16212
rect 13580 14028 13636 14084
rect 13916 14252 13972 14308
rect 13580 12572 13636 12628
rect 14140 13244 14196 13300
rect 15148 27804 15204 27860
rect 15708 31724 15764 31780
rect 15932 31388 15988 31444
rect 15820 31218 15876 31220
rect 15820 31166 15822 31218
rect 15822 31166 15874 31218
rect 15874 31166 15876 31218
rect 15820 31164 15876 31166
rect 15596 28588 15652 28644
rect 15932 30156 15988 30212
rect 15820 28476 15876 28532
rect 15596 27580 15652 27636
rect 15148 22594 15204 22596
rect 15148 22542 15150 22594
rect 15150 22542 15202 22594
rect 15202 22542 15204 22594
rect 15148 22540 15204 22542
rect 15148 21532 15204 21588
rect 15260 21474 15316 21476
rect 15260 21422 15262 21474
rect 15262 21422 15314 21474
rect 15314 21422 15316 21474
rect 15260 21420 15316 21422
rect 15148 20076 15204 20132
rect 14924 19292 14980 19348
rect 15484 23436 15540 23492
rect 17836 45612 17892 45668
rect 17052 44268 17108 44324
rect 16716 39618 16772 39620
rect 16716 39566 16718 39618
rect 16718 39566 16770 39618
rect 16770 39566 16772 39618
rect 16716 39564 16772 39566
rect 16828 35196 16884 35252
rect 16604 34076 16660 34132
rect 17724 40402 17780 40404
rect 17724 40350 17726 40402
rect 17726 40350 17778 40402
rect 17778 40350 17780 40402
rect 17724 40348 17780 40350
rect 17276 40124 17332 40180
rect 17164 37212 17220 37268
rect 17164 32620 17220 32676
rect 16828 31836 16884 31892
rect 16268 31724 16324 31780
rect 16156 28364 16212 28420
rect 16044 26572 16100 26628
rect 15708 23100 15764 23156
rect 15820 22370 15876 22372
rect 15820 22318 15822 22370
rect 15822 22318 15874 22370
rect 15874 22318 15876 22370
rect 15820 22316 15876 22318
rect 15820 21586 15876 21588
rect 15820 21534 15822 21586
rect 15822 21534 15874 21586
rect 15874 21534 15876 21586
rect 15820 21532 15876 21534
rect 15708 21362 15764 21364
rect 15708 21310 15710 21362
rect 15710 21310 15762 21362
rect 15762 21310 15764 21362
rect 15708 21308 15764 21310
rect 15596 20076 15652 20132
rect 15820 20748 15876 20804
rect 15484 20018 15540 20020
rect 15484 19966 15486 20018
rect 15486 19966 15538 20018
rect 15538 19966 15540 20018
rect 15484 19964 15540 19966
rect 16716 31666 16772 31668
rect 16716 31614 16718 31666
rect 16718 31614 16770 31666
rect 16770 31614 16772 31666
rect 16716 31612 16772 31614
rect 17948 44156 18004 44212
rect 17500 37938 17556 37940
rect 17500 37886 17502 37938
rect 17502 37886 17554 37938
rect 17554 37886 17556 37938
rect 17500 37884 17556 37886
rect 17388 36258 17444 36260
rect 17388 36206 17390 36258
rect 17390 36206 17442 36258
rect 17442 36206 17444 36258
rect 17388 36204 17444 36206
rect 17724 33516 17780 33572
rect 17612 32284 17668 32340
rect 17052 31164 17108 31220
rect 16716 30604 16772 30660
rect 16380 28476 16436 28532
rect 16828 30210 16884 30212
rect 16828 30158 16830 30210
rect 16830 30158 16882 30210
rect 16882 30158 16884 30210
rect 16828 30156 16884 30158
rect 16940 28476 16996 28532
rect 16492 27020 16548 27076
rect 18284 53116 18340 53172
rect 18508 52668 18564 52724
rect 18060 40236 18116 40292
rect 18284 46844 18340 46900
rect 18284 36652 18340 36708
rect 18284 36204 18340 36260
rect 17948 35026 18004 35028
rect 17948 34974 17950 35026
rect 17950 34974 18002 35026
rect 18002 34974 18004 35026
rect 17948 34972 18004 34974
rect 17948 33234 18004 33236
rect 17948 33182 17950 33234
rect 17950 33182 18002 33234
rect 18002 33182 18004 33234
rect 17948 33180 18004 33182
rect 18844 37772 18900 37828
rect 19404 54626 19460 54628
rect 19404 54574 19406 54626
rect 19406 54574 19458 54626
rect 19458 54574 19460 54626
rect 19404 54572 19460 54574
rect 20188 55356 20244 55412
rect 21084 55916 21140 55972
rect 19516 53228 19572 53284
rect 19964 52220 20020 52276
rect 20524 55298 20580 55300
rect 20524 55246 20526 55298
rect 20526 55246 20578 55298
rect 20578 55246 20580 55298
rect 20524 55244 20580 55246
rect 20636 54290 20692 54292
rect 20636 54238 20638 54290
rect 20638 54238 20690 54290
rect 20690 54238 20692 54290
rect 20636 54236 20692 54238
rect 20524 53730 20580 53732
rect 20524 53678 20526 53730
rect 20526 53678 20578 53730
rect 20578 53678 20580 53730
rect 20524 53676 20580 53678
rect 21980 55916 22036 55972
rect 21644 55804 21700 55860
rect 21308 53618 21364 53620
rect 21308 53566 21310 53618
rect 21310 53566 21362 53618
rect 21362 53566 21364 53618
rect 21308 53564 21364 53566
rect 21420 52946 21476 52948
rect 21420 52894 21422 52946
rect 21422 52894 21474 52946
rect 21474 52894 21476 52946
rect 21420 52892 21476 52894
rect 20860 50428 20916 50484
rect 21084 51100 21140 51156
rect 19628 40236 19684 40292
rect 18508 34130 18564 34132
rect 18508 34078 18510 34130
rect 18510 34078 18562 34130
rect 18562 34078 18564 34130
rect 18508 34076 18564 34078
rect 18396 33570 18452 33572
rect 18396 33518 18398 33570
rect 18398 33518 18450 33570
rect 18450 33518 18452 33570
rect 18396 33516 18452 33518
rect 18284 32786 18340 32788
rect 18284 32734 18286 32786
rect 18286 32734 18338 32786
rect 18338 32734 18340 32786
rect 18284 32732 18340 32734
rect 17164 26796 17220 26852
rect 16380 23436 16436 23492
rect 16940 25228 16996 25284
rect 16380 22540 16436 22596
rect 16268 21868 16324 21924
rect 16380 21586 16436 21588
rect 16380 21534 16382 21586
rect 16382 21534 16434 21586
rect 16434 21534 16436 21586
rect 16380 21532 16436 21534
rect 16156 21308 16212 21364
rect 16604 24498 16660 24500
rect 16604 24446 16606 24498
rect 16606 24446 16658 24498
rect 16658 24446 16660 24498
rect 16604 24444 16660 24446
rect 16828 23714 16884 23716
rect 16828 23662 16830 23714
rect 16830 23662 16882 23714
rect 16882 23662 16884 23714
rect 16828 23660 16884 23662
rect 17164 23772 17220 23828
rect 17836 30604 17892 30660
rect 17052 22652 17108 22708
rect 15932 20300 15988 20356
rect 16044 20524 16100 20580
rect 15596 19794 15652 19796
rect 15596 19742 15598 19794
rect 15598 19742 15650 19794
rect 15650 19742 15652 19794
rect 15596 19740 15652 19742
rect 15372 19404 15428 19460
rect 16268 20412 16324 20468
rect 16828 22092 16884 22148
rect 16716 21308 16772 21364
rect 16716 20802 16772 20804
rect 16716 20750 16718 20802
rect 16718 20750 16770 20802
rect 16770 20750 16772 20802
rect 16716 20748 16772 20750
rect 16716 20578 16772 20580
rect 16716 20526 16718 20578
rect 16718 20526 16770 20578
rect 16770 20526 16772 20578
rect 16716 20524 16772 20526
rect 16156 19292 16212 19348
rect 15148 18620 15204 18676
rect 15708 19180 15764 19236
rect 14924 17612 14980 17668
rect 15036 18396 15092 18452
rect 15260 18060 15316 18116
rect 15148 17948 15204 18004
rect 14924 17164 14980 17220
rect 14812 15820 14868 15876
rect 14924 15202 14980 15204
rect 14924 15150 14926 15202
rect 14926 15150 14978 15202
rect 14978 15150 14980 15202
rect 14924 15148 14980 15150
rect 15596 17052 15652 17108
rect 16044 19068 16100 19124
rect 15820 18674 15876 18676
rect 15820 18622 15822 18674
rect 15822 18622 15874 18674
rect 15874 18622 15876 18674
rect 15820 18620 15876 18622
rect 16268 18562 16324 18564
rect 16268 18510 16270 18562
rect 16270 18510 16322 18562
rect 16322 18510 16324 18562
rect 16268 18508 16324 18510
rect 15932 18060 15988 18116
rect 16044 18172 16100 18228
rect 15372 16604 15428 16660
rect 15260 16492 15316 16548
rect 15260 16210 15316 16212
rect 15260 16158 15262 16210
rect 15262 16158 15314 16210
rect 15314 16158 15316 16210
rect 15260 16156 15316 16158
rect 15708 16210 15764 16212
rect 15708 16158 15710 16210
rect 15710 16158 15762 16210
rect 15762 16158 15764 16210
rect 15708 16156 15764 16158
rect 15372 15932 15428 15988
rect 15372 15708 15428 15764
rect 15708 15932 15764 15988
rect 15148 15596 15204 15652
rect 15260 15426 15316 15428
rect 15260 15374 15262 15426
rect 15262 15374 15314 15426
rect 15314 15374 15316 15426
rect 15260 15372 15316 15374
rect 15484 15148 15540 15204
rect 14700 14028 14756 14084
rect 15036 14700 15092 14756
rect 14588 13244 14644 13300
rect 14252 11788 14308 11844
rect 14476 11900 14532 11956
rect 14924 13468 14980 13524
rect 15484 14924 15540 14980
rect 15148 14476 15204 14532
rect 14028 10780 14084 10836
rect 13916 8764 13972 8820
rect 15260 14812 15316 14868
rect 16044 16940 16100 16996
rect 16156 17052 16212 17108
rect 16604 19964 16660 20020
rect 17164 21474 17220 21476
rect 17164 21422 17166 21474
rect 17166 21422 17218 21474
rect 17218 21422 17220 21474
rect 17164 21420 17220 21422
rect 17052 20860 17108 20916
rect 17052 20578 17108 20580
rect 17052 20526 17054 20578
rect 17054 20526 17106 20578
rect 17106 20526 17108 20578
rect 17052 20524 17108 20526
rect 16716 19516 16772 19572
rect 16604 19404 16660 19460
rect 16492 18226 16548 18228
rect 16492 18174 16494 18226
rect 16494 18174 16546 18226
rect 16546 18174 16548 18226
rect 16492 18172 16548 18174
rect 16380 16882 16436 16884
rect 16380 16830 16382 16882
rect 16382 16830 16434 16882
rect 16434 16830 16436 16882
rect 16380 16828 16436 16830
rect 16156 15932 16212 15988
rect 16044 15874 16100 15876
rect 16044 15822 16046 15874
rect 16046 15822 16098 15874
rect 16098 15822 16100 15874
rect 16044 15820 16100 15822
rect 15932 15372 15988 15428
rect 16044 15314 16100 15316
rect 16044 15262 16046 15314
rect 16046 15262 16098 15314
rect 16098 15262 16100 15314
rect 16044 15260 16100 15262
rect 15708 14812 15764 14868
rect 16044 14812 16100 14868
rect 15932 14642 15988 14644
rect 15932 14590 15934 14642
rect 15934 14590 15986 14642
rect 15986 14590 15988 14642
rect 15932 14588 15988 14590
rect 16044 14476 16100 14532
rect 16716 19068 16772 19124
rect 16828 18620 16884 18676
rect 17052 18620 17108 18676
rect 16940 18396 16996 18452
rect 17052 18226 17108 18228
rect 17052 18174 17054 18226
rect 17054 18174 17106 18226
rect 17106 18174 17108 18226
rect 17052 18172 17108 18174
rect 17164 17948 17220 18004
rect 17500 27970 17556 27972
rect 17500 27918 17502 27970
rect 17502 27918 17554 27970
rect 17554 27918 17556 27970
rect 17500 27916 17556 27918
rect 17724 27916 17780 27972
rect 17388 27692 17444 27748
rect 17724 27074 17780 27076
rect 17724 27022 17726 27074
rect 17726 27022 17778 27074
rect 17778 27022 17780 27074
rect 17724 27020 17780 27022
rect 17500 25676 17556 25732
rect 17724 24332 17780 24388
rect 17388 22316 17444 22372
rect 17388 20748 17444 20804
rect 17388 18226 17444 18228
rect 17388 18174 17390 18226
rect 17390 18174 17442 18226
rect 17442 18174 17444 18226
rect 17388 18172 17444 18174
rect 16940 17836 16996 17892
rect 16716 16828 16772 16884
rect 16940 17612 16996 17668
rect 16940 17052 16996 17108
rect 16716 16492 16772 16548
rect 16604 16044 16660 16100
rect 16492 15426 16548 15428
rect 16492 15374 16494 15426
rect 16494 15374 16546 15426
rect 16546 15374 16548 15426
rect 16492 15372 16548 15374
rect 17276 15708 17332 15764
rect 16716 15148 16772 15204
rect 16828 15260 16884 15316
rect 16492 14588 16548 14644
rect 16268 14364 16324 14420
rect 15372 13634 15428 13636
rect 15372 13582 15374 13634
rect 15374 13582 15426 13634
rect 15426 13582 15428 13634
rect 15372 13580 15428 13582
rect 15260 13356 15316 13412
rect 15820 13356 15876 13412
rect 15148 12124 15204 12180
rect 15260 13074 15316 13076
rect 15260 13022 15262 13074
rect 15262 13022 15314 13074
rect 15314 13022 15316 13074
rect 15260 13020 15316 13022
rect 15036 12012 15092 12068
rect 14588 4844 14644 4900
rect 15148 9772 15204 9828
rect 14140 3612 14196 3668
rect 13020 2940 13076 2996
rect 13580 2492 13636 2548
rect 12124 1596 12180 1652
rect 12796 1596 12852 1652
rect 15484 12850 15540 12852
rect 15484 12798 15486 12850
rect 15486 12798 15538 12850
rect 15538 12798 15540 12850
rect 15484 12796 15540 12798
rect 16380 14028 16436 14084
rect 16156 13580 16212 13636
rect 16716 14530 16772 14532
rect 16716 14478 16718 14530
rect 16718 14478 16770 14530
rect 16770 14478 16772 14530
rect 16716 14476 16772 14478
rect 16828 14364 16884 14420
rect 17052 14924 17108 14980
rect 16940 14140 16996 14196
rect 17164 14812 17220 14868
rect 16716 13356 16772 13412
rect 16044 12796 16100 12852
rect 16156 12684 16212 12740
rect 16604 12124 16660 12180
rect 16156 10668 16212 10724
rect 16492 12012 16548 12068
rect 16492 7196 16548 7252
rect 17612 21532 17668 21588
rect 17500 14924 17556 14980
rect 17612 15820 17668 15876
rect 17388 14812 17444 14868
rect 17500 13468 17556 13524
rect 18172 31890 18228 31892
rect 18172 31838 18174 31890
rect 18174 31838 18226 31890
rect 18226 31838 18228 31890
rect 18172 31836 18228 31838
rect 18172 27916 18228 27972
rect 18172 26796 18228 26852
rect 17948 22652 18004 22708
rect 18172 25004 18228 25060
rect 18172 24332 18228 24388
rect 18172 22764 18228 22820
rect 18620 32674 18676 32676
rect 18620 32622 18622 32674
rect 18622 32622 18674 32674
rect 18674 32622 18676 32674
rect 18620 32620 18676 32622
rect 18396 29036 18452 29092
rect 18396 25676 18452 25732
rect 18732 29036 18788 29092
rect 18956 32732 19012 32788
rect 19068 32562 19124 32564
rect 19068 32510 19070 32562
rect 19070 32510 19122 32562
rect 19122 32510 19124 32562
rect 19068 32508 19124 32510
rect 19180 31724 19236 31780
rect 19068 31612 19124 31668
rect 18956 28812 19012 28868
rect 19068 27580 19124 27636
rect 18620 26012 18676 26068
rect 18508 25618 18564 25620
rect 18508 25566 18510 25618
rect 18510 25566 18562 25618
rect 18562 25566 18564 25618
rect 18508 25564 18564 25566
rect 18396 25340 18452 25396
rect 18396 25004 18452 25060
rect 18396 23548 18452 23604
rect 18508 23772 18564 23828
rect 18508 22764 18564 22820
rect 17836 21420 17892 21476
rect 17724 12796 17780 12852
rect 17836 20524 17892 20580
rect 17164 9884 17220 9940
rect 16716 9660 16772 9716
rect 16604 6524 16660 6580
rect 15932 6076 15988 6132
rect 15260 5180 15316 5236
rect 16828 4508 16884 4564
rect 15148 1372 15204 1428
rect 15484 1596 15540 1652
rect 18284 21474 18340 21476
rect 18284 21422 18286 21474
rect 18286 21422 18338 21474
rect 18338 21422 18340 21474
rect 18284 21420 18340 21422
rect 17948 16882 18004 16884
rect 17948 16830 17950 16882
rect 17950 16830 18002 16882
rect 18002 16830 18004 16882
rect 17948 16828 18004 16830
rect 17948 16492 18004 16548
rect 17948 14812 18004 14868
rect 17948 10780 18004 10836
rect 17836 4060 17892 4116
rect 18284 18844 18340 18900
rect 18732 23548 18788 23604
rect 18732 21698 18788 21700
rect 18732 21646 18734 21698
rect 18734 21646 18786 21698
rect 18786 21646 18788 21698
rect 18732 21644 18788 21646
rect 18284 18620 18340 18676
rect 18396 18396 18452 18452
rect 18956 25564 19012 25620
rect 18956 23548 19012 23604
rect 18508 18172 18564 18228
rect 18508 16492 18564 16548
rect 18956 18396 19012 18452
rect 18956 18226 19012 18228
rect 18956 18174 18958 18226
rect 18958 18174 19010 18226
rect 19010 18174 19012 18226
rect 18956 18172 19012 18174
rect 18396 14252 18452 14308
rect 18284 4284 18340 4340
rect 19516 32508 19572 32564
rect 19516 28140 19572 28196
rect 19740 35308 19796 35364
rect 19852 35026 19908 35028
rect 19852 34974 19854 35026
rect 19854 34974 19906 35026
rect 19906 34974 19908 35026
rect 19852 34972 19908 34974
rect 19852 31778 19908 31780
rect 19852 31726 19854 31778
rect 19854 31726 19906 31778
rect 19906 31726 19908 31778
rect 19852 31724 19908 31726
rect 19852 30994 19908 30996
rect 19852 30942 19854 30994
rect 19854 30942 19906 30994
rect 19906 30942 19908 30994
rect 19852 30940 19908 30942
rect 19740 29426 19796 29428
rect 19740 29374 19742 29426
rect 19742 29374 19794 29426
rect 19794 29374 19796 29426
rect 19740 29372 19796 29374
rect 19964 29372 20020 29428
rect 20076 46396 20132 46452
rect 19740 28924 19796 28980
rect 20076 28924 20132 28980
rect 20188 29372 20244 29428
rect 19292 27580 19348 27636
rect 19516 27468 19572 27524
rect 19180 26066 19236 26068
rect 19180 26014 19182 26066
rect 19182 26014 19234 26066
rect 19234 26014 19236 26066
rect 19180 26012 19236 26014
rect 19292 25676 19348 25732
rect 19628 26124 19684 26180
rect 19740 25506 19796 25508
rect 19740 25454 19742 25506
rect 19742 25454 19794 25506
rect 19794 25454 19796 25506
rect 19740 25452 19796 25454
rect 19404 24108 19460 24164
rect 19404 23772 19460 23828
rect 20076 28642 20132 28644
rect 20076 28590 20078 28642
rect 20078 28590 20130 28642
rect 20130 28590 20132 28642
rect 20076 28588 20132 28590
rect 20076 28028 20132 28084
rect 19964 25340 20020 25396
rect 19404 21868 19460 21924
rect 19180 21644 19236 21700
rect 19292 21474 19348 21476
rect 19292 21422 19294 21474
rect 19294 21422 19346 21474
rect 19346 21422 19348 21474
rect 19292 21420 19348 21422
rect 19068 8876 19124 8932
rect 19740 20860 19796 20916
rect 19516 18450 19572 18452
rect 19516 18398 19518 18450
rect 19518 18398 19570 18450
rect 19570 18398 19572 18450
rect 19516 18396 19572 18398
rect 19964 16604 20020 16660
rect 20188 25900 20244 25956
rect 20972 45836 21028 45892
rect 20412 44380 20468 44436
rect 20412 28812 20468 28868
rect 20412 20914 20468 20916
rect 20412 20862 20414 20914
rect 20414 20862 20466 20914
rect 20466 20862 20468 20914
rect 20412 20860 20468 20862
rect 20636 25452 20692 25508
rect 20524 20300 20580 20356
rect 20748 21084 20804 21140
rect 20300 12684 20356 12740
rect 20076 5068 20132 5124
rect 20972 7308 21028 7364
rect 21532 37324 21588 37380
rect 21644 53676 21700 53732
rect 21532 35420 21588 35476
rect 21308 25452 21364 25508
rect 21084 5964 21140 6020
rect 21196 20300 21252 20356
rect 20748 1148 20804 1204
rect 20860 3276 20916 3332
rect 19404 924 19460 980
rect 19180 140 19236 196
rect 19516 140 19572 196
rect 21308 9212 21364 9268
rect 21532 21532 21588 21588
rect 21420 16828 21476 16884
rect 21868 53452 21924 53508
rect 21756 53116 21812 53172
rect 23804 56474 23860 56476
rect 23804 56422 23806 56474
rect 23806 56422 23858 56474
rect 23858 56422 23860 56474
rect 23804 56420 23860 56422
rect 23908 56474 23964 56476
rect 23908 56422 23910 56474
rect 23910 56422 23962 56474
rect 23962 56422 23964 56474
rect 23908 56420 23964 56422
rect 24012 56474 24068 56476
rect 24012 56422 24014 56474
rect 24014 56422 24066 56474
rect 24066 56422 24068 56474
rect 24012 56420 24068 56422
rect 23548 56252 23604 56308
rect 24444 56306 24500 56308
rect 24444 56254 24446 56306
rect 24446 56254 24498 56306
rect 24498 56254 24500 56306
rect 24444 56252 24500 56254
rect 25452 57260 25508 57316
rect 24892 56252 24948 56308
rect 25116 57148 25172 57204
rect 23548 56028 23604 56084
rect 23436 55468 23492 55524
rect 22316 53900 22372 53956
rect 22652 53228 22708 53284
rect 22204 52722 22260 52724
rect 22204 52670 22206 52722
rect 22206 52670 22258 52722
rect 22258 52670 22260 52722
rect 22204 52668 22260 52670
rect 22764 52274 22820 52276
rect 22764 52222 22766 52274
rect 22766 52222 22818 52274
rect 22818 52222 22820 52274
rect 22764 52220 22820 52222
rect 22204 36652 22260 36708
rect 21868 27356 21924 27412
rect 21868 21644 21924 21700
rect 21644 16716 21700 16772
rect 21420 5628 21476 5684
rect 21196 2044 21252 2100
rect 22876 51436 22932 51492
rect 22652 40348 22708 40404
rect 22652 9324 22708 9380
rect 23100 51324 23156 51380
rect 22988 49868 23044 49924
rect 23884 55970 23940 55972
rect 23884 55918 23886 55970
rect 23886 55918 23938 55970
rect 23938 55918 23940 55970
rect 23884 55916 23940 55918
rect 24464 55690 24520 55692
rect 24464 55638 24466 55690
rect 24466 55638 24518 55690
rect 24518 55638 24520 55690
rect 24464 55636 24520 55638
rect 24568 55690 24624 55692
rect 24568 55638 24570 55690
rect 24570 55638 24622 55690
rect 24622 55638 24624 55690
rect 24568 55636 24624 55638
rect 24672 55690 24728 55692
rect 24672 55638 24674 55690
rect 24674 55638 24726 55690
rect 24726 55638 24728 55690
rect 24672 55636 24728 55638
rect 24780 55356 24836 55412
rect 23660 55298 23716 55300
rect 23660 55246 23662 55298
rect 23662 55246 23714 55298
rect 23714 55246 23716 55298
rect 23660 55244 23716 55246
rect 24668 55132 24724 55188
rect 24332 55020 24388 55076
rect 23804 54906 23860 54908
rect 23804 54854 23806 54906
rect 23806 54854 23858 54906
rect 23858 54854 23860 54906
rect 23804 54852 23860 54854
rect 23908 54906 23964 54908
rect 23908 54854 23910 54906
rect 23910 54854 23962 54906
rect 23962 54854 23964 54906
rect 23908 54852 23964 54854
rect 24012 54906 24068 54908
rect 24012 54854 24014 54906
rect 24014 54854 24066 54906
rect 24066 54854 24068 54906
rect 24012 54852 24068 54854
rect 24220 54908 24276 54964
rect 23660 54460 23716 54516
rect 23772 54124 23828 54180
rect 23804 53338 23860 53340
rect 23804 53286 23806 53338
rect 23806 53286 23858 53338
rect 23858 53286 23860 53338
rect 23804 53284 23860 53286
rect 23908 53338 23964 53340
rect 23908 53286 23910 53338
rect 23910 53286 23962 53338
rect 23962 53286 23964 53338
rect 23908 53284 23964 53286
rect 24012 53338 24068 53340
rect 24012 53286 24014 53338
rect 24014 53286 24066 53338
rect 24066 53286 24068 53338
rect 24012 53284 24068 53286
rect 24108 53170 24164 53172
rect 24108 53118 24110 53170
rect 24110 53118 24162 53170
rect 24162 53118 24164 53170
rect 24108 53116 24164 53118
rect 23804 51770 23860 51772
rect 23804 51718 23806 51770
rect 23806 51718 23858 51770
rect 23858 51718 23860 51770
rect 23804 51716 23860 51718
rect 23908 51770 23964 51772
rect 23908 51718 23910 51770
rect 23910 51718 23962 51770
rect 23962 51718 23964 51770
rect 23908 51716 23964 51718
rect 24012 51770 24068 51772
rect 24012 51718 24014 51770
rect 24014 51718 24066 51770
rect 24066 51718 24068 51770
rect 24012 51716 24068 51718
rect 24668 54514 24724 54516
rect 24668 54462 24670 54514
rect 24670 54462 24722 54514
rect 24722 54462 24724 54514
rect 24668 54460 24724 54462
rect 24780 54236 24836 54292
rect 25004 55244 25060 55300
rect 24464 54122 24520 54124
rect 24464 54070 24466 54122
rect 24466 54070 24518 54122
rect 24518 54070 24520 54122
rect 24464 54068 24520 54070
rect 24568 54122 24624 54124
rect 24568 54070 24570 54122
rect 24570 54070 24622 54122
rect 24622 54070 24624 54122
rect 24568 54068 24624 54070
rect 24672 54122 24728 54124
rect 24672 54070 24674 54122
rect 24674 54070 24726 54122
rect 24726 54070 24728 54122
rect 24672 54068 24728 54070
rect 24892 53730 24948 53732
rect 24892 53678 24894 53730
rect 24894 53678 24946 53730
rect 24946 53678 24948 53730
rect 24892 53676 24948 53678
rect 24668 53004 24724 53060
rect 24464 52554 24520 52556
rect 24464 52502 24466 52554
rect 24466 52502 24518 52554
rect 24518 52502 24520 52554
rect 24464 52500 24520 52502
rect 24568 52554 24624 52556
rect 24568 52502 24570 52554
rect 24570 52502 24622 52554
rect 24622 52502 24624 52554
rect 24568 52500 24624 52502
rect 24672 52554 24728 52556
rect 24672 52502 24674 52554
rect 24674 52502 24726 52554
rect 24726 52502 24728 52554
rect 24672 52500 24728 52502
rect 24668 52332 24724 52388
rect 24668 51266 24724 51268
rect 24668 51214 24670 51266
rect 24670 51214 24722 51266
rect 24722 51214 24724 51266
rect 24668 51212 24724 51214
rect 23772 51154 23828 51156
rect 23772 51102 23774 51154
rect 23774 51102 23826 51154
rect 23826 51102 23828 51154
rect 23772 51100 23828 51102
rect 24464 50986 24520 50988
rect 24464 50934 24466 50986
rect 24466 50934 24518 50986
rect 24518 50934 24520 50986
rect 24464 50932 24520 50934
rect 24568 50986 24624 50988
rect 24568 50934 24570 50986
rect 24570 50934 24622 50986
rect 24622 50934 24624 50986
rect 24568 50932 24624 50934
rect 24672 50986 24728 50988
rect 24672 50934 24674 50986
rect 24674 50934 24726 50986
rect 24726 50934 24728 50986
rect 24672 50932 24728 50934
rect 23212 39340 23268 39396
rect 22764 3612 22820 3668
rect 22876 30940 22932 30996
rect 22428 1260 22484 1316
rect 23100 29932 23156 29988
rect 22988 21308 23044 21364
rect 23100 19068 23156 19124
rect 23804 50202 23860 50204
rect 23804 50150 23806 50202
rect 23806 50150 23858 50202
rect 23858 50150 23860 50202
rect 23804 50148 23860 50150
rect 23908 50202 23964 50204
rect 23908 50150 23910 50202
rect 23910 50150 23962 50202
rect 23962 50150 23964 50202
rect 23908 50148 23964 50150
rect 24012 50202 24068 50204
rect 24012 50150 24014 50202
rect 24014 50150 24066 50202
rect 24066 50150 24068 50202
rect 24012 50148 24068 50150
rect 24220 49922 24276 49924
rect 24220 49870 24222 49922
rect 24222 49870 24274 49922
rect 24274 49870 24276 49922
rect 24220 49868 24276 49870
rect 24668 49532 24724 49588
rect 24464 49418 24520 49420
rect 24464 49366 24466 49418
rect 24466 49366 24518 49418
rect 24518 49366 24520 49418
rect 24464 49364 24520 49366
rect 24568 49418 24624 49420
rect 24568 49366 24570 49418
rect 24570 49366 24622 49418
rect 24622 49366 24624 49418
rect 24568 49364 24624 49366
rect 24672 49418 24728 49420
rect 24672 49366 24674 49418
rect 24674 49366 24726 49418
rect 24726 49366 24728 49418
rect 24672 49364 24728 49366
rect 23772 49196 23828 49252
rect 24668 48860 24724 48916
rect 23804 48634 23860 48636
rect 23804 48582 23806 48634
rect 23806 48582 23858 48634
rect 23858 48582 23860 48634
rect 23804 48580 23860 48582
rect 23908 48634 23964 48636
rect 23908 48582 23910 48634
rect 23910 48582 23962 48634
rect 23962 48582 23964 48634
rect 23908 48580 23964 48582
rect 24012 48634 24068 48636
rect 24012 48582 24014 48634
rect 24014 48582 24066 48634
rect 24066 48582 24068 48634
rect 24012 48580 24068 48582
rect 25116 53116 25172 53172
rect 25340 56700 25396 56756
rect 26236 57260 26292 57316
rect 26012 56306 26068 56308
rect 26012 56254 26014 56306
rect 26014 56254 26066 56306
rect 26066 56254 26068 56306
rect 26012 56252 26068 56254
rect 25564 54460 25620 54516
rect 25564 53618 25620 53620
rect 25564 53566 25566 53618
rect 25566 53566 25618 53618
rect 25618 53566 25620 53618
rect 25564 53564 25620 53566
rect 25452 52668 25508 52724
rect 25564 51772 25620 51828
rect 25564 50482 25620 50484
rect 25564 50430 25566 50482
rect 25566 50430 25618 50482
rect 25618 50430 25620 50482
rect 25564 50428 25620 50430
rect 27580 56028 27636 56084
rect 25676 49532 25732 49588
rect 25676 48636 25732 48692
rect 24892 48188 24948 48244
rect 25340 48018 25396 48020
rect 25340 47966 25342 48018
rect 25342 47966 25394 48018
rect 25394 47966 25396 48018
rect 25340 47964 25396 47966
rect 24464 47850 24520 47852
rect 24464 47798 24466 47850
rect 24466 47798 24518 47850
rect 24518 47798 24520 47850
rect 24464 47796 24520 47798
rect 24568 47850 24624 47852
rect 24568 47798 24570 47850
rect 24570 47798 24622 47850
rect 24622 47798 24624 47850
rect 24568 47796 24624 47798
rect 24672 47850 24728 47852
rect 24672 47798 24674 47850
rect 24674 47798 24726 47850
rect 24726 47798 24728 47850
rect 24672 47796 24728 47798
rect 24332 47180 24388 47236
rect 23804 47066 23860 47068
rect 23804 47014 23806 47066
rect 23806 47014 23858 47066
rect 23858 47014 23860 47066
rect 23804 47012 23860 47014
rect 23908 47066 23964 47068
rect 23908 47014 23910 47066
rect 23910 47014 23962 47066
rect 23962 47014 23964 47066
rect 23908 47012 23964 47014
rect 24012 47066 24068 47068
rect 24012 47014 24014 47066
rect 24014 47014 24066 47066
rect 24066 47014 24068 47066
rect 24012 47012 24068 47014
rect 25676 47346 25732 47348
rect 25676 47294 25678 47346
rect 25678 47294 25730 47346
rect 25730 47294 25732 47346
rect 25676 47292 25732 47294
rect 24668 46396 24724 46452
rect 24464 46282 24520 46284
rect 24464 46230 24466 46282
rect 24466 46230 24518 46282
rect 24518 46230 24520 46282
rect 24464 46228 24520 46230
rect 24568 46282 24624 46284
rect 24568 46230 24570 46282
rect 24570 46230 24622 46282
rect 24622 46230 24624 46282
rect 24568 46228 24624 46230
rect 24672 46282 24728 46284
rect 24672 46230 24674 46282
rect 24674 46230 24726 46282
rect 24726 46230 24728 46282
rect 24672 46228 24728 46230
rect 24668 45890 24724 45892
rect 24668 45838 24670 45890
rect 24670 45838 24722 45890
rect 24722 45838 24724 45890
rect 24668 45836 24724 45838
rect 23804 45498 23860 45500
rect 23804 45446 23806 45498
rect 23806 45446 23858 45498
rect 23858 45446 23860 45498
rect 23804 45444 23860 45446
rect 23908 45498 23964 45500
rect 23908 45446 23910 45498
rect 23910 45446 23962 45498
rect 23962 45446 23964 45498
rect 23908 45444 23964 45446
rect 24012 45498 24068 45500
rect 24012 45446 24014 45498
rect 24014 45446 24066 45498
rect 24066 45446 24068 45498
rect 24012 45444 24068 45446
rect 24464 44714 24520 44716
rect 24464 44662 24466 44714
rect 24466 44662 24518 44714
rect 24518 44662 24520 44714
rect 24464 44660 24520 44662
rect 24568 44714 24624 44716
rect 24568 44662 24570 44714
rect 24570 44662 24622 44714
rect 24622 44662 24624 44714
rect 24568 44660 24624 44662
rect 24672 44714 24728 44716
rect 24672 44662 24674 44714
rect 24674 44662 24726 44714
rect 24726 44662 24728 44714
rect 24672 44660 24728 44662
rect 25676 46396 25732 46452
rect 25676 45500 25732 45556
rect 24892 44492 24948 44548
rect 26236 54402 26292 54404
rect 26236 54350 26238 54402
rect 26238 54350 26290 54402
rect 26290 54350 26292 54402
rect 26236 54348 26292 54350
rect 26796 53676 26852 53732
rect 26236 52834 26292 52836
rect 26236 52782 26238 52834
rect 26238 52782 26290 52834
rect 26290 52782 26292 52834
rect 26236 52780 26292 52782
rect 26236 52162 26292 52164
rect 26236 52110 26238 52162
rect 26238 52110 26290 52162
rect 26290 52110 26292 52162
rect 26236 52108 26292 52110
rect 26348 51884 26404 51940
rect 26236 50764 26292 50820
rect 26236 49026 26292 49028
rect 26236 48974 26238 49026
rect 26238 48974 26290 49026
rect 26290 48974 26292 49026
rect 26236 48972 26292 48974
rect 26348 48748 26404 48804
rect 26236 48130 26292 48132
rect 26236 48078 26238 48130
rect 26238 48078 26290 48130
rect 26290 48078 26292 48130
rect 26236 48076 26292 48078
rect 26124 46060 26180 46116
rect 25900 44380 25956 44436
rect 25676 44210 25732 44212
rect 25676 44158 25678 44210
rect 25678 44158 25730 44210
rect 25730 44158 25732 44210
rect 25676 44156 25732 44158
rect 24668 44044 24724 44100
rect 23804 43930 23860 43932
rect 23804 43878 23806 43930
rect 23806 43878 23858 43930
rect 23858 43878 23860 43930
rect 23804 43876 23860 43878
rect 23908 43930 23964 43932
rect 23908 43878 23910 43930
rect 23910 43878 23962 43930
rect 23962 43878 23964 43930
rect 23908 43876 23964 43878
rect 24012 43930 24068 43932
rect 24012 43878 24014 43930
rect 24014 43878 24066 43930
rect 24066 43878 24068 43930
rect 24012 43876 24068 43878
rect 24464 43146 24520 43148
rect 24464 43094 24466 43146
rect 24466 43094 24518 43146
rect 24518 43094 24520 43146
rect 24464 43092 24520 43094
rect 24568 43146 24624 43148
rect 24568 43094 24570 43146
rect 24570 43094 24622 43146
rect 24622 43094 24624 43146
rect 24568 43092 24624 43094
rect 24672 43146 24728 43148
rect 24672 43094 24674 43146
rect 24674 43094 24726 43146
rect 24726 43094 24728 43146
rect 24672 43092 24728 43094
rect 24668 42588 24724 42644
rect 23804 42362 23860 42364
rect 23804 42310 23806 42362
rect 23806 42310 23858 42362
rect 23858 42310 23860 42362
rect 23804 42308 23860 42310
rect 23908 42362 23964 42364
rect 23908 42310 23910 42362
rect 23910 42310 23962 42362
rect 23962 42310 23964 42362
rect 23908 42308 23964 42310
rect 24012 42362 24068 42364
rect 24012 42310 24014 42362
rect 24014 42310 24066 42362
rect 24066 42310 24068 42362
rect 24012 42308 24068 42310
rect 24464 41578 24520 41580
rect 24464 41526 24466 41578
rect 24466 41526 24518 41578
rect 24518 41526 24520 41578
rect 24464 41524 24520 41526
rect 24568 41578 24624 41580
rect 24568 41526 24570 41578
rect 24570 41526 24622 41578
rect 24622 41526 24624 41578
rect 24568 41524 24624 41526
rect 24672 41578 24728 41580
rect 24672 41526 24674 41578
rect 24674 41526 24726 41578
rect 24726 41526 24728 41578
rect 24672 41524 24728 41526
rect 23804 40794 23860 40796
rect 23804 40742 23806 40794
rect 23806 40742 23858 40794
rect 23858 40742 23860 40794
rect 23804 40740 23860 40742
rect 23908 40794 23964 40796
rect 23908 40742 23910 40794
rect 23910 40742 23962 40794
rect 23962 40742 23964 40794
rect 23908 40740 23964 40742
rect 24012 40794 24068 40796
rect 24012 40742 24014 40794
rect 24014 40742 24066 40794
rect 24066 40742 24068 40794
rect 24012 40740 24068 40742
rect 24668 40402 24724 40404
rect 24668 40350 24670 40402
rect 24670 40350 24722 40402
rect 24722 40350 24724 40402
rect 24668 40348 24724 40350
rect 25676 43260 25732 43316
rect 25676 42364 25732 42420
rect 25676 41074 25732 41076
rect 25676 41022 25678 41074
rect 25678 41022 25730 41074
rect 25730 41022 25732 41074
rect 25676 41020 25732 41022
rect 24892 40572 24948 40628
rect 24780 40124 24836 40180
rect 25676 40124 25732 40180
rect 24464 40010 24520 40012
rect 24464 39958 24466 40010
rect 24466 39958 24518 40010
rect 24518 39958 24520 40010
rect 24464 39956 24520 39958
rect 24568 40010 24624 40012
rect 24568 39958 24570 40010
rect 24570 39958 24622 40010
rect 24622 39958 24624 40010
rect 24568 39956 24624 39958
rect 24672 40010 24728 40012
rect 24672 39958 24674 40010
rect 24674 39958 24726 40010
rect 24726 39958 24728 40010
rect 24672 39956 24728 39958
rect 24668 39730 24724 39732
rect 24668 39678 24670 39730
rect 24670 39678 24722 39730
rect 24722 39678 24724 39730
rect 24668 39676 24724 39678
rect 23804 39226 23860 39228
rect 23804 39174 23806 39226
rect 23806 39174 23858 39226
rect 23858 39174 23860 39226
rect 23804 39172 23860 39174
rect 23908 39226 23964 39228
rect 23908 39174 23910 39226
rect 23910 39174 23962 39226
rect 23962 39174 23964 39226
rect 23908 39172 23964 39174
rect 24012 39226 24068 39228
rect 24012 39174 24014 39226
rect 24014 39174 24066 39226
rect 24066 39174 24068 39226
rect 25676 39228 25732 39284
rect 24012 39172 24068 39174
rect 24464 38442 24520 38444
rect 24464 38390 24466 38442
rect 24466 38390 24518 38442
rect 24518 38390 24520 38442
rect 24464 38388 24520 38390
rect 24568 38442 24624 38444
rect 24568 38390 24570 38442
rect 24570 38390 24622 38442
rect 24622 38390 24624 38442
rect 24568 38388 24624 38390
rect 24672 38442 24728 38444
rect 24672 38390 24674 38442
rect 24674 38390 24726 38442
rect 24726 38390 24728 38442
rect 24672 38388 24728 38390
rect 23804 37658 23860 37660
rect 23804 37606 23806 37658
rect 23806 37606 23858 37658
rect 23858 37606 23860 37658
rect 23804 37604 23860 37606
rect 23908 37658 23964 37660
rect 23908 37606 23910 37658
rect 23910 37606 23962 37658
rect 23962 37606 23964 37658
rect 23908 37604 23964 37606
rect 24012 37658 24068 37660
rect 24012 37606 24014 37658
rect 24014 37606 24066 37658
rect 24066 37606 24068 37658
rect 24012 37604 24068 37606
rect 23660 36092 23716 36148
rect 23548 33852 23604 33908
rect 23804 36090 23860 36092
rect 23804 36038 23806 36090
rect 23806 36038 23858 36090
rect 23858 36038 23860 36090
rect 23804 36036 23860 36038
rect 23908 36090 23964 36092
rect 23908 36038 23910 36090
rect 23910 36038 23962 36090
rect 23962 36038 23964 36090
rect 23908 36036 23964 36038
rect 24012 36090 24068 36092
rect 24012 36038 24014 36090
rect 24014 36038 24066 36090
rect 24066 36038 24068 36090
rect 24012 36036 24068 36038
rect 23804 34522 23860 34524
rect 23804 34470 23806 34522
rect 23806 34470 23858 34522
rect 23858 34470 23860 34522
rect 23804 34468 23860 34470
rect 23908 34522 23964 34524
rect 23908 34470 23910 34522
rect 23910 34470 23962 34522
rect 23962 34470 23964 34522
rect 23908 34468 23964 34470
rect 24012 34522 24068 34524
rect 24012 34470 24014 34522
rect 24014 34470 24066 34522
rect 24066 34470 24068 34522
rect 24012 34468 24068 34470
rect 23804 32954 23860 32956
rect 23804 32902 23806 32954
rect 23806 32902 23858 32954
rect 23858 32902 23860 32954
rect 23804 32900 23860 32902
rect 23908 32954 23964 32956
rect 23908 32902 23910 32954
rect 23910 32902 23962 32954
rect 23962 32902 23964 32954
rect 23908 32900 23964 32902
rect 24012 32954 24068 32956
rect 24012 32902 24014 32954
rect 24014 32902 24066 32954
rect 24066 32902 24068 32954
rect 24012 32900 24068 32902
rect 24464 36874 24520 36876
rect 24464 36822 24466 36874
rect 24466 36822 24518 36874
rect 24518 36822 24520 36874
rect 24464 36820 24520 36822
rect 24568 36874 24624 36876
rect 24568 36822 24570 36874
rect 24570 36822 24622 36874
rect 24622 36822 24624 36874
rect 24568 36820 24624 36822
rect 24672 36874 24728 36876
rect 24672 36822 24674 36874
rect 24674 36822 24726 36874
rect 24726 36822 24728 36874
rect 24672 36820 24728 36822
rect 24464 35306 24520 35308
rect 24464 35254 24466 35306
rect 24466 35254 24518 35306
rect 24518 35254 24520 35306
rect 24464 35252 24520 35254
rect 24568 35306 24624 35308
rect 24568 35254 24570 35306
rect 24570 35254 24622 35306
rect 24622 35254 24624 35306
rect 24568 35252 24624 35254
rect 24672 35306 24728 35308
rect 24672 35254 24674 35306
rect 24674 35254 24726 35306
rect 24726 35254 24728 35306
rect 24672 35252 24728 35254
rect 24668 34300 24724 34356
rect 24892 34748 24948 34804
rect 24668 33852 24724 33908
rect 24464 33738 24520 33740
rect 24464 33686 24466 33738
rect 24466 33686 24518 33738
rect 24518 33686 24520 33738
rect 24464 33684 24520 33686
rect 24568 33738 24624 33740
rect 24568 33686 24570 33738
rect 24570 33686 24622 33738
rect 24622 33686 24624 33738
rect 24568 33684 24624 33686
rect 24672 33738 24728 33740
rect 24672 33686 24674 33738
rect 24674 33686 24726 33738
rect 24726 33686 24728 33738
rect 24672 33684 24728 33686
rect 24668 32284 24724 32340
rect 24464 32170 24520 32172
rect 24464 32118 24466 32170
rect 24466 32118 24518 32170
rect 24518 32118 24520 32170
rect 24464 32116 24520 32118
rect 24568 32170 24624 32172
rect 24568 32118 24570 32170
rect 24570 32118 24622 32170
rect 24622 32118 24624 32170
rect 24568 32116 24624 32118
rect 24672 32170 24728 32172
rect 24672 32118 24674 32170
rect 24674 32118 24726 32170
rect 24726 32118 24728 32170
rect 24672 32116 24728 32118
rect 24332 31948 24388 32004
rect 23804 31386 23860 31388
rect 23804 31334 23806 31386
rect 23806 31334 23858 31386
rect 23858 31334 23860 31386
rect 23804 31332 23860 31334
rect 23908 31386 23964 31388
rect 23908 31334 23910 31386
rect 23910 31334 23962 31386
rect 23962 31334 23964 31386
rect 23908 31332 23964 31334
rect 24012 31386 24068 31388
rect 24012 31334 24014 31386
rect 24014 31334 24066 31386
rect 24066 31334 24068 31386
rect 24012 31332 24068 31334
rect 23660 30716 23716 30772
rect 23804 29818 23860 29820
rect 23804 29766 23806 29818
rect 23806 29766 23858 29818
rect 23858 29766 23860 29818
rect 23804 29764 23860 29766
rect 23908 29818 23964 29820
rect 23908 29766 23910 29818
rect 23910 29766 23962 29818
rect 23962 29766 23964 29818
rect 23908 29764 23964 29766
rect 24012 29818 24068 29820
rect 24012 29766 24014 29818
rect 24014 29766 24066 29818
rect 24066 29766 24068 29818
rect 24012 29764 24068 29766
rect 23804 28250 23860 28252
rect 23804 28198 23806 28250
rect 23806 28198 23858 28250
rect 23858 28198 23860 28250
rect 23804 28196 23860 28198
rect 23908 28250 23964 28252
rect 23908 28198 23910 28250
rect 23910 28198 23962 28250
rect 23962 28198 23964 28250
rect 23908 28196 23964 28198
rect 24012 28250 24068 28252
rect 24012 28198 24014 28250
rect 24014 28198 24066 28250
rect 24066 28198 24068 28250
rect 24012 28196 24068 28198
rect 23804 26682 23860 26684
rect 23804 26630 23806 26682
rect 23806 26630 23858 26682
rect 23858 26630 23860 26682
rect 23804 26628 23860 26630
rect 23908 26682 23964 26684
rect 23908 26630 23910 26682
rect 23910 26630 23962 26682
rect 23962 26630 23964 26682
rect 23908 26628 23964 26630
rect 24012 26682 24068 26684
rect 24012 26630 24014 26682
rect 24014 26630 24066 26682
rect 24066 26630 24068 26682
rect 24012 26628 24068 26630
rect 23548 25228 23604 25284
rect 23804 25114 23860 25116
rect 23804 25062 23806 25114
rect 23806 25062 23858 25114
rect 23858 25062 23860 25114
rect 23804 25060 23860 25062
rect 23908 25114 23964 25116
rect 23908 25062 23910 25114
rect 23910 25062 23962 25114
rect 23962 25062 23964 25114
rect 23908 25060 23964 25062
rect 24012 25114 24068 25116
rect 24012 25062 24014 25114
rect 24014 25062 24066 25114
rect 24066 25062 24068 25114
rect 24012 25060 24068 25062
rect 23804 23546 23860 23548
rect 23804 23494 23806 23546
rect 23806 23494 23858 23546
rect 23858 23494 23860 23546
rect 23804 23492 23860 23494
rect 23908 23546 23964 23548
rect 23908 23494 23910 23546
rect 23910 23494 23962 23546
rect 23962 23494 23964 23546
rect 23908 23492 23964 23494
rect 24012 23546 24068 23548
rect 24012 23494 24014 23546
rect 24014 23494 24066 23546
rect 24066 23494 24068 23546
rect 24012 23492 24068 23494
rect 24892 30716 24948 30772
rect 24464 30602 24520 30604
rect 24464 30550 24466 30602
rect 24466 30550 24518 30602
rect 24518 30550 24520 30602
rect 24464 30548 24520 30550
rect 24568 30602 24624 30604
rect 24568 30550 24570 30602
rect 24570 30550 24622 30602
rect 24622 30550 24624 30602
rect 24568 30548 24624 30550
rect 24672 30602 24728 30604
rect 24672 30550 24674 30602
rect 24674 30550 24726 30602
rect 24726 30550 24728 30602
rect 24672 30548 24728 30550
rect 24464 29034 24520 29036
rect 24464 28982 24466 29034
rect 24466 28982 24518 29034
rect 24518 28982 24520 29034
rect 24464 28980 24520 28982
rect 24568 29034 24624 29036
rect 24568 28982 24570 29034
rect 24570 28982 24622 29034
rect 24622 28982 24624 29034
rect 24568 28980 24624 28982
rect 24672 29034 24728 29036
rect 24672 28982 24674 29034
rect 24674 28982 24726 29034
rect 24726 28982 24728 29034
rect 24672 28980 24728 28982
rect 24332 27804 24388 27860
rect 24668 27746 24724 27748
rect 24668 27694 24670 27746
rect 24670 27694 24722 27746
rect 24722 27694 24724 27746
rect 24668 27692 24724 27694
rect 24464 27466 24520 27468
rect 24464 27414 24466 27466
rect 24466 27414 24518 27466
rect 24518 27414 24520 27466
rect 24464 27412 24520 27414
rect 24568 27466 24624 27468
rect 24568 27414 24570 27466
rect 24570 27414 24622 27466
rect 24622 27414 24624 27466
rect 24568 27412 24624 27414
rect 24672 27466 24728 27468
rect 24672 27414 24674 27466
rect 24674 27414 24726 27466
rect 24726 27414 24728 27466
rect 24672 27412 24728 27414
rect 24668 27244 24724 27300
rect 24464 25898 24520 25900
rect 24464 25846 24466 25898
rect 24466 25846 24518 25898
rect 24518 25846 24520 25898
rect 24464 25844 24520 25846
rect 24568 25898 24624 25900
rect 24568 25846 24570 25898
rect 24570 25846 24622 25898
rect 24622 25846 24624 25898
rect 24568 25844 24624 25846
rect 24672 25898 24728 25900
rect 24672 25846 24674 25898
rect 24674 25846 24726 25898
rect 24726 25846 24728 25898
rect 24672 25844 24728 25846
rect 25004 29484 25060 29540
rect 25564 37996 25620 38052
rect 25452 36988 25508 37044
rect 25452 30716 25508 30772
rect 25116 29148 25172 29204
rect 25676 37938 25732 37940
rect 25676 37886 25678 37938
rect 25678 37886 25730 37938
rect 25730 37886 25732 37938
rect 25676 37884 25732 37886
rect 25676 36092 25732 36148
rect 25900 35532 25956 35588
rect 25676 34802 25732 34804
rect 25676 34750 25678 34802
rect 25678 34750 25730 34802
rect 25730 34750 25732 34802
rect 25676 34748 25732 34750
rect 25676 33852 25732 33908
rect 25676 32956 25732 33012
rect 25676 31666 25732 31668
rect 25676 31614 25678 31666
rect 25678 31614 25730 31666
rect 25730 31614 25732 31666
rect 25676 31612 25732 31614
rect 25900 30940 25956 30996
rect 25564 28700 25620 28756
rect 25676 30828 25732 30884
rect 25788 30380 25844 30436
rect 25788 28700 25844 28756
rect 25900 30156 25956 30212
rect 25676 28364 25732 28420
rect 25676 27132 25732 27188
rect 25676 26236 25732 26292
rect 25564 25452 25620 25508
rect 24464 24330 24520 24332
rect 24464 24278 24466 24330
rect 24466 24278 24518 24330
rect 24518 24278 24520 24330
rect 24464 24276 24520 24278
rect 24568 24330 24624 24332
rect 24568 24278 24570 24330
rect 24570 24278 24622 24330
rect 24622 24278 24624 24330
rect 24568 24276 24624 24278
rect 24672 24330 24728 24332
rect 24672 24278 24674 24330
rect 24674 24278 24726 24330
rect 24726 24278 24728 24330
rect 24672 24276 24728 24278
rect 24668 24050 24724 24052
rect 24668 23998 24670 24050
rect 24670 23998 24722 24050
rect 24722 23998 24724 24050
rect 24668 23996 24724 23998
rect 25452 23996 25508 24052
rect 24220 23212 24276 23268
rect 24464 22762 24520 22764
rect 24464 22710 24466 22762
rect 24466 22710 24518 22762
rect 24518 22710 24520 22762
rect 24464 22708 24520 22710
rect 24568 22762 24624 22764
rect 24568 22710 24570 22762
rect 24570 22710 24622 22762
rect 24622 22710 24624 22762
rect 24568 22708 24624 22710
rect 24672 22762 24728 22764
rect 24672 22710 24674 22762
rect 24674 22710 24726 22762
rect 24726 22710 24728 22762
rect 24672 22708 24728 22710
rect 23804 21978 23860 21980
rect 23804 21926 23806 21978
rect 23806 21926 23858 21978
rect 23858 21926 23860 21978
rect 23804 21924 23860 21926
rect 23908 21978 23964 21980
rect 23908 21926 23910 21978
rect 23910 21926 23962 21978
rect 23962 21926 23964 21978
rect 23908 21924 23964 21926
rect 24012 21978 24068 21980
rect 24012 21926 24014 21978
rect 24014 21926 24066 21978
rect 24066 21926 24068 21978
rect 24012 21924 24068 21926
rect 24464 21194 24520 21196
rect 24464 21142 24466 21194
rect 24466 21142 24518 21194
rect 24518 21142 24520 21194
rect 24464 21140 24520 21142
rect 24568 21194 24624 21196
rect 24568 21142 24570 21194
rect 24570 21142 24622 21194
rect 24622 21142 24624 21194
rect 24568 21140 24624 21142
rect 24672 21194 24728 21196
rect 24672 21142 24674 21194
rect 24674 21142 24726 21194
rect 24726 21142 24728 21194
rect 24672 21140 24728 21142
rect 23804 20410 23860 20412
rect 23804 20358 23806 20410
rect 23806 20358 23858 20410
rect 23858 20358 23860 20410
rect 23804 20356 23860 20358
rect 23908 20410 23964 20412
rect 23908 20358 23910 20410
rect 23910 20358 23962 20410
rect 23962 20358 23964 20410
rect 23908 20356 23964 20358
rect 24012 20410 24068 20412
rect 24012 20358 24014 20410
rect 24014 20358 24066 20410
rect 24066 20358 24068 20410
rect 24012 20356 24068 20358
rect 24464 19626 24520 19628
rect 24464 19574 24466 19626
rect 24466 19574 24518 19626
rect 24518 19574 24520 19626
rect 24464 19572 24520 19574
rect 24568 19626 24624 19628
rect 24568 19574 24570 19626
rect 24570 19574 24622 19626
rect 24622 19574 24624 19626
rect 24568 19572 24624 19574
rect 24672 19626 24728 19628
rect 24672 19574 24674 19626
rect 24674 19574 24726 19626
rect 24726 19574 24728 19626
rect 24672 19572 24728 19574
rect 23804 18842 23860 18844
rect 23804 18790 23806 18842
rect 23806 18790 23858 18842
rect 23858 18790 23860 18842
rect 23804 18788 23860 18790
rect 23908 18842 23964 18844
rect 23908 18790 23910 18842
rect 23910 18790 23962 18842
rect 23962 18790 23964 18842
rect 23908 18788 23964 18790
rect 24012 18842 24068 18844
rect 24012 18790 24014 18842
rect 24014 18790 24066 18842
rect 24066 18790 24068 18842
rect 24012 18788 24068 18790
rect 24464 18058 24520 18060
rect 24464 18006 24466 18058
rect 24466 18006 24518 18058
rect 24518 18006 24520 18058
rect 24464 18004 24520 18006
rect 24568 18058 24624 18060
rect 24568 18006 24570 18058
rect 24570 18006 24622 18058
rect 24622 18006 24624 18058
rect 24568 18004 24624 18006
rect 24672 18058 24728 18060
rect 24672 18006 24674 18058
rect 24674 18006 24726 18058
rect 24726 18006 24728 18058
rect 24672 18004 24728 18006
rect 23804 17274 23860 17276
rect 23804 17222 23806 17274
rect 23806 17222 23858 17274
rect 23858 17222 23860 17274
rect 23804 17220 23860 17222
rect 23908 17274 23964 17276
rect 23908 17222 23910 17274
rect 23910 17222 23962 17274
rect 23962 17222 23964 17274
rect 23908 17220 23964 17222
rect 24012 17274 24068 17276
rect 24012 17222 24014 17274
rect 24014 17222 24066 17274
rect 24066 17222 24068 17274
rect 24012 17220 24068 17222
rect 24464 16490 24520 16492
rect 24464 16438 24466 16490
rect 24466 16438 24518 16490
rect 24518 16438 24520 16490
rect 24464 16436 24520 16438
rect 24568 16490 24624 16492
rect 24568 16438 24570 16490
rect 24570 16438 24622 16490
rect 24622 16438 24624 16490
rect 24568 16436 24624 16438
rect 24672 16490 24728 16492
rect 24672 16438 24674 16490
rect 24674 16438 24726 16490
rect 24726 16438 24728 16490
rect 24672 16436 24728 16438
rect 23804 15706 23860 15708
rect 23804 15654 23806 15706
rect 23806 15654 23858 15706
rect 23858 15654 23860 15706
rect 23804 15652 23860 15654
rect 23908 15706 23964 15708
rect 23908 15654 23910 15706
rect 23910 15654 23962 15706
rect 23962 15654 23964 15706
rect 23908 15652 23964 15654
rect 24012 15706 24068 15708
rect 24012 15654 24014 15706
rect 24014 15654 24066 15706
rect 24066 15654 24068 15706
rect 24012 15652 24068 15654
rect 24464 14922 24520 14924
rect 24464 14870 24466 14922
rect 24466 14870 24518 14922
rect 24518 14870 24520 14922
rect 24464 14868 24520 14870
rect 24568 14922 24624 14924
rect 24568 14870 24570 14922
rect 24570 14870 24622 14922
rect 24622 14870 24624 14922
rect 24568 14868 24624 14870
rect 24672 14922 24728 14924
rect 24672 14870 24674 14922
rect 24674 14870 24726 14922
rect 24726 14870 24728 14922
rect 24672 14868 24728 14870
rect 24892 14700 24948 14756
rect 25004 22204 25060 22260
rect 23804 14138 23860 14140
rect 23804 14086 23806 14138
rect 23806 14086 23858 14138
rect 23858 14086 23860 14138
rect 23804 14084 23860 14086
rect 23908 14138 23964 14140
rect 23908 14086 23910 14138
rect 23910 14086 23962 14138
rect 23962 14086 23964 14138
rect 23908 14084 23964 14086
rect 24012 14138 24068 14140
rect 24012 14086 24014 14138
rect 24014 14086 24066 14138
rect 24066 14086 24068 14138
rect 24012 14084 24068 14086
rect 24464 13354 24520 13356
rect 24464 13302 24466 13354
rect 24466 13302 24518 13354
rect 24518 13302 24520 13354
rect 24464 13300 24520 13302
rect 24568 13354 24624 13356
rect 24568 13302 24570 13354
rect 24570 13302 24622 13354
rect 24622 13302 24624 13354
rect 24568 13300 24624 13302
rect 24672 13354 24728 13356
rect 24672 13302 24674 13354
rect 24674 13302 24726 13354
rect 24726 13302 24728 13354
rect 24672 13300 24728 13302
rect 23804 12570 23860 12572
rect 23804 12518 23806 12570
rect 23806 12518 23858 12570
rect 23858 12518 23860 12570
rect 23804 12516 23860 12518
rect 23908 12570 23964 12572
rect 23908 12518 23910 12570
rect 23910 12518 23962 12570
rect 23962 12518 23964 12570
rect 23908 12516 23964 12518
rect 24012 12570 24068 12572
rect 24012 12518 24014 12570
rect 24014 12518 24066 12570
rect 24066 12518 24068 12570
rect 24012 12516 24068 12518
rect 24464 11786 24520 11788
rect 24464 11734 24466 11786
rect 24466 11734 24518 11786
rect 24518 11734 24520 11786
rect 24464 11732 24520 11734
rect 24568 11786 24624 11788
rect 24568 11734 24570 11786
rect 24570 11734 24622 11786
rect 24622 11734 24624 11786
rect 24568 11732 24624 11734
rect 24672 11786 24728 11788
rect 24672 11734 24674 11786
rect 24674 11734 24726 11786
rect 24726 11734 24728 11786
rect 24672 11732 24728 11734
rect 23436 11228 23492 11284
rect 23804 11002 23860 11004
rect 23804 10950 23806 11002
rect 23806 10950 23858 11002
rect 23858 10950 23860 11002
rect 23804 10948 23860 10950
rect 23908 11002 23964 11004
rect 23908 10950 23910 11002
rect 23910 10950 23962 11002
rect 23962 10950 23964 11002
rect 23908 10948 23964 10950
rect 24012 11002 24068 11004
rect 24012 10950 24014 11002
rect 24014 10950 24066 11002
rect 24066 10950 24068 11002
rect 24012 10948 24068 10950
rect 25676 24892 25732 24948
rect 25676 23100 25732 23156
rect 25676 21756 25732 21812
rect 25564 13020 25620 13076
rect 26236 44994 26292 44996
rect 26236 44942 26238 44994
rect 26238 44942 26290 44994
rect 26290 44942 26292 44994
rect 26236 44940 26292 44942
rect 26236 44322 26292 44324
rect 26236 44270 26238 44322
rect 26238 44270 26290 44322
rect 26290 44270 26292 44322
rect 26236 44268 26292 44270
rect 26236 43426 26292 43428
rect 26236 43374 26238 43426
rect 26238 43374 26290 43426
rect 26290 43374 26292 43426
rect 26236 43372 26292 43374
rect 26572 44828 26628 44884
rect 27244 54012 27300 54068
rect 27020 53116 27076 53172
rect 26012 19740 26068 19796
rect 26908 52892 26964 52948
rect 25900 12908 25956 12964
rect 26012 16716 26068 16772
rect 25004 10556 25060 10612
rect 24464 10218 24520 10220
rect 24464 10166 24466 10218
rect 24466 10166 24518 10218
rect 24518 10166 24520 10218
rect 24464 10164 24520 10166
rect 24568 10218 24624 10220
rect 24568 10166 24570 10218
rect 24570 10166 24622 10218
rect 24622 10166 24624 10218
rect 24568 10164 24624 10166
rect 24672 10218 24728 10220
rect 24672 10166 24674 10218
rect 24674 10166 24726 10218
rect 24726 10166 24728 10218
rect 24672 10164 24728 10166
rect 23804 9434 23860 9436
rect 23804 9382 23806 9434
rect 23806 9382 23858 9434
rect 23858 9382 23860 9434
rect 23804 9380 23860 9382
rect 23908 9434 23964 9436
rect 23908 9382 23910 9434
rect 23910 9382 23962 9434
rect 23962 9382 23964 9434
rect 23908 9380 23964 9382
rect 24012 9434 24068 9436
rect 24012 9382 24014 9434
rect 24014 9382 24066 9434
rect 24066 9382 24068 9434
rect 24012 9380 24068 9382
rect 24464 8650 24520 8652
rect 24464 8598 24466 8650
rect 24466 8598 24518 8650
rect 24518 8598 24520 8650
rect 24464 8596 24520 8598
rect 24568 8650 24624 8652
rect 24568 8598 24570 8650
rect 24570 8598 24622 8650
rect 24622 8598 24624 8650
rect 24568 8596 24624 8598
rect 24672 8650 24728 8652
rect 24672 8598 24674 8650
rect 24674 8598 24726 8650
rect 24726 8598 24728 8650
rect 24672 8596 24728 8598
rect 23804 7866 23860 7868
rect 23804 7814 23806 7866
rect 23806 7814 23858 7866
rect 23858 7814 23860 7866
rect 23804 7812 23860 7814
rect 23908 7866 23964 7868
rect 23908 7814 23910 7866
rect 23910 7814 23962 7866
rect 23962 7814 23964 7866
rect 23908 7812 23964 7814
rect 24012 7866 24068 7868
rect 24012 7814 24014 7866
rect 24014 7814 24066 7866
rect 24066 7814 24068 7866
rect 24012 7812 24068 7814
rect 24464 7082 24520 7084
rect 24464 7030 24466 7082
rect 24466 7030 24518 7082
rect 24518 7030 24520 7082
rect 24464 7028 24520 7030
rect 24568 7082 24624 7084
rect 24568 7030 24570 7082
rect 24570 7030 24622 7082
rect 24622 7030 24624 7082
rect 24568 7028 24624 7030
rect 24672 7082 24728 7084
rect 24672 7030 24674 7082
rect 24674 7030 24726 7082
rect 24726 7030 24728 7082
rect 24672 7028 24728 7030
rect 23804 6298 23860 6300
rect 23804 6246 23806 6298
rect 23806 6246 23858 6298
rect 23858 6246 23860 6298
rect 23804 6244 23860 6246
rect 23908 6298 23964 6300
rect 23908 6246 23910 6298
rect 23910 6246 23962 6298
rect 23962 6246 23964 6298
rect 23908 6244 23964 6246
rect 24012 6298 24068 6300
rect 24012 6246 24014 6298
rect 24014 6246 24066 6298
rect 24066 6246 24068 6298
rect 24012 6244 24068 6246
rect 24464 5514 24520 5516
rect 24464 5462 24466 5514
rect 24466 5462 24518 5514
rect 24518 5462 24520 5514
rect 24464 5460 24520 5462
rect 24568 5514 24624 5516
rect 24568 5462 24570 5514
rect 24570 5462 24622 5514
rect 24622 5462 24624 5514
rect 24568 5460 24624 5462
rect 24672 5514 24728 5516
rect 24672 5462 24674 5514
rect 24674 5462 24726 5514
rect 24726 5462 24728 5514
rect 24672 5460 24728 5462
rect 23804 4730 23860 4732
rect 23804 4678 23806 4730
rect 23806 4678 23858 4730
rect 23858 4678 23860 4730
rect 23804 4676 23860 4678
rect 23908 4730 23964 4732
rect 23908 4678 23910 4730
rect 23910 4678 23962 4730
rect 23962 4678 23964 4730
rect 23908 4676 23964 4678
rect 24012 4730 24068 4732
rect 24012 4678 24014 4730
rect 24014 4678 24066 4730
rect 24066 4678 24068 4730
rect 24012 4676 24068 4678
rect 24464 3946 24520 3948
rect 24464 3894 24466 3946
rect 24466 3894 24518 3946
rect 24518 3894 24520 3946
rect 24464 3892 24520 3894
rect 24568 3946 24624 3948
rect 24568 3894 24570 3946
rect 24570 3894 24622 3946
rect 24622 3894 24624 3946
rect 24568 3892 24624 3894
rect 24672 3946 24728 3948
rect 24672 3894 24674 3946
rect 24674 3894 24726 3946
rect 24726 3894 24728 3946
rect 24672 3892 24728 3894
rect 22988 3388 23044 3444
rect 23804 3162 23860 3164
rect 23804 3110 23806 3162
rect 23806 3110 23858 3162
rect 23858 3110 23860 3162
rect 23804 3108 23860 3110
rect 23908 3162 23964 3164
rect 23908 3110 23910 3162
rect 23910 3110 23962 3162
rect 23962 3110 23964 3162
rect 23908 3108 23964 3110
rect 24012 3162 24068 3164
rect 24012 3110 24014 3162
rect 24014 3110 24066 3162
rect 24066 3110 24068 3162
rect 24012 3108 24068 3110
rect 24464 2378 24520 2380
rect 24464 2326 24466 2378
rect 24466 2326 24518 2378
rect 24518 2326 24520 2378
rect 24464 2324 24520 2326
rect 24568 2378 24624 2380
rect 24568 2326 24570 2378
rect 24570 2326 24622 2378
rect 24622 2326 24624 2378
rect 24568 2324 24624 2326
rect 24672 2378 24728 2380
rect 24672 2326 24674 2378
rect 24674 2326 24726 2378
rect 24726 2326 24728 2378
rect 24672 2324 24728 2326
rect 23804 1594 23860 1596
rect 23804 1542 23806 1594
rect 23806 1542 23858 1594
rect 23858 1542 23860 1594
rect 23804 1540 23860 1542
rect 23908 1594 23964 1596
rect 23908 1542 23910 1594
rect 23910 1542 23962 1594
rect 23962 1542 23964 1594
rect 23908 1540 23964 1542
rect 24012 1594 24068 1596
rect 24012 1542 24014 1594
rect 24014 1542 24066 1594
rect 24066 1542 24068 1594
rect 24012 1540 24068 1542
rect 24892 1596 24948 1652
rect 22876 252 22932 308
rect 23548 1260 23604 1316
rect 24464 810 24520 812
rect 24464 758 24466 810
rect 24466 758 24518 810
rect 24518 758 24520 810
rect 24464 756 24520 758
rect 24568 810 24624 812
rect 24568 758 24570 810
rect 24570 758 24622 810
rect 24622 758 24624 810
rect 24568 756 24624 758
rect 24672 810 24728 812
rect 24672 758 24674 810
rect 24674 758 24726 810
rect 24726 758 24728 810
rect 24672 756 24728 758
rect 26236 42754 26292 42756
rect 26236 42702 26238 42754
rect 26238 42702 26290 42754
rect 26290 42702 26292 42754
rect 26236 42700 26292 42702
rect 26460 42588 26516 42644
rect 26236 41858 26292 41860
rect 26236 41806 26238 41858
rect 26238 41806 26290 41858
rect 26290 41806 26292 41858
rect 26236 41804 26292 41806
rect 26236 41186 26292 41188
rect 26236 41134 26238 41186
rect 26238 41134 26290 41186
rect 26290 41134 26292 41186
rect 26236 41132 26292 41134
rect 26236 40460 26292 40516
rect 26236 39004 26292 39060
rect 26236 38834 26292 38836
rect 26236 38782 26238 38834
rect 26238 38782 26290 38834
rect 26290 38782 26292 38834
rect 26236 38780 26292 38782
rect 26348 38220 26404 38276
rect 26236 38050 26292 38052
rect 26236 37998 26238 38050
rect 26238 37998 26290 38050
rect 26290 37998 26292 38050
rect 26236 37996 26292 37998
rect 26236 37436 26292 37492
rect 26348 35868 26404 35924
rect 26236 35586 26292 35588
rect 26236 35534 26238 35586
rect 26238 35534 26290 35586
rect 26290 35534 26292 35586
rect 26236 35532 26292 35534
rect 26236 34914 26292 34916
rect 26236 34862 26238 34914
rect 26238 34862 26290 34914
rect 26290 34862 26292 34914
rect 26236 34860 26292 34862
rect 26236 34018 26292 34020
rect 26236 33966 26238 34018
rect 26238 33966 26290 34018
rect 26290 33966 26292 34018
rect 26236 33964 26292 33966
rect 26348 32396 26404 32452
rect 26236 30882 26292 30884
rect 26236 30830 26238 30882
rect 26238 30830 26290 30882
rect 26290 30830 26292 30882
rect 26236 30828 26292 30830
rect 26236 30210 26292 30212
rect 26236 30158 26238 30210
rect 26238 30158 26290 30210
rect 26290 30158 26292 30210
rect 26236 30156 26292 30158
rect 26236 29314 26292 29316
rect 26236 29262 26238 29314
rect 26238 29262 26290 29314
rect 26290 29262 26292 29314
rect 26236 29260 26292 29262
rect 26236 28754 26292 28756
rect 26236 28702 26238 28754
rect 26238 28702 26290 28754
rect 26290 28702 26292 28754
rect 26236 28700 26292 28702
rect 26348 28028 26404 28084
rect 26236 26908 26292 26964
rect 26348 26348 26404 26404
rect 26236 26178 26292 26180
rect 26236 26126 26238 26178
rect 26238 26126 26290 26178
rect 26290 26126 26292 26178
rect 26236 26124 26292 26126
rect 26236 25506 26292 25508
rect 26236 25454 26238 25506
rect 26238 25454 26290 25506
rect 26290 25454 26292 25506
rect 26236 25452 26292 25454
rect 26348 24780 26404 24836
rect 26236 24722 26292 24724
rect 26236 24670 26238 24722
rect 26238 24670 26290 24722
rect 26290 24670 26292 24722
rect 26236 24668 26292 24670
rect 26236 23938 26292 23940
rect 26236 23886 26238 23938
rect 26238 23886 26290 23938
rect 26290 23886 26292 23938
rect 26236 23884 26292 23886
rect 26236 21474 26292 21476
rect 26236 21422 26238 21474
rect 26238 21422 26290 21474
rect 26290 21422 26292 21474
rect 26236 21420 26292 21422
rect 26684 44380 26740 44436
rect 27244 52220 27300 52276
rect 27132 51324 27188 51380
rect 27244 50876 27300 50932
rect 27020 49980 27076 50036
rect 27244 49084 27300 49140
rect 27468 49196 27524 49252
rect 27132 48188 27188 48244
rect 27244 47740 27300 47796
rect 27356 47964 27412 48020
rect 27020 46844 27076 46900
rect 27244 45948 27300 46004
rect 27132 45052 27188 45108
rect 27244 44604 27300 44660
rect 27020 43820 27076 43876
rect 26908 41916 26964 41972
rect 26908 40572 26964 40628
rect 26908 39116 26964 39172
rect 26908 37436 26964 37492
rect 26908 35980 26964 36036
rect 26908 34300 26964 34356
rect 26908 32844 26964 32900
rect 26908 31836 26964 31892
rect 26684 31052 26740 31108
rect 26908 30268 26964 30324
rect 26908 29372 26964 29428
rect 26684 18396 26740 18452
rect 26572 12684 26628 12740
rect 26348 12236 26404 12292
rect 26124 8092 26180 8148
rect 26236 11228 26292 11284
rect 26012 1484 26068 1540
rect 27020 4508 27076 4564
rect 27244 42812 27300 42868
rect 27244 41468 27300 41524
rect 27244 39676 27300 39732
rect 27244 38332 27300 38388
rect 27356 39340 27412 39396
rect 27244 36540 27300 36596
rect 27244 35196 27300 35252
rect 27244 33404 27300 33460
rect 27244 32284 27300 32340
rect 28140 35084 28196 35140
rect 28028 31836 28084 31892
rect 27804 31500 27860 31556
rect 27244 31276 27300 31332
rect 27468 31164 27524 31220
rect 27244 29820 27300 29876
rect 27244 28924 27300 28980
rect 27244 28530 27300 28532
rect 27244 28478 27246 28530
rect 27246 28478 27298 28530
rect 27298 28478 27300 28530
rect 27244 28476 27300 28478
rect 27244 28082 27300 28084
rect 27244 28030 27246 28082
rect 27246 28030 27298 28082
rect 27298 28030 27300 28082
rect 27244 28028 27300 28030
rect 27244 27580 27300 27636
rect 27244 26684 27300 26740
rect 27244 25788 27300 25844
rect 27356 25340 27412 25396
rect 27244 24444 27300 24500
rect 27356 23548 27412 23604
rect 27244 22652 27300 22708
rect 27356 22204 27412 22260
rect 27468 21644 27524 21700
rect 27356 21084 27412 21140
rect 27468 16828 27524 16884
rect 27692 21084 27748 21140
rect 28028 31164 28084 31220
rect 27804 20412 27860 20468
rect 27916 21532 27972 21588
rect 27916 15484 27972 15540
rect 27580 13916 27636 13972
rect 28252 24108 28308 24164
rect 28140 11900 28196 11956
rect 28252 16268 28308 16324
rect 28364 11452 28420 11508
rect 28364 8316 28420 8372
rect 27356 3276 27412 3332
rect 27132 1596 27188 1652
rect 27580 1484 27636 1540
<< metal3 >>
rect 4722 57260 4732 57316
rect 4788 57260 5516 57316
rect 5572 57260 5582 57316
rect 25442 57260 25452 57316
rect 25508 57260 26236 57316
rect 26292 57260 26302 57316
rect 28448 57204 28560 57232
rect 25106 57148 25116 57204
rect 25172 57148 28560 57204
rect 28448 57120 28560 57148
rect 28448 56756 28560 56784
rect 25330 56700 25340 56756
rect 25396 56700 28560 56756
rect 28448 56672 28560 56700
rect 3794 56420 3804 56476
rect 3860 56420 3908 56476
rect 3964 56420 4012 56476
rect 4068 56420 4078 56476
rect 23794 56420 23804 56476
rect 23860 56420 23908 56476
rect 23964 56420 24012 56476
rect 24068 56420 24078 56476
rect 28448 56308 28560 56336
rect 15474 56252 15484 56308
rect 15540 56252 16492 56308
rect 16548 56252 16558 56308
rect 19506 56252 19516 56308
rect 19572 56252 20636 56308
rect 20692 56252 20702 56308
rect 20850 56252 20860 56308
rect 20916 56252 21868 56308
rect 21924 56252 21934 56308
rect 23538 56252 23548 56308
rect 23604 56252 24444 56308
rect 24500 56252 24510 56308
rect 24882 56252 24892 56308
rect 24948 56252 26012 56308
rect 26068 56252 26078 56308
rect 26236 56252 28560 56308
rect 26236 56196 26292 56252
rect 28448 56224 28560 56252
rect 22530 56140 22540 56196
rect 22596 56140 26292 56196
rect 23538 56028 23548 56084
rect 23604 56028 27580 56084
rect 27636 56028 27646 56084
rect 1698 55916 1708 55972
rect 1764 55916 3052 55972
rect 3108 55916 3118 55972
rect 8082 55916 8092 55972
rect 8148 55916 21084 55972
rect 21140 55916 21150 55972
rect 21970 55916 21980 55972
rect 22036 55916 23884 55972
rect 23940 55916 23950 55972
rect 28448 55860 28560 55888
rect 21634 55804 21644 55860
rect 21700 55804 28560 55860
rect 28448 55776 28560 55804
rect 4454 55636 4464 55692
rect 4520 55636 4568 55692
rect 4624 55636 4672 55692
rect 4728 55636 4738 55692
rect 24454 55636 24464 55692
rect 24520 55636 24568 55692
rect 24624 55636 24672 55692
rect 24728 55636 24738 55692
rect 15586 55468 15596 55524
rect 15652 55468 23436 55524
rect 23492 55468 23502 55524
rect 28448 55412 28560 55440
rect 11554 55356 11564 55412
rect 11620 55356 11630 55412
rect 18834 55356 18844 55412
rect 18900 55356 20188 55412
rect 20244 55356 20254 55412
rect 24770 55356 24780 55412
rect 24836 55356 28560 55412
rect 11564 55300 11620 55356
rect 28448 55328 28560 55356
rect 11564 55244 20524 55300
rect 20580 55244 20590 55300
rect 23650 55244 23660 55300
rect 23716 55244 25004 55300
rect 25060 55244 25070 55300
rect 18050 55132 18060 55188
rect 18116 55132 24668 55188
rect 24724 55132 24734 55188
rect 12898 55020 12908 55076
rect 12964 55020 24332 55076
rect 24388 55020 24398 55076
rect 28448 54964 28560 54992
rect 24210 54908 24220 54964
rect 24276 54908 28560 54964
rect 3794 54852 3804 54908
rect 3860 54852 3908 54908
rect 3964 54852 4012 54908
rect 4068 54852 4078 54908
rect 23794 54852 23804 54908
rect 23860 54852 23908 54908
rect 23964 54852 24012 54908
rect 24068 54852 24078 54908
rect 28448 54880 28560 54908
rect 9986 54572 9996 54628
rect 10052 54572 19404 54628
rect 19460 54572 19470 54628
rect 28448 54516 28560 54544
rect 23650 54460 23660 54516
rect 23716 54460 24668 54516
rect 24724 54460 24734 54516
rect 25554 54460 25564 54516
rect 25620 54460 28560 54516
rect 28448 54432 28560 54460
rect 14690 54348 14700 54404
rect 14756 54348 26236 54404
rect 26292 54348 26302 54404
rect 8642 54236 8652 54292
rect 8708 54236 20636 54292
rect 20692 54236 20702 54292
rect 23772 54236 24780 54292
rect 24836 54236 24846 54292
rect 23772 54180 23828 54236
rect 23762 54124 23772 54180
rect 23828 54124 23838 54180
rect 4454 54068 4464 54124
rect 4520 54068 4568 54124
rect 4624 54068 4672 54124
rect 4728 54068 4738 54124
rect 24454 54068 24464 54124
rect 24520 54068 24568 54124
rect 24624 54068 24672 54124
rect 24728 54068 24738 54124
rect 28448 54068 28560 54096
rect 27234 54012 27244 54068
rect 27300 54012 28560 54068
rect 28448 53984 28560 54012
rect 14018 53900 14028 53956
rect 14084 53900 22316 53956
rect 22372 53900 22382 53956
rect 20514 53676 20524 53732
rect 20580 53676 21644 53732
rect 21700 53676 21710 53732
rect 24882 53676 24892 53732
rect 24948 53676 26796 53732
rect 26852 53676 26862 53732
rect 0 53620 112 53648
rect 28448 53620 28560 53648
rect 0 53564 364 53620
rect 420 53564 430 53620
rect 17490 53564 17500 53620
rect 17556 53564 21308 53620
rect 21364 53564 21374 53620
rect 25554 53564 25564 53620
rect 25620 53564 28560 53620
rect 0 53536 112 53564
rect 28448 53536 28560 53564
rect 14242 53452 14252 53508
rect 14308 53452 21868 53508
rect 21924 53452 21934 53508
rect 3794 53284 3804 53340
rect 3860 53284 3908 53340
rect 3964 53284 4012 53340
rect 4068 53284 4078 53340
rect 23794 53284 23804 53340
rect 23860 53284 23908 53340
rect 23964 53284 24012 53340
rect 24068 53284 24078 53340
rect 19506 53228 19516 53284
rect 19572 53228 22652 53284
rect 22708 53228 22718 53284
rect 28448 53172 28560 53200
rect 18274 53116 18284 53172
rect 18340 53116 21756 53172
rect 21812 53116 21822 53172
rect 24098 53116 24108 53172
rect 24164 53116 25116 53172
rect 25172 53116 25182 53172
rect 27010 53116 27020 53172
rect 27076 53116 28560 53172
rect 28448 53088 28560 53116
rect 6290 53004 6300 53060
rect 6356 53004 24668 53060
rect 24724 53004 24734 53060
rect 1362 52892 1372 52948
rect 1428 52892 15148 52948
rect 15204 52892 15214 52948
rect 21410 52892 21420 52948
rect 21476 52892 26908 52948
rect 26964 52892 26974 52948
rect 22194 52780 22204 52836
rect 22260 52780 26236 52836
rect 26292 52780 26302 52836
rect 28448 52724 28560 52752
rect 18498 52668 18508 52724
rect 18564 52668 22204 52724
rect 22260 52668 22270 52724
rect 25442 52668 25452 52724
rect 25508 52668 28560 52724
rect 28448 52640 28560 52668
rect 4454 52500 4464 52556
rect 4520 52500 4568 52556
rect 4624 52500 4672 52556
rect 4728 52500 4738 52556
rect 24454 52500 24464 52556
rect 24520 52500 24568 52556
rect 24624 52500 24672 52556
rect 24728 52500 24738 52556
rect 12674 52444 12684 52500
rect 12740 52444 22484 52500
rect 22428 52388 22484 52444
rect 10098 52332 10108 52388
rect 10164 52332 22204 52388
rect 22260 52332 22270 52388
rect 22428 52332 24668 52388
rect 24724 52332 24734 52388
rect 0 52276 112 52304
rect 28448 52276 28560 52304
rect 0 52220 1820 52276
rect 1876 52220 1886 52276
rect 19954 52220 19964 52276
rect 20020 52220 22764 52276
rect 22820 52220 22830 52276
rect 27234 52220 27244 52276
rect 27300 52220 28560 52276
rect 0 52192 112 52220
rect 28448 52192 28560 52220
rect 17602 52108 17612 52164
rect 17668 52108 26236 52164
rect 26292 52108 26302 52164
rect 5954 51884 5964 51940
rect 6020 51884 26348 51940
rect 26404 51884 26414 51940
rect 28448 51828 28560 51856
rect 25554 51772 25564 51828
rect 25620 51772 28560 51828
rect 3794 51716 3804 51772
rect 3860 51716 3908 51772
rect 3964 51716 4012 51772
rect 4068 51716 4078 51772
rect 23794 51716 23804 51772
rect 23860 51716 23908 51772
rect 23964 51716 24012 51772
rect 24068 51716 24078 51772
rect 28448 51744 28560 51772
rect 6626 51436 6636 51492
rect 6692 51436 22876 51492
rect 22932 51436 22942 51492
rect 28448 51380 28560 51408
rect 4162 51324 4172 51380
rect 4228 51324 23100 51380
rect 23156 51324 23166 51380
rect 27122 51324 27132 51380
rect 27188 51324 28560 51380
rect 28448 51296 28560 51324
rect 16706 51212 16716 51268
rect 16772 51212 24668 51268
rect 24724 51212 24734 51268
rect 21074 51100 21084 51156
rect 21140 51100 23772 51156
rect 23828 51100 23838 51156
rect 0 50932 112 50960
rect 4454 50932 4464 50988
rect 4520 50932 4568 50988
rect 4624 50932 4672 50988
rect 4728 50932 4738 50988
rect 24454 50932 24464 50988
rect 24520 50932 24568 50988
rect 24624 50932 24672 50988
rect 24728 50932 24738 50988
rect 28448 50932 28560 50960
rect 0 50876 1932 50932
rect 1988 50876 1998 50932
rect 27234 50876 27244 50932
rect 27300 50876 28560 50932
rect 0 50848 112 50876
rect 28448 50848 28560 50876
rect 10882 50764 10892 50820
rect 10948 50764 26236 50820
rect 26292 50764 26302 50820
rect 28448 50484 28560 50512
rect 15474 50428 15484 50484
rect 15540 50428 20860 50484
rect 20916 50428 20926 50484
rect 25554 50428 25564 50484
rect 25620 50428 28560 50484
rect 28448 50400 28560 50428
rect 3794 50148 3804 50204
rect 3860 50148 3908 50204
rect 3964 50148 4012 50204
rect 4068 50148 4078 50204
rect 23794 50148 23804 50204
rect 23860 50148 23908 50204
rect 23964 50148 24012 50204
rect 24068 50148 24078 50204
rect 28448 50036 28560 50064
rect 27010 49980 27020 50036
rect 27076 49980 28560 50036
rect 28448 49952 28560 49980
rect 22978 49868 22988 49924
rect 23044 49868 24220 49924
rect 24276 49868 24286 49924
rect 0 49588 112 49616
rect 28448 49588 28560 49616
rect 0 49532 5740 49588
rect 5796 49532 5806 49588
rect 7410 49532 7420 49588
rect 7476 49532 24668 49588
rect 24724 49532 24734 49588
rect 25666 49532 25676 49588
rect 25732 49532 28560 49588
rect 0 49504 112 49532
rect 28448 49504 28560 49532
rect 4454 49364 4464 49420
rect 4520 49364 4568 49420
rect 4624 49364 4672 49420
rect 4728 49364 4738 49420
rect 24454 49364 24464 49420
rect 24520 49364 24568 49420
rect 24624 49364 24672 49420
rect 24728 49364 24738 49420
rect 23762 49196 23772 49252
rect 23828 49196 27468 49252
rect 27524 49196 27534 49252
rect 28448 49140 28560 49168
rect 27234 49084 27244 49140
rect 27300 49084 28560 49140
rect 28448 49056 28560 49084
rect 7186 48972 7196 49028
rect 7252 48972 26236 49028
rect 26292 48972 26302 49028
rect 11778 48860 11788 48916
rect 11844 48860 24668 48916
rect 24724 48860 24734 48916
rect 9090 48748 9100 48804
rect 9156 48748 26348 48804
rect 26404 48748 26414 48804
rect 28448 48692 28560 48720
rect 25666 48636 25676 48692
rect 25732 48636 28560 48692
rect 3794 48580 3804 48636
rect 3860 48580 3908 48636
rect 3964 48580 4012 48636
rect 4068 48580 4078 48636
rect 23794 48580 23804 48636
rect 23860 48580 23908 48636
rect 23964 48580 24012 48636
rect 24068 48580 24078 48636
rect 28448 48608 28560 48636
rect 0 48244 112 48272
rect 28448 48244 28560 48272
rect 0 48188 6076 48244
rect 6132 48188 6142 48244
rect 14354 48188 14364 48244
rect 14420 48188 24892 48244
rect 24948 48188 24958 48244
rect 27122 48188 27132 48244
rect 27188 48188 28560 48244
rect 0 48160 112 48188
rect 28448 48160 28560 48188
rect 16370 48076 16380 48132
rect 16436 48076 26236 48132
rect 26292 48076 26302 48132
rect 25330 47964 25340 48020
rect 25396 47964 27356 48020
rect 27412 47964 27422 48020
rect 14914 47852 14924 47908
rect 14980 47852 17612 47908
rect 17668 47852 17678 47908
rect 4454 47796 4464 47852
rect 4520 47796 4568 47852
rect 4624 47796 4672 47852
rect 4728 47796 4738 47852
rect 24454 47796 24464 47852
rect 24520 47796 24568 47852
rect 24624 47796 24672 47852
rect 24728 47796 24738 47852
rect 28448 47796 28560 47824
rect 27234 47740 27244 47796
rect 27300 47740 28560 47796
rect 28448 47712 28560 47740
rect 28448 47348 28560 47376
rect 25666 47292 25676 47348
rect 25732 47292 28560 47348
rect 28448 47264 28560 47292
rect 18284 47180 24332 47236
rect 24388 47180 24398 47236
rect 3794 47012 3804 47068
rect 3860 47012 3908 47068
rect 3964 47012 4012 47068
rect 4068 47012 4078 47068
rect 0 46900 112 46928
rect 18284 46900 18340 47180
rect 23794 47012 23804 47068
rect 23860 47012 23908 47068
rect 23964 47012 24012 47068
rect 24068 47012 24078 47068
rect 28448 46900 28560 46928
rect 0 46844 3276 46900
rect 3332 46844 3342 46900
rect 18274 46844 18284 46900
rect 18340 46844 18350 46900
rect 27010 46844 27020 46900
rect 27076 46844 28560 46900
rect 0 46816 112 46844
rect 28448 46816 28560 46844
rect 28448 46452 28560 46480
rect 20066 46396 20076 46452
rect 20132 46396 24668 46452
rect 24724 46396 24734 46452
rect 25666 46396 25676 46452
rect 25732 46396 28560 46452
rect 28448 46368 28560 46396
rect 4454 46228 4464 46284
rect 4520 46228 4568 46284
rect 4624 46228 4672 46284
rect 4728 46228 4738 46284
rect 24454 46228 24464 46284
rect 24520 46228 24568 46284
rect 24624 46228 24672 46284
rect 24728 46228 24738 46284
rect 26086 46060 26124 46116
rect 26180 46060 26190 46116
rect 28448 46004 28560 46032
rect 27234 45948 27244 46004
rect 27300 45948 28560 46004
rect 28448 45920 28560 45948
rect 20962 45836 20972 45892
rect 21028 45836 24668 45892
rect 24724 45836 24734 45892
rect 3332 45612 17836 45668
rect 17892 45612 17902 45668
rect 0 45556 112 45584
rect 3332 45556 3388 45612
rect 28448 45556 28560 45584
rect 0 45500 3388 45556
rect 25666 45500 25676 45556
rect 25732 45500 28560 45556
rect 0 45472 112 45500
rect 3794 45444 3804 45500
rect 3860 45444 3908 45500
rect 3964 45444 4012 45500
rect 4068 45444 4078 45500
rect 23794 45444 23804 45500
rect 23860 45444 23908 45500
rect 23964 45444 24012 45500
rect 24068 45444 24078 45500
rect 28448 45472 28560 45500
rect 28448 45108 28560 45136
rect 27122 45052 27132 45108
rect 27188 45052 28560 45108
rect 28448 45024 28560 45052
rect 2258 44940 2268 44996
rect 2324 44940 26236 44996
rect 26292 44940 26302 44996
rect 26562 44828 26572 44884
rect 26628 44828 26740 44884
rect 4454 44660 4464 44716
rect 4520 44660 4568 44716
rect 4624 44660 4672 44716
rect 4728 44660 4738 44716
rect 24454 44660 24464 44716
rect 24520 44660 24568 44716
rect 24624 44660 24672 44716
rect 24728 44660 24738 44716
rect 12002 44492 12012 44548
rect 12068 44492 24892 44548
rect 24948 44492 24958 44548
rect 26684 44436 26740 44828
rect 28448 44660 28560 44688
rect 27234 44604 27244 44660
rect 27300 44604 28560 44660
rect 28448 44576 28560 44604
rect 20402 44380 20412 44436
rect 20468 44380 25900 44436
rect 25956 44380 25966 44436
rect 26674 44380 26684 44436
rect 26740 44380 26750 44436
rect 17042 44268 17052 44324
rect 17108 44268 26236 44324
rect 26292 44268 26302 44324
rect 0 44212 112 44240
rect 28448 44212 28560 44240
rect 0 44156 17948 44212
rect 18004 44156 18014 44212
rect 25666 44156 25676 44212
rect 25732 44156 28560 44212
rect 0 44128 112 44156
rect 28448 44128 28560 44156
rect 7970 44044 7980 44100
rect 8036 44044 24668 44100
rect 24724 44044 24734 44100
rect 3794 43876 3804 43932
rect 3860 43876 3908 43932
rect 3964 43876 4012 43932
rect 4068 43876 4078 43932
rect 23794 43876 23804 43932
rect 23860 43876 23908 43932
rect 23964 43876 24012 43932
rect 24068 43876 24078 43932
rect 27010 43820 27020 43876
rect 27076 43820 27086 43876
rect 27020 43764 27076 43820
rect 28448 43764 28560 43792
rect 27020 43708 28560 43764
rect 28448 43680 28560 43708
rect 3490 43596 3500 43652
rect 3556 43596 11340 43652
rect 11396 43596 11406 43652
rect 7746 43372 7756 43428
rect 7812 43372 26236 43428
rect 26292 43372 26302 43428
rect 28448 43316 28560 43344
rect 25666 43260 25676 43316
rect 25732 43260 28560 43316
rect 28448 43232 28560 43260
rect 4454 43092 4464 43148
rect 4520 43092 4568 43148
rect 4624 43092 4672 43148
rect 4728 43092 4738 43148
rect 24454 43092 24464 43148
rect 24520 43092 24568 43148
rect 24624 43092 24672 43148
rect 24728 43092 24738 43148
rect 1474 42924 1484 42980
rect 1540 42924 11788 42980
rect 11844 42924 11854 42980
rect 0 42868 112 42896
rect 28448 42868 28560 42896
rect 0 42812 13916 42868
rect 13972 42812 13982 42868
rect 27234 42812 27244 42868
rect 27300 42812 28560 42868
rect 0 42784 112 42812
rect 28448 42784 28560 42812
rect 9762 42700 9772 42756
rect 9828 42700 26236 42756
rect 26292 42700 26302 42756
rect 13122 42588 13132 42644
rect 13188 42588 24668 42644
rect 24724 42588 24734 42644
rect 26114 42588 26124 42644
rect 26180 42588 26460 42644
rect 26516 42588 26526 42644
rect 28448 42420 28560 42448
rect 25666 42364 25676 42420
rect 25732 42364 28560 42420
rect 3794 42308 3804 42364
rect 3860 42308 3908 42364
rect 3964 42308 4012 42364
rect 4068 42308 4078 42364
rect 23794 42308 23804 42364
rect 23860 42308 23908 42364
rect 23964 42308 24012 42364
rect 24068 42308 24078 42364
rect 28448 42336 28560 42364
rect 2034 42028 2044 42084
rect 2100 42028 10892 42084
rect 10948 42028 10958 42084
rect 28448 41972 28560 42000
rect 26898 41916 26908 41972
rect 26964 41916 28560 41972
rect 28448 41888 28560 41916
rect 12226 41804 12236 41860
rect 12292 41804 26236 41860
rect 26292 41804 26302 41860
rect 0 41524 112 41552
rect 4454 41524 4464 41580
rect 4520 41524 4568 41580
rect 4624 41524 4672 41580
rect 4728 41524 4738 41580
rect 24454 41524 24464 41580
rect 24520 41524 24568 41580
rect 24624 41524 24672 41580
rect 24728 41524 24738 41580
rect 28448 41524 28560 41552
rect 0 41468 3388 41524
rect 27234 41468 27244 41524
rect 27300 41468 28560 41524
rect 0 41440 112 41468
rect 3332 41412 3388 41468
rect 28448 41440 28560 41468
rect 3332 41356 4564 41412
rect 5282 41356 5292 41412
rect 5348 41356 6076 41412
rect 6132 41356 6142 41412
rect 4508 41300 4564 41356
rect 1698 41244 1708 41300
rect 1764 41244 4284 41300
rect 4340 41244 4350 41300
rect 4508 41244 12124 41300
rect 12180 41244 12190 41300
rect 3266 41132 3276 41188
rect 3332 41132 10556 41188
rect 10612 41132 10622 41188
rect 16034 41132 16044 41188
rect 16100 41132 26236 41188
rect 26292 41132 26302 41188
rect 28448 41076 28560 41104
rect 9538 41020 9548 41076
rect 9604 41020 10220 41076
rect 10276 41020 10286 41076
rect 25666 41020 25676 41076
rect 25732 41020 28560 41076
rect 28448 40992 28560 41020
rect 3794 40740 3804 40796
rect 3860 40740 3908 40796
rect 3964 40740 4012 40796
rect 4068 40740 4078 40796
rect 23794 40740 23804 40796
rect 23860 40740 23908 40796
rect 23964 40740 24012 40796
rect 24068 40740 24078 40796
rect 28448 40628 28560 40656
rect 1922 40572 1932 40628
rect 1988 40572 1998 40628
rect 2146 40572 2156 40628
rect 2212 40572 24892 40628
rect 24948 40572 24958 40628
rect 26898 40572 26908 40628
rect 26964 40572 28560 40628
rect 1932 40516 1988 40572
rect 28448 40544 28560 40572
rect 1932 40460 2212 40516
rect 7858 40460 7868 40516
rect 7924 40460 26236 40516
rect 26292 40460 26302 40516
rect 1698 40348 1708 40404
rect 1764 40348 1932 40404
rect 1988 40348 1998 40404
rect 2156 40292 2212 40460
rect 4274 40348 4284 40404
rect 4340 40348 8764 40404
rect 8820 40348 8830 40404
rect 15362 40348 15372 40404
rect 15428 40348 17724 40404
rect 17780 40348 17790 40404
rect 22642 40348 22652 40404
rect 22708 40348 24668 40404
rect 24724 40348 24734 40404
rect 2146 40236 2156 40292
rect 2212 40236 2222 40292
rect 8194 40236 8204 40292
rect 8260 40236 9324 40292
rect 9380 40236 9996 40292
rect 10052 40236 10062 40292
rect 18050 40236 18060 40292
rect 18116 40236 19628 40292
rect 19684 40236 19694 40292
rect 0 40180 112 40208
rect 28448 40180 28560 40208
rect 0 40124 812 40180
rect 868 40124 878 40180
rect 5058 40124 5068 40180
rect 5124 40124 8092 40180
rect 8148 40124 8158 40180
rect 17266 40124 17276 40180
rect 17332 40124 24780 40180
rect 24836 40124 24846 40180
rect 25666 40124 25676 40180
rect 25732 40124 28560 40180
rect 0 40096 112 40124
rect 28448 40096 28560 40124
rect 4454 39956 4464 40012
rect 4520 39956 4568 40012
rect 4624 39956 4672 40012
rect 4728 39956 4738 40012
rect 24454 39956 24464 40012
rect 24520 39956 24568 40012
rect 24624 39956 24672 40012
rect 24728 39956 24738 40012
rect 5282 39900 5292 39956
rect 5348 39900 9884 39956
rect 9940 39900 9950 39956
rect 6962 39788 6972 39844
rect 7028 39788 15148 39844
rect 15092 39732 15148 39788
rect 28448 39732 28560 39760
rect 3154 39676 3164 39732
rect 3220 39676 5964 39732
rect 6020 39676 6030 39732
rect 11890 39676 11900 39732
rect 11956 39676 12908 39732
rect 12964 39676 12974 39732
rect 15092 39676 24668 39732
rect 24724 39676 24734 39732
rect 27234 39676 27244 39732
rect 27300 39676 28560 39732
rect 28448 39648 28560 39676
rect 6626 39564 6636 39620
rect 6692 39564 15820 39620
rect 15876 39564 16716 39620
rect 16772 39564 16782 39620
rect 10994 39452 11004 39508
rect 11060 39452 11788 39508
rect 11844 39452 11854 39508
rect 12114 39340 12124 39396
rect 12180 39340 12348 39396
rect 12404 39340 12414 39396
rect 23202 39340 23212 39396
rect 23268 39340 27356 39396
rect 27412 39340 27422 39396
rect 28448 39284 28560 39312
rect 25666 39228 25676 39284
rect 25732 39228 28560 39284
rect 3794 39172 3804 39228
rect 3860 39172 3908 39228
rect 3964 39172 4012 39228
rect 4068 39172 4078 39228
rect 23794 39172 23804 39228
rect 23860 39172 23908 39228
rect 23964 39172 24012 39228
rect 24068 39172 24078 39228
rect 28448 39200 28560 39228
rect 26898 39116 26908 39172
rect 26964 39116 26974 39172
rect 6738 39004 6748 39060
rect 6804 39004 7196 39060
rect 7252 39004 7262 39060
rect 11218 39004 11228 39060
rect 11284 39004 26236 39060
rect 26292 39004 26302 39060
rect 2706 38892 2716 38948
rect 2772 38892 3612 38948
rect 3668 38892 5180 38948
rect 5236 38892 5628 38948
rect 5684 38892 5694 38948
rect 6178 38892 6188 38948
rect 6244 38892 7644 38948
rect 7700 38892 7710 38948
rect 0 38836 112 38864
rect 26908 38836 26964 39116
rect 28448 38836 28560 38864
rect 0 38780 588 38836
rect 644 38780 654 38836
rect 4274 38780 4284 38836
rect 4340 38780 8988 38836
rect 9044 38780 9054 38836
rect 15026 38780 15036 38836
rect 15092 38780 26236 38836
rect 26292 38780 26302 38836
rect 26908 38780 28560 38836
rect 0 38752 112 38780
rect 28448 38752 28560 38780
rect 1698 38668 1708 38724
rect 1764 38668 5964 38724
rect 6020 38668 6030 38724
rect 1698 38556 1708 38612
rect 1764 38556 1774 38612
rect 7634 38556 7644 38612
rect 7700 38556 12460 38612
rect 12516 38556 12526 38612
rect 1708 38052 1764 38556
rect 4454 38388 4464 38444
rect 4520 38388 4568 38444
rect 4624 38388 4672 38444
rect 4728 38388 4738 38444
rect 24454 38388 24464 38444
rect 24520 38388 24568 38444
rect 24624 38388 24672 38444
rect 24728 38388 24738 38444
rect 28448 38388 28560 38416
rect 27234 38332 27244 38388
rect 27300 38332 28560 38388
rect 28448 38304 28560 38332
rect 12562 38220 12572 38276
rect 12628 38220 12908 38276
rect 12964 38220 12974 38276
rect 13346 38220 13356 38276
rect 13412 38220 26348 38276
rect 26404 38220 26414 38276
rect 2370 38108 2380 38164
rect 2436 38108 2604 38164
rect 2660 38108 2670 38164
rect 1586 37996 1596 38052
rect 1652 37996 1764 38052
rect 9202 37996 9212 38052
rect 9268 37996 9548 38052
rect 9604 37996 10556 38052
rect 10612 37996 10622 38052
rect 11106 37996 11116 38052
rect 11172 37996 11900 38052
rect 11956 37996 11966 38052
rect 12114 37996 12124 38052
rect 12180 37996 13132 38052
rect 13188 37996 13198 38052
rect 25554 37996 25564 38052
rect 25620 37996 26236 38052
rect 26292 37996 26302 38052
rect 28448 37940 28560 37968
rect 3154 37884 3164 37940
rect 3220 37884 6748 37940
rect 6804 37884 11004 37940
rect 11060 37884 11070 37940
rect 12450 37884 12460 37940
rect 12516 37884 17500 37940
rect 17556 37884 17566 37940
rect 25666 37884 25676 37940
rect 25732 37884 28560 37940
rect 28448 37856 28560 37884
rect 2706 37772 2716 37828
rect 2772 37772 6356 37828
rect 7522 37772 7532 37828
rect 7588 37772 18844 37828
rect 18900 37772 18910 37828
rect 6300 37716 6356 37772
rect 6300 37660 9212 37716
rect 9268 37660 9278 37716
rect 3794 37604 3804 37660
rect 3860 37604 3908 37660
rect 3964 37604 4012 37660
rect 4068 37604 4078 37660
rect 23794 37604 23804 37660
rect 23860 37604 23908 37660
rect 23964 37604 24012 37660
rect 24068 37604 24078 37660
rect 1250 37548 1260 37604
rect 1316 37548 2716 37604
rect 2772 37548 2782 37604
rect 9314 37548 9324 37604
rect 9380 37548 9772 37604
rect 9828 37548 9838 37604
rect 0 37492 112 37520
rect 28448 37492 28560 37520
rect 0 37436 924 37492
rect 980 37436 990 37492
rect 6738 37436 6748 37492
rect 6804 37436 7756 37492
rect 7812 37436 7822 37492
rect 8194 37436 8204 37492
rect 8260 37436 26236 37492
rect 26292 37436 26302 37492
rect 26898 37436 26908 37492
rect 26964 37436 28560 37492
rect 0 37408 112 37436
rect 28448 37408 28560 37436
rect 2482 37324 2492 37380
rect 2548 37324 21532 37380
rect 21588 37324 21598 37380
rect 1922 37212 1932 37268
rect 1988 37212 2268 37268
rect 2324 37212 2334 37268
rect 3490 37212 3500 37268
rect 3556 37212 8316 37268
rect 8372 37212 15596 37268
rect 15652 37212 17164 37268
rect 17220 37212 17230 37268
rect 7522 37100 7532 37156
rect 7588 37100 13580 37156
rect 13636 37100 13646 37156
rect 28448 37044 28560 37072
rect 466 36988 476 37044
rect 532 36988 1036 37044
rect 1092 36988 5068 37044
rect 5124 36988 5628 37044
rect 5684 36988 5694 37044
rect 25442 36988 25452 37044
rect 25508 36988 28560 37044
rect 1596 36932 1652 36988
rect 28448 36960 28560 36988
rect 1586 36876 1596 36932
rect 1652 36876 1662 36932
rect 12786 36876 12796 36932
rect 12852 36876 14252 36932
rect 14308 36876 14318 36932
rect 4454 36820 4464 36876
rect 4520 36820 4568 36876
rect 4624 36820 4672 36876
rect 4728 36820 4738 36876
rect 24454 36820 24464 36876
rect 24520 36820 24568 36876
rect 24624 36820 24672 36876
rect 24728 36820 24738 36876
rect 14690 36764 14700 36820
rect 14756 36764 14766 36820
rect 1922 36652 1932 36708
rect 1988 36652 3052 36708
rect 3108 36652 4844 36708
rect 4900 36652 10108 36708
rect 10164 36652 10174 36708
rect 12786 36652 12796 36708
rect 12852 36652 13244 36708
rect 13300 36652 13310 36708
rect 14700 36596 14756 36764
rect 18274 36652 18284 36708
rect 18340 36652 22204 36708
rect 22260 36652 22270 36708
rect 28448 36596 28560 36624
rect 1698 36540 1708 36596
rect 1764 36540 2044 36596
rect 2100 36540 3948 36596
rect 4004 36540 9996 36596
rect 10052 36540 12124 36596
rect 12180 36540 12190 36596
rect 14690 36540 14700 36596
rect 14756 36540 14766 36596
rect 27234 36540 27244 36596
rect 27300 36540 28560 36596
rect 28448 36512 28560 36540
rect 2594 36428 2604 36484
rect 2660 36428 3388 36484
rect 3444 36428 3454 36484
rect 9314 36428 9324 36484
rect 9380 36428 9548 36484
rect 9604 36428 9614 36484
rect 14354 36428 14364 36484
rect 14420 36428 14812 36484
rect 14868 36428 14878 36484
rect 690 36316 700 36372
rect 756 36316 6636 36372
rect 6692 36316 6702 36372
rect 10546 36316 10556 36372
rect 10612 36316 17444 36372
rect 17388 36260 17444 36316
rect 8978 36204 8988 36260
rect 9044 36204 9324 36260
rect 9380 36204 9390 36260
rect 17378 36204 17388 36260
rect 17444 36204 18284 36260
rect 18340 36204 18350 36260
rect 0 36148 112 36176
rect 28448 36148 28560 36176
rect 0 36092 252 36148
rect 308 36092 318 36148
rect 7858 36092 7868 36148
rect 7924 36092 23660 36148
rect 23716 36092 23726 36148
rect 25666 36092 25676 36148
rect 25732 36092 28560 36148
rect 0 36064 112 36092
rect 3794 36036 3804 36092
rect 3860 36036 3908 36092
rect 3964 36036 4012 36092
rect 4068 36036 4078 36092
rect 23794 36036 23804 36092
rect 23860 36036 23908 36092
rect 23964 36036 24012 36092
rect 24068 36036 24078 36092
rect 28448 36064 28560 36092
rect 6850 35980 6860 36036
rect 6916 35980 8092 36036
rect 8148 35980 8158 36036
rect 8306 35980 8316 36036
rect 8372 35980 9100 36036
rect 9156 35980 9166 36036
rect 26898 35980 26908 36036
rect 26964 35980 26974 36036
rect 6738 35868 6748 35924
rect 6804 35868 26348 35924
rect 26404 35868 26414 35924
rect 5842 35756 5852 35812
rect 5908 35756 10556 35812
rect 10612 35756 10622 35812
rect 26908 35700 26964 35980
rect 28448 35700 28560 35728
rect 7634 35644 7644 35700
rect 7700 35644 8316 35700
rect 8372 35644 8382 35700
rect 26908 35644 28560 35700
rect 28448 35616 28560 35644
rect 5394 35532 5404 35588
rect 5460 35532 5852 35588
rect 5908 35532 5918 35588
rect 7074 35532 7084 35588
rect 7140 35532 7868 35588
rect 7924 35532 15148 35588
rect 25890 35532 25900 35588
rect 25956 35532 26236 35588
rect 26292 35532 26302 35588
rect 15092 35476 15148 35532
rect 5730 35420 5740 35476
rect 5796 35420 6300 35476
rect 6356 35420 6366 35476
rect 8866 35420 8876 35476
rect 8932 35420 9100 35476
rect 9156 35420 9166 35476
rect 15092 35420 21532 35476
rect 21588 35420 21598 35476
rect 8082 35308 8092 35364
rect 8148 35308 8652 35364
rect 8708 35308 9324 35364
rect 9380 35308 9390 35364
rect 13122 35308 13132 35364
rect 13188 35308 19740 35364
rect 19796 35308 19806 35364
rect 4454 35252 4464 35308
rect 4520 35252 4568 35308
rect 4624 35252 4672 35308
rect 4728 35252 4738 35308
rect 24454 35252 24464 35308
rect 24520 35252 24568 35308
rect 24624 35252 24672 35308
rect 24728 35252 24738 35308
rect 28448 35252 28560 35280
rect 12086 35196 12124 35252
rect 12180 35196 12190 35252
rect 15922 35196 15932 35252
rect 15988 35196 16828 35252
rect 16884 35196 16894 35252
rect 27234 35196 27244 35252
rect 27300 35196 28560 35252
rect 28448 35168 28560 35196
rect 9986 35084 9996 35140
rect 10052 35084 28140 35140
rect 28196 35084 28206 35140
rect 13234 34972 13244 35028
rect 13300 34972 14028 35028
rect 14084 34972 14094 35028
rect 17910 34972 17948 35028
rect 18004 34972 19852 35028
rect 19908 34972 19918 35028
rect 4274 34860 4284 34916
rect 4340 34860 5404 34916
rect 5460 34860 5470 34916
rect 12114 34860 12124 34916
rect 12180 34860 12908 34916
rect 12964 34860 12974 34916
rect 14578 34860 14588 34916
rect 14644 34860 26236 34916
rect 26292 34860 26302 34916
rect 0 34804 112 34832
rect 28448 34804 28560 34832
rect 0 34748 6076 34804
rect 6132 34748 6142 34804
rect 13010 34748 13020 34804
rect 13076 34748 24892 34804
rect 24948 34748 24958 34804
rect 25666 34748 25676 34804
rect 25732 34748 28560 34804
rect 0 34720 112 34748
rect 28448 34720 28560 34748
rect 12562 34636 12572 34692
rect 12628 34636 13692 34692
rect 13748 34636 13758 34692
rect 3794 34468 3804 34524
rect 3860 34468 3908 34524
rect 3964 34468 4012 34524
rect 4068 34468 4078 34524
rect 23794 34468 23804 34524
rect 23860 34468 23908 34524
rect 23964 34468 24012 34524
rect 24068 34468 24078 34524
rect 5954 34412 5964 34468
rect 6020 34412 7084 34468
rect 7140 34412 15148 34468
rect 15204 34412 15214 34468
rect 28448 34356 28560 34384
rect 1698 34300 1708 34356
rect 1764 34300 24668 34356
rect 24724 34300 24734 34356
rect 26898 34300 26908 34356
rect 26964 34300 28560 34356
rect 28448 34272 28560 34300
rect 2482 34188 2492 34244
rect 2548 34188 5180 34244
rect 5236 34188 5246 34244
rect 12226 34188 12236 34244
rect 12292 34188 13356 34244
rect 13412 34188 13422 34244
rect 4274 34076 4284 34132
rect 4340 34076 5404 34132
rect 5460 34076 12572 34132
rect 12628 34076 12638 34132
rect 16594 34076 16604 34132
rect 16660 34076 18508 34132
rect 18564 34076 18574 34132
rect 11890 33964 11900 34020
rect 11956 33964 26236 34020
rect 26292 33964 26302 34020
rect 28448 33908 28560 33936
rect 5730 33852 5740 33908
rect 5796 33852 7420 33908
rect 7476 33852 7486 33908
rect 23538 33852 23548 33908
rect 23604 33852 24668 33908
rect 24724 33852 24734 33908
rect 25666 33852 25676 33908
rect 25732 33852 28560 33908
rect 28448 33824 28560 33852
rect 7298 33740 7308 33796
rect 7364 33740 7868 33796
rect 7924 33740 7934 33796
rect 4454 33684 4464 33740
rect 4520 33684 4568 33740
rect 4624 33684 4672 33740
rect 4728 33684 4738 33740
rect 24454 33684 24464 33740
rect 24520 33684 24568 33740
rect 24624 33684 24672 33740
rect 24728 33684 24738 33740
rect 5170 33628 5180 33684
rect 5236 33628 8540 33684
rect 8596 33628 9548 33684
rect 9604 33628 9614 33684
rect 3266 33516 3276 33572
rect 3332 33516 4172 33572
rect 4228 33516 4238 33572
rect 6066 33516 6076 33572
rect 6132 33516 9996 33572
rect 10052 33516 10062 33572
rect 15092 33516 15596 33572
rect 15652 33516 15662 33572
rect 17714 33516 17724 33572
rect 17780 33516 18396 33572
rect 18452 33516 18462 33572
rect 0 33460 112 33488
rect 9996 33460 10052 33516
rect 15092 33460 15148 33516
rect 28448 33460 28560 33488
rect 0 33404 3388 33460
rect 7186 33404 7196 33460
rect 7252 33404 8316 33460
rect 8372 33404 8382 33460
rect 9996 33404 14588 33460
rect 14644 33404 15148 33460
rect 27234 33404 27244 33460
rect 27300 33404 28560 33460
rect 0 33376 112 33404
rect 3332 33348 3388 33404
rect 28448 33376 28560 33404
rect 3332 33292 8652 33348
rect 8708 33292 8718 33348
rect 1698 33180 1708 33236
rect 1764 33180 1932 33236
rect 1988 33180 1998 33236
rect 5170 33180 5180 33236
rect 5236 33180 5628 33236
rect 5684 33180 9212 33236
rect 9268 33180 9278 33236
rect 10882 33180 10892 33236
rect 10948 33180 17948 33236
rect 18004 33180 18014 33236
rect 10658 33068 10668 33124
rect 10724 33068 11452 33124
rect 11508 33068 11518 33124
rect 28448 33012 28560 33040
rect 10546 32956 10556 33012
rect 10612 32956 10622 33012
rect 25666 32956 25676 33012
rect 25732 32956 28560 33012
rect 3794 32900 3804 32956
rect 3860 32900 3908 32956
rect 3964 32900 4012 32956
rect 4068 32900 4078 32956
rect 7410 32732 7420 32788
rect 7476 32732 7980 32788
rect 8036 32732 8046 32788
rect 10556 32564 10612 32956
rect 23794 32900 23804 32956
rect 23860 32900 23908 32956
rect 23964 32900 24012 32956
rect 24068 32900 24078 32956
rect 28448 32928 28560 32956
rect 26898 32844 26908 32900
rect 26964 32844 26974 32900
rect 18274 32732 18284 32788
rect 18340 32732 18956 32788
rect 19012 32732 19022 32788
rect 17154 32620 17164 32676
rect 17220 32620 18620 32676
rect 18676 32620 18686 32676
rect 26908 32564 26964 32844
rect 28448 32564 28560 32592
rect 1250 32508 1260 32564
rect 1316 32508 1596 32564
rect 1652 32508 1662 32564
rect 6738 32508 6748 32564
rect 6804 32508 7196 32564
rect 7252 32508 7262 32564
rect 9202 32508 9212 32564
rect 9268 32508 10444 32564
rect 10500 32508 11788 32564
rect 11844 32508 11854 32564
rect 19058 32508 19068 32564
rect 19124 32508 19516 32564
rect 19572 32508 19582 32564
rect 26908 32508 28560 32564
rect 28448 32480 28560 32508
rect 2258 32396 2268 32452
rect 2324 32396 2604 32452
rect 2660 32396 2670 32452
rect 4274 32396 4284 32452
rect 4340 32396 26348 32452
rect 26404 32396 26414 32452
rect 8642 32284 8652 32340
rect 8708 32284 13804 32340
rect 13860 32284 13870 32340
rect 17602 32284 17612 32340
rect 17668 32284 24668 32340
rect 24724 32284 24734 32340
rect 27234 32284 27244 32340
rect 27300 32284 27310 32340
rect 9314 32172 9324 32228
rect 9380 32172 9996 32228
rect 10052 32172 10062 32228
rect 0 32116 112 32144
rect 4454 32116 4464 32172
rect 4520 32116 4568 32172
rect 4624 32116 4672 32172
rect 4728 32116 4738 32172
rect 24454 32116 24464 32172
rect 24520 32116 24568 32172
rect 24624 32116 24672 32172
rect 24728 32116 24738 32172
rect 27244 32116 27300 32284
rect 28448 32116 28560 32144
rect 0 32060 2044 32116
rect 2100 32060 2110 32116
rect 2258 32060 2268 32116
rect 2324 32060 2828 32116
rect 2884 32060 2894 32116
rect 27244 32060 28560 32116
rect 0 32032 112 32060
rect 28448 32032 28560 32060
rect 15362 31948 15372 32004
rect 15428 31948 24332 32004
rect 24388 31948 24398 32004
rect 2818 31836 2828 31892
rect 2884 31836 3724 31892
rect 3780 31836 3790 31892
rect 5058 31836 5068 31892
rect 5124 31836 6300 31892
rect 6356 31836 6366 31892
rect 16818 31836 16828 31892
rect 16884 31836 18172 31892
rect 18228 31836 18238 31892
rect 26898 31836 26908 31892
rect 26964 31836 28028 31892
rect 28084 31836 28094 31892
rect 2706 31724 2716 31780
rect 2772 31724 3500 31780
rect 3556 31724 3566 31780
rect 4050 31724 4060 31780
rect 4116 31724 4284 31780
rect 4340 31724 4350 31780
rect 7298 31724 7308 31780
rect 7364 31724 7644 31780
rect 7700 31724 8876 31780
rect 8932 31724 8942 31780
rect 12786 31724 12796 31780
rect 12852 31724 13244 31780
rect 13300 31724 13310 31780
rect 15026 31724 15036 31780
rect 15092 31724 15708 31780
rect 15764 31724 16268 31780
rect 16324 31724 16334 31780
rect 19170 31724 19180 31780
rect 19236 31724 19852 31780
rect 19908 31724 19918 31780
rect 28448 31668 28560 31696
rect 1250 31612 1260 31668
rect 1316 31612 1708 31668
rect 1764 31612 4844 31668
rect 4900 31612 4910 31668
rect 5282 31612 5292 31668
rect 5348 31612 5964 31668
rect 6020 31612 6030 31668
rect 8082 31612 8092 31668
rect 8148 31612 8540 31668
rect 8596 31612 8606 31668
rect 14802 31612 14812 31668
rect 14868 31612 16716 31668
rect 16772 31612 19068 31668
rect 19124 31612 19134 31668
rect 25666 31612 25676 31668
rect 25732 31612 28560 31668
rect 28448 31584 28560 31612
rect 4386 31500 4396 31556
rect 4452 31500 12012 31556
rect 12068 31500 27804 31556
rect 27860 31500 27870 31556
rect 10668 31388 10892 31444
rect 10948 31388 10958 31444
rect 13878 31388 13916 31444
rect 13972 31388 13982 31444
rect 14242 31388 14252 31444
rect 14308 31388 15148 31444
rect 15204 31388 15932 31444
rect 15988 31388 15998 31444
rect 3794 31332 3804 31388
rect 3860 31332 3908 31388
rect 3964 31332 4012 31388
rect 4068 31332 4078 31388
rect 10668 31332 10724 31388
rect 23794 31332 23804 31388
rect 23860 31332 23908 31388
rect 23964 31332 24012 31388
rect 24068 31332 24078 31388
rect 10658 31276 10668 31332
rect 10724 31276 10734 31332
rect 27234 31276 27244 31332
rect 27300 31276 27310 31332
rect 27244 31220 27300 31276
rect 28448 31220 28560 31248
rect 1810 31164 1820 31220
rect 1876 31164 4396 31220
rect 4452 31164 4462 31220
rect 15810 31164 15820 31220
rect 15876 31164 17052 31220
rect 17108 31164 17118 31220
rect 27244 31164 27468 31220
rect 27524 31164 27534 31220
rect 28018 31164 28028 31220
rect 28084 31164 28560 31220
rect 28448 31136 28560 31164
rect 10994 31052 11004 31108
rect 11060 31052 11340 31108
rect 11396 31052 11676 31108
rect 11732 31052 11742 31108
rect 11890 31052 11900 31108
rect 11956 31052 26684 31108
rect 26740 31052 26750 31108
rect 690 30940 700 30996
rect 756 30940 1260 30996
rect 1316 30940 1326 30996
rect 7970 30940 7980 30996
rect 8036 30940 14252 30996
rect 14308 30940 14318 30996
rect 19842 30940 19852 30996
rect 19908 30940 22876 30996
rect 22932 30940 22942 30996
rect 23100 30940 25900 30996
rect 25956 30940 25966 30996
rect 23100 30884 23156 30940
rect 2156 30828 2828 30884
rect 2884 30828 2894 30884
rect 6626 30828 6636 30884
rect 6692 30828 23156 30884
rect 25666 30828 25676 30884
rect 25732 30828 26236 30884
rect 26292 30828 26302 30884
rect 0 30772 112 30800
rect 2156 30772 2212 30828
rect 28448 30772 28560 30800
rect 0 30716 2212 30772
rect 2370 30716 2380 30772
rect 2436 30716 4284 30772
rect 4340 30716 4844 30772
rect 4900 30716 4910 30772
rect 13794 30716 13804 30772
rect 13860 30716 14700 30772
rect 14756 30716 14766 30772
rect 23650 30716 23660 30772
rect 23716 30716 24892 30772
rect 24948 30716 24958 30772
rect 25442 30716 25452 30772
rect 25508 30716 28560 30772
rect 0 30688 112 30716
rect 28448 30688 28560 30716
rect 6290 30604 6300 30660
rect 6356 30604 16716 30660
rect 16772 30604 16782 30660
rect 17826 30604 17836 30660
rect 17892 30604 17948 30660
rect 18004 30604 18014 30660
rect 4454 30548 4464 30604
rect 4520 30548 4568 30604
rect 4624 30548 4672 30604
rect 4728 30548 4738 30604
rect 7084 30548 7140 30604
rect 24454 30548 24464 30604
rect 24520 30548 24568 30604
rect 24624 30548 24672 30604
rect 24728 30548 24738 30604
rect 7074 30492 7084 30548
rect 7140 30492 7150 30548
rect 5394 30380 5404 30436
rect 5460 30380 5628 30436
rect 5684 30380 5694 30436
rect 5842 30380 5852 30436
rect 5908 30380 5918 30436
rect 10882 30380 10892 30436
rect 10948 30380 25788 30436
rect 25844 30380 25854 30436
rect 5852 30324 5908 30380
rect 28448 30324 28560 30352
rect 3378 30268 3388 30324
rect 3444 30268 7980 30324
rect 8036 30268 8046 30324
rect 26898 30268 26908 30324
rect 26964 30268 28560 30324
rect 28448 30240 28560 30268
rect 1138 30156 1148 30212
rect 1204 30156 2156 30212
rect 2212 30156 2222 30212
rect 5842 30156 5852 30212
rect 5908 30156 5918 30212
rect 8194 30156 8204 30212
rect 8260 30156 10220 30212
rect 10276 30156 15148 30212
rect 15922 30156 15932 30212
rect 15988 30156 16828 30212
rect 16884 30156 16894 30212
rect 25890 30156 25900 30212
rect 25956 30156 26236 30212
rect 26292 30156 26302 30212
rect 5852 30100 5908 30156
rect 15092 30100 15148 30156
rect 2818 30044 2828 30100
rect 2884 30044 3948 30100
rect 4004 30044 4014 30100
rect 5852 30044 7756 30100
rect 7812 30044 8316 30100
rect 8372 30044 8382 30100
rect 9986 30044 9996 30100
rect 10052 30044 13188 30100
rect 15092 30044 28364 30100
rect 28420 30044 28430 30100
rect 13132 29988 13188 30044
rect 3332 29932 12908 29988
rect 12964 29932 12974 29988
rect 13132 29932 23100 29988
rect 23156 29932 23166 29988
rect 1820 29820 2268 29876
rect 2324 29820 2334 29876
rect 0 29428 112 29456
rect 1820 29428 1876 29820
rect 3332 29652 3388 29932
rect 28448 29876 28560 29904
rect 5058 29820 5068 29876
rect 5124 29820 9996 29876
rect 10052 29820 10062 29876
rect 27234 29820 27244 29876
rect 27300 29820 28560 29876
rect 3794 29764 3804 29820
rect 3860 29764 3908 29820
rect 3964 29764 4012 29820
rect 4068 29764 4078 29820
rect 23794 29764 23804 29820
rect 23860 29764 23908 29820
rect 23964 29764 24012 29820
rect 24068 29764 24078 29820
rect 28448 29792 28560 29820
rect 2258 29596 2268 29652
rect 2324 29596 3388 29652
rect 3500 29596 5180 29652
rect 5236 29596 5246 29652
rect 12086 29596 12124 29652
rect 12180 29596 12190 29652
rect 3500 29540 3556 29596
rect 2034 29484 2044 29540
rect 2100 29484 2604 29540
rect 2660 29484 3500 29540
rect 3556 29484 3566 29540
rect 4050 29484 4060 29540
rect 4116 29484 25004 29540
rect 25060 29484 25070 29540
rect 28448 29428 28560 29456
rect 0 29372 1876 29428
rect 9762 29372 9772 29428
rect 9828 29372 10220 29428
rect 10276 29372 10286 29428
rect 11778 29372 11788 29428
rect 11844 29372 12460 29428
rect 12516 29372 12526 29428
rect 19702 29372 19740 29428
rect 19796 29372 19806 29428
rect 19954 29372 19964 29428
rect 20020 29372 20188 29428
rect 20244 29372 20254 29428
rect 26898 29372 26908 29428
rect 26964 29372 28560 29428
rect 0 29344 112 29372
rect 28448 29344 28560 29372
rect 802 29260 812 29316
rect 868 29260 1596 29316
rect 1652 29260 1662 29316
rect 9538 29260 9548 29316
rect 9604 29260 26236 29316
rect 26292 29260 26302 29316
rect 130 29148 140 29204
rect 196 29148 1484 29204
rect 1540 29148 8988 29204
rect 9044 29148 9054 29204
rect 15092 29148 25116 29204
rect 25172 29148 25182 29204
rect 15092 29092 15148 29148
rect 5506 29036 5516 29092
rect 5572 29036 15148 29092
rect 18386 29036 18396 29092
rect 18452 29036 18732 29092
rect 18788 29036 18798 29092
rect 4454 28980 4464 29036
rect 4520 28980 4568 29036
rect 4624 28980 4672 29036
rect 4728 28980 4738 29036
rect 24454 28980 24464 29036
rect 24520 28980 24568 29036
rect 24624 28980 24672 29036
rect 24728 28980 24738 29036
rect 28448 28980 28560 29008
rect 6738 28924 6748 28980
rect 6804 28924 6972 28980
rect 7028 28924 7038 28980
rect 19730 28924 19740 28980
rect 19796 28924 20076 28980
rect 20132 28924 20142 28980
rect 27234 28924 27244 28980
rect 27300 28924 28560 28980
rect 28448 28896 28560 28924
rect 10994 28812 11004 28868
rect 11060 28812 11340 28868
rect 11396 28812 11788 28868
rect 11844 28812 11854 28868
rect 12898 28812 12908 28868
rect 12964 28812 13580 28868
rect 13636 28812 14364 28868
rect 14420 28812 14430 28868
rect 18946 28812 18956 28868
rect 19012 28812 20412 28868
rect 20468 28812 20478 28868
rect 578 28700 588 28756
rect 644 28700 1596 28756
rect 1652 28700 1662 28756
rect 2706 28700 2716 28756
rect 2772 28700 25564 28756
rect 25620 28700 25630 28756
rect 25778 28700 25788 28756
rect 25844 28700 26236 28756
rect 26292 28700 26302 28756
rect 1810 28588 1820 28644
rect 1876 28588 2492 28644
rect 2548 28588 6972 28644
rect 7028 28588 7038 28644
rect 11862 28588 11900 28644
rect 11956 28588 11966 28644
rect 12450 28588 12460 28644
rect 12516 28588 14364 28644
rect 14420 28588 14430 28644
rect 14578 28588 14588 28644
rect 14644 28588 14924 28644
rect 14980 28588 15596 28644
rect 15652 28588 15662 28644
rect 19730 28588 19740 28644
rect 19796 28588 20076 28644
rect 20132 28588 20142 28644
rect 28448 28532 28560 28560
rect 3462 28476 3500 28532
rect 3556 28476 3566 28532
rect 6626 28476 6636 28532
rect 6692 28476 8652 28532
rect 8708 28476 8718 28532
rect 10882 28476 10892 28532
rect 10948 28476 11340 28532
rect 11396 28476 11406 28532
rect 15810 28476 15820 28532
rect 15876 28476 16380 28532
rect 16436 28476 16940 28532
rect 16996 28476 17006 28532
rect 27234 28476 27244 28532
rect 27300 28476 28560 28532
rect 28448 28448 28560 28476
rect 5058 28364 5068 28420
rect 5124 28364 5740 28420
rect 5796 28364 5806 28420
rect 16146 28364 16156 28420
rect 16212 28364 25676 28420
rect 25732 28364 25742 28420
rect 3794 28196 3804 28252
rect 3860 28196 3908 28252
rect 3964 28196 4012 28252
rect 4068 28196 4078 28252
rect 23794 28196 23804 28252
rect 23860 28196 23908 28252
rect 23964 28196 24012 28252
rect 24068 28196 24078 28252
rect 19478 28140 19516 28196
rect 19572 28140 19582 28196
rect 0 28084 112 28112
rect 28448 28084 28560 28112
rect 0 28028 476 28084
rect 532 28028 542 28084
rect 3378 28028 3388 28084
rect 3444 28028 3482 28084
rect 4946 28028 4956 28084
rect 5012 28028 19908 28084
rect 20066 28028 20076 28084
rect 20132 28028 26348 28084
rect 26404 28028 26414 28084
rect 27234 28028 27244 28084
rect 27300 28028 28560 28084
rect 0 28000 112 28028
rect 19852 27972 19908 28028
rect 28448 28000 28560 28028
rect 2594 27916 2604 27972
rect 2660 27916 4844 27972
rect 4900 27916 4910 27972
rect 8978 27916 8988 27972
rect 9044 27916 9436 27972
rect 9492 27916 9502 27972
rect 10882 27916 10892 27972
rect 10948 27916 17332 27972
rect 17490 27916 17500 27972
rect 17556 27916 17724 27972
rect 17780 27916 18172 27972
rect 18228 27916 18238 27972
rect 19852 27916 25676 27972
rect 25732 27916 25742 27972
rect 17276 27860 17332 27916
rect 4274 27804 4284 27860
rect 4340 27804 5292 27860
rect 5348 27804 5358 27860
rect 5702 27804 5740 27860
rect 5796 27804 7084 27860
rect 7140 27804 7150 27860
rect 8194 27804 8204 27860
rect 8260 27804 9324 27860
rect 9380 27804 9390 27860
rect 14018 27804 14028 27860
rect 14084 27804 15148 27860
rect 15204 27804 15214 27860
rect 17276 27804 24332 27860
rect 24388 27804 24398 27860
rect 914 27692 924 27748
rect 980 27692 1484 27748
rect 1540 27692 1550 27748
rect 17378 27692 17388 27748
rect 17444 27692 24668 27748
rect 24724 27692 24734 27748
rect 28448 27636 28560 27664
rect 14578 27580 14588 27636
rect 14644 27580 15596 27636
rect 15652 27580 15662 27636
rect 19058 27580 19068 27636
rect 19124 27580 19292 27636
rect 19348 27580 19358 27636
rect 27234 27580 27244 27636
rect 27300 27580 28560 27636
rect 28448 27552 28560 27580
rect 19478 27468 19516 27524
rect 19572 27468 19582 27524
rect 4454 27412 4464 27468
rect 4520 27412 4568 27468
rect 4624 27412 4672 27468
rect 4728 27412 4738 27468
rect 24454 27412 24464 27468
rect 24520 27412 24568 27468
rect 24624 27412 24672 27468
rect 24728 27412 24738 27468
rect 10770 27356 10780 27412
rect 10836 27356 10846 27412
rect 13682 27356 13692 27412
rect 13748 27356 14476 27412
rect 14532 27356 21868 27412
rect 21924 27356 21934 27412
rect 10780 27300 10836 27356
rect 5506 27244 5516 27300
rect 5572 27244 5852 27300
rect 5908 27244 5918 27300
rect 10546 27244 10556 27300
rect 10612 27244 10836 27300
rect 14690 27244 14700 27300
rect 14756 27244 24668 27300
rect 24724 27244 24734 27300
rect 28448 27188 28560 27216
rect 25666 27132 25676 27188
rect 25732 27132 28560 27188
rect 28448 27104 28560 27132
rect 1250 27020 1260 27076
rect 1316 27020 1708 27076
rect 1764 27020 1774 27076
rect 8306 27020 8316 27076
rect 8372 27020 8652 27076
rect 8708 27020 11340 27076
rect 11396 27020 16492 27076
rect 16548 27020 17724 27076
rect 17780 27020 17790 27076
rect 914 26908 924 26964
rect 980 26908 6748 26964
rect 6804 26908 6814 26964
rect 9874 26908 9884 26964
rect 9940 26908 26236 26964
rect 26292 26908 26302 26964
rect 2482 26796 2492 26852
rect 2548 26796 2828 26852
rect 2884 26796 2894 26852
rect 12898 26796 12908 26852
rect 12964 26796 13916 26852
rect 13972 26796 13982 26852
rect 17154 26796 17164 26852
rect 17220 26796 18172 26852
rect 18228 26796 18238 26852
rect 0 26740 112 26768
rect 28448 26740 28560 26768
rect 0 26684 3612 26740
rect 3668 26684 3678 26740
rect 27234 26684 27244 26740
rect 27300 26684 28560 26740
rect 0 26656 112 26684
rect 3794 26628 3804 26684
rect 3860 26628 3908 26684
rect 3964 26628 4012 26684
rect 4068 26628 4078 26684
rect 23794 26628 23804 26684
rect 23860 26628 23908 26684
rect 23964 26628 24012 26684
rect 24068 26628 24078 26684
rect 28448 26656 28560 26684
rect 5842 26572 5852 26628
rect 5908 26572 16044 26628
rect 16100 26572 16110 26628
rect 3490 26460 3500 26516
rect 3556 26460 3836 26516
rect 3892 26460 6300 26516
rect 6356 26460 7644 26516
rect 7700 26460 13468 26516
rect 13524 26460 13534 26516
rect 14550 26460 14588 26516
rect 14644 26460 14654 26516
rect 13346 26348 13356 26404
rect 13412 26348 14700 26404
rect 14756 26348 14766 26404
rect 15092 26348 26348 26404
rect 26404 26348 26414 26404
rect 15092 26292 15148 26348
rect 28448 26292 28560 26320
rect 6178 26236 6188 26292
rect 6244 26236 15148 26292
rect 25666 26236 25676 26292
rect 25732 26236 28560 26292
rect 28448 26208 28560 26236
rect 242 26124 252 26180
rect 308 26124 1036 26180
rect 1092 26124 2044 26180
rect 2100 26124 2110 26180
rect 2818 26124 2828 26180
rect 2884 26124 13244 26180
rect 13300 26124 15148 26180
rect 19618 26124 19628 26180
rect 19684 26124 26236 26180
rect 26292 26124 26302 26180
rect 1474 26012 1484 26068
rect 1540 26012 8092 26068
rect 8148 26012 9324 26068
rect 9380 26012 9390 26068
rect 15092 25956 15148 26124
rect 18610 26012 18620 26068
rect 18676 26012 19180 26068
rect 19236 26012 19246 26068
rect 15092 25900 20188 25956
rect 20244 25900 20254 25956
rect 4454 25844 4464 25900
rect 4520 25844 4568 25900
rect 4624 25844 4672 25900
rect 4728 25844 4738 25900
rect 24454 25844 24464 25900
rect 24520 25844 24568 25900
rect 24624 25844 24672 25900
rect 24728 25844 24738 25900
rect 28448 25844 28560 25872
rect 3266 25788 3276 25844
rect 3332 25788 3500 25844
rect 3556 25788 3566 25844
rect 27234 25788 27244 25844
rect 27300 25788 28560 25844
rect 28448 25760 28560 25788
rect 3042 25676 3052 25732
rect 3108 25676 3724 25732
rect 3780 25676 3790 25732
rect 12002 25676 12012 25732
rect 12068 25676 14924 25732
rect 14980 25676 14990 25732
rect 17490 25676 17500 25732
rect 17556 25676 18396 25732
rect 18452 25676 18462 25732
rect 19282 25676 19292 25732
rect 19348 25676 19358 25732
rect 2034 25564 2044 25620
rect 2100 25564 6636 25620
rect 6692 25564 10332 25620
rect 10388 25564 10398 25620
rect 18498 25564 18508 25620
rect 18564 25564 18956 25620
rect 19012 25564 19022 25620
rect 1698 25452 1708 25508
rect 1764 25452 3836 25508
rect 3892 25452 3902 25508
rect 0 25396 112 25424
rect 19292 25396 19348 25676
rect 19730 25452 19740 25508
rect 19796 25452 20636 25508
rect 20692 25452 21308 25508
rect 21364 25452 21374 25508
rect 25554 25452 25564 25508
rect 25620 25452 26236 25508
rect 26292 25452 26302 25508
rect 28448 25396 28560 25424
rect 0 25340 2716 25396
rect 2772 25340 5292 25396
rect 5348 25340 5358 25396
rect 18386 25340 18396 25396
rect 18452 25340 19964 25396
rect 20020 25340 20030 25396
rect 27346 25340 27356 25396
rect 27412 25340 28560 25396
rect 0 25312 112 25340
rect 28448 25312 28560 25340
rect 2818 25228 2828 25284
rect 2884 25228 3500 25284
rect 3556 25228 3566 25284
rect 16930 25228 16940 25284
rect 16996 25228 23548 25284
rect 23604 25228 23614 25284
rect 8726 25116 8764 25172
rect 8820 25116 8830 25172
rect 10434 25116 10444 25172
rect 10500 25116 10780 25172
rect 10836 25116 12684 25172
rect 12740 25116 15148 25172
rect 3794 25060 3804 25116
rect 3860 25060 3908 25116
rect 3964 25060 4012 25116
rect 4068 25060 4078 25116
rect 15092 25060 15148 25116
rect 23794 25060 23804 25116
rect 23860 25060 23908 25116
rect 23964 25060 24012 25116
rect 24068 25060 24078 25116
rect 6738 25004 6748 25060
rect 6804 25004 8316 25060
rect 8372 25004 8382 25060
rect 10658 25004 10668 25060
rect 10724 25004 13804 25060
rect 13860 25004 13870 25060
rect 15092 25004 18172 25060
rect 18228 25004 18396 25060
rect 18452 25004 18462 25060
rect 28448 24948 28560 24976
rect 1138 24892 1148 24948
rect 1204 24892 9660 24948
rect 9716 24892 9726 24948
rect 25666 24892 25676 24948
rect 25732 24892 28560 24948
rect 28448 24864 28560 24892
rect 7186 24780 7196 24836
rect 7252 24780 7532 24836
rect 7588 24780 7598 24836
rect 13906 24780 13916 24836
rect 13972 24780 26348 24836
rect 26404 24780 26414 24836
rect 1250 24668 1260 24724
rect 1316 24668 6692 24724
rect 9314 24668 9324 24724
rect 9380 24668 26236 24724
rect 26292 24668 26302 24724
rect 4454 24276 4464 24332
rect 4520 24276 4568 24332
rect 4624 24276 4672 24332
rect 4728 24276 4738 24332
rect 6636 24276 6692 24668
rect 13906 24556 13916 24612
rect 13972 24556 14700 24612
rect 14756 24556 14766 24612
rect 28448 24500 28560 24528
rect 8726 24444 8764 24500
rect 8820 24444 8830 24500
rect 12002 24444 12012 24500
rect 12068 24444 12460 24500
rect 12516 24444 12526 24500
rect 13346 24444 13356 24500
rect 13412 24444 16604 24500
rect 16660 24444 16670 24500
rect 27234 24444 27244 24500
rect 27300 24444 28560 24500
rect 28448 24416 28560 24444
rect 7522 24332 7532 24388
rect 7588 24332 8876 24388
rect 8932 24332 8942 24388
rect 10994 24332 11004 24388
rect 11060 24332 11564 24388
rect 11620 24332 11630 24388
rect 12338 24332 12348 24388
rect 12404 24332 13132 24388
rect 13188 24332 13198 24388
rect 14130 24332 14140 24388
rect 14196 24332 17724 24388
rect 17780 24332 18172 24388
rect 18228 24332 18238 24388
rect 24454 24276 24464 24332
rect 24520 24276 24568 24332
rect 24624 24276 24672 24332
rect 24728 24276 24738 24332
rect 6626 24220 6636 24276
rect 6692 24220 21028 24276
rect 20972 24164 21028 24220
rect 2006 24108 2044 24164
rect 2100 24108 2110 24164
rect 6178 24108 6188 24164
rect 6244 24108 15148 24164
rect 19394 24108 19404 24164
rect 19460 24108 19470 24164
rect 20972 24108 28252 24164
rect 28308 24108 28318 24164
rect 0 24052 112 24080
rect 0 23996 9268 24052
rect 13570 23996 13580 24052
rect 13636 23996 14140 24052
rect 14196 23996 14206 24052
rect 0 23968 112 23996
rect 4834 23884 4844 23940
rect 4900 23884 5404 23940
rect 5460 23884 5470 23940
rect 9212 23828 9268 23996
rect 15092 23940 15148 24108
rect 19404 24052 19460 24108
rect 28448 24052 28560 24080
rect 19404 23996 24668 24052
rect 24724 23996 24734 24052
rect 25442 23996 25452 24052
rect 25508 23996 28560 24052
rect 28448 23968 28560 23996
rect 12338 23884 12348 23940
rect 12404 23884 14252 23940
rect 14308 23884 14318 23940
rect 15092 23884 26236 23940
rect 26292 23884 26302 23940
rect 2258 23772 2268 23828
rect 2324 23772 4620 23828
rect 4676 23772 4686 23828
rect 9212 23772 17164 23828
rect 17220 23772 18508 23828
rect 18564 23772 19404 23828
rect 19460 23772 19470 23828
rect 2146 23660 2156 23716
rect 2212 23660 3052 23716
rect 3108 23660 4060 23716
rect 4116 23660 4126 23716
rect 4274 23660 4284 23716
rect 4340 23660 10780 23716
rect 10836 23660 10846 23716
rect 14690 23660 14700 23716
rect 14756 23660 16828 23716
rect 16884 23660 16894 23716
rect 28448 23604 28560 23632
rect 2006 23548 2044 23604
rect 2100 23548 2110 23604
rect 5618 23548 5628 23604
rect 5684 23548 5852 23604
rect 5908 23548 5918 23604
rect 6066 23548 6076 23604
rect 6132 23548 6972 23604
rect 7028 23548 7038 23604
rect 18386 23548 18396 23604
rect 18452 23548 18732 23604
rect 18788 23548 18956 23604
rect 19012 23548 19022 23604
rect 27346 23548 27356 23604
rect 27412 23548 28560 23604
rect 3794 23492 3804 23548
rect 3860 23492 3908 23548
rect 3964 23492 4012 23548
rect 4068 23492 4078 23548
rect 23794 23492 23804 23548
rect 23860 23492 23908 23548
rect 23964 23492 24012 23548
rect 24068 23492 24078 23548
rect 28448 23520 28560 23548
rect 5506 23436 5516 23492
rect 5572 23436 5628 23492
rect 5684 23436 5694 23492
rect 10658 23436 10668 23492
rect 10724 23436 14140 23492
rect 14196 23436 14206 23492
rect 15474 23436 15484 23492
rect 15540 23436 16380 23492
rect 16436 23436 16446 23492
rect 5058 23324 5068 23380
rect 5124 23324 6412 23380
rect 6468 23324 6478 23380
rect 6626 23324 6636 23380
rect 6692 23324 6972 23380
rect 7028 23324 7038 23380
rect 8642 23324 8652 23380
rect 8708 23324 8988 23380
rect 9044 23324 9054 23380
rect 12226 23324 12236 23380
rect 12292 23324 13804 23380
rect 13860 23324 13870 23380
rect 1698 23212 1708 23268
rect 1764 23212 24220 23268
rect 24276 23212 24286 23268
rect 28448 23156 28560 23184
rect 1586 23100 1596 23156
rect 1652 23100 3276 23156
rect 3332 23100 3342 23156
rect 5814 23100 5852 23156
rect 5908 23100 5918 23156
rect 6486 23100 6524 23156
rect 6580 23100 6590 23156
rect 14802 23100 14812 23156
rect 14868 23100 15708 23156
rect 15764 23100 15774 23156
rect 25666 23100 25676 23156
rect 25732 23100 28560 23156
rect 28448 23072 28560 23100
rect 10546 22988 10556 23044
rect 10612 22988 12012 23044
rect 12068 22988 14364 23044
rect 14420 22988 14430 23044
rect 6514 22876 6524 22932
rect 6580 22876 7196 22932
rect 7252 22876 7262 22932
rect 8306 22876 8316 22932
rect 8372 22876 10332 22932
rect 10388 22876 10398 22932
rect 11106 22764 11116 22820
rect 11172 22764 11340 22820
rect 11396 22764 11406 22820
rect 18162 22764 18172 22820
rect 18228 22764 18508 22820
rect 18564 22764 18574 22820
rect 0 22708 112 22736
rect 4454 22708 4464 22764
rect 4520 22708 4568 22764
rect 4624 22708 4672 22764
rect 4728 22708 4738 22764
rect 24454 22708 24464 22764
rect 24520 22708 24568 22764
rect 24624 22708 24672 22764
rect 24728 22708 24738 22764
rect 28448 22708 28560 22736
rect 0 22652 3388 22708
rect 0 22624 112 22652
rect 3332 22596 3388 22652
rect 5068 22652 17052 22708
rect 17108 22652 17948 22708
rect 18004 22652 18014 22708
rect 27234 22652 27244 22708
rect 27300 22652 28560 22708
rect 5068 22596 5124 22652
rect 28448 22624 28560 22652
rect 1922 22540 1932 22596
rect 1988 22540 2716 22596
rect 2772 22540 3052 22596
rect 3108 22540 3118 22596
rect 3332 22540 5124 22596
rect 5282 22540 5292 22596
rect 5348 22540 5852 22596
rect 5908 22540 5918 22596
rect 6860 22540 10220 22596
rect 10276 22540 10286 22596
rect 12226 22540 12236 22596
rect 12292 22540 12908 22596
rect 12964 22540 12974 22596
rect 15138 22540 15148 22596
rect 15204 22540 16380 22596
rect 16436 22540 16446 22596
rect 6860 22484 6916 22540
rect 1586 22428 1596 22484
rect 1652 22428 6916 22484
rect 8530 22428 8540 22484
rect 8596 22428 9772 22484
rect 9828 22428 11116 22484
rect 11172 22428 15148 22484
rect 4274 22316 4284 22372
rect 4340 22316 5292 22372
rect 5348 22316 5358 22372
rect 8194 22316 8204 22372
rect 8260 22316 9212 22372
rect 9268 22316 9278 22372
rect 11890 22316 11900 22372
rect 11956 22316 13692 22372
rect 13748 22316 13758 22372
rect 15092 22260 15148 22428
rect 15810 22316 15820 22372
rect 15876 22316 17388 22372
rect 17444 22316 17454 22372
rect 28448 22260 28560 22288
rect 8082 22204 8092 22260
rect 8148 22204 13916 22260
rect 13972 22204 14476 22260
rect 14532 22204 14542 22260
rect 15092 22204 25004 22260
rect 25060 22204 25070 22260
rect 27346 22204 27356 22260
rect 27412 22204 28560 22260
rect 14476 22148 14532 22204
rect 28448 22176 28560 22204
rect 13010 22092 13020 22148
rect 13076 22092 13086 22148
rect 14476 22092 16828 22148
rect 16884 22092 16894 22148
rect 5478 21980 5516 22036
rect 5572 21980 5582 22036
rect 12226 21980 12236 22036
rect 12292 21980 12460 22036
rect 12516 21980 12526 22036
rect 3794 21924 3804 21980
rect 3860 21924 3908 21980
rect 3964 21924 4012 21980
rect 4068 21924 4078 21980
rect 13020 21924 13076 22092
rect 23794 21924 23804 21980
rect 23860 21924 23908 21980
rect 23964 21924 24012 21980
rect 24068 21924 24078 21980
rect 7634 21868 7644 21924
rect 7700 21868 7710 21924
rect 13020 21868 13580 21924
rect 13636 21868 14812 21924
rect 14868 21868 14878 21924
rect 16258 21868 16268 21924
rect 16324 21868 19404 21924
rect 19460 21868 19470 21924
rect 7644 21812 7700 21868
rect 28448 21812 28560 21840
rect 6850 21756 6860 21812
rect 6916 21756 7196 21812
rect 7252 21756 7262 21812
rect 7644 21756 8092 21812
rect 8148 21756 8158 21812
rect 11228 21756 11452 21812
rect 11508 21756 11518 21812
rect 11666 21756 11676 21812
rect 11732 21756 13132 21812
rect 13188 21756 13198 21812
rect 25666 21756 25676 21812
rect 25732 21756 28560 21812
rect 2258 21644 2268 21700
rect 2324 21644 5740 21700
rect 5796 21644 5806 21700
rect 7046 21532 7084 21588
rect 7140 21532 7150 21588
rect 7298 21532 7308 21588
rect 7364 21532 7402 21588
rect 8418 21532 8428 21588
rect 8484 21532 9436 21588
rect 9492 21532 9502 21588
rect 3332 21420 10892 21476
rect 10948 21420 10958 21476
rect 0 21364 112 21392
rect 3332 21364 3388 21420
rect 11228 21364 11284 21756
rect 28448 21728 28560 21756
rect 18722 21644 18732 21700
rect 18788 21644 19180 21700
rect 19236 21644 19246 21700
rect 21858 21644 21868 21700
rect 21924 21644 27468 21700
rect 27524 21644 27534 21700
rect 11442 21532 11452 21588
rect 11508 21532 12124 21588
rect 12180 21532 12190 21588
rect 15138 21532 15148 21588
rect 15204 21532 15820 21588
rect 15876 21532 15886 21588
rect 16370 21532 16380 21588
rect 16436 21532 17612 21588
rect 17668 21532 17678 21588
rect 21522 21532 21532 21588
rect 21588 21532 27916 21588
rect 27972 21532 27982 21588
rect 12908 21420 14924 21476
rect 14980 21420 14990 21476
rect 15250 21420 15260 21476
rect 15316 21420 17164 21476
rect 17220 21420 17230 21476
rect 17826 21420 17836 21476
rect 17892 21420 18284 21476
rect 18340 21420 18350 21476
rect 19282 21420 19292 21476
rect 19348 21420 26236 21476
rect 26292 21420 26302 21476
rect 12908 21364 12964 21420
rect 28448 21364 28560 21392
rect 0 21308 3388 21364
rect 5954 21308 5964 21364
rect 6020 21308 7308 21364
rect 7364 21308 7374 21364
rect 9762 21308 9772 21364
rect 9828 21308 12124 21364
rect 12180 21308 12190 21364
rect 12898 21308 12908 21364
rect 12964 21308 12974 21364
rect 13682 21308 13692 21364
rect 13748 21308 13758 21364
rect 14690 21308 14700 21364
rect 14756 21308 15708 21364
rect 15764 21308 15774 21364
rect 16146 21308 16156 21364
rect 16212 21308 16716 21364
rect 16772 21308 22988 21364
rect 23044 21308 23054 21364
rect 25666 21308 25676 21364
rect 25732 21308 28560 21364
rect 0 21280 112 21308
rect 13692 21252 13748 21308
rect 16156 21252 16212 21308
rect 28448 21280 28560 21308
rect 3042 21196 3052 21252
rect 3108 21196 3276 21252
rect 3332 21196 3342 21252
rect 4946 21196 4956 21252
rect 5012 21196 12572 21252
rect 12628 21196 12638 21252
rect 13692 21196 14252 21252
rect 14308 21196 16212 21252
rect 4454 21140 4464 21196
rect 4520 21140 4568 21196
rect 4624 21140 4672 21196
rect 4728 21140 4738 21196
rect 24454 21140 24464 21196
rect 24520 21140 24568 21196
rect 24624 21140 24672 21196
rect 24728 21140 24738 21196
rect 8866 21084 8876 21140
rect 8932 21084 15148 21140
rect 15810 21084 15820 21140
rect 15876 21084 20748 21140
rect 20804 21084 20814 21140
rect 27346 21084 27356 21140
rect 27412 21084 27692 21140
rect 27748 21084 27758 21140
rect 15092 21028 15148 21084
rect 2146 20972 2156 21028
rect 2212 20972 3276 21028
rect 3332 20972 3342 21028
rect 5730 20972 5740 21028
rect 5796 20972 6300 21028
rect 6356 20972 8316 21028
rect 8372 20972 9660 21028
rect 9716 20972 9726 21028
rect 14914 20972 14924 21028
rect 14980 20972 14990 21028
rect 15092 20972 28028 21028
rect 28084 20972 28094 21028
rect 14924 20916 14980 20972
rect 28448 20916 28560 20944
rect 1698 20860 1708 20916
rect 1764 20860 1932 20916
rect 1988 20860 1998 20916
rect 5618 20860 5628 20916
rect 5684 20860 6524 20916
rect 6580 20860 6748 20916
rect 6804 20860 6814 20916
rect 13794 20860 13804 20916
rect 13860 20860 14252 20916
rect 14308 20860 14318 20916
rect 14924 20860 17052 20916
rect 17108 20860 17118 20916
rect 19730 20860 19740 20916
rect 19796 20860 20412 20916
rect 20468 20860 20478 20916
rect 26852 20860 28560 20916
rect 2146 20748 2156 20804
rect 2212 20748 2940 20804
rect 2996 20748 3006 20804
rect 5730 20748 5740 20804
rect 5796 20748 6412 20804
rect 6468 20748 6478 20804
rect 7858 20748 7868 20804
rect 7924 20748 8092 20804
rect 8148 20748 9716 20804
rect 9874 20748 9884 20804
rect 9940 20748 10444 20804
rect 10500 20748 10510 20804
rect 13346 20748 13356 20804
rect 13412 20748 14476 20804
rect 14532 20748 15820 20804
rect 15876 20748 16716 20804
rect 16772 20748 17388 20804
rect 17444 20748 17454 20804
rect 9660 20692 9716 20748
rect 26852 20692 26908 20860
rect 28448 20832 28560 20860
rect 9426 20636 9436 20692
rect 9492 20636 9604 20692
rect 9660 20636 26908 20692
rect 9548 20580 9604 20636
rect 802 20524 812 20580
rect 868 20524 9324 20580
rect 9380 20524 9390 20580
rect 9548 20524 15820 20580
rect 15876 20524 15886 20580
rect 16034 20524 16044 20580
rect 16100 20524 16716 20580
rect 16772 20524 16782 20580
rect 17042 20524 17052 20580
rect 17108 20524 17836 20580
rect 17892 20524 17902 20580
rect 28448 20468 28560 20496
rect 4498 20412 4508 20468
rect 4564 20412 5852 20468
rect 5908 20412 12180 20468
rect 12870 20412 12908 20468
rect 12964 20412 12974 20468
rect 14578 20412 14588 20468
rect 14644 20412 16268 20468
rect 16324 20412 16334 20468
rect 27794 20412 27804 20468
rect 27860 20412 28560 20468
rect 3794 20356 3804 20412
rect 3860 20356 3908 20412
rect 3964 20356 4012 20412
rect 4068 20356 4078 20412
rect 12124 20356 12180 20412
rect 23794 20356 23804 20412
rect 23860 20356 23908 20412
rect 23964 20356 24012 20412
rect 24068 20356 24078 20412
rect 28448 20384 28560 20412
rect 9538 20300 9548 20356
rect 9604 20300 10556 20356
rect 10612 20300 11900 20356
rect 11956 20300 11966 20356
rect 12124 20300 15148 20356
rect 15922 20300 15932 20356
rect 15988 20300 20524 20356
rect 20580 20300 21196 20356
rect 21252 20300 21262 20356
rect 15092 20244 15148 20300
rect 2370 20188 2380 20244
rect 2436 20188 2828 20244
rect 2884 20188 2894 20244
rect 11732 20188 12236 20244
rect 12292 20188 12796 20244
rect 12852 20188 12862 20244
rect 15092 20188 27916 20244
rect 27972 20188 27982 20244
rect 11732 20132 11788 20188
rect 5282 20076 5292 20132
rect 5348 20076 6748 20132
rect 6804 20076 8148 20132
rect 8306 20076 8316 20132
rect 8372 20076 11788 20132
rect 13234 20076 13244 20132
rect 13300 20076 15148 20132
rect 15204 20076 15214 20132
rect 15586 20076 15596 20132
rect 15652 20076 26908 20132
rect 0 20020 112 20048
rect 8092 20020 8148 20076
rect 26852 20020 26908 20076
rect 28448 20020 28560 20048
rect 0 19964 4788 20020
rect 4946 19964 4956 20020
rect 5012 19964 7196 20020
rect 7252 19964 7262 20020
rect 8092 19964 8876 20020
rect 8932 19964 8942 20020
rect 11442 19964 11452 20020
rect 11508 19964 12124 20020
rect 12180 19964 13132 20020
rect 13188 19964 13468 20020
rect 13524 19964 13534 20020
rect 15474 19964 15484 20020
rect 15540 19964 16604 20020
rect 16660 19964 16670 20020
rect 26852 19964 28560 20020
rect 0 19936 112 19964
rect 4732 19908 4788 19964
rect 15484 19908 15540 19964
rect 28448 19936 28560 19964
rect 1698 19852 1708 19908
rect 1764 19852 3500 19908
rect 3556 19852 4172 19908
rect 4228 19852 4238 19908
rect 4732 19852 11228 19908
rect 11284 19852 11294 19908
rect 11666 19852 11676 19908
rect 11732 19852 15540 19908
rect 578 19740 588 19796
rect 644 19740 7196 19796
rect 7252 19740 7262 19796
rect 9538 19740 9548 19796
rect 9604 19740 12348 19796
rect 12404 19740 13356 19796
rect 13412 19740 13422 19796
rect 14242 19740 14252 19796
rect 14308 19740 15596 19796
rect 15652 19740 15662 19796
rect 20524 19740 26012 19796
rect 26068 19740 26078 19796
rect 20524 19684 20580 19740
rect 6178 19628 6188 19684
rect 6244 19628 20580 19684
rect 4454 19572 4464 19628
rect 4520 19572 4568 19628
rect 4624 19572 4672 19628
rect 4728 19572 4738 19628
rect 24454 19572 24464 19628
rect 24520 19572 24568 19628
rect 24624 19572 24672 19628
rect 24728 19572 24738 19628
rect 28448 19572 28560 19600
rect 10882 19516 10892 19572
rect 10948 19516 11676 19572
rect 11732 19516 12572 19572
rect 12628 19516 12638 19572
rect 13906 19516 13916 19572
rect 13972 19516 16716 19572
rect 16772 19516 16782 19572
rect 24882 19516 24892 19572
rect 24948 19516 28560 19572
rect 28448 19488 28560 19516
rect 1586 19404 1596 19460
rect 1652 19404 2604 19460
rect 2660 19404 2670 19460
rect 2930 19404 2940 19460
rect 2996 19404 7644 19460
rect 7700 19404 7710 19460
rect 9986 19404 9996 19460
rect 10052 19404 11564 19460
rect 11620 19404 11630 19460
rect 11890 19404 11900 19460
rect 11956 19404 14364 19460
rect 14420 19404 14430 19460
rect 15362 19404 15372 19460
rect 15428 19404 16604 19460
rect 16660 19404 16670 19460
rect 11900 19348 11956 19404
rect 354 19292 364 19348
rect 420 19292 2716 19348
rect 2772 19292 3052 19348
rect 3108 19292 4508 19348
rect 4564 19292 4574 19348
rect 11106 19292 11116 19348
rect 11172 19292 11956 19348
rect 13794 19292 13804 19348
rect 13860 19292 14140 19348
rect 14196 19292 14206 19348
rect 14914 19292 14924 19348
rect 14980 19292 16156 19348
rect 16212 19292 16222 19348
rect 6626 19180 6636 19236
rect 6692 19180 7420 19236
rect 7476 19180 7486 19236
rect 7746 19180 7756 19236
rect 7812 19180 10332 19236
rect 10388 19180 10398 19236
rect 11778 19180 11788 19236
rect 11844 19180 14700 19236
rect 14756 19180 14766 19236
rect 15092 19180 15708 19236
rect 15764 19180 15774 19236
rect 10332 19124 10388 19180
rect 15092 19124 15148 19180
rect 28448 19124 28560 19152
rect 10332 19068 13244 19124
rect 13300 19068 13310 19124
rect 14130 19068 14140 19124
rect 14196 19068 15148 19124
rect 16034 19068 16044 19124
rect 16100 19068 16716 19124
rect 16772 19068 16782 19124
rect 23090 19068 23100 19124
rect 23156 19068 28560 19124
rect 28448 19040 28560 19068
rect 2930 18956 2940 19012
rect 2996 18956 10780 19012
rect 10836 18956 10846 19012
rect 5618 18844 5628 18900
rect 5684 18844 6300 18900
rect 6356 18844 6366 18900
rect 13346 18844 13356 18900
rect 13412 18844 18284 18900
rect 18340 18844 18350 18900
rect 3794 18788 3804 18844
rect 3860 18788 3908 18844
rect 3964 18788 4012 18844
rect 4068 18788 4078 18844
rect 23794 18788 23804 18844
rect 23860 18788 23908 18844
rect 23964 18788 24012 18844
rect 24068 18788 24078 18844
rect 2258 18732 2268 18788
rect 2324 18732 2716 18788
rect 2772 18732 3164 18788
rect 3220 18732 3612 18788
rect 3668 18732 3678 18788
rect 4274 18732 4284 18788
rect 4340 18732 4956 18788
rect 5012 18732 5022 18788
rect 10994 18732 11004 18788
rect 11060 18732 12796 18788
rect 12852 18732 12862 18788
rect 0 18676 112 18704
rect 28448 18676 28560 18704
rect 0 18620 9436 18676
rect 9492 18620 9502 18676
rect 13794 18620 13804 18676
rect 13860 18620 15148 18676
rect 15204 18620 15242 18676
rect 15810 18620 15820 18676
rect 15876 18620 16828 18676
rect 16884 18620 16894 18676
rect 17042 18620 17052 18676
rect 17108 18620 18284 18676
rect 18340 18620 18350 18676
rect 27906 18620 27916 18676
rect 27972 18620 28560 18676
rect 0 18592 112 18620
rect 28448 18592 28560 18620
rect 3154 18508 3164 18564
rect 3220 18508 6524 18564
rect 6580 18508 6590 18564
rect 8866 18508 8876 18564
rect 8932 18508 9548 18564
rect 9604 18508 10332 18564
rect 10388 18508 10398 18564
rect 14130 18508 14140 18564
rect 14196 18508 16268 18564
rect 16324 18508 16334 18564
rect 2482 18396 2492 18452
rect 2548 18396 9268 18452
rect 10098 18396 10108 18452
rect 10164 18396 13692 18452
rect 13748 18396 14364 18452
rect 14420 18396 14430 18452
rect 14578 18396 14588 18452
rect 14644 18396 15036 18452
rect 15092 18396 15102 18452
rect 16044 18396 16940 18452
rect 16996 18396 17006 18452
rect 18386 18396 18396 18452
rect 18452 18396 18956 18452
rect 19012 18396 19022 18452
rect 19506 18396 19516 18452
rect 19572 18396 26684 18452
rect 26740 18396 26750 18452
rect 3938 18284 3948 18340
rect 4004 18284 5964 18340
rect 6020 18284 6972 18340
rect 7028 18284 7038 18340
rect 4454 18004 4464 18060
rect 4520 18004 4568 18060
rect 4624 18004 4672 18060
rect 4728 18004 4738 18060
rect 2034 17836 2044 17892
rect 2100 17836 2828 17892
rect 2884 17836 4284 17892
rect 4340 17836 4350 17892
rect 4834 17836 4844 17892
rect 4900 17836 5852 17892
rect 5908 17836 9156 17892
rect 2146 17724 2156 17780
rect 2212 17724 2604 17780
rect 2660 17724 2670 17780
rect 9100 17668 9156 17836
rect 9212 17780 9268 18396
rect 16044 18228 16100 18396
rect 28448 18228 28560 18256
rect 11890 18172 11900 18228
rect 11956 18172 13804 18228
rect 13860 18172 13870 18228
rect 14018 18172 14028 18228
rect 14084 18172 14588 18228
rect 14644 18172 14654 18228
rect 15260 18172 16044 18228
rect 16100 18172 16110 18228
rect 16482 18172 16492 18228
rect 16548 18172 17052 18228
rect 17108 18172 17118 18228
rect 17378 18172 17388 18228
rect 17444 18172 17454 18228
rect 18498 18172 18508 18228
rect 18564 18172 18956 18228
rect 19012 18172 19022 18228
rect 28354 18172 28364 18228
rect 28420 18172 28560 18228
rect 15260 18116 15316 18172
rect 17388 18116 17444 18172
rect 28448 18144 28560 18172
rect 11218 18060 11228 18116
rect 11284 18060 15260 18116
rect 15316 18060 15326 18116
rect 15922 18060 15932 18116
rect 15988 18060 17444 18116
rect 24454 18004 24464 18060
rect 24520 18004 24568 18060
rect 24624 18004 24672 18060
rect 24728 18004 24738 18060
rect 14354 17948 14364 18004
rect 14420 17948 15148 18004
rect 15204 17948 17164 18004
rect 17220 17948 17230 18004
rect 14466 17836 14476 17892
rect 14532 17836 16940 17892
rect 16996 17836 17006 17892
rect 28448 17780 28560 17808
rect 9212 17724 16716 17780
rect 16772 17724 16782 17780
rect 26852 17724 28560 17780
rect 3714 17612 3724 17668
rect 3780 17612 4844 17668
rect 4900 17612 4910 17668
rect 6626 17612 6636 17668
rect 6692 17612 8092 17668
rect 8148 17612 8158 17668
rect 9100 17612 9996 17668
rect 10052 17612 10062 17668
rect 10770 17612 10780 17668
rect 10836 17612 10846 17668
rect 13458 17612 13468 17668
rect 13524 17612 13692 17668
rect 13748 17612 13758 17668
rect 14914 17612 14924 17668
rect 14980 17612 16940 17668
rect 16996 17612 17006 17668
rect 10780 17556 10836 17612
rect 26852 17556 26908 17724
rect 28448 17696 28560 17724
rect 2594 17500 2604 17556
rect 2660 17500 10836 17556
rect 10892 17500 26908 17556
rect 10892 17444 10948 17500
rect 3332 17388 6972 17444
rect 7028 17388 7038 17444
rect 9874 17388 9884 17444
rect 9940 17388 10948 17444
rect 11302 17388 11340 17444
rect 11396 17388 26908 17444
rect 0 17332 112 17360
rect 3332 17332 3388 17388
rect 26852 17332 26908 17388
rect 28448 17332 28560 17360
rect 0 17276 3388 17332
rect 3574 17276 3612 17332
rect 3668 17276 3678 17332
rect 4498 17276 4508 17332
rect 4564 17276 13356 17332
rect 13412 17276 13422 17332
rect 26852 17276 28560 17332
rect 0 17248 112 17276
rect 3794 17220 3804 17276
rect 3860 17220 3908 17276
rect 3964 17220 4012 17276
rect 4068 17220 4078 17276
rect 23794 17220 23804 17276
rect 23860 17220 23908 17276
rect 23964 17220 24012 17276
rect 24068 17220 24078 17276
rect 28448 17248 28560 17276
rect 5394 17164 5404 17220
rect 5460 17164 6188 17220
rect 6244 17164 7084 17220
rect 7140 17164 7150 17220
rect 13010 17164 13020 17220
rect 13076 17164 14924 17220
rect 14980 17164 14990 17220
rect 1586 17052 1596 17108
rect 1652 17052 3500 17108
rect 3556 17052 6636 17108
rect 6692 17052 6702 17108
rect 13122 17052 13132 17108
rect 13188 17052 13916 17108
rect 13972 17052 13982 17108
rect 14578 17052 14588 17108
rect 14644 17052 15596 17108
rect 15652 17052 15662 17108
rect 16146 17052 16156 17108
rect 16212 17052 16940 17108
rect 16996 17052 17006 17108
rect 8306 16940 8316 16996
rect 8372 16940 16044 16996
rect 16100 16940 16110 16996
rect 28448 16884 28560 16912
rect 3826 16828 3836 16884
rect 3892 16828 4956 16884
rect 5012 16828 5740 16884
rect 5796 16828 6636 16884
rect 6692 16828 7868 16884
rect 7924 16828 7934 16884
rect 9650 16828 9660 16884
rect 9716 16828 10164 16884
rect 13122 16828 13132 16884
rect 13188 16828 13356 16884
rect 13412 16828 13422 16884
rect 14018 16828 14028 16884
rect 14084 16828 16380 16884
rect 16436 16828 16446 16884
rect 16706 16828 16716 16884
rect 16772 16828 17948 16884
rect 18004 16828 21420 16884
rect 21476 16828 21486 16884
rect 27458 16828 27468 16884
rect 27524 16828 28560 16884
rect 10108 16772 10164 16828
rect 28448 16800 28560 16828
rect 10108 16716 13916 16772
rect 13972 16716 13982 16772
rect 21634 16716 21644 16772
rect 21700 16716 26012 16772
rect 26068 16716 26078 16772
rect 4386 16604 4396 16660
rect 4452 16604 4956 16660
rect 5012 16604 5628 16660
rect 5684 16604 5694 16660
rect 5842 16604 5852 16660
rect 5908 16604 8428 16660
rect 8484 16604 8494 16660
rect 10322 16604 10332 16660
rect 10388 16604 10892 16660
rect 10948 16604 10958 16660
rect 14326 16604 14364 16660
rect 14420 16604 14430 16660
rect 15092 16604 15372 16660
rect 15428 16604 15438 16660
rect 19954 16604 19964 16660
rect 20020 16604 26908 16660
rect 4454 16436 4464 16492
rect 4520 16436 4568 16492
rect 4624 16436 4672 16492
rect 4728 16436 4738 16492
rect 10098 16380 10108 16436
rect 10164 16380 11676 16436
rect 11732 16380 11742 16436
rect 13570 16380 13580 16436
rect 13636 16380 13804 16436
rect 13860 16380 13870 16436
rect 11676 16324 11732 16380
rect 15092 16324 15148 16604
rect 15250 16492 15260 16548
rect 15316 16492 16716 16548
rect 16772 16492 16782 16548
rect 17938 16492 17948 16548
rect 18004 16492 18508 16548
rect 18564 16492 18574 16548
rect 24454 16436 24464 16492
rect 24520 16436 24568 16492
rect 24624 16436 24672 16492
rect 24728 16436 24738 16492
rect 26852 16436 26908 16604
rect 28448 16436 28560 16464
rect 26852 16380 28560 16436
rect 28448 16352 28560 16380
rect 4722 16268 4732 16324
rect 4788 16268 4844 16324
rect 4900 16268 8036 16324
rect 8194 16268 8204 16324
rect 8260 16268 11116 16324
rect 11172 16268 11182 16324
rect 11676 16268 28252 16324
rect 28308 16268 28318 16324
rect 7980 16212 8036 16268
rect 1922 16156 1932 16212
rect 1988 16156 3164 16212
rect 3220 16156 6860 16212
rect 6916 16156 6926 16212
rect 7980 16156 8316 16212
rect 8372 16156 8382 16212
rect 9762 16156 9772 16212
rect 9828 16156 12236 16212
rect 12292 16156 12302 16212
rect 13906 16156 13916 16212
rect 13972 16156 15260 16212
rect 15316 16156 15326 16212
rect 15670 16156 15708 16212
rect 15764 16156 15774 16212
rect 16380 16156 24892 16212
rect 24948 16156 24958 16212
rect 16380 16100 16436 16156
rect 5842 16044 5852 16100
rect 5908 16044 5918 16100
rect 9314 16044 9324 16100
rect 9380 16044 9996 16100
rect 10052 16044 10062 16100
rect 10220 16044 16436 16100
rect 16594 16044 16604 16100
rect 16660 16044 16716 16100
rect 16772 16044 16782 16100
rect 0 15988 112 16016
rect 5852 15988 5908 16044
rect 0 15932 5908 15988
rect 8082 15932 8092 15988
rect 8148 15932 9884 15988
rect 9940 15932 9950 15988
rect 0 15904 112 15932
rect 10220 15876 10276 16044
rect 28448 15988 28560 16016
rect 10994 15932 11004 15988
rect 11060 15932 15372 15988
rect 15428 15932 15438 15988
rect 15698 15932 15708 15988
rect 15764 15932 16156 15988
rect 16212 15932 16222 15988
rect 26852 15932 28560 15988
rect 5282 15820 5292 15876
rect 5348 15820 10276 15876
rect 10770 15820 10780 15876
rect 10836 15820 12012 15876
rect 12068 15820 12348 15876
rect 12404 15820 12414 15876
rect 13570 15820 13580 15876
rect 13636 15820 14812 15876
rect 14868 15820 14878 15876
rect 16034 15820 16044 15876
rect 16100 15820 17612 15876
rect 17668 15820 17678 15876
rect 17948 15820 26348 15876
rect 26404 15820 26414 15876
rect 3462 15708 3500 15764
rect 3556 15708 3566 15764
rect 4946 15708 4956 15764
rect 5012 15708 12180 15764
rect 3794 15652 3804 15708
rect 3860 15652 3908 15708
rect 3964 15652 4012 15708
rect 4068 15652 4078 15708
rect 3574 15596 3612 15652
rect 3668 15596 3678 15652
rect 9650 15596 9660 15652
rect 9716 15596 10556 15652
rect 10612 15596 10622 15652
rect 12124 15540 12180 15708
rect 12348 15652 12404 15820
rect 15362 15708 15372 15764
rect 15428 15708 17276 15764
rect 17332 15708 17342 15764
rect 17948 15652 18004 15820
rect 23794 15652 23804 15708
rect 23860 15652 23908 15708
rect 23964 15652 24012 15708
rect 24068 15652 24078 15708
rect 12348 15596 15148 15652
rect 15204 15596 18004 15652
rect 26852 15540 26908 15932
rect 28448 15904 28560 15932
rect 28448 15540 28560 15568
rect 9090 15484 9100 15540
rect 9156 15484 11900 15540
rect 11956 15484 11966 15540
rect 12124 15484 26908 15540
rect 27906 15484 27916 15540
rect 27972 15484 28560 15540
rect 28448 15456 28560 15484
rect 7746 15372 7756 15428
rect 7812 15372 7980 15428
rect 8036 15372 8046 15428
rect 9538 15372 9548 15428
rect 9604 15372 11004 15428
rect 11060 15372 11070 15428
rect 15250 15372 15260 15428
rect 15316 15372 15932 15428
rect 15988 15372 15998 15428
rect 16454 15372 16492 15428
rect 16548 15372 16558 15428
rect 10070 15260 10108 15316
rect 10164 15260 10174 15316
rect 11330 15260 11340 15316
rect 11396 15260 11788 15316
rect 11844 15260 11854 15316
rect 15260 15260 16044 15316
rect 16100 15260 16828 15316
rect 16884 15260 16894 15316
rect 3042 15148 3052 15204
rect 3108 15148 6076 15204
rect 6132 15148 6142 15204
rect 11732 15092 11788 15260
rect 15260 15204 15316 15260
rect 14914 15148 14924 15204
rect 14980 15148 15316 15204
rect 15474 15148 15484 15204
rect 15540 15148 15932 15204
rect 15988 15148 16716 15204
rect 16772 15148 16782 15204
rect 28448 15092 28560 15120
rect 1586 15036 1596 15092
rect 1652 15036 1932 15092
rect 1988 15036 1998 15092
rect 3332 15036 4396 15092
rect 4452 15036 4462 15092
rect 10098 15036 10108 15092
rect 10164 15036 11788 15092
rect 12450 15036 12460 15092
rect 12516 15036 28560 15092
rect 3332 14980 3388 15036
rect 28448 15008 28560 15036
rect 1708 14924 3388 14980
rect 15474 14924 15484 14980
rect 15540 14924 15708 14980
rect 15764 14924 16884 14980
rect 17042 14924 17052 14980
rect 17108 14924 17500 14980
rect 17556 14924 17566 14980
rect 0 14644 112 14672
rect 1708 14644 1764 14924
rect 4454 14868 4464 14924
rect 4520 14868 4568 14924
rect 4624 14868 4672 14924
rect 4728 14868 4738 14924
rect 16828 14868 16884 14924
rect 24454 14868 24464 14924
rect 24520 14868 24568 14924
rect 24624 14868 24672 14924
rect 24728 14868 24738 14924
rect 1922 14812 1932 14868
rect 1988 14812 3052 14868
rect 3108 14812 3118 14868
rect 3378 14812 3388 14868
rect 3444 14812 3454 14868
rect 7298 14812 7308 14868
rect 7364 14812 10220 14868
rect 10276 14812 11228 14868
rect 11284 14812 11294 14868
rect 15250 14812 15260 14868
rect 15316 14812 15708 14868
rect 15764 14812 15774 14868
rect 16006 14812 16044 14868
rect 16100 14812 16110 14868
rect 16828 14812 17164 14868
rect 17220 14812 17230 14868
rect 17378 14812 17388 14868
rect 17444 14812 17948 14868
rect 18004 14812 18014 14868
rect 3388 14756 3444 14812
rect 2818 14700 2828 14756
rect 2884 14700 5628 14756
rect 5684 14700 5694 14756
rect 7634 14700 7644 14756
rect 7700 14700 9436 14756
rect 9492 14700 10724 14756
rect 15026 14700 15036 14756
rect 15092 14700 24892 14756
rect 24948 14700 24958 14756
rect 10668 14644 10724 14700
rect 28448 14644 28560 14672
rect 0 14588 1764 14644
rect 3378 14588 3388 14644
rect 3444 14588 4508 14644
rect 4564 14588 4956 14644
rect 5012 14588 5022 14644
rect 9538 14588 9548 14644
rect 9604 14588 10108 14644
rect 10164 14588 10174 14644
rect 10668 14588 15260 14644
rect 15316 14588 15326 14644
rect 15894 14588 15932 14644
rect 15988 14588 16492 14644
rect 16548 14588 16558 14644
rect 27804 14588 28560 14644
rect 0 14560 112 14588
rect 4946 14476 4956 14532
rect 5012 14476 7532 14532
rect 7588 14476 7598 14532
rect 9986 14476 9996 14532
rect 10052 14476 13244 14532
rect 13300 14476 13310 14532
rect 15138 14476 15148 14532
rect 15204 14476 16044 14532
rect 16100 14476 16110 14532
rect 16482 14476 16492 14532
rect 16548 14476 16716 14532
rect 16772 14476 16782 14532
rect 3266 14364 3276 14420
rect 3332 14364 8988 14420
rect 9044 14364 9054 14420
rect 16258 14364 16268 14420
rect 16324 14364 16828 14420
rect 16884 14364 16894 14420
rect 2902 14252 2940 14308
rect 2996 14252 3006 14308
rect 7298 14252 7308 14308
rect 7364 14252 7644 14308
rect 7700 14252 7710 14308
rect 9426 14252 9436 14308
rect 9492 14252 11004 14308
rect 11060 14252 11070 14308
rect 13878 14252 13916 14308
rect 13972 14252 18396 14308
rect 18452 14252 18462 14308
rect 16930 14140 16940 14196
rect 16996 14140 17006 14196
rect 3794 14084 3804 14140
rect 3860 14084 3908 14140
rect 3964 14084 4012 14140
rect 4068 14084 4078 14140
rect 16940 14084 16996 14140
rect 23794 14084 23804 14140
rect 23860 14084 23908 14140
rect 23964 14084 24012 14140
rect 24068 14084 24078 14140
rect 13570 14028 13580 14084
rect 13636 14028 14700 14084
rect 14756 14028 14766 14084
rect 16370 14028 16380 14084
rect 16436 14028 16996 14084
rect 2482 13916 2492 13972
rect 2548 13916 27580 13972
rect 27636 13916 27646 13972
rect 27804 13860 27860 14588
rect 28448 14560 28560 14588
rect 28448 14196 28560 14224
rect 28018 14140 28028 14196
rect 28084 14140 28560 14196
rect 28448 14112 28560 14140
rect 690 13804 700 13860
rect 756 13804 1148 13860
rect 1204 13804 4956 13860
rect 5012 13804 5292 13860
rect 5348 13804 5358 13860
rect 8642 13804 8652 13860
rect 8708 13804 27860 13860
rect 28448 13748 28560 13776
rect 5842 13692 5852 13748
rect 5908 13692 8316 13748
rect 8372 13692 8382 13748
rect 9874 13692 9884 13748
rect 9940 13692 28560 13748
rect 28448 13664 28560 13692
rect 5058 13580 5068 13636
rect 5124 13580 5292 13636
rect 5348 13580 5358 13636
rect 9762 13580 9772 13636
rect 9828 13580 10556 13636
rect 10612 13580 10622 13636
rect 10770 13580 10780 13636
rect 10836 13580 11340 13636
rect 11396 13580 11406 13636
rect 15362 13580 15372 13636
rect 15428 13580 16156 13636
rect 16212 13580 16222 13636
rect 1922 13468 1932 13524
rect 1988 13468 3052 13524
rect 3108 13468 5012 13524
rect 5842 13468 5852 13524
rect 5908 13468 6748 13524
rect 6804 13468 6814 13524
rect 14914 13468 14924 13524
rect 14980 13468 17500 13524
rect 17556 13468 17566 13524
rect 0 13300 112 13328
rect 4454 13300 4464 13356
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4728 13300 4738 13356
rect 4956 13300 5012 13468
rect 5170 13356 5180 13412
rect 5236 13356 7756 13412
rect 7812 13356 7822 13412
rect 15250 13356 15260 13412
rect 15316 13356 15820 13412
rect 15876 13356 15886 13412
rect 16678 13356 16716 13412
rect 16772 13356 16782 13412
rect 24454 13300 24464 13356
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24728 13300 24738 13356
rect 28448 13300 28560 13328
rect 0 13244 140 13300
rect 196 13244 206 13300
rect 4274 13244 4284 13300
rect 4340 13244 4350 13300
rect 4956 13244 7084 13300
rect 7140 13244 14140 13300
rect 14196 13244 14206 13300
rect 14578 13244 14588 13300
rect 14644 13244 21028 13300
rect 0 13216 112 13244
rect 4284 13188 4340 13244
rect 20972 13188 21028 13244
rect 26852 13244 28560 13300
rect 26852 13188 26908 13244
rect 28448 13216 28560 13244
rect 1138 13132 1148 13188
rect 1204 13132 2604 13188
rect 2660 13132 2670 13188
rect 4284 13132 6412 13188
rect 6468 13132 6478 13188
rect 11890 13132 11900 13188
rect 11956 13132 20356 13188
rect 20972 13132 26908 13188
rect 20300 13076 20356 13132
rect 2034 13020 2044 13076
rect 2100 13020 9212 13076
rect 9268 13020 9436 13076
rect 9492 13020 9502 13076
rect 15250 13020 15260 13076
rect 15316 13020 15354 13076
rect 20300 13020 25564 13076
rect 25620 13020 25630 13076
rect 1698 12908 1708 12964
rect 1764 12908 2156 12964
rect 2212 12908 5068 12964
rect 5124 12908 5134 12964
rect 10098 12908 10108 12964
rect 10164 12908 12236 12964
rect 12292 12908 12302 12964
rect 12786 12908 12796 12964
rect 12852 12908 25900 12964
rect 25956 12908 25966 12964
rect 28448 12852 28560 12880
rect 3378 12796 3388 12852
rect 3444 12796 4172 12852
rect 4228 12796 4238 12852
rect 6850 12796 6860 12852
rect 6916 12796 8204 12852
rect 8260 12796 9100 12852
rect 9156 12796 9166 12852
rect 15474 12796 15484 12852
rect 15540 12796 16044 12852
rect 16100 12796 16110 12852
rect 17714 12796 17724 12852
rect 17780 12796 28560 12852
rect 28448 12768 28560 12796
rect 3154 12684 3164 12740
rect 3220 12684 15148 12740
rect 16146 12684 16156 12740
rect 16212 12684 20300 12740
rect 20356 12684 20366 12740
rect 20524 12684 26572 12740
rect 26628 12684 26638 12740
rect 15092 12628 15148 12684
rect 20524 12628 20580 12684
rect 7186 12572 7196 12628
rect 7252 12572 13580 12628
rect 13636 12572 13646 12628
rect 15092 12572 20580 12628
rect 3794 12516 3804 12572
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 4068 12516 4078 12572
rect 23794 12516 23804 12572
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 24068 12516 24078 12572
rect 5954 12460 5964 12516
rect 6020 12460 20804 12516
rect 2146 12348 2156 12404
rect 2212 12348 13356 12404
rect 13412 12348 13422 12404
rect 20748 12292 20804 12460
rect 28448 12404 28560 12432
rect 26852 12348 28560 12404
rect 914 12236 924 12292
rect 980 12236 1596 12292
rect 1652 12236 1662 12292
rect 2482 12236 2492 12292
rect 2548 12236 5292 12292
rect 5348 12236 5358 12292
rect 6402 12236 6412 12292
rect 6468 12236 20692 12292
rect 20748 12236 26348 12292
rect 26404 12236 26414 12292
rect 20636 12180 20692 12236
rect 26852 12180 26908 12348
rect 28448 12320 28560 12348
rect 8530 12124 8540 12180
rect 8596 12124 9324 12180
rect 9380 12124 9390 12180
rect 12114 12124 12124 12180
rect 12180 12124 15148 12180
rect 15204 12124 16604 12180
rect 16660 12124 16670 12180
rect 20636 12124 26908 12180
rect 9874 12012 9884 12068
rect 9940 12012 10220 12068
rect 10276 12012 10780 12068
rect 10836 12012 10846 12068
rect 15026 12012 15036 12068
rect 15092 12012 16044 12068
rect 16100 12012 16492 12068
rect 16548 12012 16558 12068
rect 0 11956 112 11984
rect 28448 11956 28560 11984
rect 0 11900 1932 11956
rect 1988 11900 1998 11956
rect 2370 11900 2380 11956
rect 2436 11900 14476 11956
rect 14532 11900 14542 11956
rect 28130 11900 28140 11956
rect 28196 11900 28560 11956
rect 0 11872 112 11900
rect 28448 11872 28560 11900
rect 6178 11788 6188 11844
rect 6244 11788 10892 11844
rect 10948 11788 10958 11844
rect 12114 11788 12124 11844
rect 12180 11788 14252 11844
rect 14308 11788 14318 11844
rect 4454 11732 4464 11788
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4728 11732 4738 11788
rect 24454 11732 24464 11788
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24728 11732 24738 11788
rect 2258 11564 2268 11620
rect 2324 11564 10444 11620
rect 10500 11564 10510 11620
rect 28448 11508 28560 11536
rect 2594 11452 2604 11508
rect 2660 11452 7308 11508
rect 7364 11452 7374 11508
rect 28354 11452 28364 11508
rect 28420 11452 28560 11508
rect 28448 11424 28560 11452
rect 3490 11340 3500 11396
rect 3556 11340 4284 11396
rect 4340 11340 4350 11396
rect 4834 11340 4844 11396
rect 4900 11340 5404 11396
rect 5460 11340 6076 11396
rect 6132 11340 6142 11396
rect 8194 11340 8204 11396
rect 8260 11340 10220 11396
rect 10276 11340 10286 11396
rect 11218 11340 11228 11396
rect 11284 11340 12012 11396
rect 12068 11340 24892 11396
rect 24948 11340 24958 11396
rect 23426 11228 23436 11284
rect 23492 11228 26236 11284
rect 26292 11228 26302 11284
rect 11554 11116 11564 11172
rect 11620 11116 26908 11172
rect 26852 11060 26908 11116
rect 28448 11060 28560 11088
rect 26852 11004 28560 11060
rect 3794 10948 3804 11004
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 4068 10948 4078 11004
rect 23794 10948 23804 11004
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 24068 10948 24078 11004
rect 28448 10976 28560 11004
rect 6738 10780 6748 10836
rect 6804 10780 7980 10836
rect 8036 10780 8046 10836
rect 14018 10780 14028 10836
rect 14084 10780 17948 10836
rect 18004 10780 18014 10836
rect 5842 10668 5852 10724
rect 5908 10668 16156 10724
rect 16212 10668 16222 10724
rect 0 10612 112 10640
rect 28448 10612 28560 10640
rect 0 10556 1260 10612
rect 1316 10556 1326 10612
rect 5954 10556 5964 10612
rect 6020 10556 7084 10612
rect 7140 10556 7150 10612
rect 24994 10556 25004 10612
rect 25060 10556 28560 10612
rect 0 10528 112 10556
rect 28448 10528 28560 10556
rect 4274 10444 4284 10500
rect 4340 10444 9548 10500
rect 9604 10444 10444 10500
rect 10500 10444 10510 10500
rect 11218 10444 11228 10500
rect 11284 10444 13132 10500
rect 13188 10444 13198 10500
rect 4454 10164 4464 10220
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4728 10164 4738 10220
rect 24454 10164 24464 10220
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24728 10164 24738 10220
rect 28448 10164 28560 10192
rect 24882 10108 24892 10164
rect 24948 10108 28560 10164
rect 28448 10080 28560 10108
rect 7410 9996 7420 10052
rect 7476 9996 10892 10052
rect 10948 9996 10958 10052
rect 4722 9884 4732 9940
rect 4788 9884 17164 9940
rect 17220 9884 17230 9940
rect 9874 9772 9884 9828
rect 9940 9772 13132 9828
rect 13188 9772 15148 9828
rect 15204 9772 15214 9828
rect 28448 9716 28560 9744
rect 6962 9660 6972 9716
rect 7028 9660 11228 9716
rect 11284 9660 11294 9716
rect 16706 9660 16716 9716
rect 16772 9660 28560 9716
rect 28448 9632 28560 9660
rect 3794 9380 3804 9436
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 4068 9380 4078 9436
rect 23794 9380 23804 9436
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 24068 9380 24078 9436
rect 11666 9324 11676 9380
rect 11732 9324 22652 9380
rect 22708 9324 22718 9380
rect 0 9268 112 9296
rect 28448 9268 28560 9296
rect 0 9212 1260 9268
rect 1316 9212 1326 9268
rect 8866 9212 8876 9268
rect 8932 9212 10444 9268
rect 10500 9212 10510 9268
rect 21298 9212 21308 9268
rect 21364 9212 28560 9268
rect 0 9184 112 9212
rect 28448 9184 28560 9212
rect 7298 9100 7308 9156
rect 7364 9100 9660 9156
rect 9716 9100 9726 9156
rect 7074 8876 7084 8932
rect 7140 8876 7644 8932
rect 7700 8876 9884 8932
rect 9940 8876 9950 8932
rect 12114 8876 12124 8932
rect 12180 8876 19068 8932
rect 19124 8876 19134 8932
rect 28448 8820 28560 8848
rect 13906 8764 13916 8820
rect 13972 8764 28560 8820
rect 28448 8736 28560 8764
rect 4454 8596 4464 8652
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4728 8596 4738 8652
rect 24454 8596 24464 8652
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24728 8596 24738 8652
rect 28448 8372 28560 8400
rect 28354 8316 28364 8372
rect 28420 8316 28560 8372
rect 28448 8288 28560 8316
rect 8306 8092 8316 8148
rect 8372 8092 26124 8148
rect 26180 8092 26190 8148
rect 3332 7980 7420 8036
rect 7476 7980 7486 8036
rect 13234 7980 13244 8036
rect 13300 7980 26908 8036
rect 0 7924 112 7952
rect 3332 7924 3388 7980
rect 0 7868 3388 7924
rect 26852 7924 26908 7980
rect 28448 7924 28560 7952
rect 26852 7868 28560 7924
rect 0 7840 112 7868
rect 3794 7812 3804 7868
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 4068 7812 4078 7868
rect 23794 7812 23804 7868
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 24068 7812 24078 7868
rect 28448 7840 28560 7868
rect 28448 7476 28560 7504
rect 26338 7420 26348 7476
rect 26404 7420 28560 7476
rect 28448 7392 28560 7420
rect 10658 7308 10668 7364
rect 10724 7308 20972 7364
rect 21028 7308 21038 7364
rect 16482 7196 16492 7252
rect 16548 7196 26908 7252
rect 4454 7028 4464 7084
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4728 7028 4738 7084
rect 24454 7028 24464 7084
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 24728 7028 24738 7084
rect 26852 7028 26908 7196
rect 28448 7028 28560 7056
rect 26852 6972 28560 7028
rect 28448 6944 28560 6972
rect 0 6580 112 6608
rect 28448 6580 28560 6608
rect 0 6524 1260 6580
rect 1316 6524 1326 6580
rect 16594 6524 16604 6580
rect 16660 6524 28560 6580
rect 0 6496 112 6524
rect 28448 6496 28560 6524
rect 3794 6244 3804 6300
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 4068 6244 4078 6300
rect 23794 6244 23804 6300
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 24068 6244 24078 6300
rect 28448 6132 28560 6160
rect 15922 6076 15932 6132
rect 15988 6076 28560 6132
rect 28448 6048 28560 6076
rect 11442 5964 11452 6020
rect 11508 5964 21084 6020
rect 21140 5964 21150 6020
rect 28448 5684 28560 5712
rect 21410 5628 21420 5684
rect 21476 5628 28560 5684
rect 28448 5600 28560 5628
rect 4454 5460 4464 5516
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4728 5460 4738 5516
rect 24454 5460 24464 5516
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24728 5460 24738 5516
rect 0 5236 112 5264
rect 28448 5236 28560 5264
rect 0 5180 1260 5236
rect 1316 5180 1326 5236
rect 15250 5180 15260 5236
rect 15316 5180 28560 5236
rect 0 5152 112 5180
rect 28448 5152 28560 5180
rect 10098 5068 10108 5124
rect 10164 5068 20076 5124
rect 20132 5068 20142 5124
rect 14578 4844 14588 4900
rect 14644 4844 26908 4900
rect 26852 4788 26908 4844
rect 28448 4788 28560 4816
rect 26852 4732 28560 4788
rect 3794 4676 3804 4732
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 4068 4676 4078 4732
rect 23794 4676 23804 4732
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 24068 4676 24078 4732
rect 28448 4704 28560 4732
rect 16818 4508 16828 4564
rect 16884 4508 27020 4564
rect 27076 4508 27086 4564
rect 28448 4340 28560 4368
rect 18274 4284 18284 4340
rect 18340 4284 28560 4340
rect 28448 4256 28560 4284
rect 17826 4060 17836 4116
rect 17892 4060 26908 4116
rect 0 3892 112 3920
rect 4454 3892 4464 3948
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4728 3892 4738 3948
rect 24454 3892 24464 3948
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24728 3892 24738 3948
rect 26852 3892 26908 4060
rect 28448 3892 28560 3920
rect 0 3836 3052 3892
rect 3108 3836 3118 3892
rect 26852 3836 28560 3892
rect 0 3808 112 3836
rect 28448 3808 28560 3836
rect 14130 3612 14140 3668
rect 14196 3612 22764 3668
rect 22820 3612 22830 3668
rect 28448 3444 28560 3472
rect 22978 3388 22988 3444
rect 23044 3388 28560 3444
rect 28448 3360 28560 3388
rect 20850 3276 20860 3332
rect 20916 3276 27356 3332
rect 27412 3276 27422 3332
rect 3794 3108 3804 3164
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 4068 3108 4078 3164
rect 23794 3108 23804 3164
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 24068 3108 24078 3164
rect 7410 3052 7420 3108
rect 7476 3052 8764 3108
rect 8820 3052 8830 3108
rect 28448 2996 28560 3024
rect 13010 2940 13020 2996
rect 13076 2940 28560 2996
rect 28448 2912 28560 2940
rect 28448 2548 28560 2576
rect 13570 2492 13580 2548
rect 13636 2492 28560 2548
rect 28448 2464 28560 2492
rect 1362 2380 1372 2436
rect 1428 2380 3388 2436
rect 3444 2380 3454 2436
rect 4454 2324 4464 2380
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4728 2324 4738 2380
rect 24454 2324 24464 2380
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24728 2324 24738 2380
rect 28448 2100 28560 2128
rect 21186 2044 21196 2100
rect 21252 2044 28560 2100
rect 28448 2016 28560 2044
rect 28448 1652 28560 1680
rect 662 1596 700 1652
rect 756 1596 766 1652
rect 8754 1596 8764 1652
rect 8820 1596 12124 1652
rect 12180 1596 12190 1652
rect 12758 1596 12796 1652
rect 12852 1596 12862 1652
rect 15446 1596 15484 1652
rect 15540 1596 15550 1652
rect 24882 1596 24892 1652
rect 24948 1596 27132 1652
rect 27188 1596 27198 1652
rect 28252 1596 28560 1652
rect 3794 1540 3804 1596
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 4068 1540 4078 1596
rect 23794 1540 23804 1596
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 24068 1540 24078 1596
rect 26002 1484 26012 1540
rect 26068 1484 27580 1540
rect 27636 1484 27646 1540
rect 28252 1428 28308 1596
rect 28448 1568 28560 1596
rect 2034 1372 2044 1428
rect 2100 1372 7980 1428
rect 8036 1372 8046 1428
rect 15138 1372 15148 1428
rect 15204 1372 28308 1428
rect 22418 1260 22428 1316
rect 22484 1260 23548 1316
rect 23604 1260 23614 1316
rect 28448 1204 28560 1232
rect 20738 1148 20748 1204
rect 20804 1148 28560 1204
rect 28448 1120 28560 1148
rect 19394 924 19404 980
rect 19460 924 24948 980
rect 4454 756 4464 812
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4728 756 4738 812
rect 24454 756 24464 812
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24728 756 24738 812
rect 24892 756 24948 924
rect 28448 756 28560 784
rect 24892 700 28560 756
rect 28448 672 28560 700
rect 28448 308 28560 336
rect 22866 252 22876 308
rect 22932 252 28560 308
rect 28448 224 28560 252
rect 3602 140 3612 196
rect 3668 140 4732 196
rect 4788 140 4798 196
rect 19170 140 19180 196
rect 19236 140 19516 196
rect 19572 140 19582 196
<< via3 >>
rect 3804 56420 3860 56476
rect 3908 56420 3964 56476
rect 4012 56420 4068 56476
rect 23804 56420 23860 56476
rect 23908 56420 23964 56476
rect 24012 56420 24068 56476
rect 1708 55916 1764 55972
rect 4464 55636 4520 55692
rect 4568 55636 4624 55692
rect 4672 55636 4728 55692
rect 24464 55636 24520 55692
rect 24568 55636 24624 55692
rect 24672 55636 24728 55692
rect 3804 54852 3860 54908
rect 3908 54852 3964 54908
rect 4012 54852 4068 54908
rect 23804 54852 23860 54908
rect 23908 54852 23964 54908
rect 24012 54852 24068 54908
rect 4464 54068 4520 54124
rect 4568 54068 4624 54124
rect 4672 54068 4728 54124
rect 24464 54068 24520 54124
rect 24568 54068 24624 54124
rect 24672 54068 24728 54124
rect 3804 53284 3860 53340
rect 3908 53284 3964 53340
rect 4012 53284 4068 53340
rect 23804 53284 23860 53340
rect 23908 53284 23964 53340
rect 24012 53284 24068 53340
rect 22204 52780 22260 52836
rect 4464 52500 4520 52556
rect 4568 52500 4624 52556
rect 4672 52500 4728 52556
rect 24464 52500 24520 52556
rect 24568 52500 24624 52556
rect 24672 52500 24728 52556
rect 22204 52332 22260 52388
rect 3804 51716 3860 51772
rect 3908 51716 3964 51772
rect 4012 51716 4068 51772
rect 23804 51716 23860 51772
rect 23908 51716 23964 51772
rect 24012 51716 24068 51772
rect 16716 51212 16772 51268
rect 4464 50932 4520 50988
rect 4568 50932 4624 50988
rect 4672 50932 4728 50988
rect 24464 50932 24520 50988
rect 24568 50932 24624 50988
rect 24672 50932 24728 50988
rect 15484 50428 15540 50484
rect 3804 50148 3860 50204
rect 3908 50148 3964 50204
rect 4012 50148 4068 50204
rect 23804 50148 23860 50204
rect 23908 50148 23964 50204
rect 24012 50148 24068 50204
rect 4464 49364 4520 49420
rect 4568 49364 4624 49420
rect 4672 49364 4728 49420
rect 24464 49364 24520 49420
rect 24568 49364 24624 49420
rect 24672 49364 24728 49420
rect 3804 48580 3860 48636
rect 3908 48580 3964 48636
rect 4012 48580 4068 48636
rect 23804 48580 23860 48636
rect 23908 48580 23964 48636
rect 24012 48580 24068 48636
rect 4464 47796 4520 47852
rect 4568 47796 4624 47852
rect 4672 47796 4728 47852
rect 24464 47796 24520 47852
rect 24568 47796 24624 47852
rect 24672 47796 24728 47852
rect 3804 47012 3860 47068
rect 3908 47012 3964 47068
rect 4012 47012 4068 47068
rect 23804 47012 23860 47068
rect 23908 47012 23964 47068
rect 24012 47012 24068 47068
rect 4464 46228 4520 46284
rect 4568 46228 4624 46284
rect 4672 46228 4728 46284
rect 24464 46228 24520 46284
rect 24568 46228 24624 46284
rect 24672 46228 24728 46284
rect 26124 46060 26180 46116
rect 3804 45444 3860 45500
rect 3908 45444 3964 45500
rect 4012 45444 4068 45500
rect 23804 45444 23860 45500
rect 23908 45444 23964 45500
rect 24012 45444 24068 45500
rect 4464 44660 4520 44716
rect 4568 44660 4624 44716
rect 4672 44660 4728 44716
rect 24464 44660 24520 44716
rect 24568 44660 24624 44716
rect 24672 44660 24728 44716
rect 3804 43876 3860 43932
rect 3908 43876 3964 43932
rect 4012 43876 4068 43932
rect 23804 43876 23860 43932
rect 23908 43876 23964 43932
rect 24012 43876 24068 43932
rect 4464 43092 4520 43148
rect 4568 43092 4624 43148
rect 4672 43092 4728 43148
rect 24464 43092 24520 43148
rect 24568 43092 24624 43148
rect 24672 43092 24728 43148
rect 26124 42588 26180 42644
rect 3804 42308 3860 42364
rect 3908 42308 3964 42364
rect 4012 42308 4068 42364
rect 23804 42308 23860 42364
rect 23908 42308 23964 42364
rect 24012 42308 24068 42364
rect 4464 41524 4520 41580
rect 4568 41524 4624 41580
rect 4672 41524 4728 41580
rect 24464 41524 24520 41580
rect 24568 41524 24624 41580
rect 24672 41524 24728 41580
rect 3804 40740 3860 40796
rect 3908 40740 3964 40796
rect 4012 40740 4068 40796
rect 23804 40740 23860 40796
rect 23908 40740 23964 40796
rect 24012 40740 24068 40796
rect 4464 39956 4520 40012
rect 4568 39956 4624 40012
rect 4672 39956 4728 40012
rect 24464 39956 24520 40012
rect 24568 39956 24624 40012
rect 24672 39956 24728 40012
rect 3804 39172 3860 39228
rect 3908 39172 3964 39228
rect 4012 39172 4068 39228
rect 23804 39172 23860 39228
rect 23908 39172 23964 39228
rect 24012 39172 24068 39228
rect 11228 39004 11284 39060
rect 4464 38388 4520 38444
rect 4568 38388 4624 38444
rect 4672 38388 4728 38444
rect 24464 38388 24520 38444
rect 24568 38388 24624 38444
rect 24672 38388 24728 38444
rect 3804 37604 3860 37660
rect 3908 37604 3964 37660
rect 4012 37604 4068 37660
rect 23804 37604 23860 37660
rect 23908 37604 23964 37660
rect 24012 37604 24068 37660
rect 12796 36876 12852 36932
rect 4464 36820 4520 36876
rect 4568 36820 4624 36876
rect 4672 36820 4728 36876
rect 24464 36820 24520 36876
rect 24568 36820 24624 36876
rect 24672 36820 24728 36876
rect 4844 36652 4900 36708
rect 700 36316 756 36372
rect 3804 36036 3860 36092
rect 3908 36036 3964 36092
rect 4012 36036 4068 36092
rect 23804 36036 23860 36092
rect 23908 36036 23964 36092
rect 24012 36036 24068 36092
rect 4464 35252 4520 35308
rect 4568 35252 4624 35308
rect 4672 35252 4728 35308
rect 24464 35252 24520 35308
rect 24568 35252 24624 35308
rect 24672 35252 24728 35308
rect 12124 35196 12180 35252
rect 17948 34972 18004 35028
rect 14588 34860 14644 34916
rect 3804 34468 3860 34524
rect 3908 34468 3964 34524
rect 4012 34468 4068 34524
rect 23804 34468 23860 34524
rect 23908 34468 23964 34524
rect 24012 34468 24068 34524
rect 11900 33964 11956 34020
rect 5740 33852 5796 33908
rect 4464 33684 4520 33740
rect 4568 33684 4624 33740
rect 4672 33684 4728 33740
rect 24464 33684 24520 33740
rect 24568 33684 24624 33740
rect 24672 33684 24728 33740
rect 10892 33180 10948 33236
rect 3804 32900 3860 32956
rect 3908 32900 3964 32956
rect 4012 32900 4068 32956
rect 23804 32900 23860 32956
rect 23908 32900 23964 32956
rect 24012 32900 24068 32956
rect 4464 32116 4520 32172
rect 4568 32116 4624 32172
rect 4672 32116 4728 32172
rect 24464 32116 24520 32172
rect 24568 32116 24624 32172
rect 24672 32116 24728 32172
rect 13916 31388 13972 31444
rect 3804 31332 3860 31388
rect 3908 31332 3964 31388
rect 4012 31332 4068 31388
rect 23804 31332 23860 31388
rect 23908 31332 23964 31388
rect 24012 31332 24068 31388
rect 17948 30604 18004 30660
rect 4464 30548 4520 30604
rect 4568 30548 4624 30604
rect 4672 30548 4728 30604
rect 24464 30548 24520 30604
rect 24568 30548 24624 30604
rect 24672 30548 24728 30604
rect 3388 30268 3444 30324
rect 28364 30044 28420 30100
rect 3804 29764 3860 29820
rect 3908 29764 3964 29820
rect 4012 29764 4068 29820
rect 23804 29764 23860 29820
rect 23908 29764 23964 29820
rect 24012 29764 24068 29820
rect 12124 29596 12180 29652
rect 3500 29484 3556 29540
rect 19740 29372 19796 29428
rect 4464 28980 4520 29036
rect 4568 28980 4624 29036
rect 4672 28980 4728 29036
rect 24464 28980 24520 29036
rect 24568 28980 24624 29036
rect 24672 28980 24728 29036
rect 11900 28588 11956 28644
rect 19740 28588 19796 28644
rect 3500 28476 3556 28532
rect 3804 28196 3860 28252
rect 3908 28196 3964 28252
rect 4012 28196 4068 28252
rect 23804 28196 23860 28252
rect 23908 28196 23964 28252
rect 24012 28196 24068 28252
rect 19516 28140 19572 28196
rect 3388 28028 3444 28084
rect 25676 27916 25732 27972
rect 5740 27804 5796 27860
rect 19516 27468 19572 27524
rect 4464 27412 4520 27468
rect 4568 27412 4624 27468
rect 4672 27412 4728 27468
rect 24464 27412 24520 27468
rect 24568 27412 24624 27468
rect 24672 27412 24728 27468
rect 3804 26628 3860 26684
rect 3908 26628 3964 26684
rect 4012 26628 4068 26684
rect 23804 26628 23860 26684
rect 23908 26628 23964 26684
rect 24012 26628 24068 26684
rect 14588 26460 14644 26516
rect 4464 25844 4520 25900
rect 4568 25844 4624 25900
rect 4672 25844 4728 25900
rect 24464 25844 24520 25900
rect 24568 25844 24624 25900
rect 24672 25844 24728 25900
rect 8764 25116 8820 25172
rect 3804 25060 3860 25116
rect 3908 25060 3964 25116
rect 4012 25060 4068 25116
rect 23804 25060 23860 25116
rect 23908 25060 23964 25116
rect 24012 25060 24068 25116
rect 13916 24780 13972 24836
rect 4464 24276 4520 24332
rect 4568 24276 4624 24332
rect 4672 24276 4728 24332
rect 8764 24444 8820 24500
rect 24464 24276 24520 24332
rect 24568 24276 24624 24332
rect 24672 24276 24728 24332
rect 2044 24108 2100 24164
rect 2044 23548 2100 23604
rect 3804 23492 3860 23548
rect 3908 23492 3964 23548
rect 4012 23492 4068 23548
rect 23804 23492 23860 23548
rect 23908 23492 23964 23548
rect 24012 23492 24068 23548
rect 5516 23436 5572 23492
rect 5852 23100 5908 23156
rect 6524 23100 6580 23156
rect 4464 22708 4520 22764
rect 4568 22708 4624 22764
rect 4672 22708 4728 22764
rect 24464 22708 24520 22764
rect 24568 22708 24624 22764
rect 24672 22708 24728 22764
rect 12908 22540 12964 22596
rect 5516 21980 5572 22036
rect 3804 21924 3860 21980
rect 3908 21924 3964 21980
rect 4012 21924 4068 21980
rect 23804 21924 23860 21980
rect 23908 21924 23964 21980
rect 24012 21924 24068 21980
rect 7084 21532 7140 21588
rect 7308 21532 7364 21588
rect 25676 21308 25732 21364
rect 4464 21140 4520 21196
rect 4568 21140 4624 21196
rect 4672 21140 4728 21196
rect 24464 21140 24520 21196
rect 24568 21140 24624 21196
rect 24672 21140 24728 21196
rect 15820 21084 15876 21140
rect 28028 20972 28084 21028
rect 1708 20860 1764 20916
rect 15820 20524 15876 20580
rect 12908 20412 12964 20468
rect 3804 20356 3860 20412
rect 3908 20356 3964 20412
rect 4012 20356 4068 20412
rect 23804 20356 23860 20412
rect 23908 20356 23964 20412
rect 24012 20356 24068 20412
rect 27916 20188 27972 20244
rect 4464 19572 4520 19628
rect 4568 19572 4624 19628
rect 4672 19572 4728 19628
rect 24464 19572 24520 19628
rect 24568 19572 24624 19628
rect 24672 19572 24728 19628
rect 24892 19516 24948 19572
rect 2940 18956 2996 19012
rect 3804 18788 3860 18844
rect 3908 18788 3964 18844
rect 4012 18788 4068 18844
rect 23804 18788 23860 18844
rect 23908 18788 23964 18844
rect 24012 18788 24068 18844
rect 15148 18620 15204 18676
rect 27916 18620 27972 18676
rect 6524 18508 6580 18564
rect 14364 18396 14420 18452
rect 4464 18004 4520 18060
rect 4568 18004 4624 18060
rect 4672 18004 4728 18060
rect 5852 17836 5908 17892
rect 28364 18172 28420 18228
rect 24464 18004 24520 18060
rect 24568 18004 24624 18060
rect 24672 18004 24728 18060
rect 16716 17724 16772 17780
rect 11340 17388 11396 17444
rect 3612 17276 3668 17332
rect 3804 17220 3860 17276
rect 3908 17220 3964 17276
rect 4012 17220 4068 17276
rect 23804 17220 23860 17276
rect 23908 17220 23964 17276
rect 24012 17220 24068 17276
rect 3500 17052 3556 17108
rect 13916 16716 13972 16772
rect 4956 16604 5012 16660
rect 14364 16604 14420 16660
rect 4464 16436 4520 16492
rect 4568 16436 4624 16492
rect 4672 16436 4728 16492
rect 24464 16436 24520 16492
rect 24568 16436 24624 16492
rect 24672 16436 24728 16492
rect 4844 16268 4900 16324
rect 15708 16156 15764 16212
rect 24892 16156 24948 16212
rect 16716 16044 16772 16100
rect 26348 15820 26404 15876
rect 3500 15708 3556 15764
rect 3804 15652 3860 15708
rect 3908 15652 3964 15708
rect 4012 15652 4068 15708
rect 3612 15596 3668 15652
rect 23804 15652 23860 15708
rect 23908 15652 23964 15708
rect 24012 15652 24068 15708
rect 16492 15372 16548 15428
rect 10108 15260 10164 15316
rect 15932 15148 15988 15204
rect 10108 15036 10164 15092
rect 15708 14924 15764 14980
rect 4464 14868 4520 14924
rect 4568 14868 4624 14924
rect 4672 14868 4728 14924
rect 24464 14868 24520 14924
rect 24568 14868 24624 14924
rect 24672 14868 24728 14924
rect 16044 14812 16100 14868
rect 15260 14588 15316 14644
rect 15932 14588 15988 14644
rect 4956 14476 5012 14532
rect 16492 14476 16548 14532
rect 2940 14252 2996 14308
rect 7308 14252 7364 14308
rect 13916 14252 13972 14308
rect 3804 14084 3860 14140
rect 3908 14084 3964 14140
rect 4012 14084 4068 14140
rect 23804 14084 23860 14140
rect 23908 14084 23964 14140
rect 24012 14084 24068 14140
rect 28028 14140 28084 14196
rect 11340 13580 11396 13636
rect 4464 13300 4520 13356
rect 4568 13300 4624 13356
rect 4672 13300 4728 13356
rect 16716 13356 16772 13412
rect 24464 13300 24520 13356
rect 24568 13300 24624 13356
rect 24672 13300 24728 13356
rect 7084 13244 7140 13300
rect 15260 13020 15316 13076
rect 3804 12516 3860 12572
rect 3908 12516 3964 12572
rect 4012 12516 4068 12572
rect 23804 12516 23860 12572
rect 23908 12516 23964 12572
rect 24012 12516 24068 12572
rect 16044 12012 16100 12068
rect 10892 11788 10948 11844
rect 4464 11732 4520 11788
rect 4568 11732 4624 11788
rect 4672 11732 4728 11788
rect 24464 11732 24520 11788
rect 24568 11732 24624 11788
rect 24672 11732 24728 11788
rect 24892 11340 24948 11396
rect 3804 10948 3860 11004
rect 3908 10948 3964 11004
rect 4012 10948 4068 11004
rect 23804 10948 23860 11004
rect 23908 10948 23964 11004
rect 24012 10948 24068 11004
rect 4464 10164 4520 10220
rect 4568 10164 4624 10220
rect 4672 10164 4728 10220
rect 24464 10164 24520 10220
rect 24568 10164 24624 10220
rect 24672 10164 24728 10220
rect 24892 10108 24948 10164
rect 11228 9660 11284 9716
rect 3804 9380 3860 9436
rect 3908 9380 3964 9436
rect 4012 9380 4068 9436
rect 23804 9380 23860 9436
rect 23908 9380 23964 9436
rect 24012 9380 24068 9436
rect 4464 8596 4520 8652
rect 4568 8596 4624 8652
rect 4672 8596 4728 8652
rect 24464 8596 24520 8652
rect 24568 8596 24624 8652
rect 24672 8596 24728 8652
rect 3804 7812 3860 7868
rect 3908 7812 3964 7868
rect 4012 7812 4068 7868
rect 23804 7812 23860 7868
rect 23908 7812 23964 7868
rect 24012 7812 24068 7868
rect 26348 7420 26404 7476
rect 4464 7028 4520 7084
rect 4568 7028 4624 7084
rect 4672 7028 4728 7084
rect 24464 7028 24520 7084
rect 24568 7028 24624 7084
rect 24672 7028 24728 7084
rect 3804 6244 3860 6300
rect 3908 6244 3964 6300
rect 4012 6244 4068 6300
rect 23804 6244 23860 6300
rect 23908 6244 23964 6300
rect 24012 6244 24068 6300
rect 4464 5460 4520 5516
rect 4568 5460 4624 5516
rect 4672 5460 4728 5516
rect 24464 5460 24520 5516
rect 24568 5460 24624 5516
rect 24672 5460 24728 5516
rect 3804 4676 3860 4732
rect 3908 4676 3964 4732
rect 4012 4676 4068 4732
rect 23804 4676 23860 4732
rect 23908 4676 23964 4732
rect 24012 4676 24068 4732
rect 4464 3892 4520 3948
rect 4568 3892 4624 3948
rect 4672 3892 4728 3948
rect 24464 3892 24520 3948
rect 24568 3892 24624 3948
rect 24672 3892 24728 3948
rect 3804 3108 3860 3164
rect 3908 3108 3964 3164
rect 4012 3108 4068 3164
rect 23804 3108 23860 3164
rect 23908 3108 23964 3164
rect 24012 3108 24068 3164
rect 4464 2324 4520 2380
rect 4568 2324 4624 2380
rect 4672 2324 4728 2380
rect 24464 2324 24520 2380
rect 24568 2324 24624 2380
rect 24672 2324 24728 2380
rect 700 1596 756 1652
rect 12796 1596 12852 1652
rect 15484 1596 15540 1652
rect 3804 1540 3860 1596
rect 3908 1540 3964 1596
rect 4012 1540 4068 1596
rect 23804 1540 23860 1596
rect 23908 1540 23964 1596
rect 24012 1540 24068 1596
rect 4464 756 4520 812
rect 4568 756 4624 812
rect 4672 756 4728 812
rect 24464 756 24520 812
rect 24568 756 24624 812
rect 24672 756 24728 812
<< metal4 >>
rect 3776 56476 4096 57456
rect 3776 56420 3804 56476
rect 3860 56420 3908 56476
rect 3964 56420 4012 56476
rect 4068 56420 4096 56476
rect 1708 55972 1764 55982
rect 700 36372 756 36382
rect 700 1652 756 36316
rect 1708 20916 1764 55916
rect 3776 54908 4096 56420
rect 3776 54852 3804 54908
rect 3860 54852 3908 54908
rect 3964 54852 4012 54908
rect 4068 54852 4096 54908
rect 3776 53340 4096 54852
rect 3776 53284 3804 53340
rect 3860 53284 3908 53340
rect 3964 53284 4012 53340
rect 4068 53284 4096 53340
rect 3776 51772 4096 53284
rect 3776 51716 3804 51772
rect 3860 51716 3908 51772
rect 3964 51716 4012 51772
rect 4068 51716 4096 51772
rect 3776 50204 4096 51716
rect 3776 50148 3804 50204
rect 3860 50148 3908 50204
rect 3964 50148 4012 50204
rect 4068 50148 4096 50204
rect 3776 48636 4096 50148
rect 3776 48580 3804 48636
rect 3860 48580 3908 48636
rect 3964 48580 4012 48636
rect 4068 48580 4096 48636
rect 3776 47068 4096 48580
rect 3776 47012 3804 47068
rect 3860 47012 3908 47068
rect 3964 47012 4012 47068
rect 4068 47012 4096 47068
rect 3776 45500 4096 47012
rect 3776 45444 3804 45500
rect 3860 45444 3908 45500
rect 3964 45444 4012 45500
rect 4068 45444 4096 45500
rect 3776 43932 4096 45444
rect 3776 43876 3804 43932
rect 3860 43876 3908 43932
rect 3964 43876 4012 43932
rect 4068 43876 4096 43932
rect 3776 42364 4096 43876
rect 3776 42308 3804 42364
rect 3860 42308 3908 42364
rect 3964 42308 4012 42364
rect 4068 42308 4096 42364
rect 3776 40796 4096 42308
rect 3776 40740 3804 40796
rect 3860 40740 3908 40796
rect 3964 40740 4012 40796
rect 4068 40740 4096 40796
rect 3776 39228 4096 40740
rect 3776 39172 3804 39228
rect 3860 39172 3908 39228
rect 3964 39172 4012 39228
rect 4068 39172 4096 39228
rect 3776 37660 4096 39172
rect 3776 37604 3804 37660
rect 3860 37604 3908 37660
rect 3964 37604 4012 37660
rect 4068 37604 4096 37660
rect 3776 36092 4096 37604
rect 3776 36036 3804 36092
rect 3860 36036 3908 36092
rect 3964 36036 4012 36092
rect 4068 36036 4096 36092
rect 3776 34524 4096 36036
rect 3776 34468 3804 34524
rect 3860 34468 3908 34524
rect 3964 34468 4012 34524
rect 4068 34468 4096 34524
rect 3776 32956 4096 34468
rect 3776 32900 3804 32956
rect 3860 32900 3908 32956
rect 3964 32900 4012 32956
rect 4068 32900 4096 32956
rect 3776 31388 4096 32900
rect 3776 31332 3804 31388
rect 3860 31332 3908 31388
rect 3964 31332 4012 31388
rect 4068 31332 4096 31388
rect 3388 30324 3444 30334
rect 3388 28084 3444 30268
rect 3776 29820 4096 31332
rect 3776 29764 3804 29820
rect 3860 29764 3908 29820
rect 3964 29764 4012 29820
rect 4068 29764 4096 29820
rect 3500 29540 3556 29550
rect 3500 28532 3556 29484
rect 3500 28466 3556 28476
rect 3388 28018 3444 28028
rect 3776 28252 4096 29764
rect 3776 28196 3804 28252
rect 3860 28196 3908 28252
rect 3964 28196 4012 28252
rect 4068 28196 4096 28252
rect 3776 26684 4096 28196
rect 3776 26628 3804 26684
rect 3860 26628 3908 26684
rect 3964 26628 4012 26684
rect 4068 26628 4096 26684
rect 3776 25116 4096 26628
rect 3776 25060 3804 25116
rect 3860 25060 3908 25116
rect 3964 25060 4012 25116
rect 4068 25060 4096 25116
rect 2044 24164 2100 24174
rect 2044 23604 2100 24108
rect 2044 23538 2100 23548
rect 3776 23548 4096 25060
rect 1708 20850 1764 20860
rect 3776 23492 3804 23548
rect 3860 23492 3908 23548
rect 3964 23492 4012 23548
rect 4068 23492 4096 23548
rect 3776 21980 4096 23492
rect 3776 21924 3804 21980
rect 3860 21924 3908 21980
rect 3964 21924 4012 21980
rect 4068 21924 4096 21980
rect 3776 20412 4096 21924
rect 3776 20356 3804 20412
rect 3860 20356 3908 20412
rect 3964 20356 4012 20412
rect 4068 20356 4096 20412
rect 2940 19012 2996 19022
rect 2940 14308 2996 18956
rect 3776 18844 4096 20356
rect 3776 18788 3804 18844
rect 3860 18788 3908 18844
rect 3964 18788 4012 18844
rect 4068 18788 4096 18844
rect 3612 17332 3668 17342
rect 3500 17108 3556 17118
rect 3500 15764 3556 17052
rect 3500 15698 3556 15708
rect 3612 15652 3668 17276
rect 3612 15586 3668 15596
rect 3776 17276 4096 18788
rect 3776 17220 3804 17276
rect 3860 17220 3908 17276
rect 3964 17220 4012 17276
rect 4068 17220 4096 17276
rect 3776 15708 4096 17220
rect 3776 15652 3804 15708
rect 3860 15652 3908 15708
rect 3964 15652 4012 15708
rect 4068 15652 4096 15708
rect 2940 14242 2996 14252
rect 700 1586 756 1596
rect 3776 14140 4096 15652
rect 3776 14084 3804 14140
rect 3860 14084 3908 14140
rect 3964 14084 4012 14140
rect 4068 14084 4096 14140
rect 3776 12572 4096 14084
rect 3776 12516 3804 12572
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 4068 12516 4096 12572
rect 3776 11004 4096 12516
rect 3776 10948 3804 11004
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 4068 10948 4096 11004
rect 3776 9436 4096 10948
rect 3776 9380 3804 9436
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 4068 9380 4096 9436
rect 3776 7868 4096 9380
rect 3776 7812 3804 7868
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 4068 7812 4096 7868
rect 3776 6300 4096 7812
rect 3776 6244 3804 6300
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 4068 6244 4096 6300
rect 3776 4732 4096 6244
rect 3776 4676 3804 4732
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 4068 4676 4096 4732
rect 3776 3164 4096 4676
rect 3776 3108 3804 3164
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 4068 3108 4096 3164
rect 3776 1596 4096 3108
rect 3776 1540 3804 1596
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 4068 1540 4096 1596
rect 3776 0 4096 1540
rect 4436 55692 4756 57456
rect 4436 55636 4464 55692
rect 4520 55636 4568 55692
rect 4624 55636 4672 55692
rect 4728 55636 4756 55692
rect 4436 54124 4756 55636
rect 4436 54068 4464 54124
rect 4520 54068 4568 54124
rect 4624 54068 4672 54124
rect 4728 54068 4756 54124
rect 4436 52556 4756 54068
rect 23776 56476 24096 57456
rect 23776 56420 23804 56476
rect 23860 56420 23908 56476
rect 23964 56420 24012 56476
rect 24068 56420 24096 56476
rect 23776 54908 24096 56420
rect 23776 54852 23804 54908
rect 23860 54852 23908 54908
rect 23964 54852 24012 54908
rect 24068 54852 24096 54908
rect 23776 53340 24096 54852
rect 23776 53284 23804 53340
rect 23860 53284 23908 53340
rect 23964 53284 24012 53340
rect 24068 53284 24096 53340
rect 4436 52500 4464 52556
rect 4520 52500 4568 52556
rect 4624 52500 4672 52556
rect 4728 52500 4756 52556
rect 4436 50988 4756 52500
rect 22204 52836 22260 52846
rect 22204 52388 22260 52780
rect 22204 52322 22260 52332
rect 23776 51772 24096 53284
rect 23776 51716 23804 51772
rect 23860 51716 23908 51772
rect 23964 51716 24012 51772
rect 24068 51716 24096 51772
rect 4436 50932 4464 50988
rect 4520 50932 4568 50988
rect 4624 50932 4672 50988
rect 4728 50932 4756 50988
rect 4436 49420 4756 50932
rect 16716 51268 16772 51278
rect 4436 49364 4464 49420
rect 4520 49364 4568 49420
rect 4624 49364 4672 49420
rect 4728 49364 4756 49420
rect 4436 47852 4756 49364
rect 4436 47796 4464 47852
rect 4520 47796 4568 47852
rect 4624 47796 4672 47852
rect 4728 47796 4756 47852
rect 4436 46284 4756 47796
rect 4436 46228 4464 46284
rect 4520 46228 4568 46284
rect 4624 46228 4672 46284
rect 4728 46228 4756 46284
rect 4436 44716 4756 46228
rect 4436 44660 4464 44716
rect 4520 44660 4568 44716
rect 4624 44660 4672 44716
rect 4728 44660 4756 44716
rect 4436 43148 4756 44660
rect 4436 43092 4464 43148
rect 4520 43092 4568 43148
rect 4624 43092 4672 43148
rect 4728 43092 4756 43148
rect 4436 41580 4756 43092
rect 4436 41524 4464 41580
rect 4520 41524 4568 41580
rect 4624 41524 4672 41580
rect 4728 41524 4756 41580
rect 4436 40012 4756 41524
rect 4436 39956 4464 40012
rect 4520 39956 4568 40012
rect 4624 39956 4672 40012
rect 4728 39956 4756 40012
rect 4436 38444 4756 39956
rect 15484 50484 15540 50494
rect 4436 38388 4464 38444
rect 4520 38388 4568 38444
rect 4624 38388 4672 38444
rect 4728 38388 4756 38444
rect 4436 36876 4756 38388
rect 4436 36820 4464 36876
rect 4520 36820 4568 36876
rect 4624 36820 4672 36876
rect 4728 36820 4756 36876
rect 4436 35308 4756 36820
rect 11228 39060 11284 39070
rect 4436 35252 4464 35308
rect 4520 35252 4568 35308
rect 4624 35252 4672 35308
rect 4728 35252 4756 35308
rect 4436 33740 4756 35252
rect 4436 33684 4464 33740
rect 4520 33684 4568 33740
rect 4624 33684 4672 33740
rect 4728 33684 4756 33740
rect 4436 32172 4756 33684
rect 4436 32116 4464 32172
rect 4520 32116 4568 32172
rect 4624 32116 4672 32172
rect 4728 32116 4756 32172
rect 4436 30604 4756 32116
rect 4436 30548 4464 30604
rect 4520 30548 4568 30604
rect 4624 30548 4672 30604
rect 4728 30548 4756 30604
rect 4436 29036 4756 30548
rect 4436 28980 4464 29036
rect 4520 28980 4568 29036
rect 4624 28980 4672 29036
rect 4728 28980 4756 29036
rect 4436 27468 4756 28980
rect 4436 27412 4464 27468
rect 4520 27412 4568 27468
rect 4624 27412 4672 27468
rect 4728 27412 4756 27468
rect 4436 25900 4756 27412
rect 4436 25844 4464 25900
rect 4520 25844 4568 25900
rect 4624 25844 4672 25900
rect 4728 25844 4756 25900
rect 4436 24332 4756 25844
rect 4436 24276 4464 24332
rect 4520 24276 4568 24332
rect 4624 24276 4672 24332
rect 4728 24276 4756 24332
rect 4436 22764 4756 24276
rect 4436 22708 4464 22764
rect 4520 22708 4568 22764
rect 4624 22708 4672 22764
rect 4728 22708 4756 22764
rect 4436 21196 4756 22708
rect 4436 21140 4464 21196
rect 4520 21140 4568 21196
rect 4624 21140 4672 21196
rect 4728 21140 4756 21196
rect 4436 19628 4756 21140
rect 4436 19572 4464 19628
rect 4520 19572 4568 19628
rect 4624 19572 4672 19628
rect 4728 19572 4756 19628
rect 4436 18060 4756 19572
rect 4436 18004 4464 18060
rect 4520 18004 4568 18060
rect 4624 18004 4672 18060
rect 4728 18004 4756 18060
rect 4436 16492 4756 18004
rect 4436 16436 4464 16492
rect 4520 16436 4568 16492
rect 4624 16436 4672 16492
rect 4728 16436 4756 16492
rect 4436 14924 4756 16436
rect 4844 36708 4900 36718
rect 4844 16324 4900 36652
rect 5740 33908 5796 33918
rect 5740 27860 5796 33852
rect 5740 27794 5796 27804
rect 10892 33236 10948 33246
rect 8764 25172 8820 25182
rect 8764 24500 8820 25116
rect 8764 24434 8820 24444
rect 5516 23492 5572 23502
rect 5516 22036 5572 23436
rect 5516 21970 5572 21980
rect 5852 23156 5908 23166
rect 5852 17892 5908 23100
rect 6524 23156 6580 23166
rect 6524 18564 6580 23100
rect 6524 18498 6580 18508
rect 7084 21588 7140 21598
rect 5852 17826 5908 17836
rect 4844 16258 4900 16268
rect 4956 16660 5012 16670
rect 4436 14868 4464 14924
rect 4520 14868 4568 14924
rect 4624 14868 4672 14924
rect 4728 14868 4756 14924
rect 4436 13356 4756 14868
rect 4956 14532 5012 16604
rect 4956 14466 5012 14476
rect 4436 13300 4464 13356
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4728 13300 4756 13356
rect 4436 11788 4756 13300
rect 7084 13300 7140 21532
rect 7308 21588 7364 21598
rect 7308 14308 7364 21532
rect 10108 15316 10164 15326
rect 10108 15092 10164 15260
rect 10108 15026 10164 15036
rect 7308 14242 7364 14252
rect 7084 13234 7140 13244
rect 4436 11732 4464 11788
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4728 11732 4756 11788
rect 10892 11844 10948 33180
rect 10892 11778 10948 11788
rect 4436 10220 4756 11732
rect 4436 10164 4464 10220
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4728 10164 4756 10220
rect 4436 8652 4756 10164
rect 11228 9716 11284 39004
rect 12796 36932 12852 36942
rect 12124 35252 12180 35262
rect 11900 34020 11956 34030
rect 11900 28644 11956 33964
rect 12124 29652 12180 35196
rect 12124 29586 12180 29596
rect 11900 28578 11956 28588
rect 11340 17444 11396 17454
rect 11340 13636 11396 17388
rect 11340 13570 11396 13580
rect 11228 9650 11284 9660
rect 4436 8596 4464 8652
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4728 8596 4756 8652
rect 4436 7084 4756 8596
rect 4436 7028 4464 7084
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4728 7028 4756 7084
rect 4436 5516 4756 7028
rect 4436 5460 4464 5516
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4728 5460 4756 5516
rect 4436 3948 4756 5460
rect 4436 3892 4464 3948
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4728 3892 4756 3948
rect 4436 2380 4756 3892
rect 4436 2324 4464 2380
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4728 2324 4756 2380
rect 4436 812 4756 2324
rect 12796 1652 12852 36876
rect 14588 34916 14644 34926
rect 13916 31444 13972 31454
rect 13916 24836 13972 31388
rect 14588 26516 14644 34860
rect 14588 26450 14644 26460
rect 13916 24770 13972 24780
rect 12908 22596 12964 22606
rect 12908 20468 12964 22540
rect 12908 20402 12964 20412
rect 15148 18676 15204 18686
rect 15204 18620 15316 18658
rect 15148 18602 15316 18620
rect 14364 18452 14420 18462
rect 13916 16772 13972 16782
rect 13916 14308 13972 16716
rect 14364 16660 14420 18396
rect 14364 16594 14420 16604
rect 13916 14242 13972 14252
rect 15260 14644 15316 18602
rect 15260 13076 15316 14588
rect 15260 13010 15316 13020
rect 12796 1586 12852 1596
rect 15484 1652 15540 50428
rect 15820 21140 15876 21150
rect 15820 20580 15876 21084
rect 15820 20514 15876 20524
rect 16716 17780 16772 51212
rect 23776 50204 24096 51716
rect 23776 50148 23804 50204
rect 23860 50148 23908 50204
rect 23964 50148 24012 50204
rect 24068 50148 24096 50204
rect 23776 48636 24096 50148
rect 23776 48580 23804 48636
rect 23860 48580 23908 48636
rect 23964 48580 24012 48636
rect 24068 48580 24096 48636
rect 23776 47068 24096 48580
rect 23776 47012 23804 47068
rect 23860 47012 23908 47068
rect 23964 47012 24012 47068
rect 24068 47012 24096 47068
rect 23776 45500 24096 47012
rect 23776 45444 23804 45500
rect 23860 45444 23908 45500
rect 23964 45444 24012 45500
rect 24068 45444 24096 45500
rect 23776 43932 24096 45444
rect 23776 43876 23804 43932
rect 23860 43876 23908 43932
rect 23964 43876 24012 43932
rect 24068 43876 24096 43932
rect 23776 42364 24096 43876
rect 23776 42308 23804 42364
rect 23860 42308 23908 42364
rect 23964 42308 24012 42364
rect 24068 42308 24096 42364
rect 23776 40796 24096 42308
rect 23776 40740 23804 40796
rect 23860 40740 23908 40796
rect 23964 40740 24012 40796
rect 24068 40740 24096 40796
rect 23776 39228 24096 40740
rect 23776 39172 23804 39228
rect 23860 39172 23908 39228
rect 23964 39172 24012 39228
rect 24068 39172 24096 39228
rect 23776 37660 24096 39172
rect 23776 37604 23804 37660
rect 23860 37604 23908 37660
rect 23964 37604 24012 37660
rect 24068 37604 24096 37660
rect 23776 36092 24096 37604
rect 23776 36036 23804 36092
rect 23860 36036 23908 36092
rect 23964 36036 24012 36092
rect 24068 36036 24096 36092
rect 17948 35028 18004 35038
rect 17948 30660 18004 34972
rect 17948 30594 18004 30604
rect 23776 34524 24096 36036
rect 23776 34468 23804 34524
rect 23860 34468 23908 34524
rect 23964 34468 24012 34524
rect 24068 34468 24096 34524
rect 23776 32956 24096 34468
rect 23776 32900 23804 32956
rect 23860 32900 23908 32956
rect 23964 32900 24012 32956
rect 24068 32900 24096 32956
rect 23776 31388 24096 32900
rect 23776 31332 23804 31388
rect 23860 31332 23908 31388
rect 23964 31332 24012 31388
rect 24068 31332 24096 31388
rect 23776 29820 24096 31332
rect 23776 29764 23804 29820
rect 23860 29764 23908 29820
rect 23964 29764 24012 29820
rect 24068 29764 24096 29820
rect 19740 29428 19796 29438
rect 19740 28644 19796 29372
rect 19740 28578 19796 28588
rect 23776 28252 24096 29764
rect 19516 28196 19572 28206
rect 19516 27524 19572 28140
rect 19516 27458 19572 27468
rect 23776 28196 23804 28252
rect 23860 28196 23908 28252
rect 23964 28196 24012 28252
rect 24068 28196 24096 28252
rect 16716 17714 16772 17724
rect 23776 26684 24096 28196
rect 23776 26628 23804 26684
rect 23860 26628 23908 26684
rect 23964 26628 24012 26684
rect 24068 26628 24096 26684
rect 23776 25116 24096 26628
rect 23776 25060 23804 25116
rect 23860 25060 23908 25116
rect 23964 25060 24012 25116
rect 24068 25060 24096 25116
rect 23776 23548 24096 25060
rect 23776 23492 23804 23548
rect 23860 23492 23908 23548
rect 23964 23492 24012 23548
rect 24068 23492 24096 23548
rect 23776 21980 24096 23492
rect 23776 21924 23804 21980
rect 23860 21924 23908 21980
rect 23964 21924 24012 21980
rect 24068 21924 24096 21980
rect 23776 20412 24096 21924
rect 23776 20356 23804 20412
rect 23860 20356 23908 20412
rect 23964 20356 24012 20412
rect 24068 20356 24096 20412
rect 23776 18844 24096 20356
rect 23776 18788 23804 18844
rect 23860 18788 23908 18844
rect 23964 18788 24012 18844
rect 24068 18788 24096 18844
rect 23776 17276 24096 18788
rect 23776 17220 23804 17276
rect 23860 17220 23908 17276
rect 23964 17220 24012 17276
rect 24068 17220 24096 17276
rect 15708 16212 15764 16222
rect 15708 14980 15764 16156
rect 16716 16100 16772 16110
rect 16492 15428 16548 15438
rect 15708 14914 15764 14924
rect 15932 15204 15988 15214
rect 15932 14644 15988 15148
rect 15932 14578 15988 14588
rect 16044 14868 16100 14878
rect 16044 12068 16100 14812
rect 16492 14532 16548 15372
rect 16492 14466 16548 14476
rect 16716 13412 16772 16044
rect 16716 13346 16772 13356
rect 23776 15708 24096 17220
rect 23776 15652 23804 15708
rect 23860 15652 23908 15708
rect 23964 15652 24012 15708
rect 24068 15652 24096 15708
rect 23776 14140 24096 15652
rect 23776 14084 23804 14140
rect 23860 14084 23908 14140
rect 23964 14084 24012 14140
rect 24068 14084 24096 14140
rect 16044 12002 16100 12012
rect 23776 12572 24096 14084
rect 23776 12516 23804 12572
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 24068 12516 24096 12572
rect 15484 1586 15540 1596
rect 23776 11004 24096 12516
rect 23776 10948 23804 11004
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 24068 10948 24096 11004
rect 23776 9436 24096 10948
rect 23776 9380 23804 9436
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 24068 9380 24096 9436
rect 23776 7868 24096 9380
rect 23776 7812 23804 7868
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 24068 7812 24096 7868
rect 23776 6300 24096 7812
rect 23776 6244 23804 6300
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 24068 6244 24096 6300
rect 23776 4732 24096 6244
rect 23776 4676 23804 4732
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 24068 4676 24096 4732
rect 23776 3164 24096 4676
rect 23776 3108 23804 3164
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 24068 3108 24096 3164
rect 23776 1596 24096 3108
rect 4436 756 4464 812
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4728 756 4756 812
rect 4436 0 4756 756
rect 23776 1540 23804 1596
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 24068 1540 24096 1596
rect 23776 0 24096 1540
rect 24436 55692 24756 57456
rect 24436 55636 24464 55692
rect 24520 55636 24568 55692
rect 24624 55636 24672 55692
rect 24728 55636 24756 55692
rect 24436 54124 24756 55636
rect 24436 54068 24464 54124
rect 24520 54068 24568 54124
rect 24624 54068 24672 54124
rect 24728 54068 24756 54124
rect 24436 52556 24756 54068
rect 24436 52500 24464 52556
rect 24520 52500 24568 52556
rect 24624 52500 24672 52556
rect 24728 52500 24756 52556
rect 24436 50988 24756 52500
rect 24436 50932 24464 50988
rect 24520 50932 24568 50988
rect 24624 50932 24672 50988
rect 24728 50932 24756 50988
rect 24436 49420 24756 50932
rect 24436 49364 24464 49420
rect 24520 49364 24568 49420
rect 24624 49364 24672 49420
rect 24728 49364 24756 49420
rect 24436 47852 24756 49364
rect 24436 47796 24464 47852
rect 24520 47796 24568 47852
rect 24624 47796 24672 47852
rect 24728 47796 24756 47852
rect 24436 46284 24756 47796
rect 24436 46228 24464 46284
rect 24520 46228 24568 46284
rect 24624 46228 24672 46284
rect 24728 46228 24756 46284
rect 24436 44716 24756 46228
rect 24436 44660 24464 44716
rect 24520 44660 24568 44716
rect 24624 44660 24672 44716
rect 24728 44660 24756 44716
rect 24436 43148 24756 44660
rect 24436 43092 24464 43148
rect 24520 43092 24568 43148
rect 24624 43092 24672 43148
rect 24728 43092 24756 43148
rect 24436 41580 24756 43092
rect 26124 46116 26180 46126
rect 26124 42644 26180 46060
rect 26124 42578 26180 42588
rect 24436 41524 24464 41580
rect 24520 41524 24568 41580
rect 24624 41524 24672 41580
rect 24728 41524 24756 41580
rect 24436 40012 24756 41524
rect 24436 39956 24464 40012
rect 24520 39956 24568 40012
rect 24624 39956 24672 40012
rect 24728 39956 24756 40012
rect 24436 38444 24756 39956
rect 24436 38388 24464 38444
rect 24520 38388 24568 38444
rect 24624 38388 24672 38444
rect 24728 38388 24756 38444
rect 24436 36876 24756 38388
rect 24436 36820 24464 36876
rect 24520 36820 24568 36876
rect 24624 36820 24672 36876
rect 24728 36820 24756 36876
rect 24436 35308 24756 36820
rect 24436 35252 24464 35308
rect 24520 35252 24568 35308
rect 24624 35252 24672 35308
rect 24728 35252 24756 35308
rect 24436 33740 24756 35252
rect 24436 33684 24464 33740
rect 24520 33684 24568 33740
rect 24624 33684 24672 33740
rect 24728 33684 24756 33740
rect 24436 32172 24756 33684
rect 24436 32116 24464 32172
rect 24520 32116 24568 32172
rect 24624 32116 24672 32172
rect 24728 32116 24756 32172
rect 24436 30604 24756 32116
rect 24436 30548 24464 30604
rect 24520 30548 24568 30604
rect 24624 30548 24672 30604
rect 24728 30548 24756 30604
rect 24436 29036 24756 30548
rect 24436 28980 24464 29036
rect 24520 28980 24568 29036
rect 24624 28980 24672 29036
rect 24728 28980 24756 29036
rect 24436 27468 24756 28980
rect 28364 30100 28420 30110
rect 24436 27412 24464 27468
rect 24520 27412 24568 27468
rect 24624 27412 24672 27468
rect 24728 27412 24756 27468
rect 24436 25900 24756 27412
rect 24436 25844 24464 25900
rect 24520 25844 24568 25900
rect 24624 25844 24672 25900
rect 24728 25844 24756 25900
rect 24436 24332 24756 25844
rect 24436 24276 24464 24332
rect 24520 24276 24568 24332
rect 24624 24276 24672 24332
rect 24728 24276 24756 24332
rect 24436 22764 24756 24276
rect 24436 22708 24464 22764
rect 24520 22708 24568 22764
rect 24624 22708 24672 22764
rect 24728 22708 24756 22764
rect 24436 21196 24756 22708
rect 25676 27972 25732 27982
rect 25676 21364 25732 27916
rect 25676 21298 25732 21308
rect 24436 21140 24464 21196
rect 24520 21140 24568 21196
rect 24624 21140 24672 21196
rect 24728 21140 24756 21196
rect 24436 19628 24756 21140
rect 28028 21028 28084 21038
rect 24436 19572 24464 19628
rect 24520 19572 24568 19628
rect 24624 19572 24672 19628
rect 24728 19572 24756 19628
rect 27916 20244 27972 20254
rect 24436 18060 24756 19572
rect 24436 18004 24464 18060
rect 24520 18004 24568 18060
rect 24624 18004 24672 18060
rect 24728 18004 24756 18060
rect 24436 16492 24756 18004
rect 24436 16436 24464 16492
rect 24520 16436 24568 16492
rect 24624 16436 24672 16492
rect 24728 16436 24756 16492
rect 24436 14924 24756 16436
rect 24892 19572 24948 19582
rect 24892 16212 24948 19516
rect 27916 18676 27972 20188
rect 27916 18610 27972 18620
rect 24892 16146 24948 16156
rect 24436 14868 24464 14924
rect 24520 14868 24568 14924
rect 24624 14868 24672 14924
rect 24728 14868 24756 14924
rect 24436 13356 24756 14868
rect 24436 13300 24464 13356
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24728 13300 24756 13356
rect 24436 11788 24756 13300
rect 24436 11732 24464 11788
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24728 11732 24756 11788
rect 24436 10220 24756 11732
rect 26348 15876 26404 15886
rect 24436 10164 24464 10220
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24728 10164 24756 10220
rect 24436 8652 24756 10164
rect 24892 11396 24948 11406
rect 24892 10164 24948 11340
rect 24892 10098 24948 10108
rect 24436 8596 24464 8652
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24728 8596 24756 8652
rect 24436 7084 24756 8596
rect 26348 7476 26404 15820
rect 28028 14196 28084 20972
rect 28364 18228 28420 30044
rect 28364 18162 28420 18172
rect 28028 14130 28084 14140
rect 26348 7410 26404 7420
rect 24436 7028 24464 7084
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 24728 7028 24756 7084
rect 24436 5516 24756 7028
rect 24436 5460 24464 5516
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24728 5460 24756 5516
rect 24436 3948 24756 5460
rect 24436 3892 24464 3948
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24728 3892 24756 3948
rect 24436 2380 24756 3892
rect 24436 2324 24464 2380
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24728 2324 24756 2380
rect 24436 812 24756 2324
rect 24436 756 24464 812
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24728 756 24756 812
rect 24436 0 24756 756
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _042_
timestamp 1486834041
transform -1 0 17024 0 -1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _043_
timestamp 1486834041
transform -1 0 15456 0 1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _044_
timestamp 1486834041
transform 1 0 15120 0 -1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _045_
timestamp 1486834041
transform 1 0 15120 0 1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _046_
timestamp 1486834041
transform -1 0 12432 0 1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _047_
timestamp 1486834041
transform -1 0 16352 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _048_
timestamp 1486834041
transform -1 0 10304 0 1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _049_
timestamp 1486834041
transform 1 0 14784 0 1 16464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _050_
timestamp 1486834041
transform 1 0 15680 0 -1 18032
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _051_
timestamp 1486834041
transform -1 0 15680 0 -1 18032
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _052_
timestamp 1486834041
transform 1 0 16800 0 1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _053_
timestamp 1486834041
transform 1 0 12768 0 -1 21168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _054_
timestamp 1486834041
transform 1 0 16576 0 -1 19600
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _055_
timestamp 1486834041
transform 1 0 13216 0 1 18032
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _056_
timestamp 1486834041
transform -1 0 17248 0 -1 21168
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _057_
timestamp 1486834041
transform 1 0 15344 0 1 19600
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _058_
timestamp 1486834041
transform 1 0 13664 0 1 16464
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _059_
timestamp 1486834041
transform 1 0 15456 0 1 18032
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _060_
timestamp 1486834041
transform 1 0 12768 0 -1 19600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _061_
timestamp 1486834041
transform -1 0 13328 0 1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _062_
timestamp 1486834041
transform -1 0 12768 0 -1 19600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _063_
timestamp 1486834041
transform -1 0 10192 0 -1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _064_
timestamp 1486834041
transform 1 0 12656 0 1 22736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _065_
timestamp 1486834041
transform -1 0 12432 0 1 24304
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _066_
timestamp 1486834041
transform 1 0 12656 0 1 19600
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _067_
timestamp 1486834041
transform -1 0 13328 0 1 21168
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _068_
timestamp 1486834041
transform 1 0 11312 0 1 19600
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _069_
timestamp 1486834041
transform -1 0 12432 0 1 22736
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _070_
timestamp 1486834041
transform -1 0 12768 0 -1 21168
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _071_
timestamp 1486834041
transform 1 0 16576 0 -1 32144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _072_
timestamp 1486834041
transform 1 0 12432 0 -1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _073_
timestamp 1486834041
transform 1 0 7392 0 1 36848
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _074_
timestamp 1486834041
transform -1 0 4592 0 1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _075_
timestamp 1486834041
transform 1 0 16576 0 1 30576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _076_
timestamp 1486834041
transform 1 0 11872 0 -1 32144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _077_
timestamp 1486834041
transform 1 0 9968 0 -1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _078_
timestamp 1486834041
transform 1 0 6160 0 1 21168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _079_
timestamp 1486834041
transform 1 0 4928 0 -1 39984
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _080_
timestamp 1486834041
transform 1 0 1008 0 1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _081_
timestamp 1486834041
transform 1 0 6608 0 1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _082_
timestamp 1486834041
transform 1 0 4816 0 1 27440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _083_
timestamp 1486834041
transform -1 0 16912 0 1 21168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _084_
timestamp 1486834041
transform 1 0 12768 0 1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _085_
timestamp 1486834041
transform -1 0 4592 0 1 30576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _086_
timestamp 1486834041
transform 1 0 1904 0 -1 25872
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _087_
timestamp 1486834041
transform 1 0 6160 0 1 32144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _088_
timestamp 1486834041
transform 1 0 11424 0 -1 38416
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _089_
timestamp 1486834041
transform 1 0 1008 0 1 33712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _090_
timestamp 1486834041
transform 1 0 4928 0 -1 30576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _091_
timestamp 1486834041
transform -1 0 16352 0 -1 22736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _092_
timestamp 1486834041
transform 1 0 12656 0 -1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _093_
timestamp 1486834041
transform 1 0 12656 0 1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _094_
timestamp 1486834041
transform 1 0 10640 0 -1 16464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _095_
timestamp 1486834041
transform 1 0 1680 0 -1 32144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _096_
timestamp 1486834041
transform 1 0 2128 0 -1 21168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _097_
timestamp 1486834041
transform 1 0 4928 0 -1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _098_
timestamp 1486834041
transform 1 0 11312 0 -1 39984
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _099_
timestamp 1486834041
transform 1 0 18256 0 -1 29008
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _100_
timestamp 1486834041
transform 1 0 13440 0 1 27440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _101_
timestamp 1486834041
transform 1 0 8848 0 1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _102_
timestamp 1486834041
transform 1 0 7392 0 1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _103_
timestamp 1486834041
transform 1 0 9296 0 -1 30576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _104_
timestamp 1486834041
transform 1 0 4480 0 -1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _105_
timestamp 1486834041
transform 1 0 7168 0 1 39984
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _106_
timestamp 1486834041
transform 1 0 4032 0 -1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _107_
timestamp 1486834041
transform 1 0 17360 0 -1 25872
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _108_
timestamp 1486834041
transform 1 0 12768 0 -1 29008
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _109_
timestamp 1486834041
transform 1 0 9744 0 -1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _110_
timestamp 1486834041
transform 1 0 8736 0 -1 22736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _111_
timestamp 1486834041
transform 1 0 8848 0 1 27440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _112_
timestamp 1486834041
transform 1 0 4816 0 -1 22736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _113_
timestamp 1486834041
transform 1 0 7728 0 1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _114_
timestamp 1486834041
transform 1 0 4368 0 -1 14896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _115_
timestamp 1486834041
transform 1 0 18032 0 1 32144
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _116_
timestamp 1486834041
transform 1 0 14560 0 -1 36848
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _117_
timestamp 1486834041
transform 1 0 19600 0 -1 21168
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _118_
timestamp 1486834041
transform 1 0 13888 0 -1 11760
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _119_
timestamp 1486834041
transform -1 0 15680 0 -1 13328
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _120_
timestamp 1486834041
transform -1 0 16688 0 1 13328
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _121_
timestamp 1486834041
transform 1 0 15568 0 1 14896
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _122_
timestamp 1486834041
transform 1 0 16688 0 1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _123_
timestamp 1486834041
transform -1 0 15568 0 1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _124_
timestamp 1486834041
transform 1 0 15792 0 -1 14896
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _125_
timestamp 1486834041
transform -1 0 16352 0 -1 16464
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _126_
timestamp 1486834041
transform 1 0 16576 0 -1 14896
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _127_
timestamp 1486834041
transform 1 0 9744 0 1 16464
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _128_
timestamp 1486834041
transform -1 0 11536 0 1 16464
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _129_
timestamp 1486834041
transform 1 0 9744 0 -1 14896
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _130_
timestamp 1486834041
transform -1 0 9744 0 -1 14896
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _131_
timestamp 1486834041
transform 1 0 10864 0 -1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _132_
timestamp 1486834041
transform 1 0 9744 0 -1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _133_
timestamp 1486834041
transform 1 0 11648 0 1 14896
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _134_
timestamp 1486834041
transform 1 0 8960 0 -1 16464
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _135_
timestamp 1486834041
transform -1 0 11648 0 1 14896
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _136_
timestamp 1486834041
transform 1 0 12880 0 1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _137_
timestamp 1486834041
transform 1 0 17808 0 1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _138_
timestamp 1486834041
transform -1 0 18816 0 -1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _139_
timestamp 1486834041
transform 1 0 17584 0 -1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _140_
timestamp 1486834041
transform 1 0 1792 0 -1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _141_
timestamp 1486834041
transform 1 0 4032 0 -1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _142_
timestamp 1486834041
transform 1 0 5488 0 1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _143_
timestamp 1486834041
transform -1 0 10976 0 -1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _144_
timestamp 1486834041
transform 1 0 2352 0 1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _145_
timestamp 1486834041
transform 1 0 3808 0 -1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _146_
timestamp 1486834041
transform 1 0 6272 0 -1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _147_
timestamp 1486834041
transform 1 0 8176 0 1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _148_
timestamp 1486834041
transform 1 0 6272 0 -1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _149_
timestamp 1486834041
transform 1 0 6384 0 1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _150_
timestamp 1486834041
transform 1 0 6272 0 -1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _151_
timestamp 1486834041
transform 1 0 9072 0 1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _152_
timestamp 1486834041
transform 1 0 10976 0 -1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _153_
timestamp 1486834041
transform 1 0 10528 0 -1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _154_
timestamp 1486834041
transform 1 0 16128 0 1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _155_
timestamp 1486834041
transform 1 0 17472 0 -1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _156_
timestamp 1486834041
transform 1 0 1792 0 -1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _157_
timestamp 1486834041
transform 1 0 4816 0 1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _158_
timestamp 1486834041
transform 1 0 4368 0 -1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _159_
timestamp 1486834041
transform 1 0 2352 0 1 39984
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _160_
timestamp 1486834041
transform 1 0 2352 0 1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _161_
timestamp 1486834041
transform 1 0 3136 0 -1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _162_
timestamp 1486834041
transform 1 0 7840 0 1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _163_
timestamp 1486834041
transform 1 0 9184 0 -1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _164_
timestamp 1486834041
transform 1 0 5936 0 -1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _165_
timestamp 1486834041
transform 1 0 7280 0 1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _166_
timestamp 1486834041
transform 1 0 6608 0 1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _167_
timestamp 1486834041
transform 1 0 8736 0 -1 13328
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _168_
timestamp 1486834041
transform 1 0 13216 0 -1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _169_
timestamp 1486834041
transform 1 0 13328 0 1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _170_
timestamp 1486834041
transform 1 0 17136 0 1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _171_
timestamp 1486834041
transform 1 0 17808 0 1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _172_
timestamp 1486834041
transform 1 0 9856 0 -1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _173_
timestamp 1486834041
transform 1 0 9072 0 -1 39984
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _174_
timestamp 1486834041
transform 1 0 4816 0 1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _175_
timestamp 1486834041
transform 1 0 2352 0 -1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _176_
timestamp 1486834041
transform 1 0 1904 0 -1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _177_
timestamp 1486834041
transform -1 0 3584 0 -1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _178_
timestamp 1486834041
transform 1 0 1344 0 1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _179_
timestamp 1486834041
transform 1 0 896 0 -1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _180_
timestamp 1486834041
transform 1 0 6272 0 -1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _181_
timestamp 1486834041
transform 1 0 7728 0 1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _182_
timestamp 1486834041
transform 1 0 9184 0 1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _183_
timestamp 1486834041
transform 1 0 10192 0 1 10192
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _184_
timestamp 1486834041
transform 1 0 10416 0 -1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _185_
timestamp 1486834041
transform 1 0 10080 0 -1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _186_
timestamp 1486834041
transform -1 0 18816 0 -1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _187_
timestamp 1486834041
transform -1 0 19376 0 1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _188_
timestamp 1486834041
transform 1 0 4816 0 1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _189_
timestamp 1486834041
transform 1 0 3136 0 -1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _190_
timestamp 1486834041
transform 1 0 896 0 -1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _191_
timestamp 1486834041
transform -1 0 3136 0 -1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _192_
timestamp 1486834041
transform 1 0 10192 0 1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _193_
timestamp 1486834041
transform 1 0 9184 0 -1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _194_
timestamp 1486834041
transform -1 0 9520 0 1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _195_
timestamp 1486834041
transform 1 0 5264 0 -1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _196_
timestamp 1486834041
transform 1 0 1344 0 1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _197_
timestamp 1486834041
transform 1 0 896 0 -1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _198_
timestamp 1486834041
transform 1 0 896 0 -1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _199_
timestamp 1486834041
transform 1 0 896 0 1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _200_
timestamp 1486834041
transform 1 0 12320 0 -1 25872
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _201_
timestamp 1486834041
transform -1 0 18592 0 1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _202_
timestamp 1486834041
transform -1 0 19152 0 1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _203_
timestamp 1486834041
transform -1 0 19600 0 -1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _204_
timestamp 1486834041
transform 1 0 2352 0 1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _205_
timestamp 1486834041
transform 1 0 4592 0 -1 27440
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _206_
timestamp 1486834041
transform 1 0 4032 0 -1 11760
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _207_
timestamp 1486834041
transform 1 0 3920 0 -1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _208_
timestamp 1486834041
transform -1 0 3920 0 1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _209_
timestamp 1486834041
transform -1 0 3920 0 -1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _210_
timestamp 1486834041
transform 1 0 3584 0 -1 41552
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _211_
timestamp 1486834041
transform 1 0 5264 0 1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _212_
timestamp 1486834041
transform 1 0 5264 0 1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _213_
timestamp 1486834041
transform 1 0 5936 0 -1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _214_
timestamp 1486834041
transform 1 0 6944 0 1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _215_
timestamp 1486834041
transform 1 0 9408 0 -1 8624
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _216_
timestamp 1486834041
transform 1 0 10192 0 1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _217_
timestamp 1486834041
transform 1 0 11536 0 -1 33712
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _218_
timestamp 1486834041
transform 1 0 15568 0 1 29008
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _219_
timestamp 1486834041
transform 1 0 16576 0 -1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _220_
timestamp 1486834041
transform 1 0 1904 0 1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _221_
timestamp 1486834041
transform -1 0 4480 0 -1 24304
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _222_
timestamp 1486834041
transform 1 0 4816 0 1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _223_
timestamp 1486834041
transform 1 0 2352 0 1 38416
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _224_
timestamp 1486834041
transform 1 0 10192 0 -1 35280
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _225_
timestamp 1486834041
transform 1 0 11424 0 -1 36848
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _226_
timestamp 1486834041
transform 1 0 13888 0 1 30576
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _227_
timestamp 1486834041
transform 1 0 14896 0 1 32144
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _228_
timestamp 1486834041
transform 1 0 9744 0 1 21168
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _229_
timestamp 1486834041
transform 1 0 8624 0 1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _230_
timestamp 1486834041
transform 1 0 6384 0 1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _231_
timestamp 1486834041
transform 1 0 8624 0 1 19600
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _232_
timestamp 1486834041
transform 1 0 13552 0 -1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _233_
timestamp 1486834041
transform -1 0 18816 0 -1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _234_
timestamp 1486834041
transform -1 0 18928 0 1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _235_
timestamp 1486834041
transform -1 0 19376 0 -1 22736
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _236_
timestamp 1486834041
transform 1 0 9968 0 1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _237_
timestamp 1486834041
transform 1 0 9296 0 -1 18032
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _238_
timestamp 1486834041
transform 1 0 6384 0 1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _239_
timestamp 1486834041
transform 1 0 7616 0 1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _240_
timestamp 1486834041
transform 1 0 6160 0 -1 16464
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__latq_1  _241_
timestamp 1486834041
transform 1 0 5376 0 1 14896
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_4  _242_
timestamp 1486834041
transform 1 0 16576 0 -1 38416
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_4  _243_
timestamp 1486834041
transform -1 0 18704 0 1 39984
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _244_
timestamp 1486834041
transform -1 0 2352 0 1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _245_
timestamp 1486834041
transform 1 0 3584 0 1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _246_
timestamp 1486834041
transform 1 0 11536 0 1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _247_
timestamp 1486834041
transform 1 0 13328 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _248_
timestamp 1486834041
transform 1 0 13888 0 1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _249_
timestamp 1486834041
transform 1 0 16240 0 1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _250_
timestamp 1486834041
transform 1 0 6048 0 1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _251_
timestamp 1486834041
transform -1 0 2352 0 -1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _252_
timestamp 1486834041
transform 1 0 12768 0 1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _253_
timestamp 1486834041
transform 1 0 7504 0 -1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _254_
timestamp 1486834041
transform 1 0 3584 0 1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _255_
timestamp 1486834041
transform -1 0 3360 0 -1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _256_
timestamp 1486834041
transform 1 0 14560 0 -1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _257_
timestamp 1486834041
transform 1 0 14448 0 1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _258_
timestamp 1486834041
transform 1 0 1456 0 1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _259_
timestamp 1486834041
transform 1 0 1568 0 -1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _260_
timestamp 1486834041
transform 1 0 3696 0 1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _261_
timestamp 1486834041
transform 1 0 5488 0 1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _262_
timestamp 1486834041
transform 1 0 7616 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _263_
timestamp 1486834041
transform 1 0 9968 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _264_
timestamp 1486834041
transform 1 0 11200 0 1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _265_
timestamp 1486834041
transform 1 0 11536 0 1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _266_
timestamp 1486834041
transform 1 0 15456 0 -1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _267_
timestamp 1486834041
transform 1 0 19264 0 -1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _268_
timestamp 1486834041
transform 1 0 896 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _269_
timestamp 1486834041
transform 1 0 2688 0 -1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _270_
timestamp 1486834041
transform 1 0 896 0 1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _271_
timestamp 1486834041
transform 1 0 2464 0 -1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _272_
timestamp 1486834041
transform 1 0 6608 0 -1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _273_
timestamp 1486834041
transform 1 0 1456 0 1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _274_
timestamp 1486834041
transform 1 0 13664 0 1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _275_
timestamp 1486834041
transform 1 0 14448 0 -1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _276_
timestamp 1486834041
transform 1 0 1008 0 -1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _277_
timestamp 1486834041
transform 1 0 1344 0 -1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _278_
timestamp 1486834041
transform 1 0 2464 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _279_
timestamp 1486834041
transform 1 0 1792 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _280_
timestamp 1486834041
transform 1 0 12656 0 1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _281_
timestamp 1486834041
transform 1 0 18816 0 1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _282_
timestamp 1486834041
transform 1 0 19712 0 -1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _283_
timestamp 1486834041
transform 1 0 19040 0 1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _284_
timestamp 1486834041
transform 1 0 3472 0 1 41552
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _285_
timestamp 1486834041
transform 1 0 5936 0 -1 41552
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _286_
timestamp 1486834041
transform 1 0 5152 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _287_
timestamp 1486834041
transform 1 0 1792 0 1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _288_
timestamp 1486834041
transform 1 0 1792 0 1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _289_
timestamp 1486834041
transform 1 0 1792 0 -1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _290_
timestamp 1486834041
transform -1 0 12208 0 1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _291_
timestamp 1486834041
transform 1 0 1232 0 -1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _292_
timestamp 1486834041
transform 1 0 2464 0 1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _293_
timestamp 1486834041
transform 1 0 18144 0 -1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _294_
timestamp 1486834041
transform 1 0 20496 0 1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _295_
timestamp 1486834041
transform 1 0 18816 0 1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _296_
timestamp 1486834041
transform 1 0 19824 0 -1 55664
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _297_
timestamp 1486834041
transform 1 0 23632 0 1 50960
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _298_
timestamp 1486834041
transform 1 0 21616 0 -1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _299_
timestamp 1486834041
transform 1 0 22624 0 1 50960
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _300_
timestamp 1486834041
transform 1 0 20720 0 -1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _301_
timestamp 1486834041
transform 1 0 21168 0 1 52528
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _302_
timestamp 1486834041
transform 1 0 22064 0 1 52528
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _303_
timestamp 1486834041
transform -1 0 19600 0 -1 55664
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _304_
timestamp 1486834041
transform 1 0 23632 0 1 49392
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _305_
timestamp 1486834041
transform 1 0 24304 0 1 47824
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _306_
timestamp 1486834041
transform -1 0 22624 0 -1 52528
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _307_
timestamp 1486834041
transform 1 0 25200 0 1 47824
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _308_
timestamp 1486834041
transform -1 0 24192 0 -1 50960
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _309_
timestamp 1486834041
transform -1 0 20720 0 -1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _310_
timestamp 1486834041
transform -1 0 15680 0 -1 38416
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _311_
timestamp 1486834041
transform 1 0 14224 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _312_
timestamp 1486834041
transform -1 0 20048 0 1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _313_
timestamp 1486834041
transform -1 0 14560 0 -1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _314_
timestamp 1486834041
transform 1 0 18816 0 -1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _315_
timestamp 1486834041
transform 1 0 5264 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _316_
timestamp 1486834041
transform -1 0 8512 0 -1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _317_
timestamp 1486834041
transform 1 0 5488 0 1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _318_
timestamp 1486834041
transform 1 0 10080 0 -1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _319_
timestamp 1486834041
transform -1 0 10080 0 -1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _320_
timestamp 1486834041
transform 1 0 11200 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _321_
timestamp 1486834041
transform 1 0 14000 0 -1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _322_
timestamp 1486834041
transform 1 0 18816 0 1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _323_
timestamp 1486834041
transform -1 0 5488 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _324_
timestamp 1486834041
transform 1 0 8736 0 -1 41552
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _325_
timestamp 1486834041
transform 1 0 5488 0 1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _326_
timestamp 1486834041
transform 1 0 10192 0 1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _327_
timestamp 1486834041
transform 1 0 8736 0 -1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _328_
timestamp 1486834041
transform 1 0 12096 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _329_
timestamp 1486834041
transform 1 0 15456 0 -1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _330_
timestamp 1486834041
transform 1 0 19376 0 1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _331_
timestamp 1486834041
transform -1 0 6272 0 -1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _332_
timestamp 1486834041
transform -1 0 7728 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _333_
timestamp 1486834041
transform 1 0 2688 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _334_
timestamp 1486834041
transform 1 0 6272 0 1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _335_
timestamp 1486834041
transform -1 0 6160 0 1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _336_
timestamp 1486834041
transform 1 0 10864 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _337_
timestamp 1486834041
transform 1 0 12768 0 1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _338_
timestamp 1486834041
transform -1 0 18032 0 1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _339_
timestamp 1486834041
transform -1 0 1904 0 1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _340_
timestamp 1486834041
transform -1 0 8512 0 -1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _341_
timestamp 1486834041
transform -1 0 13552 0 1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _342_
timestamp 1486834041
transform -1 0 17584 0 -1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _343_
timestamp 1486834041
transform 1 0 12768 0 1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _344_
timestamp 1486834041
transform 1 0 6048 0 -1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_UserCLK
timestamp 1486834041
transform 1 0 16576 0 -1 39984
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_UserCLK_regs
timestamp 1486834041
transform -1 0 20272 0 1 36848
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_UserCLK
timestamp 1486834041
transform -1 0 19152 0 1 35280
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_UserCLK_regs
timestamp 1486834041
transform -1 0 20160 0 1 33712
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_UserCLK_regs
timestamp 1486834041
transform 1 0 14672 0 1 41552
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_regs_0_UserCLK
timestamp 1486834041
transform 1 0 14672 0 1 38416
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout27
timestamp 1486834041
transform -1 0 18144 0 -1 36848
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout28
timestamp 1486834041
transform -1 0 8624 0 1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout29
timestamp 1486834041
transform 1 0 7616 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout30
timestamp 1486834041
transform -1 0 2464 0 1 18032
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout31
timestamp 1486834041
transform -1 0 4032 0 1 19600
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout32
timestamp 1486834041
transform 1 0 896 0 1 19600
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout33
timestamp 1486834041
transform 1 0 896 0 -1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout34
timestamp 1486834041
transform 1 0 896 0 -1 30576
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout35
timestamp 1486834041
transform 1 0 896 0 1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout36
timestamp 1486834041
transform -1 0 1792 0 1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout37
timestamp 1486834041
transform 1 0 4816 0 1 16464
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout38
timestamp 1486834041
transform -1 0 4592 0 1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout39
timestamp 1486834041
transform -1 0 7840 0 1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout40
timestamp 1486834041
transform 1 0 6944 0 -1 32144
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout41
timestamp 1486834041
transform 1 0 8736 0 -1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2
timestamp 1486834041
transform 1 0 896 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36
timestamp 1486834041
transform 1 0 4704 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_70
timestamp 1486834041
transform 1 0 8512 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_104
timestamp 1486834041
transform 1 0 12320 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_138
timestamp 1486834041
transform 1 0 16128 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_172
timestamp 1486834041
transform 1 0 19936 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_206
timestamp 1486834041
transform 1 0 23744 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_240
timestamp 1486834041
transform 1 0 27552 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_2
timestamp 1486834041
transform 1 0 896 0 -1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_66
timestamp 1486834041
transform 1 0 8064 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_72
timestamp 1486834041
transform 1 0 8736 0 -1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_136
timestamp 1486834041
transform 1 0 15904 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_142
timestamp 1486834041
transform 1 0 16576 0 -1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_206
timestamp 1486834041
transform 1 0 23744 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_212
timestamp 1486834041
transform 1 0 24416 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_228
timestamp 1486834041
transform 1 0 26208 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_236
timestamp 1486834041
transform 1 0 27104 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_240
timestamp 1486834041
transform 1 0 27552 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_2
timestamp 1486834041
transform 1 0 896 0 1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1486834041
transform 1 0 4480 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_37
timestamp 1486834041
transform 1 0 4816 0 1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_101
timestamp 1486834041
transform 1 0 11984 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_107
timestamp 1486834041
transform 1 0 12656 0 1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_171
timestamp 1486834041
transform 1 0 19824 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_177
timestamp 1486834041
transform 1 0 20496 0 1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_2
timestamp 1486834041
transform 1 0 896 0 -1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_66
timestamp 1486834041
transform 1 0 8064 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_72
timestamp 1486834041
transform 1 0 8736 0 -1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_136
timestamp 1486834041
transform 1 0 15904 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_142
timestamp 1486834041
transform 1 0 16576 0 -1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_206
timestamp 1486834041
transform 1 0 23744 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_212
timestamp 1486834041
transform 1 0 24416 0 -1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_228
timestamp 1486834041
transform 1 0 26208 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_236
timestamp 1486834041
transform 1 0 27104 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_240
timestamp 1486834041
transform 1 0 27552 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_2
timestamp 1486834041
transform 1 0 896 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1486834041
transform 1 0 4480 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_37
timestamp 1486834041
transform 1 0 4816 0 1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_101
timestamp 1486834041
transform 1 0 11984 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_107
timestamp 1486834041
transform 1 0 12656 0 1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_171
timestamp 1486834041
transform 1 0 19824 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_177
timestamp 1486834041
transform 1 0 20496 0 1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_2
timestamp 1486834041
transform 1 0 896 0 -1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_66
timestamp 1486834041
transform 1 0 8064 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_72
timestamp 1486834041
transform 1 0 8736 0 -1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_136
timestamp 1486834041
transform 1 0 15904 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_142
timestamp 1486834041
transform 1 0 16576 0 -1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_206
timestamp 1486834041
transform 1 0 23744 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_212
timestamp 1486834041
transform 1 0 24416 0 -1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_228
timestamp 1486834041
transform 1 0 26208 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_236
timestamp 1486834041
transform 1 0 27104 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_240
timestamp 1486834041
transform 1 0 27552 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_16
timestamp 1486834041
transform 1 0 2464 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_32
timestamp 1486834041
transform 1 0 4256 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1486834041
transform 1 0 4480 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_37
timestamp 1486834041
transform 1 0 4816 0 1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_101
timestamp 1486834041
transform 1 0 11984 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_107
timestamp 1486834041
transform 1 0 12656 0 1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_171
timestamp 1486834041
transform 1 0 19824 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_177
timestamp 1486834041
transform 1 0 20496 0 1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_16
timestamp 1486834041
transform 1 0 2464 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_48
timestamp 1486834041
transform 1 0 6048 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_64
timestamp 1486834041
transform 1 0 7840 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_68
timestamp 1486834041
transform 1 0 8288 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_72
timestamp 1486834041
transform 1 0 8736 0 -1 7056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_136
timestamp 1486834041
transform 1 0 15904 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_142
timestamp 1486834041
transform 1 0 16576 0 -1 7056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_206
timestamp 1486834041
transform 1 0 23744 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_212
timestamp 1486834041
transform 1 0 24416 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_228
timestamp 1486834041
transform 1 0 26208 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_236
timestamp 1486834041
transform 1 0 27104 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_240
timestamp 1486834041
transform 1 0 27552 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1486834041
transform 1 0 896 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1486834041
transform 1 0 4480 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_37
timestamp 1486834041
transform 1 0 4816 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_69
timestamp 1486834041
transform 1 0 8400 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_77
timestamp 1486834041
transform 1 0 9296 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_81
timestamp 1486834041
transform 1 0 9744 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_99
timestamp 1486834041
transform 1 0 11760 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_103
timestamp 1486834041
transform 1 0 12208 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_107
timestamp 1486834041
transform 1 0 12656 0 1 7056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_171
timestamp 1486834041
transform 1 0 19824 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_177
timestamp 1486834041
transform 1 0 20496 0 1 7056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_2
timestamp 1486834041
transform 1 0 896 0 -1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_34
timestamp 1486834041
transform 1 0 4480 0 -1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_50
timestamp 1486834041
transform 1 0 6272 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_58
timestamp 1486834041
transform 1 0 7168 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_72
timestamp 1486834041
transform 1 0 8736 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_76
timestamp 1486834041
transform 1 0 9184 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_98
timestamp 1486834041
transform 1 0 11648 0 -1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_130
timestamp 1486834041
transform 1 0 15232 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_138
timestamp 1486834041
transform 1 0 16128 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_142
timestamp 1486834041
transform 1 0 16576 0 -1 8624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_206
timestamp 1486834041
transform 1 0 23744 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_212
timestamp 1486834041
transform 1 0 24416 0 -1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_228
timestamp 1486834041
transform 1 0 26208 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_236
timestamp 1486834041
transform 1 0 27104 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_240
timestamp 1486834041
transform 1 0 27552 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_2
timestamp 1486834041
transform 1 0 896 0 1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1486834041
transform 1 0 4480 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_37
timestamp 1486834041
transform 1 0 4816 0 1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_53
timestamp 1486834041
transform 1 0 6608 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_55
timestamp 1486834041
transform 1 0 6832 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_96
timestamp 1486834041
transform 1 0 11424 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_104
timestamp 1486834041
transform 1 0 12320 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_107
timestamp 1486834041
transform 1 0 12656 0 1 8624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_171
timestamp 1486834041
transform 1 0 19824 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_177
timestamp 1486834041
transform 1 0 20496 0 1 8624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_16
timestamp 1486834041
transform 1 0 2464 0 -1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_32
timestamp 1486834041
transform 1 0 4256 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_34
timestamp 1486834041
transform 1 0 4480 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_43
timestamp 1486834041
transform 1 0 5488 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_51
timestamp 1486834041
transform 1 0 6384 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_63
timestamp 1486834041
transform 1 0 7728 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_67
timestamp 1486834041
transform 1 0 8176 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_69
timestamp 1486834041
transform 1 0 8400 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_72
timestamp 1486834041
transform 1 0 8736 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_80
timestamp 1486834041
transform 1 0 9632 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_82
timestamp 1486834041
transform 1 0 9856 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_115
timestamp 1486834041
transform 1 0 13552 0 -1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_131
timestamp 1486834041
transform 1 0 15344 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_139
timestamp 1486834041
transform 1 0 16240 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_142
timestamp 1486834041
transform 1 0 16576 0 -1 10192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_206
timestamp 1486834041
transform 1 0 23744 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_212
timestamp 1486834041
transform 1 0 24416 0 -1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_228
timestamp 1486834041
transform 1 0 26208 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_236
timestamp 1486834041
transform 1 0 27104 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_240
timestamp 1486834041
transform 1 0 27552 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_2
timestamp 1486834041
transform 1 0 896 0 1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1486834041
transform 1 0 4480 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_37
timestamp 1486834041
transform 1 0 4816 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_39
timestamp 1486834041
transform 1 0 5040 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_48
timestamp 1486834041
transform 1 0 6048 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_52
timestamp 1486834041
transform 1 0 6496 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_107
timestamp 1486834041
transform 1 0 12656 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_111
timestamp 1486834041
transform 1 0 13104 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_129
timestamp 1486834041
transform 1 0 15120 0 1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_161
timestamp 1486834041
transform 1 0 18704 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_169
timestamp 1486834041
transform 1 0 19600 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_173
timestamp 1486834041
transform 1 0 20048 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_177
timestamp 1486834041
transform 1 0 20496 0 1 10192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_24
timestamp 1486834041
transform 1 0 3360 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_28
timestamp 1486834041
transform 1 0 3808 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_72
timestamp 1486834041
transform 1 0 8736 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_80
timestamp 1486834041
transform 1 0 9632 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_113
timestamp 1486834041
transform 1 0 13328 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_117
timestamp 1486834041
transform 1 0 13776 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_133
timestamp 1486834041
transform 1 0 15568 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_137
timestamp 1486834041
transform 1 0 16016 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_139
timestamp 1486834041
transform 1 0 16240 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_142
timestamp 1486834041
transform 1 0 16576 0 -1 11760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_206
timestamp 1486834041
transform 1 0 23744 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_212
timestamp 1486834041
transform 1 0 24416 0 -1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_228
timestamp 1486834041
transform 1 0 26208 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_236
timestamp 1486834041
transform 1 0 27104 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_240
timestamp 1486834041
transform 1 0 27552 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_26
timestamp 1486834041
transform 1 0 3584 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1486834041
transform 1 0 4480 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_37
timestamp 1486834041
transform 1 0 4816 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_49
timestamp 1486834041
transform 1 0 6160 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_139
timestamp 1486834041
transform 1 0 16240 0 1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_171
timestamp 1486834041
transform 1 0 19824 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_177
timestamp 1486834041
transform 1 0 20496 0 1 11760
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_2
timestamp 1486834041
transform 1 0 896 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_92
timestamp 1486834041
transform 1 0 10976 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_110
timestamp 1486834041
transform 1 0 12992 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_118
timestamp 1486834041
transform 1 0 13888 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_134
timestamp 1486834041
transform 1 0 15680 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_142
timestamp 1486834041
transform 1 0 16576 0 -1 13328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_206
timestamp 1486834041
transform 1 0 23744 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_212
timestamp 1486834041
transform 1 0 24416 0 -1 13328
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_228
timestamp 1486834041
transform 1 0 26208 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_236
timestamp 1486834041
transform 1 0 27104 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_240
timestamp 1486834041
transform 1 0 27552 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_2
timestamp 1486834041
transform 1 0 896 0 1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_71
timestamp 1486834041
transform 1 0 8624 0 1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_95
timestamp 1486834041
transform 1 0 11312 0 1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_103
timestamp 1486834041
transform 1 0 12208 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_107
timestamp 1486834041
transform 1 0 12656 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_151
timestamp 1486834041
transform 1 0 17584 0 1 13328
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_167
timestamp 1486834041
transform 1 0 19376 0 1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_177
timestamp 1486834041
transform 1 0 20496 0 1 13328
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_2
timestamp 1486834041
transform 1 0 896 0 -1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_26
timestamp 1486834041
transform 1 0 3584 0 -1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_30
timestamp 1486834041
transform 1 0 4032 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_32
timestamp 1486834041
transform 1 0 4256 0 -1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_65
timestamp 1486834041
transform 1 0 7952 0 -1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_69
timestamp 1486834041
transform 1 0 8400 0 -1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_72
timestamp 1486834041
transform 1 0 8736 0 -1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_97
timestamp 1486834041
transform 1 0 11536 0 -1 14896
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_113
timestamp 1486834041
transform 1 0 13328 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_17_154
timestamp 1486834041
transform 1 0 17920 0 -1 14896
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_186
timestamp 1486834041
transform 1 0 21504 0 -1 14896
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_202
timestamp 1486834041
transform 1 0 23296 0 -1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_212
timestamp 1486834041
transform 1 0 24416 0 -1 14896
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_228
timestamp 1486834041
transform 1 0 26208 0 -1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_236
timestamp 1486834041
transform 1 0 27104 0 -1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_240
timestamp 1486834041
transform 1 0 27552 0 -1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_2
timestamp 1486834041
transform 1 0 896 0 1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_6
timestamp 1486834041
transform 1 0 1344 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_8
timestamp 1486834041
transform 1 0 1568 0 1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_29
timestamp 1486834041
transform 1 0 3920 0 1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_33
timestamp 1486834041
transform 1 0 4368 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_37
timestamp 1486834041
transform 1 0 4816 0 1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_41
timestamp 1486834041
transform 1 0 5264 0 1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_103
timestamp 1486834041
transform 1 0 12208 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_107
timestamp 1486834041
transform 1 0 12656 0 1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_111
timestamp 1486834041
transform 1 0 13104 0 1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_118
timestamp 1486834041
transform 1 0 13888 0 1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_122
timestamp 1486834041
transform 1 0 14336 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_124
timestamp 1486834041
transform 1 0 14560 0 1 14896
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_163
timestamp 1486834041
transform 1 0 18928 0 1 14896
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_171
timestamp 1486834041
transform 1 0 19824 0 1 14896
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_177
timestamp 1486834041
transform 1 0 20496 0 1 14896
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_2
timestamp 1486834041
transform 1 0 896 0 -1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_6
timestamp 1486834041
transform 1 0 1344 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_8
timestamp 1486834041
transform 1 0 1568 0 -1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_69
timestamp 1486834041
transform 1 0 8400 0 -1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_72
timestamp 1486834041
transform 1 0 8736 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_121
timestamp 1486834041
transform 1 0 14224 0 -1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_19_162
timestamp 1486834041
transform 1 0 18816 0 -1 16464
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_194
timestamp 1486834041
transform 1 0 22400 0 -1 16464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_212
timestamp 1486834041
transform 1 0 24416 0 -1 16464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_228
timestamp 1486834041
transform 1 0 26208 0 -1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_236
timestamp 1486834041
transform 1 0 27104 0 -1 16464
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_240
timestamp 1486834041
transform 1 0 27552 0 -1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_18
timestamp 1486834041
transform 1 0 2688 0 1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_26
timestamp 1486834041
transform 1 0 3584 0 1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_71
timestamp 1486834041
transform 1 0 8624 0 1 16464
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_79
timestamp 1486834041
transform 1 0 9520 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_113
timestamp 1486834041
transform 1 0 13328 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_115
timestamp 1486834041
transform 1 0 13552 0 1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_158
timestamp 1486834041
transform 1 0 18368 0 1 16464
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_174
timestamp 1486834041
transform 1 0 20160 0 1 16464
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_177
timestamp 1486834041
transform 1 0 20496 0 1 16464
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_72
timestamp 1486834041
transform 1 0 8736 0 -1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_76
timestamp 1486834041
transform 1 0 9184 0 -1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_97
timestamp 1486834041
transform 1 0 11536 0 -1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_101
timestamp 1486834041
transform 1 0 11984 0 -1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_142
timestamp 1486834041
transform 1 0 16576 0 -1 18032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_206
timestamp 1486834041
transform 1 0 23744 0 -1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_212
timestamp 1486834041
transform 1 0 24416 0 -1 18032
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_228
timestamp 1486834041
transform 1 0 26208 0 -1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_236
timestamp 1486834041
transform 1 0 27104 0 -1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_240
timestamp 1486834041
transform 1 0 27552 0 -1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_24
timestamp 1486834041
transform 1 0 3360 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_26
timestamp 1486834041
transform 1 0 3584 0 1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_37
timestamp 1486834041
transform 1 0 4816 0 1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_61
timestamp 1486834041
transform 1 0 7504 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_103
timestamp 1486834041
transform 1 0 12208 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_107
timestamp 1486834041
transform 1 0 12656 0 1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_111
timestamp 1486834041
transform 1 0 13104 0 1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_127
timestamp 1486834041
transform 1 0 14896 0 1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_152
timestamp 1486834041
transform 1 0 17696 0 1 18032
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_160
timestamp 1486834041
transform 1 0 18592 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_170
timestamp 1486834041
transform 1 0 19712 0 1 18032
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_174
timestamp 1486834041
transform 1 0 20160 0 1 18032
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_177
timestamp 1486834041
transform 1 0 20496 0 1 18032
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_2
timestamp 1486834041
transform 1 0 896 0 -1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_26
timestamp 1486834041
transform 1 0 3584 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_48
timestamp 1486834041
transform 1 0 6048 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_72
timestamp 1486834041
transform 1 0 8736 0 -1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_23_148
timestamp 1486834041
transform 1 0 17248 0 -1 19600
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_180
timestamp 1486834041
transform 1 0 20832 0 -1 19600
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_196
timestamp 1486834041
transform 1 0 22624 0 -1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_204
timestamp 1486834041
transform 1 0 23520 0 -1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_208
timestamp 1486834041
transform 1 0 23968 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_212
timestamp 1486834041
transform 1 0 24416 0 -1 19600
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_228
timestamp 1486834041
transform 1 0 26208 0 -1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_236
timestamp 1486834041
transform 1 0 27104 0 -1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_240
timestamp 1486834041
transform 1 0 27552 0 -1 19600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_30
timestamp 1486834041
transform 1 0 4032 0 1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_34
timestamp 1486834041
transform 1 0 4480 0 1 19600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_37
timestamp 1486834041
transform 1 0 4816 0 1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_41
timestamp 1486834041
transform 1 0 5264 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_91
timestamp 1486834041
transform 1 0 10864 0 1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_122
timestamp 1486834041
transform 1 0 14336 0 1 19600
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_141
timestamp 1486834041
transform 1 0 16464 0 1 19600
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_149
timestamp 1486834041
transform 1 0 17360 0 1 19600
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_173
timestamp 1486834041
transform 1 0 20048 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_177
timestamp 1486834041
transform 1 0 20496 0 1 19600
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_2
timestamp 1486834041
transform 1 0 896 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_4
timestamp 1486834041
transform 1 0 1120 0 -1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_45
timestamp 1486834041
transform 1 0 5712 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_67
timestamp 1486834041
transform 1 0 8176 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_69
timestamp 1486834041
transform 1 0 8400 0 -1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_72
timestamp 1486834041
transform 1 0 8736 0 -1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_76
timestamp 1486834041
transform 1 0 9184 0 -1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_148
timestamp 1486834041
transform 1 0 17248 0 -1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_184
timestamp 1486834041
transform 1 0 21280 0 -1 21168
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_200
timestamp 1486834041
transform 1 0 23072 0 -1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_208
timestamp 1486834041
transform 1 0 23968 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_212
timestamp 1486834041
transform 1 0 24416 0 -1 21168
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_228
timestamp 1486834041
transform 1 0 26208 0 -1 21168
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_236
timestamp 1486834041
transform 1 0 27104 0 -1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_240
timestamp 1486834041
transform 1 0 27552 0 -1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_2
timestamp 1486834041
transform 1 0 896 0 1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_6
timestamp 1486834041
transform 1 0 1344 0 1 21168
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_37
timestamp 1486834041
transform 1 0 4816 0 1 21168
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_173
timestamp 1486834041
transform 1 0 20048 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_177
timestamp 1486834041
transform 1 0 20496 0 1 21168
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_209
timestamp 1486834041
transform 1 0 24080 0 1 21168
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_225
timestamp 1486834041
transform 1 0 25872 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_2
timestamp 1486834041
transform 1 0 896 0 -1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_31
timestamp 1486834041
transform 1 0 4144 0 -1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_35
timestamp 1486834041
transform 1 0 4592 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_69
timestamp 1486834041
transform 1 0 8400 0 -1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_104
timestamp 1486834041
transform 1 0 12320 0 -1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_146
timestamp 1486834041
transform 1 0 17024 0 -1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_27_167
timestamp 1486834041
transform 1 0 19376 0 -1 22736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_199
timestamp 1486834041
transform 1 0 22960 0 -1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_207
timestamp 1486834041
transform 1 0 23856 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_209
timestamp 1486834041
transform 1 0 24080 0 -1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_212
timestamp 1486834041
transform 1 0 24416 0 -1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_2
timestamp 1486834041
transform 1 0 896 0 1 22736
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_31
timestamp 1486834041
transform 1 0 4144 0 1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_37
timestamp 1486834041
transform 1 0 4816 0 1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_41
timestamp 1486834041
transform 1 0 5264 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_91
timestamp 1486834041
transform 1 0 10864 0 1 22736
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_167
timestamp 1486834041
transform 1 0 19376 0 1 22736
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_177
timestamp 1486834041
transform 1 0 20496 0 1 22736
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_209
timestamp 1486834041
transform 1 0 24080 0 1 22736
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_225
timestamp 1486834041
transform 1 0 25872 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_2
timestamp 1486834041
transform 1 0 896 0 -1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_66
timestamp 1486834041
transform 1 0 8064 0 -1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_72
timestamp 1486834041
transform 1 0 8736 0 -1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_84
timestamp 1486834041
transform 1 0 10080 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_86
timestamp 1486834041
transform 1 0 10304 0 -1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_139
timestamp 1486834041
transform 1 0 16240 0 -1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_162
timestamp 1486834041
transform 1 0 18816 0 -1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_29_174
timestamp 1486834041
transform 1 0 20160 0 -1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_206
timestamp 1486834041
transform 1 0 23744 0 -1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_212
timestamp 1486834041
transform 1 0 24416 0 -1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_2
timestamp 1486834041
transform 1 0 896 0 1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_37
timestamp 1486834041
transform 1 0 4816 0 1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_41
timestamp 1486834041
transform 1 0 5264 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_51
timestamp 1486834041
transform 1 0 6384 0 1 24304
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_59
timestamp 1486834041
transform 1 0 7280 0 1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_92
timestamp 1486834041
transform 1 0 10976 0 1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_96
timestamp 1486834041
transform 1 0 11424 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_98
timestamp 1486834041
transform 1 0 11648 0 1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_107
timestamp 1486834041
transform 1 0 12656 0 1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_160
timestamp 1486834041
transform 1 0 18592 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_170
timestamp 1486834041
transform 1 0 19712 0 1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_174
timestamp 1486834041
transform 1 0 20160 0 1 24304
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_177
timestamp 1486834041
transform 1 0 20496 0 1 24304
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_209
timestamp 1486834041
transform 1 0 24080 0 1 24304
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_2
timestamp 1486834041
transform 1 0 896 0 -1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_10
timestamp 1486834041
transform 1 0 1792 0 -1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_43
timestamp 1486834041
transform 1 0 5488 0 -1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_67
timestamp 1486834041
transform 1 0 8176 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_69
timestamp 1486834041
transform 1 0 8400 0 -1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_80
timestamp 1486834041
transform 1 0 9632 0 -1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_132
timestamp 1486834041
transform 1 0 15456 0 -1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_142
timestamp 1486834041
transform 1 0 16576 0 -1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_146
timestamp 1486834041
transform 1 0 17024 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_148
timestamp 1486834041
transform 1 0 17248 0 -1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_181
timestamp 1486834041
transform 1 0 20944 0 -1 25872
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_197
timestamp 1486834041
transform 1 0 22736 0 -1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_205
timestamp 1486834041
transform 1 0 23632 0 -1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_209
timestamp 1486834041
transform 1 0 24080 0 -1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_212
timestamp 1486834041
transform 1 0 24416 0 -1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_2
timestamp 1486834041
transform 1 0 896 0 1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_34
timestamp 1486834041
transform 1 0 4480 0 1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_37
timestamp 1486834041
transform 1 0 4816 0 1 25872
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_53
timestamp 1486834041
transform 1 0 6608 0 1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_57
timestamp 1486834041
transform 1 0 7056 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_79
timestamp 1486834041
transform 1 0 9520 0 1 25872
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_95
timestamp 1486834041
transform 1 0 11312 0 1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_103
timestamp 1486834041
transform 1 0 12208 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_115
timestamp 1486834041
transform 1 0 13552 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_117
timestamp 1486834041
transform 1 0 13776 0 1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_126
timestamp 1486834041
transform 1 0 14784 0 1 25872
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_134
timestamp 1486834041
transform 1 0 15680 0 1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_158
timestamp 1486834041
transform 1 0 18368 0 1 25872
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_162
timestamp 1486834041
transform 1 0 18816 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_172
timestamp 1486834041
transform 1 0 19936 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_174
timestamp 1486834041
transform 1 0 20160 0 1 25872
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_177
timestamp 1486834041
transform 1 0 20496 0 1 25872
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_209
timestamp 1486834041
transform 1 0 24080 0 1 25872
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_225
timestamp 1486834041
transform 1 0 25872 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_22
timestamp 1486834041
transform 1 0 3136 0 -1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_30
timestamp 1486834041
transform 1 0 4032 0 -1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_34
timestamp 1486834041
transform 1 0 4480 0 -1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_55
timestamp 1486834041
transform 1 0 6832 0 -1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_63
timestamp 1486834041
transform 1 0 7728 0 -1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_67
timestamp 1486834041
transform 1 0 8176 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_69
timestamp 1486834041
transform 1 0 8400 0 -1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_72
timestamp 1486834041
transform 1 0 8736 0 -1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_80
timestamp 1486834041
transform 1 0 9632 0 -1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_142
timestamp 1486834041
transform 1 0 16576 0 -1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_33_170
timestamp 1486834041
transform 1 0 19712 0 -1 27440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_202
timestamp 1486834041
transform 1 0 23296 0 -1 27440
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_212
timestamp 1486834041
transform 1 0 24416 0 -1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_10
timestamp 1486834041
transform 1 0 1792 0 1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_14
timestamp 1486834041
transform 1 0 2240 0 1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_69
timestamp 1486834041
transform 1 0 8400 0 1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_107
timestamp 1486834041
transform 1 0 12656 0 1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_111
timestamp 1486834041
transform 1 0 13104 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_113
timestamp 1486834041
transform 1 0 13328 0 1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_146
timestamp 1486834041
transform 1 0 17024 0 1 27440
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_177
timestamp 1486834041
transform 1 0 20496 0 1 27440
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_209
timestamp 1486834041
transform 1 0 24080 0 1 27440
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_72
timestamp 1486834041
transform 1 0 8736 0 -1 29008
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_142
timestamp 1486834041
transform 1 0 16576 0 -1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_150
timestamp 1486834041
transform 1 0 17472 0 -1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_154
timestamp 1486834041
transform 1 0 17920 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_156
timestamp 1486834041
transform 1 0 18144 0 -1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_189
timestamp 1486834041
transform 1 0 21840 0 -1 29008
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_205
timestamp 1486834041
transform 1 0 23632 0 -1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_209
timestamp 1486834041
transform 1 0 24080 0 -1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_212
timestamp 1486834041
transform 1 0 24416 0 -1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_220
timestamp 1486834041
transform 1 0 25312 0 -1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_224
timestamp 1486834041
transform 1 0 25760 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_226
timestamp 1486834041
transform 1 0 25984 0 -1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_22
timestamp 1486834041
transform 1 0 3136 0 1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_30
timestamp 1486834041
transform 1 0 4032 0 1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_34
timestamp 1486834041
transform 1 0 4480 0 1 29008
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_57
timestamp 1486834041
transform 1 0 7056 0 1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_65
timestamp 1486834041
transform 1 0 7952 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_87
timestamp 1486834041
transform 1 0 10416 0 1 29008
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_95
timestamp 1486834041
transform 1 0 11312 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_107
timestamp 1486834041
transform 1 0 12656 0 1 29008
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_111
timestamp 1486834041
transform 1 0 13104 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_173
timestamp 1486834041
transform 1 0 20048 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_177
timestamp 1486834041
transform 1 0 20496 0 1 29008
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_209
timestamp 1486834041
transform 1 0 24080 0 1 29008
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_225
timestamp 1486834041
transform 1 0 25872 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_24
timestamp 1486834041
transform 1 0 3360 0 -1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_32
timestamp 1486834041
transform 1 0 4256 0 -1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_36
timestamp 1486834041
transform 1 0 4704 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_72
timestamp 1486834041
transform 1 0 8736 0 -1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_76
timestamp 1486834041
transform 1 0 9184 0 -1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_109
timestamp 1486834041
transform 1 0 12880 0 -1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_117
timestamp 1486834041
transform 1 0 13776 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_127
timestamp 1486834041
transform 1 0 14896 0 -1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_131
timestamp 1486834041
transform 1 0 15344 0 -1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_162
timestamp 1486834041
transform 1 0 18816 0 -1 30576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_194
timestamp 1486834041
transform 1 0 22400 0 -1 30576
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_212
timestamp 1486834041
transform 1 0 24416 0 -1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_220
timestamp 1486834041
transform 1 0 25312 0 -1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_224
timestamp 1486834041
transform 1 0 25760 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_226
timestamp 1486834041
transform 1 0 25984 0 -1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_2
timestamp 1486834041
transform 1 0 896 0 1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_37
timestamp 1486834041
transform 1 0 4816 0 1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_45
timestamp 1486834041
transform 1 0 5712 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_47
timestamp 1486834041
transform 1 0 5936 0 1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_84
timestamp 1486834041
transform 1 0 10080 0 1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_93
timestamp 1486834041
transform 1 0 11088 0 1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_102
timestamp 1486834041
transform 1 0 12096 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_104
timestamp 1486834041
transform 1 0 12320 0 1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_107
timestamp 1486834041
transform 1 0 12656 0 1 30576
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_115
timestamp 1486834041
transform 1 0 13552 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_117
timestamp 1486834041
transform 1 0 13776 0 1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_138
timestamp 1486834041
transform 1 0 16128 0 1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_174
timestamp 1486834041
transform 1 0 20160 0 1 30576
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_177
timestamp 1486834041
transform 1 0 20496 0 1 30576
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_209
timestamp 1486834041
transform 1 0 24080 0 1 30576
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_2
timestamp 1486834041
transform 1 0 896 0 -1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_6
timestamp 1486834041
transform 1 0 1344 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_8
timestamp 1486834041
transform 1 0 1568 0 -1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_41
timestamp 1486834041
transform 1 0 5264 0 -1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_49
timestamp 1486834041
transform 1 0 6160 0 -1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_53
timestamp 1486834041
transform 1 0 6608 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_55
timestamp 1486834041
transform 1 0 6832 0 -1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_80
timestamp 1486834041
transform 1 0 9632 0 -1 32144
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_96
timestamp 1486834041
transform 1 0 11424 0 -1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_132
timestamp 1486834041
transform 1 0 15456 0 -1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_39_174
timestamp 1486834041
transform 1 0 20160 0 -1 32144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_206
timestamp 1486834041
transform 1 0 23744 0 -1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_212
timestamp 1486834041
transform 1 0 24416 0 -1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_2
timestamp 1486834041
transform 1 0 896 0 1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_34
timestamp 1486834041
transform 1 0 4480 0 1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_37
timestamp 1486834041
transform 1 0 4816 0 1 32144
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_45
timestamp 1486834041
transform 1 0 5712 0 1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_81
timestamp 1486834041
transform 1 0 9744 0 1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_107
timestamp 1486834041
transform 1 0 12656 0 1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_124
timestamp 1486834041
transform 1 0 14560 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_126
timestamp 1486834041
transform 1 0 14784 0 1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_170
timestamp 1486834041
transform 1 0 19712 0 1 32144
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_174
timestamp 1486834041
transform 1 0 20160 0 1 32144
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_177
timestamp 1486834041
transform 1 0 20496 0 1 32144
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_209
timestamp 1486834041
transform 1 0 24080 0 1 32144
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_225
timestamp 1486834041
transform 1 0 25872 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_22
timestamp 1486834041
transform 1 0 3136 0 -1 33712
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_38
timestamp 1486834041
transform 1 0 4928 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_40
timestamp 1486834041
transform 1 0 5152 0 -1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_69
timestamp 1486834041
transform 1 0 8400 0 -1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_72
timestamp 1486834041
transform 1 0 8736 0 -1 33712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_96
timestamp 1486834041
transform 1 0 11424 0 -1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_117
timestamp 1486834041
transform 1 0 13776 0 -1 33712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_121
timestamp 1486834041
transform 1 0 14224 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_131
timestamp 1486834041
transform 1 0 15344 0 -1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_139
timestamp 1486834041
transform 1 0 16240 0 -1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_142
timestamp 1486834041
transform 1 0 16576 0 -1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_41_171
timestamp 1486834041
transform 1 0 19824 0 -1 33712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_203
timestamp 1486834041
transform 1 0 23408 0 -1 33712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_207
timestamp 1486834041
transform 1 0 23856 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_209
timestamp 1486834041
transform 1 0 24080 0 -1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_212
timestamp 1486834041
transform 1 0 24416 0 -1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_2
timestamp 1486834041
transform 1 0 896 0 1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_57
timestamp 1486834041
transform 1 0 7056 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_79
timestamp 1486834041
transform 1 0 9520 0 1 33712
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_95
timestamp 1486834041
transform 1 0 11312 0 1 33712
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_103
timestamp 1486834041
transform 1 0 12208 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_107
timestamp 1486834041
transform 1 0 12656 0 1 33712
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_123
timestamp 1486834041
transform 1 0 14448 0 1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_174
timestamp 1486834041
transform 1 0 20160 0 1 33712
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_177
timestamp 1486834041
transform 1 0 20496 0 1 33712
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_209
timestamp 1486834041
transform 1 0 24080 0 1 33712
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_2
timestamp 1486834041
transform 1 0 896 0 -1 35280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_6
timestamp 1486834041
transform 1 0 1344 0 -1 35280
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_35
timestamp 1486834041
transform 1 0 4592 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_37
timestamp 1486834041
transform 1 0 4816 0 -1 35280
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_72
timestamp 1486834041
transform 1 0 8736 0 -1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_80
timestamp 1486834041
transform 1 0 9632 0 -1 35280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_84
timestamp 1486834041
transform 1 0 10080 0 -1 35280
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_137
timestamp 1486834041
transform 1 0 16016 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_139
timestamp 1486834041
transform 1 0 16240 0 -1 35280
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_43_178
timestamp 1486834041
transform 1 0 20608 0 -1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_212
timestamp 1486834041
transform 1 0 24416 0 -1 35280
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_2
timestamp 1486834041
transform 1 0 896 0 1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_10
timestamp 1486834041
transform 1 0 1792 0 1 35280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_14
timestamp 1486834041
transform 1 0 2240 0 1 35280
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_37
timestamp 1486834041
transform 1 0 4816 0 1 35280
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_41
timestamp 1486834041
transform 1 0 5264 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_103
timestamp 1486834041
transform 1 0 12208 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_165
timestamp 1486834041
transform 1 0 19152 0 1 35280
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_173
timestamp 1486834041
transform 1 0 20048 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_177
timestamp 1486834041
transform 1 0 20496 0 1 35280
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_209
timestamp 1486834041
transform 1 0 24080 0 1 35280
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_225
timestamp 1486834041
transform 1 0 25872 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_42
timestamp 1486834041
transform 1 0 5376 0 -1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_46
timestamp 1486834041
transform 1 0 5824 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_56
timestamp 1486834041
transform 1 0 6944 0 -1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_60
timestamp 1486834041
transform 1 0 7392 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_92
timestamp 1486834041
transform 1 0 10976 0 -1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_139
timestamp 1486834041
transform 1 0 16240 0 -1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_45_164
timestamp 1486834041
transform 1 0 19040 0 -1 36848
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_196
timestamp 1486834041
transform 1 0 22624 0 -1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_204
timestamp 1486834041
transform 1 0 23520 0 -1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_208
timestamp 1486834041
transform 1 0 23968 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_212
timestamp 1486834041
transform 1 0 24416 0 -1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_18
timestamp 1486834041
transform 1 0 2688 0 1 36848
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_34
timestamp 1486834041
transform 1 0 4480 0 1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_57
timestamp 1486834041
transform 1 0 7056 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_59
timestamp 1486834041
transform 1 0 7280 0 1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_92
timestamp 1486834041
transform 1 0 10976 0 1 36848
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_100
timestamp 1486834041
transform 1 0 11872 0 1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_104
timestamp 1486834041
transform 1 0 12320 0 1 36848
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_107
timestamp 1486834041
transform 1 0 12656 0 1 36848
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_123
timestamp 1486834041
transform 1 0 14448 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_46_177
timestamp 1486834041
transform 1 0 20496 0 1 36848
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_209
timestamp 1486834041
transform 1 0 24080 0 1 36848
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_22
timestamp 1486834041
transform 1 0 3136 0 -1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_30
timestamp 1486834041
transform 1 0 4032 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_32
timestamp 1486834041
transform 1 0 4256 0 -1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_61
timestamp 1486834041
transform 1 0 7504 0 -1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_72
timestamp 1486834041
transform 1 0 8736 0 -1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_134
timestamp 1486834041
transform 1 0 15680 0 -1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_138
timestamp 1486834041
transform 1 0 16128 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_178
timestamp 1486834041
transform 1 0 20608 0 -1 38416
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_212
timestamp 1486834041
transform 1 0 24416 0 -1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_2
timestamp 1486834041
transform 1 0 896 0 1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_6
timestamp 1486834041
transform 1 0 1344 0 1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_37
timestamp 1486834041
transform 1 0 4816 0 1 38416
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_61
timestamp 1486834041
transform 1 0 7504 0 1 38416
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_77
timestamp 1486834041
transform 1 0 9296 0 1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_107
timestamp 1486834041
transform 1 0 12656 0 1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_116
timestamp 1486834041
transform 1 0 13664 0 1 38416
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_124
timestamp 1486834041
transform 1 0 14560 0 1 38416
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_48_177
timestamp 1486834041
transform 1 0 20496 0 1 38416
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_209
timestamp 1486834041
transform 1 0 24080 0 1 38416
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_225
timestamp 1486834041
transform 1 0 25872 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_2
timestamp 1486834041
transform 1 0 896 0 -1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_6
timestamp 1486834041
transform 1 0 1344 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_24
timestamp 1486834041
transform 1 0 3360 0 -1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_32
timestamp 1486834041
transform 1 0 4256 0 -1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_36
timestamp 1486834041
transform 1 0 4704 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_72
timestamp 1486834041
transform 1 0 8736 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_74
timestamp 1486834041
transform 1 0 8960 0 -1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_127
timestamp 1486834041
transform 1 0 14896 0 -1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_135
timestamp 1486834041
transform 1 0 15792 0 -1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_139
timestamp 1486834041
transform 1 0 16240 0 -1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_192
timestamp 1486834041
transform 1 0 22176 0 -1 39984
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_208
timestamp 1486834041
transform 1 0 23968 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_212
timestamp 1486834041
transform 1 0 24416 0 -1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_2
timestamp 1486834041
transform 1 0 896 0 1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_6
timestamp 1486834041
transform 1 0 1344 0 1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_37
timestamp 1486834041
transform 1 0 4816 0 1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_45
timestamp 1486834041
transform 1 0 5712 0 1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_49
timestamp 1486834041
transform 1 0 6160 0 1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_90
timestamp 1486834041
transform 1 0 10752 0 1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_98
timestamp 1486834041
transform 1 0 11648 0 1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_102
timestamp 1486834041
transform 1 0 12096 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_104
timestamp 1486834041
transform 1 0 12320 0 1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_107
timestamp 1486834041
transform 1 0 12656 0 1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_116
timestamp 1486834041
transform 1 0 13664 0 1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_124
timestamp 1486834041
transform 1 0 14560 0 1 39984
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_161
timestamp 1486834041
transform 1 0 18704 0 1 39984
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_169
timestamp 1486834041
transform 1 0 19600 0 1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_173
timestamp 1486834041
transform 1 0 20048 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_177
timestamp 1486834041
transform 1 0 20496 0 1 39984
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_209
timestamp 1486834041
transform 1 0 24080 0 1 39984
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_2
timestamp 1486834041
transform 1 0 896 0 -1 41552
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_18
timestamp 1486834041
transform 1 0 2688 0 -1 41552
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_46
timestamp 1486834041
transform 1 0 5824 0 -1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_55
timestamp 1486834041
transform 1 0 6832 0 -1 41552
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_63
timestamp 1486834041
transform 1 0 7728 0 -1 41552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_67
timestamp 1486834041
transform 1 0 8176 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_69
timestamp 1486834041
transform 1 0 8400 0 -1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_80
timestamp 1486834041
transform 1 0 9632 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_51_102
timestamp 1486834041
transform 1 0 12096 0 -1 41552
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_134
timestamp 1486834041
transform 1 0 15680 0 -1 41552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_138
timestamp 1486834041
transform 1 0 16128 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_142
timestamp 1486834041
transform 1 0 16576 0 -1 41552
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_206
timestamp 1486834041
transform 1 0 23744 0 -1 41552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_212
timestamp 1486834041
transform 1 0 24416 0 -1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_2
timestamp 1486834041
transform 1 0 896 0 1 41552
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_18
timestamp 1486834041
transform 1 0 2688 0 1 41552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_22
timestamp 1486834041
transform 1 0 3136 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_24
timestamp 1486834041
transform 1 0 3360 0 1 41552
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_33
timestamp 1486834041
transform 1 0 4368 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_37
timestamp 1486834041
transform 1 0 4816 0 1 41552
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_101
timestamp 1486834041
transform 1 0 11984 0 1 41552
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_107
timestamp 1486834041
transform 1 0 12656 0 1 41552
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_123
timestamp 1486834041
transform 1 0 14448 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_52_177
timestamp 1486834041
transform 1 0 20496 0 1 41552
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_209
timestamp 1486834041
transform 1 0 24080 0 1 41552
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_225
timestamp 1486834041
transform 1 0 25872 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_2
timestamp 1486834041
transform 1 0 896 0 -1 43120
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_66
timestamp 1486834041
transform 1 0 8064 0 -1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_72
timestamp 1486834041
transform 1 0 8736 0 -1 43120
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_136
timestamp 1486834041
transform 1 0 15904 0 -1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_142
timestamp 1486834041
transform 1 0 16576 0 -1 43120
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_206
timestamp 1486834041
transform 1 0 23744 0 -1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_212
timestamp 1486834041
transform 1 0 24416 0 -1 43120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_2
timestamp 1486834041
transform 1 0 896 0 1 43120
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_34
timestamp 1486834041
transform 1 0 4480 0 1 43120
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_37
timestamp 1486834041
transform 1 0 4816 0 1 43120
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_101
timestamp 1486834041
transform 1 0 11984 0 1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_107
timestamp 1486834041
transform 1 0 12656 0 1 43120
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_171
timestamp 1486834041
transform 1 0 19824 0 1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_177
timestamp 1486834041
transform 1 0 20496 0 1 43120
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_209
timestamp 1486834041
transform 1 0 24080 0 1 43120
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_2
timestamp 1486834041
transform 1 0 896 0 -1 44688
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_66
timestamp 1486834041
transform 1 0 8064 0 -1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_72
timestamp 1486834041
transform 1 0 8736 0 -1 44688
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_136
timestamp 1486834041
transform 1 0 15904 0 -1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_142
timestamp 1486834041
transform 1 0 16576 0 -1 44688
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_206
timestamp 1486834041
transform 1 0 23744 0 -1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_212
timestamp 1486834041
transform 1 0 24416 0 -1 44688
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_56_2
timestamp 1486834041
transform 1 0 896 0 1 44688
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_34
timestamp 1486834041
transform 1 0 4480 0 1 44688
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_37
timestamp 1486834041
transform 1 0 4816 0 1 44688
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_101
timestamp 1486834041
transform 1 0 11984 0 1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_107
timestamp 1486834041
transform 1 0 12656 0 1 44688
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_171
timestamp 1486834041
transform 1 0 19824 0 1 44688
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_56_177
timestamp 1486834041
transform 1 0 20496 0 1 44688
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_56_209
timestamp 1486834041
transform 1 0 24080 0 1 44688
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_225
timestamp 1486834041
transform 1 0 25872 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_2
timestamp 1486834041
transform 1 0 896 0 -1 46256
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_66
timestamp 1486834041
transform 1 0 8064 0 -1 46256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_72
timestamp 1486834041
transform 1 0 8736 0 -1 46256
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_136
timestamp 1486834041
transform 1 0 15904 0 -1 46256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_142
timestamp 1486834041
transform 1 0 16576 0 -1 46256
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_206
timestamp 1486834041
transform 1 0 23744 0 -1 46256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_212
timestamp 1486834041
transform 1 0 24416 0 -1 46256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_58_2
timestamp 1486834041
transform 1 0 896 0 1 46256
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_34
timestamp 1486834041
transform 1 0 4480 0 1 46256
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_37
timestamp 1486834041
transform 1 0 4816 0 1 46256
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_101
timestamp 1486834041
transform 1 0 11984 0 1 46256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_107
timestamp 1486834041
transform 1 0 12656 0 1 46256
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_171
timestamp 1486834041
transform 1 0 19824 0 1 46256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_58_177
timestamp 1486834041
transform 1 0 20496 0 1 46256
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_209
timestamp 1486834041
transform 1 0 24080 0 1 46256
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_2
timestamp 1486834041
transform 1 0 896 0 -1 47824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_66
timestamp 1486834041
transform 1 0 8064 0 -1 47824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_72
timestamp 1486834041
transform 1 0 8736 0 -1 47824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_136
timestamp 1486834041
transform 1 0 15904 0 -1 47824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_142
timestamp 1486834041
transform 1 0 16576 0 -1 47824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_206
timestamp 1486834041
transform 1 0 23744 0 -1 47824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_212
timestamp 1486834041
transform 1 0 24416 0 -1 47824
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_2
timestamp 1486834041
transform 1 0 896 0 1 47824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_34
timestamp 1486834041
transform 1 0 4480 0 1 47824
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_37
timestamp 1486834041
transform 1 0 4816 0 1 47824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_101
timestamp 1486834041
transform 1 0 11984 0 1 47824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_107
timestamp 1486834041
transform 1 0 12656 0 1 47824
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_171
timestamp 1486834041
transform 1 0 19824 0 1 47824
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_177
timestamp 1486834041
transform 1 0 20496 0 1 47824
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_209
timestamp 1486834041
transform 1 0 24080 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_2
timestamp 1486834041
transform 1 0 896 0 -1 49392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_66
timestamp 1486834041
transform 1 0 8064 0 -1 49392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_72
timestamp 1486834041
transform 1 0 8736 0 -1 49392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_136
timestamp 1486834041
transform 1 0 15904 0 -1 49392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_142
timestamp 1486834041
transform 1 0 16576 0 -1 49392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_206
timestamp 1486834041
transform 1 0 23744 0 -1 49392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_212
timestamp 1486834041
transform 1 0 24416 0 -1 49392
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_62_2
timestamp 1486834041
transform 1 0 896 0 1 49392
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_34
timestamp 1486834041
transform 1 0 4480 0 1 49392
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_37
timestamp 1486834041
transform 1 0 4816 0 1 49392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_101
timestamp 1486834041
transform 1 0 11984 0 1 49392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_107
timestamp 1486834041
transform 1 0 12656 0 1 49392
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_171
timestamp 1486834041
transform 1 0 19824 0 1 49392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_62_177
timestamp 1486834041
transform 1 0 20496 0 1 49392
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_193
timestamp 1486834041
transform 1 0 22288 0 1 49392
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_201
timestamp 1486834041
transform 1 0 23184 0 1 49392
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_2
timestamp 1486834041
transform 1 0 896 0 -1 50960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_66
timestamp 1486834041
transform 1 0 8064 0 -1 50960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_72
timestamp 1486834041
transform 1 0 8736 0 -1 50960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_136
timestamp 1486834041
transform 1 0 15904 0 -1 50960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_63_142
timestamp 1486834041
transform 1 0 16576 0 -1 50960
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_63_174
timestamp 1486834041
transform 1 0 20160 0 -1 50960
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_190
timestamp 1486834041
transform 1 0 21952 0 -1 50960
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_198
timestamp 1486834041
transform 1 0 22848 0 -1 50960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_212
timestamp 1486834041
transform 1 0 24416 0 -1 50960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_64_2
timestamp 1486834041
transform 1 0 896 0 1 50960
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_34
timestamp 1486834041
transform 1 0 4480 0 1 50960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_37
timestamp 1486834041
transform 1 0 4816 0 1 50960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_101
timestamp 1486834041
transform 1 0 11984 0 1 50960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_107
timestamp 1486834041
transform 1 0 12656 0 1 50960
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_171
timestamp 1486834041
transform 1 0 19824 0 1 50960
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_64_177
timestamp 1486834041
transform 1 0 20496 0 1 50960
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_193
timestamp 1486834041
transform 1 0 22288 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_195
timestamp 1486834041
transform 1 0 22512 0 1 50960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_204
timestamp 1486834041
transform 1 0 23520 0 1 50960
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_2
timestamp 1486834041
transform 1 0 896 0 -1 52528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_66
timestamp 1486834041
transform 1 0 8064 0 -1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_72
timestamp 1486834041
transform 1 0 8736 0 -1 52528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_136
timestamp 1486834041
transform 1 0 15904 0 -1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_65_142
timestamp 1486834041
transform 1 0 16576 0 -1 52528
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_174
timestamp 1486834041
transform 1 0 20160 0 -1 52528
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_182
timestamp 1486834041
transform 1 0 21056 0 -1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_186
timestamp 1486834041
transform 1 0 21504 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_212
timestamp 1486834041
transform 1 0 24416 0 -1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_66_2
timestamp 1486834041
transform 1 0 896 0 1 52528
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_34
timestamp 1486834041
transform 1 0 4480 0 1 52528
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_37
timestamp 1486834041
transform 1 0 4816 0 1 52528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_101
timestamp 1486834041
transform 1 0 11984 0 1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_107
timestamp 1486834041
transform 1 0 12656 0 1 52528
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_171
timestamp 1486834041
transform 1 0 19824 0 1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_177
timestamp 1486834041
transform 1 0 20496 0 1 52528
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_181
timestamp 1486834041
transform 1 0 20944 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_2
timestamp 1486834041
transform 1 0 896 0 -1 54096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_66
timestamp 1486834041
transform 1 0 8064 0 -1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_72
timestamp 1486834041
transform 1 0 8736 0 -1 54096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_136
timestamp 1486834041
transform 1 0 15904 0 -1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_142
timestamp 1486834041
transform 1 0 16576 0 -1 54096
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_158
timestamp 1486834041
transform 1 0 18368 0 -1 54096
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_166
timestamp 1486834041
transform 1 0 19264 0 -1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_170
timestamp 1486834041
transform 1 0 19712 0 -1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_195
timestamp 1486834041
transform 1 0 22512 0 -1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_212
timestamp 1486834041
transform 1 0 24416 0 -1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_68_2
timestamp 1486834041
transform 1 0 896 0 1 54096
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_34
timestamp 1486834041
transform 1 0 4480 0 1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_37
timestamp 1486834041
transform 1 0 4816 0 1 54096
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_101
timestamp 1486834041
transform 1 0 11984 0 1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_68_107
timestamp 1486834041
transform 1 0 12656 0 1 54096
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_68_139
timestamp 1486834041
transform 1 0 16240 0 1 54096
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_155
timestamp 1486834041
transform 1 0 18032 0 1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_159
timestamp 1486834041
transform 1 0 18480 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_161
timestamp 1486834041
transform 1 0 18704 0 1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_170
timestamp 1486834041
transform 1 0 19712 0 1 54096
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_174
timestamp 1486834041
transform 1 0 20160 0 1 54096
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_69_2
timestamp 1486834041
transform 1 0 896 0 -1 55664
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_10
timestamp 1486834041
transform 1 0 1792 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_12
timestamp 1486834041
transform 1 0 2016 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_69_27
timestamp 1486834041
transform 1 0 3696 0 -1 55664
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_43
timestamp 1486834041
transform 1 0 5488 0 -1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_47
timestamp 1486834041
transform 1 0 5936 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_63
timestamp 1486834041
transform 1 0 7728 0 -1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_67
timestamp 1486834041
transform 1 0 8176 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_69
timestamp 1486834041
transform 1 0 8400 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_69_72
timestamp 1486834041
transform 1 0 8736 0 -1 55664
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_69_88
timestamp 1486834041
transform 1 0 10528 0 -1 55664
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_96
timestamp 1486834041
transform 1 0 11424 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_69_111
timestamp 1486834041
transform 1 0 13104 0 -1 55664
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_69_127
timestamp 1486834041
transform 1 0 14896 0 -1 55664
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_135
timestamp 1486834041
transform 1 0 15792 0 -1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_139
timestamp 1486834041
transform 1 0 16240 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_142
timestamp 1486834041
transform 1 0 16576 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_144
timestamp 1486834041
transform 1 0 16800 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_159
timestamp 1486834041
transform 1 0 18480 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_169
timestamp 1486834041
transform 1 0 19600 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_207
timestamp 1486834041
transform 1 0 23856 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_209
timestamp 1486834041
transform 1 0 24080 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_212
timestamp 1486834041
transform 1 0 24416 0 -1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_70_8
timestamp 1486834041
transform 1 0 1568 0 1 55664
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_16
timestamp 1486834041
transform 1 0 2464 0 1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_36
timestamp 1486834041
transform 1 0 4704 0 1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_51
timestamp 1486834041
transform 1 0 6384 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_53
timestamp 1486834041
transform 1 0 6608 0 1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_70
timestamp 1486834041
transform 1 0 8512 0 1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_99
timestamp 1486834041
transform 1 0 11760 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_101
timestamp 1486834041
transform 1 0 11984 0 1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_104
timestamp 1486834041
transform 1 0 12320 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_106
timestamp 1486834041
transform 1 0 12544 0 1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_135
timestamp 1486834041
transform 1 0 15792 0 1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_152
timestamp 1486834041
transform 1 0 17696 0 1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_200
timestamp 1486834041
transform 1 0 23072 0 1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_234
timestamp 1486834041
transform 1 0 26880 0 1 55664
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_240
timestamp 1486834041
transform 1 0 27552 0 1 55664
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output1
timestamp 1486834041
transform -1 0 2464 0 1 5488
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output2
timestamp 1486834041
transform -1 0 2464 0 -1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output3
timestamp 1486834041
transform -1 0 2464 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output4
timestamp 1486834041
transform -1 0 2464 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output5
timestamp 1486834041
transform 1 0 24528 0 -1 22736
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output6
timestamp 1486834041
transform 1 0 26096 0 1 21168
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output7
timestamp 1486834041
transform 1 0 26096 0 -1 22736
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output8
timestamp 1486834041
transform 1 0 24528 0 -1 24304
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output9
timestamp 1486834041
transform 1 0 26096 0 1 22736
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output10
timestamp 1486834041
transform 1 0 24528 0 1 24304
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output11
timestamp 1486834041
transform 1 0 26096 0 -1 24304
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output12
timestamp 1486834041
transform 1 0 24528 0 -1 25872
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output13
timestamp 1486834041
transform 1 0 26096 0 1 24304
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output14
timestamp 1486834041
transform 1 0 26096 0 -1 25872
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output15
timestamp 1486834041
transform 1 0 24528 0 -1 27440
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output16
timestamp 1486834041
transform 1 0 26096 0 1 25872
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output17
timestamp 1486834041
transform 1 0 24528 0 1 27440
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output18
timestamp 1486834041
transform 1 0 26096 0 -1 27440
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output19
timestamp 1486834041
transform 1 0 26096 0 1 27440
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output20
timestamp 1486834041
transform 1 0 26096 0 -1 29008
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output21
timestamp 1486834041
transform 1 0 26096 0 1 29008
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output22
timestamp 1486834041
transform 1 0 26096 0 -1 30576
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output23
timestamp 1486834041
transform 1 0 26096 0 1 30576
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output24
timestamp 1486834041
transform 1 0 26096 0 -1 32144
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output25
timestamp 1486834041
transform 1 0 24528 0 -1 38416
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output26
timestamp 1486834041
transform 1 0 24528 0 -1 43120
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output27
timestamp 1486834041
transform 1 0 26096 0 -1 44688
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output28
timestamp 1486834041
transform 1 0 26096 0 -1 39984
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output29
timestamp 1486834041
transform 1 0 26096 0 1 39984
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output30
timestamp 1486834041
transform 1 0 24528 0 -1 39984
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output31
timestamp 1486834041
transform 1 0 26096 0 -1 41552
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output32
timestamp 1486834041
transform 1 0 24528 0 1 39984
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output33
timestamp 1486834041
transform 1 0 26096 0 1 41552
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output34
timestamp 1486834041
transform 1 0 24528 0 -1 41552
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output35
timestamp 1486834041
transform 1 0 26096 0 -1 43120
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output36
timestamp 1486834041
transform 1 0 26096 0 1 43120
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output37
timestamp 1486834041
transform 1 0 24528 0 1 30576
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output38
timestamp 1486834041
transform 1 0 26096 0 -1 36848
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output39
timestamp 1486834041
transform 1 0 26096 0 1 36848
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output40
timestamp 1486834041
transform 1 0 24528 0 -1 36848
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output41
timestamp 1486834041
transform 1 0 26096 0 -1 38416
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output42
timestamp 1486834041
transform 1 0 24528 0 1 36848
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output43
timestamp 1486834041
transform 1 0 26096 0 1 38416
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output44
timestamp 1486834041
transform 1 0 26096 0 1 32144
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output45
timestamp 1486834041
transform 1 0 24528 0 -1 32144
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output46
timestamp 1486834041
transform 1 0 26096 0 -1 33712
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output47
timestamp 1486834041
transform 1 0 26096 0 1 33712
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output48
timestamp 1486834041
transform 1 0 24528 0 -1 33712
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output49
timestamp 1486834041
transform 1 0 26096 0 -1 35280
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output50
timestamp 1486834041
transform 1 0 24528 0 1 33712
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output51
timestamp 1486834041
transform 1 0 26096 0 1 35280
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output52
timestamp 1486834041
transform 1 0 24528 0 -1 35280
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output53
timestamp 1486834041
transform 1 0 24528 0 1 43120
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output54
timestamp 1486834041
transform 1 0 26096 0 -1 49392
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output55
timestamp 1486834041
transform 1 0 26096 0 1 49392
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output56
timestamp 1486834041
transform 1 0 24528 0 -1 49392
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output57
timestamp 1486834041
transform 1 0 26096 0 -1 50960
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output58
timestamp 1486834041
transform 1 0 24528 0 1 49392
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output59
timestamp 1486834041
transform 1 0 26096 0 1 50960
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output60
timestamp 1486834041
transform 1 0 24528 0 -1 50960
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output61
timestamp 1486834041
transform 1 0 26096 0 -1 52528
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output62
timestamp 1486834041
transform 1 0 26096 0 1 52528
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output63
timestamp 1486834041
transform 1 0 24528 0 -1 52528
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output64
timestamp 1486834041
transform 1 0 26096 0 1 44688
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output65
timestamp 1486834041
transform 1 0 26096 0 -1 54096
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output66
timestamp 1486834041
transform 1 0 24528 0 1 52528
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output67
timestamp 1486834041
transform 1 0 26096 0 1 54096
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output68
timestamp 1486834041
transform 1 0 24528 0 -1 54096
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output69
timestamp 1486834041
transform 1 0 26096 0 -1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output70
timestamp 1486834041
transform 1 0 24528 0 -1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output71
timestamp 1486834041
transform 1 0 22960 0 1 54096
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output72
timestamp 1486834041
transform 1 0 22624 0 -1 54096
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output73
timestamp 1486834041
transform 1 0 20720 0 -1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output74
timestamp 1486834041
transform 1 0 21392 0 1 54096
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output75
timestamp 1486834041
transform 1 0 24528 0 -1 44688
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output76
timestamp 1486834041
transform 1 0 24528 0 1 50960
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output77
timestamp 1486834041
transform 1 0 22960 0 1 52528
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output78
timestamp 1486834041
transform 1 0 26096 0 -1 46256
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output79
timestamp 1486834041
transform 1 0 26096 0 1 46256
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output80
timestamp 1486834041
transform 1 0 24528 0 -1 46256
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output81
timestamp 1486834041
transform 1 0 26096 0 -1 47824
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output82
timestamp 1486834041
transform 1 0 24528 0 1 46256
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output83
timestamp 1486834041
transform 1 0 26096 0 1 47824
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output84
timestamp 1486834041
transform 1 0 24528 0 -1 47824
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output85
timestamp 1486834041
transform -1 0 3696 0 -1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output86
timestamp 1486834041
transform -1 0 17696 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output87
timestamp 1486834041
transform -1 0 18480 0 -1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output88
timestamp 1486834041
transform -1 0 19712 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output89
timestamp 1486834041
transform 1 0 19936 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output90
timestamp 1486834041
transform -1 0 23072 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output91
timestamp 1486834041
transform -1 0 23856 0 -1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output92
timestamp 1486834041
transform 1 0 23744 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output93
timestamp 1486834041
transform 1 0 25312 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output94
timestamp 1486834041
transform 1 0 24528 0 1 54096
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output95
timestamp 1486834041
transform 1 0 22624 0 -1 52528
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output96
timestamp 1486834041
transform 1 0 2912 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output97
timestamp 1486834041
transform 1 0 4816 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output98
timestamp 1486834041
transform -1 0 7728 0 -1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output99
timestamp 1486834041
transform -1 0 8288 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output100
timestamp 1486834041
transform -1 0 10192 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output101
timestamp 1486834041
transform -1 0 11760 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output102
timestamp 1486834041
transform -1 0 13104 0 -1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output103
timestamp 1486834041
transform -1 0 14224 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output104
timestamp 1486834041
transform -1 0 15792 0 1 55664
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output105
timestamp 1486834041
transform -1 0 1568 0 1 55664
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_71
timestamp 1486834041
transform 1 0 672 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1486834041
transform -1 0 27888 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_72
timestamp 1486834041
transform 1 0 672 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1486834041
transform -1 0 27888 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_73
timestamp 1486834041
transform 1 0 672 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1486834041
transform -1 0 27888 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_74
timestamp 1486834041
transform 1 0 672 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1486834041
transform -1 0 27888 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_75
timestamp 1486834041
transform 1 0 672 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1486834041
transform -1 0 27888 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_76
timestamp 1486834041
transform 1 0 672 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1486834041
transform -1 0 27888 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_77
timestamp 1486834041
transform 1 0 672 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1486834041
transform -1 0 27888 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_78
timestamp 1486834041
transform 1 0 672 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1486834041
transform -1 0 27888 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_79
timestamp 1486834041
transform 1 0 672 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1486834041
transform -1 0 27888 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_80
timestamp 1486834041
transform 1 0 672 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1486834041
transform -1 0 27888 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_81
timestamp 1486834041
transform 1 0 672 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1486834041
transform -1 0 27888 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_82
timestamp 1486834041
transform 1 0 672 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1486834041
transform -1 0 27888 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_83
timestamp 1486834041
transform 1 0 672 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1486834041
transform -1 0 27888 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_84
timestamp 1486834041
transform 1 0 672 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1486834041
transform -1 0 27888 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_85
timestamp 1486834041
transform 1 0 672 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1486834041
transform -1 0 27888 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_86
timestamp 1486834041
transform 1 0 672 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1486834041
transform -1 0 27888 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_87
timestamp 1486834041
transform 1 0 672 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1486834041
transform -1 0 27888 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_88
timestamp 1486834041
transform 1 0 672 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1486834041
transform -1 0 27888 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_89
timestamp 1486834041
transform 1 0 672 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1486834041
transform -1 0 27888 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_90
timestamp 1486834041
transform 1 0 672 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1486834041
transform -1 0 27888 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_91
timestamp 1486834041
transform 1 0 672 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1486834041
transform -1 0 27888 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_92
timestamp 1486834041
transform 1 0 672 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1486834041
transform -1 0 27888 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_93
timestamp 1486834041
transform 1 0 672 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1486834041
transform -1 0 27888 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_94
timestamp 1486834041
transform 1 0 672 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1486834041
transform -1 0 27888 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_95
timestamp 1486834041
transform 1 0 672 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1486834041
transform -1 0 27888 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_96
timestamp 1486834041
transform 1 0 672 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1486834041
transform -1 0 27888 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_97
timestamp 1486834041
transform 1 0 672 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1486834041
transform -1 0 27888 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_98
timestamp 1486834041
transform 1 0 672 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1486834041
transform -1 0 27888 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_99
timestamp 1486834041
transform 1 0 672 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1486834041
transform -1 0 27888 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_100
timestamp 1486834041
transform 1 0 672 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1486834041
transform -1 0 27888 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_101
timestamp 1486834041
transform 1 0 672 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1486834041
transform -1 0 27888 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_102
timestamp 1486834041
transform 1 0 672 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1486834041
transform -1 0 27888 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_103
timestamp 1486834041
transform 1 0 672 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1486834041
transform -1 0 27888 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_104
timestamp 1486834041
transform 1 0 672 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1486834041
transform -1 0 27888 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_105
timestamp 1486834041
transform 1 0 672 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1486834041
transform -1 0 27888 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_106
timestamp 1486834041
transform 1 0 672 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1486834041
transform -1 0 27888 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_107
timestamp 1486834041
transform 1 0 672 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1486834041
transform -1 0 27888 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_108
timestamp 1486834041
transform 1 0 672 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1486834041
transform -1 0 27888 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_109
timestamp 1486834041
transform 1 0 672 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1486834041
transform -1 0 27888 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_110
timestamp 1486834041
transform 1 0 672 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1486834041
transform -1 0 27888 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_111
timestamp 1486834041
transform 1 0 672 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1486834041
transform -1 0 27888 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_112
timestamp 1486834041
transform 1 0 672 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1486834041
transform -1 0 27888 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_113
timestamp 1486834041
transform 1 0 672 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1486834041
transform -1 0 27888 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_114
timestamp 1486834041
transform 1 0 672 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1486834041
transform -1 0 27888 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_115
timestamp 1486834041
transform 1 0 672 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1486834041
transform -1 0 27888 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_116
timestamp 1486834041
transform 1 0 672 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1486834041
transform -1 0 27888 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_117
timestamp 1486834041
transform 1 0 672 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1486834041
transform -1 0 27888 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_118
timestamp 1486834041
transform 1 0 672 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1486834041
transform -1 0 27888 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_119
timestamp 1486834041
transform 1 0 672 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1486834041
transform -1 0 27888 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_120
timestamp 1486834041
transform 1 0 672 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1486834041
transform -1 0 27888 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_121
timestamp 1486834041
transform 1 0 672 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1486834041
transform -1 0 27888 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_122
timestamp 1486834041
transform 1 0 672 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1486834041
transform -1 0 27888 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_123
timestamp 1486834041
transform 1 0 672 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1486834041
transform -1 0 27888 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_124
timestamp 1486834041
transform 1 0 672 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1486834041
transform -1 0 27888 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_125
timestamp 1486834041
transform 1 0 672 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1486834041
transform -1 0 27888 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_126
timestamp 1486834041
transform 1 0 672 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1486834041
transform -1 0 27888 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_127
timestamp 1486834041
transform 1 0 672 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1486834041
transform -1 0 27888 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_128
timestamp 1486834041
transform 1 0 672 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1486834041
transform -1 0 27888 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_129
timestamp 1486834041
transform 1 0 672 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1486834041
transform -1 0 27888 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_130
timestamp 1486834041
transform 1 0 672 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1486834041
transform -1 0 27888 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_131
timestamp 1486834041
transform 1 0 672 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1486834041
transform -1 0 27888 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_132
timestamp 1486834041
transform 1 0 672 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1486834041
transform -1 0 27888 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Left_133
timestamp 1486834041
transform 1 0 672 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Right_62
timestamp 1486834041
transform -1 0 27888 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Left_134
timestamp 1486834041
transform 1 0 672 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Right_63
timestamp 1486834041
transform -1 0 27888 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Left_135
timestamp 1486834041
transform 1 0 672 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Right_64
timestamp 1486834041
transform -1 0 27888 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Left_136
timestamp 1486834041
transform 1 0 672 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Right_65
timestamp 1486834041
transform -1 0 27888 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Left_137
timestamp 1486834041
transform 1 0 672 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Right_66
timestamp 1486834041
transform -1 0 27888 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Left_138
timestamp 1486834041
transform 1 0 672 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Right_67
timestamp 1486834041
transform -1 0 27888 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Left_139
timestamp 1486834041
transform 1 0 672 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Right_68
timestamp 1486834041
transform -1 0 27888 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Left_140
timestamp 1486834041
transform 1 0 672 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Right_69
timestamp 1486834041
transform -1 0 27888 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Left_141
timestamp 1486834041
transform 1 0 672 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Right_70
timestamp 1486834041
transform -1 0 27888 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_142
timestamp 1486834041
transform 1 0 4480 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_143
timestamp 1486834041
transform 1 0 8288 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_144
timestamp 1486834041
transform 1 0 12096 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_145
timestamp 1486834041
transform 1 0 15904 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_146
timestamp 1486834041
transform 1 0 19712 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_147
timestamp 1486834041
transform 1 0 23520 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_148
timestamp 1486834041
transform 1 0 27328 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_149
timestamp 1486834041
transform 1 0 8512 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_150
timestamp 1486834041
transform 1 0 16352 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_151
timestamp 1486834041
transform 1 0 24192 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_152
timestamp 1486834041
transform 1 0 4592 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_153
timestamp 1486834041
transform 1 0 12432 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_154
timestamp 1486834041
transform 1 0 20272 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_155
timestamp 1486834041
transform 1 0 8512 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_156
timestamp 1486834041
transform 1 0 16352 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_157
timestamp 1486834041
transform 1 0 24192 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_158
timestamp 1486834041
transform 1 0 4592 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_159
timestamp 1486834041
transform 1 0 12432 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_160
timestamp 1486834041
transform 1 0 20272 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_161
timestamp 1486834041
transform 1 0 8512 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_162
timestamp 1486834041
transform 1 0 16352 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_163
timestamp 1486834041
transform 1 0 24192 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_164
timestamp 1486834041
transform 1 0 4592 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_165
timestamp 1486834041
transform 1 0 12432 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_166
timestamp 1486834041
transform 1 0 20272 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_167
timestamp 1486834041
transform 1 0 8512 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_168
timestamp 1486834041
transform 1 0 16352 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_169
timestamp 1486834041
transform 1 0 24192 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_170
timestamp 1486834041
transform 1 0 4592 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_171
timestamp 1486834041
transform 1 0 12432 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_172
timestamp 1486834041
transform 1 0 20272 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_173
timestamp 1486834041
transform 1 0 8512 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_174
timestamp 1486834041
transform 1 0 16352 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_175
timestamp 1486834041
transform 1 0 24192 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_176
timestamp 1486834041
transform 1 0 4592 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_177
timestamp 1486834041
transform 1 0 12432 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_178
timestamp 1486834041
transform 1 0 20272 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_179
timestamp 1486834041
transform 1 0 8512 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_180
timestamp 1486834041
transform 1 0 16352 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_181
timestamp 1486834041
transform 1 0 24192 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_182
timestamp 1486834041
transform 1 0 4592 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_183
timestamp 1486834041
transform 1 0 12432 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_184
timestamp 1486834041
transform 1 0 20272 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_185
timestamp 1486834041
transform 1 0 8512 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_186
timestamp 1486834041
transform 1 0 16352 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_187
timestamp 1486834041
transform 1 0 24192 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_188
timestamp 1486834041
transform 1 0 4592 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_189
timestamp 1486834041
transform 1 0 12432 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_190
timestamp 1486834041
transform 1 0 20272 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_191
timestamp 1486834041
transform 1 0 8512 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_192
timestamp 1486834041
transform 1 0 16352 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_193
timestamp 1486834041
transform 1 0 24192 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_194
timestamp 1486834041
transform 1 0 4592 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_195
timestamp 1486834041
transform 1 0 12432 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_196
timestamp 1486834041
transform 1 0 20272 0 1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_197
timestamp 1486834041
transform 1 0 8512 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_198
timestamp 1486834041
transform 1 0 16352 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_199
timestamp 1486834041
transform 1 0 24192 0 -1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_200
timestamp 1486834041
transform 1 0 4592 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_201
timestamp 1486834041
transform 1 0 12432 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_202
timestamp 1486834041
transform 1 0 20272 0 1 14896
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_203
timestamp 1486834041
transform 1 0 8512 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_204
timestamp 1486834041
transform 1 0 16352 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_205
timestamp 1486834041
transform 1 0 24192 0 -1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_206
timestamp 1486834041
transform 1 0 4592 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_207
timestamp 1486834041
transform 1 0 12432 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_208
timestamp 1486834041
transform 1 0 20272 0 1 16464
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_209
timestamp 1486834041
transform 1 0 8512 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_210
timestamp 1486834041
transform 1 0 16352 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_211
timestamp 1486834041
transform 1 0 24192 0 -1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_212
timestamp 1486834041
transform 1 0 4592 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_213
timestamp 1486834041
transform 1 0 12432 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_214
timestamp 1486834041
transform 1 0 20272 0 1 18032
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_215
timestamp 1486834041
transform 1 0 8512 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_216
timestamp 1486834041
transform 1 0 16352 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_217
timestamp 1486834041
transform 1 0 24192 0 -1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_218
timestamp 1486834041
transform 1 0 4592 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_219
timestamp 1486834041
transform 1 0 12432 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_220
timestamp 1486834041
transform 1 0 20272 0 1 19600
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_221
timestamp 1486834041
transform 1 0 8512 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_222
timestamp 1486834041
transform 1 0 16352 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_223
timestamp 1486834041
transform 1 0 24192 0 -1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_224
timestamp 1486834041
transform 1 0 4592 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_225
timestamp 1486834041
transform 1 0 12432 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_226
timestamp 1486834041
transform 1 0 20272 0 1 21168
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_227
timestamp 1486834041
transform 1 0 8512 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_228
timestamp 1486834041
transform 1 0 16352 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_229
timestamp 1486834041
transform 1 0 24192 0 -1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_230
timestamp 1486834041
transform 1 0 4592 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_231
timestamp 1486834041
transform 1 0 12432 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_232
timestamp 1486834041
transform 1 0 20272 0 1 22736
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_233
timestamp 1486834041
transform 1 0 8512 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_234
timestamp 1486834041
transform 1 0 16352 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_235
timestamp 1486834041
transform 1 0 24192 0 -1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_236
timestamp 1486834041
transform 1 0 4592 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_237
timestamp 1486834041
transform 1 0 12432 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_238
timestamp 1486834041
transform 1 0 20272 0 1 24304
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_239
timestamp 1486834041
transform 1 0 8512 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_240
timestamp 1486834041
transform 1 0 16352 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_241
timestamp 1486834041
transform 1 0 24192 0 -1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1486834041
transform 1 0 4592 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1486834041
transform 1 0 12432 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_244
timestamp 1486834041
transform 1 0 20272 0 1 25872
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1486834041
transform 1 0 8512 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1486834041
transform 1 0 16352 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1486834041
transform 1 0 24192 0 -1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1486834041
transform 1 0 4592 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1486834041
transform 1 0 12432 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1486834041
transform 1 0 20272 0 1 27440
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_251
timestamp 1486834041
transform 1 0 8512 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_252
timestamp 1486834041
transform 1 0 16352 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1486834041
transform 1 0 24192 0 -1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_254
timestamp 1486834041
transform 1 0 4592 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_255
timestamp 1486834041
transform 1 0 12432 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_256
timestamp 1486834041
transform 1 0 20272 0 1 29008
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_257
timestamp 1486834041
transform 1 0 8512 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_258
timestamp 1486834041
transform 1 0 16352 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_259
timestamp 1486834041
transform 1 0 24192 0 -1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_260
timestamp 1486834041
transform 1 0 4592 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_261
timestamp 1486834041
transform 1 0 12432 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_262
timestamp 1486834041
transform 1 0 20272 0 1 30576
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_263
timestamp 1486834041
transform 1 0 8512 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_264
timestamp 1486834041
transform 1 0 16352 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_265
timestamp 1486834041
transform 1 0 24192 0 -1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_266
timestamp 1486834041
transform 1 0 4592 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_267
timestamp 1486834041
transform 1 0 12432 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_268
timestamp 1486834041
transform 1 0 20272 0 1 32144
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_269
timestamp 1486834041
transform 1 0 8512 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_270
timestamp 1486834041
transform 1 0 16352 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_271
timestamp 1486834041
transform 1 0 24192 0 -1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_272
timestamp 1486834041
transform 1 0 4592 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_273
timestamp 1486834041
transform 1 0 12432 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_274
timestamp 1486834041
transform 1 0 20272 0 1 33712
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_275
timestamp 1486834041
transform 1 0 8512 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_276
timestamp 1486834041
transform 1 0 16352 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_277
timestamp 1486834041
transform 1 0 24192 0 -1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_278
timestamp 1486834041
transform 1 0 4592 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_279
timestamp 1486834041
transform 1 0 12432 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_280
timestamp 1486834041
transform 1 0 20272 0 1 35280
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_281
timestamp 1486834041
transform 1 0 8512 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_282
timestamp 1486834041
transform 1 0 16352 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_283
timestamp 1486834041
transform 1 0 24192 0 -1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_284
timestamp 1486834041
transform 1 0 4592 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_285
timestamp 1486834041
transform 1 0 12432 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_286
timestamp 1486834041
transform 1 0 20272 0 1 36848
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_287
timestamp 1486834041
transform 1 0 8512 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_288
timestamp 1486834041
transform 1 0 16352 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_289
timestamp 1486834041
transform 1 0 24192 0 -1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_290
timestamp 1486834041
transform 1 0 4592 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_291
timestamp 1486834041
transform 1 0 12432 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_292
timestamp 1486834041
transform 1 0 20272 0 1 38416
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_293
timestamp 1486834041
transform 1 0 8512 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_294
timestamp 1486834041
transform 1 0 16352 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_295
timestamp 1486834041
transform 1 0 24192 0 -1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_296
timestamp 1486834041
transform 1 0 4592 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_297
timestamp 1486834041
transform 1 0 12432 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_298
timestamp 1486834041
transform 1 0 20272 0 1 39984
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_299
timestamp 1486834041
transform 1 0 8512 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_300
timestamp 1486834041
transform 1 0 16352 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_301
timestamp 1486834041
transform 1 0 24192 0 -1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_302
timestamp 1486834041
transform 1 0 4592 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_303
timestamp 1486834041
transform 1 0 12432 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_304
timestamp 1486834041
transform 1 0 20272 0 1 41552
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_305
timestamp 1486834041
transform 1 0 8512 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_306
timestamp 1486834041
transform 1 0 16352 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_307
timestamp 1486834041
transform 1 0 24192 0 -1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_308
timestamp 1486834041
transform 1 0 4592 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_309
timestamp 1486834041
transform 1 0 12432 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_310
timestamp 1486834041
transform 1 0 20272 0 1 43120
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_311
timestamp 1486834041
transform 1 0 8512 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_312
timestamp 1486834041
transform 1 0 16352 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_313
timestamp 1486834041
transform 1 0 24192 0 -1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_314
timestamp 1486834041
transform 1 0 4592 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_315
timestamp 1486834041
transform 1 0 12432 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_316
timestamp 1486834041
transform 1 0 20272 0 1 44688
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_317
timestamp 1486834041
transform 1 0 8512 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_318
timestamp 1486834041
transform 1 0 16352 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_319
timestamp 1486834041
transform 1 0 24192 0 -1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_320
timestamp 1486834041
transform 1 0 4592 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_321
timestamp 1486834041
transform 1 0 12432 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_322
timestamp 1486834041
transform 1 0 20272 0 1 46256
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_323
timestamp 1486834041
transform 1 0 8512 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_324
timestamp 1486834041
transform 1 0 16352 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_325
timestamp 1486834041
transform 1 0 24192 0 -1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_326
timestamp 1486834041
transform 1 0 4592 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_327
timestamp 1486834041
transform 1 0 12432 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_328
timestamp 1486834041
transform 1 0 20272 0 1 47824
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_329
timestamp 1486834041
transform 1 0 8512 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_330
timestamp 1486834041
transform 1 0 16352 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_331
timestamp 1486834041
transform 1 0 24192 0 -1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_332
timestamp 1486834041
transform 1 0 4592 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_333
timestamp 1486834041
transform 1 0 12432 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_334
timestamp 1486834041
transform 1 0 20272 0 1 49392
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_335
timestamp 1486834041
transform 1 0 8512 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_336
timestamp 1486834041
transform 1 0 16352 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_337
timestamp 1486834041
transform 1 0 24192 0 -1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_338
timestamp 1486834041
transform 1 0 4592 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_339
timestamp 1486834041
transform 1 0 12432 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_340
timestamp 1486834041
transform 1 0 20272 0 1 50960
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_341
timestamp 1486834041
transform 1 0 8512 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_342
timestamp 1486834041
transform 1 0 16352 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_343
timestamp 1486834041
transform 1 0 24192 0 -1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_344
timestamp 1486834041
transform 1 0 4592 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_345
timestamp 1486834041
transform 1 0 12432 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_346
timestamp 1486834041
transform 1 0 20272 0 1 52528
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_347
timestamp 1486834041
transform 1 0 8512 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_348
timestamp 1486834041
transform 1 0 16352 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_349
timestamp 1486834041
transform 1 0 24192 0 -1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_350
timestamp 1486834041
transform 1 0 4592 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_351
timestamp 1486834041
transform 1 0 12432 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_352
timestamp 1486834041
transform 1 0 20272 0 1 54096
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_353
timestamp 1486834041
transform 1 0 8512 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_354
timestamp 1486834041
transform 1 0 16352 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_355
timestamp 1486834041
transform 1 0 24192 0 -1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_356
timestamp 1486834041
transform 1 0 4480 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_357
timestamp 1486834041
transform 1 0 8288 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_358
timestamp 1486834041
transform 1 0 12096 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_359
timestamp 1486834041
transform 1 0 15904 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_360
timestamp 1486834041
transform 1 0 19712 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_361
timestamp 1486834041
transform 1 0 23520 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_362
timestamp 1486834041
transform 1 0 27328 0 1 55664
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  wire106
timestamp 1486834041
transform -1 0 13888 0 1 14896
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  wire107
timestamp 1486834041
transform -1 0 15008 0 -1 13328
box -86 -86 758 870
<< labels >>
flabel metal3 s 0 5152 112 5264 0 FreeSans 448 0 0 0 A_I_top
port 0 nsew signal output
flabel metal3 s 0 3808 112 3920 0 FreeSans 448 0 0 0 A_O_top
port 1 nsew signal input
flabel metal3 s 0 6496 112 6608 0 FreeSans 448 0 0 0 A_T_top
port 2 nsew signal output
flabel metal3 s 0 9184 112 9296 0 FreeSans 448 0 0 0 B_I_top
port 3 nsew signal output
flabel metal3 s 0 7840 112 7952 0 FreeSans 448 0 0 0 B_O_top
port 4 nsew signal input
flabel metal3 s 0 10528 112 10640 0 FreeSans 448 0 0 0 B_T_top
port 5 nsew signal output
flabel metal3 s 28448 21728 28560 21840 0 FreeSans 448 0 0 0 E1BEG[0]
port 6 nsew signal output
flabel metal3 s 28448 22176 28560 22288 0 FreeSans 448 0 0 0 E1BEG[1]
port 7 nsew signal output
flabel metal3 s 28448 22624 28560 22736 0 FreeSans 448 0 0 0 E1BEG[2]
port 8 nsew signal output
flabel metal3 s 28448 23072 28560 23184 0 FreeSans 448 0 0 0 E1BEG[3]
port 9 nsew signal output
flabel metal3 s 28448 23520 28560 23632 0 FreeSans 448 0 0 0 E2BEG[0]
port 10 nsew signal output
flabel metal3 s 28448 23968 28560 24080 0 FreeSans 448 0 0 0 E2BEG[1]
port 11 nsew signal output
flabel metal3 s 28448 24416 28560 24528 0 FreeSans 448 0 0 0 E2BEG[2]
port 12 nsew signal output
flabel metal3 s 28448 24864 28560 24976 0 FreeSans 448 0 0 0 E2BEG[3]
port 13 nsew signal output
flabel metal3 s 28448 25312 28560 25424 0 FreeSans 448 0 0 0 E2BEG[4]
port 14 nsew signal output
flabel metal3 s 28448 25760 28560 25872 0 FreeSans 448 0 0 0 E2BEG[5]
port 15 nsew signal output
flabel metal3 s 28448 26208 28560 26320 0 FreeSans 448 0 0 0 E2BEG[6]
port 16 nsew signal output
flabel metal3 s 28448 26656 28560 26768 0 FreeSans 448 0 0 0 E2BEG[7]
port 17 nsew signal output
flabel metal3 s 28448 27104 28560 27216 0 FreeSans 448 0 0 0 E2BEGb[0]
port 18 nsew signal output
flabel metal3 s 28448 27552 28560 27664 0 FreeSans 448 0 0 0 E2BEGb[1]
port 19 nsew signal output
flabel metal3 s 28448 28000 28560 28112 0 FreeSans 448 0 0 0 E2BEGb[2]
port 20 nsew signal output
flabel metal3 s 28448 28448 28560 28560 0 FreeSans 448 0 0 0 E2BEGb[3]
port 21 nsew signal output
flabel metal3 s 28448 28896 28560 29008 0 FreeSans 448 0 0 0 E2BEGb[4]
port 22 nsew signal output
flabel metal3 s 28448 29344 28560 29456 0 FreeSans 448 0 0 0 E2BEGb[5]
port 23 nsew signal output
flabel metal3 s 28448 29792 28560 29904 0 FreeSans 448 0 0 0 E2BEGb[6]
port 24 nsew signal output
flabel metal3 s 28448 30240 28560 30352 0 FreeSans 448 0 0 0 E2BEGb[7]
port 25 nsew signal output
flabel metal3 s 28448 37856 28560 37968 0 FreeSans 448 0 0 0 E6BEG[0]
port 26 nsew signal output
flabel metal3 s 28448 42336 28560 42448 0 FreeSans 448 0 0 0 E6BEG[10]
port 27 nsew signal output
flabel metal3 s 28448 42784 28560 42896 0 FreeSans 448 0 0 0 E6BEG[11]
port 28 nsew signal output
flabel metal3 s 28448 38304 28560 38416 0 FreeSans 448 0 0 0 E6BEG[1]
port 29 nsew signal output
flabel metal3 s 28448 38752 28560 38864 0 FreeSans 448 0 0 0 E6BEG[2]
port 30 nsew signal output
flabel metal3 s 28448 39200 28560 39312 0 FreeSans 448 0 0 0 E6BEG[3]
port 31 nsew signal output
flabel metal3 s 28448 39648 28560 39760 0 FreeSans 448 0 0 0 E6BEG[4]
port 32 nsew signal output
flabel metal3 s 28448 40096 28560 40208 0 FreeSans 448 0 0 0 E6BEG[5]
port 33 nsew signal output
flabel metal3 s 28448 40544 28560 40656 0 FreeSans 448 0 0 0 E6BEG[6]
port 34 nsew signal output
flabel metal3 s 28448 40992 28560 41104 0 FreeSans 448 0 0 0 E6BEG[7]
port 35 nsew signal output
flabel metal3 s 28448 41440 28560 41552 0 FreeSans 448 0 0 0 E6BEG[8]
port 36 nsew signal output
flabel metal3 s 28448 41888 28560 42000 0 FreeSans 448 0 0 0 E6BEG[9]
port 37 nsew signal output
flabel metal3 s 28448 30688 28560 30800 0 FreeSans 448 0 0 0 EE4BEG[0]
port 38 nsew signal output
flabel metal3 s 28448 35168 28560 35280 0 FreeSans 448 0 0 0 EE4BEG[10]
port 39 nsew signal output
flabel metal3 s 28448 35616 28560 35728 0 FreeSans 448 0 0 0 EE4BEG[11]
port 40 nsew signal output
flabel metal3 s 28448 36064 28560 36176 0 FreeSans 448 0 0 0 EE4BEG[12]
port 41 nsew signal output
flabel metal3 s 28448 36512 28560 36624 0 FreeSans 448 0 0 0 EE4BEG[13]
port 42 nsew signal output
flabel metal3 s 28448 36960 28560 37072 0 FreeSans 448 0 0 0 EE4BEG[14]
port 43 nsew signal output
flabel metal3 s 28448 37408 28560 37520 0 FreeSans 448 0 0 0 EE4BEG[15]
port 44 nsew signal output
flabel metal3 s 28448 31136 28560 31248 0 FreeSans 448 0 0 0 EE4BEG[1]
port 45 nsew signal output
flabel metal3 s 28448 31584 28560 31696 0 FreeSans 448 0 0 0 EE4BEG[2]
port 46 nsew signal output
flabel metal3 s 28448 32032 28560 32144 0 FreeSans 448 0 0 0 EE4BEG[3]
port 47 nsew signal output
flabel metal3 s 28448 32480 28560 32592 0 FreeSans 448 0 0 0 EE4BEG[4]
port 48 nsew signal output
flabel metal3 s 28448 32928 28560 33040 0 FreeSans 448 0 0 0 EE4BEG[5]
port 49 nsew signal output
flabel metal3 s 28448 33376 28560 33488 0 FreeSans 448 0 0 0 EE4BEG[6]
port 50 nsew signal output
flabel metal3 s 28448 33824 28560 33936 0 FreeSans 448 0 0 0 EE4BEG[7]
port 51 nsew signal output
flabel metal3 s 28448 34272 28560 34384 0 FreeSans 448 0 0 0 EE4BEG[8]
port 52 nsew signal output
flabel metal3 s 28448 34720 28560 34832 0 FreeSans 448 0 0 0 EE4BEG[9]
port 53 nsew signal output
flabel metal3 s 0 11872 112 11984 0 FreeSans 448 0 0 0 FrameData[0]
port 54 nsew signal input
flabel metal3 s 0 25312 112 25424 0 FreeSans 448 0 0 0 FrameData[10]
port 55 nsew signal input
flabel metal3 s 0 26656 112 26768 0 FreeSans 448 0 0 0 FrameData[11]
port 56 nsew signal input
flabel metal3 s 0 28000 112 28112 0 FreeSans 448 0 0 0 FrameData[12]
port 57 nsew signal input
flabel metal3 s 0 29344 112 29456 0 FreeSans 448 0 0 0 FrameData[13]
port 58 nsew signal input
flabel metal3 s 0 30688 112 30800 0 FreeSans 448 0 0 0 FrameData[14]
port 59 nsew signal input
flabel metal3 s 0 32032 112 32144 0 FreeSans 448 0 0 0 FrameData[15]
port 60 nsew signal input
flabel metal3 s 0 33376 112 33488 0 FreeSans 448 0 0 0 FrameData[16]
port 61 nsew signal input
flabel metal3 s 0 34720 112 34832 0 FreeSans 448 0 0 0 FrameData[17]
port 62 nsew signal input
flabel metal3 s 0 36064 112 36176 0 FreeSans 448 0 0 0 FrameData[18]
port 63 nsew signal input
flabel metal3 s 0 37408 112 37520 0 FreeSans 448 0 0 0 FrameData[19]
port 64 nsew signal input
flabel metal3 s 0 13216 112 13328 0 FreeSans 448 0 0 0 FrameData[1]
port 65 nsew signal input
flabel metal3 s 0 38752 112 38864 0 FreeSans 448 0 0 0 FrameData[20]
port 66 nsew signal input
flabel metal3 s 0 40096 112 40208 0 FreeSans 448 0 0 0 FrameData[21]
port 67 nsew signal input
flabel metal3 s 0 41440 112 41552 0 FreeSans 448 0 0 0 FrameData[22]
port 68 nsew signal input
flabel metal3 s 0 42784 112 42896 0 FreeSans 448 0 0 0 FrameData[23]
port 69 nsew signal input
flabel metal3 s 0 44128 112 44240 0 FreeSans 448 0 0 0 FrameData[24]
port 70 nsew signal input
flabel metal3 s 0 45472 112 45584 0 FreeSans 448 0 0 0 FrameData[25]
port 71 nsew signal input
flabel metal3 s 0 46816 112 46928 0 FreeSans 448 0 0 0 FrameData[26]
port 72 nsew signal input
flabel metal3 s 0 48160 112 48272 0 FreeSans 448 0 0 0 FrameData[27]
port 73 nsew signal input
flabel metal3 s 0 49504 112 49616 0 FreeSans 448 0 0 0 FrameData[28]
port 74 nsew signal input
flabel metal3 s 0 50848 112 50960 0 FreeSans 448 0 0 0 FrameData[29]
port 75 nsew signal input
flabel metal3 s 0 14560 112 14672 0 FreeSans 448 0 0 0 FrameData[2]
port 76 nsew signal input
flabel metal3 s 0 52192 112 52304 0 FreeSans 448 0 0 0 FrameData[30]
port 77 nsew signal input
flabel metal3 s 0 53536 112 53648 0 FreeSans 448 0 0 0 FrameData[31]
port 78 nsew signal input
flabel metal3 s 0 15904 112 16016 0 FreeSans 448 0 0 0 FrameData[3]
port 79 nsew signal input
flabel metal3 s 0 17248 112 17360 0 FreeSans 448 0 0 0 FrameData[4]
port 80 nsew signal input
flabel metal3 s 0 18592 112 18704 0 FreeSans 448 0 0 0 FrameData[5]
port 81 nsew signal input
flabel metal3 s 0 19936 112 20048 0 FreeSans 448 0 0 0 FrameData[6]
port 82 nsew signal input
flabel metal3 s 0 21280 112 21392 0 FreeSans 448 0 0 0 FrameData[7]
port 83 nsew signal input
flabel metal3 s 0 22624 112 22736 0 FreeSans 448 0 0 0 FrameData[8]
port 84 nsew signal input
flabel metal3 s 0 23968 112 24080 0 FreeSans 448 0 0 0 FrameData[9]
port 85 nsew signal input
flabel metal3 s 28448 43232 28560 43344 0 FreeSans 448 0 0 0 FrameData_O[0]
port 86 nsew signal output
flabel metal3 s 28448 47712 28560 47824 0 FreeSans 448 0 0 0 FrameData_O[10]
port 87 nsew signal output
flabel metal3 s 28448 48160 28560 48272 0 FreeSans 448 0 0 0 FrameData_O[11]
port 88 nsew signal output
flabel metal3 s 28448 48608 28560 48720 0 FreeSans 448 0 0 0 FrameData_O[12]
port 89 nsew signal output
flabel metal3 s 28448 49056 28560 49168 0 FreeSans 448 0 0 0 FrameData_O[13]
port 90 nsew signal output
flabel metal3 s 28448 49504 28560 49616 0 FreeSans 448 0 0 0 FrameData_O[14]
port 91 nsew signal output
flabel metal3 s 28448 49952 28560 50064 0 FreeSans 448 0 0 0 FrameData_O[15]
port 92 nsew signal output
flabel metal3 s 28448 50400 28560 50512 0 FreeSans 448 0 0 0 FrameData_O[16]
port 93 nsew signal output
flabel metal3 s 28448 50848 28560 50960 0 FreeSans 448 0 0 0 FrameData_O[17]
port 94 nsew signal output
flabel metal3 s 28448 51296 28560 51408 0 FreeSans 448 0 0 0 FrameData_O[18]
port 95 nsew signal output
flabel metal3 s 28448 51744 28560 51856 0 FreeSans 448 0 0 0 FrameData_O[19]
port 96 nsew signal output
flabel metal3 s 28448 43680 28560 43792 0 FreeSans 448 0 0 0 FrameData_O[1]
port 97 nsew signal output
flabel metal3 s 28448 52192 28560 52304 0 FreeSans 448 0 0 0 FrameData_O[20]
port 98 nsew signal output
flabel metal3 s 28448 52640 28560 52752 0 FreeSans 448 0 0 0 FrameData_O[21]
port 99 nsew signal output
flabel metal3 s 28448 53088 28560 53200 0 FreeSans 448 0 0 0 FrameData_O[22]
port 100 nsew signal output
flabel metal3 s 28448 53536 28560 53648 0 FreeSans 448 0 0 0 FrameData_O[23]
port 101 nsew signal output
flabel metal3 s 28448 53984 28560 54096 0 FreeSans 448 0 0 0 FrameData_O[24]
port 102 nsew signal output
flabel metal3 s 28448 54432 28560 54544 0 FreeSans 448 0 0 0 FrameData_O[25]
port 103 nsew signal output
flabel metal3 s 28448 54880 28560 54992 0 FreeSans 448 0 0 0 FrameData_O[26]
port 104 nsew signal output
flabel metal3 s 28448 55328 28560 55440 0 FreeSans 448 0 0 0 FrameData_O[27]
port 105 nsew signal output
flabel metal3 s 28448 55776 28560 55888 0 FreeSans 448 0 0 0 FrameData_O[28]
port 106 nsew signal output
flabel metal3 s 28448 56224 28560 56336 0 FreeSans 448 0 0 0 FrameData_O[29]
port 107 nsew signal output
flabel metal3 s 28448 44128 28560 44240 0 FreeSans 448 0 0 0 FrameData_O[2]
port 108 nsew signal output
flabel metal3 s 28448 56672 28560 56784 0 FreeSans 448 0 0 0 FrameData_O[30]
port 109 nsew signal output
flabel metal3 s 28448 57120 28560 57232 0 FreeSans 448 0 0 0 FrameData_O[31]
port 110 nsew signal output
flabel metal3 s 28448 44576 28560 44688 0 FreeSans 448 0 0 0 FrameData_O[3]
port 111 nsew signal output
flabel metal3 s 28448 45024 28560 45136 0 FreeSans 448 0 0 0 FrameData_O[4]
port 112 nsew signal output
flabel metal3 s 28448 45472 28560 45584 0 FreeSans 448 0 0 0 FrameData_O[5]
port 113 nsew signal output
flabel metal3 s 28448 45920 28560 46032 0 FreeSans 448 0 0 0 FrameData_O[6]
port 114 nsew signal output
flabel metal3 s 28448 46368 28560 46480 0 FreeSans 448 0 0 0 FrameData_O[7]
port 115 nsew signal output
flabel metal3 s 28448 46816 28560 46928 0 FreeSans 448 0 0 0 FrameData_O[8]
port 116 nsew signal output
flabel metal3 s 28448 47264 28560 47376 0 FreeSans 448 0 0 0 FrameData_O[9]
port 117 nsew signal output
flabel metal2 s 2016 0 2128 112 0 FreeSans 448 0 0 0 FrameStrobe[0]
port 118 nsew signal input
flabel metal2 s 15456 0 15568 112 0 FreeSans 448 0 0 0 FrameStrobe[10]
port 119 nsew signal input
flabel metal2 s 16800 0 16912 112 0 FreeSans 448 0 0 0 FrameStrobe[11]
port 120 nsew signal input
flabel metal2 s 18144 0 18256 112 0 FreeSans 448 0 0 0 FrameStrobe[12]
port 121 nsew signal input
flabel metal2 s 19488 0 19600 112 0 FreeSans 448 0 0 0 FrameStrobe[13]
port 122 nsew signal input
flabel metal2 s 20832 0 20944 112 0 FreeSans 448 0 0 0 FrameStrobe[14]
port 123 nsew signal input
flabel metal2 s 22176 0 22288 112 0 FreeSans 448 0 0 0 FrameStrobe[15]
port 124 nsew signal input
flabel metal2 s 23520 0 23632 112 0 FreeSans 448 0 0 0 FrameStrobe[16]
port 125 nsew signal input
flabel metal2 s 24864 0 24976 112 0 FreeSans 448 0 0 0 FrameStrobe[17]
port 126 nsew signal input
flabel metal2 s 26208 0 26320 112 0 FreeSans 448 0 0 0 FrameStrobe[18]
port 127 nsew signal input
flabel metal2 s 27552 0 27664 112 0 FreeSans 448 0 0 0 FrameStrobe[19]
port 128 nsew signal input
flabel metal2 s 3360 0 3472 112 0 FreeSans 448 0 0 0 FrameStrobe[1]
port 129 nsew signal input
flabel metal2 s 4704 0 4816 112 0 FreeSans 448 0 0 0 FrameStrobe[2]
port 130 nsew signal input
flabel metal2 s 6048 0 6160 112 0 FreeSans 448 0 0 0 FrameStrobe[3]
port 131 nsew signal input
flabel metal2 s 7392 0 7504 112 0 FreeSans 448 0 0 0 FrameStrobe[4]
port 132 nsew signal input
flabel metal2 s 8736 0 8848 112 0 FreeSans 448 0 0 0 FrameStrobe[5]
port 133 nsew signal input
flabel metal2 s 10080 0 10192 112 0 FreeSans 448 0 0 0 FrameStrobe[6]
port 134 nsew signal input
flabel metal2 s 11424 0 11536 112 0 FreeSans 448 0 0 0 FrameStrobe[7]
port 135 nsew signal input
flabel metal2 s 12768 0 12880 112 0 FreeSans 448 0 0 0 FrameStrobe[8]
port 136 nsew signal input
flabel metal2 s 14112 0 14224 112 0 FreeSans 448 0 0 0 FrameStrobe[9]
port 137 nsew signal input
flabel metal2 s 2016 57344 2128 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[0]
port 138 nsew signal output
flabel metal2 s 15456 57344 15568 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[10]
port 139 nsew signal output
flabel metal2 s 16800 57344 16912 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[11]
port 140 nsew signal output
flabel metal2 s 18144 57344 18256 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[12]
port 141 nsew signal output
flabel metal2 s 19488 57344 19600 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[13]
port 142 nsew signal output
flabel metal2 s 20832 57344 20944 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[14]
port 143 nsew signal output
flabel metal2 s 22176 57344 22288 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[15]
port 144 nsew signal output
flabel metal2 s 23520 57344 23632 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[16]
port 145 nsew signal output
flabel metal2 s 24864 57344 24976 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[17]
port 146 nsew signal output
flabel metal2 s 26208 57344 26320 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[18]
port 147 nsew signal output
flabel metal2 s 27552 57344 27664 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[19]
port 148 nsew signal output
flabel metal2 s 3360 57344 3472 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[1]
port 149 nsew signal output
flabel metal2 s 4704 57344 4816 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[2]
port 150 nsew signal output
flabel metal2 s 6048 57344 6160 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[3]
port 151 nsew signal output
flabel metal2 s 7392 57344 7504 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[4]
port 152 nsew signal output
flabel metal2 s 8736 57344 8848 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[5]
port 153 nsew signal output
flabel metal2 s 10080 57344 10192 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[6]
port 154 nsew signal output
flabel metal2 s 11424 57344 11536 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[7]
port 155 nsew signal output
flabel metal2 s 12768 57344 12880 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[8]
port 156 nsew signal output
flabel metal2 s 14112 57344 14224 57456 0 FreeSans 448 0 0 0 FrameStrobe_O[9]
port 157 nsew signal output
flabel metal2 s 672 0 784 112 0 FreeSans 448 0 0 0 UserCLK
port 158 nsew signal input
flabel metal2 s 672 57344 784 57456 0 FreeSans 448 0 0 0 UserCLKo
port 159 nsew signal output
flabel metal4 s 3776 0 4096 57456 0 FreeSans 1472 90 0 0 VDD
port 160 nsew power bidirectional
flabel metal4 s 3776 0 4096 56 0 FreeSans 368 0 0 0 VDD
port 160 nsew power bidirectional
flabel metal4 s 3776 57400 4096 57456 0 FreeSans 368 0 0 0 VDD
port 160 nsew power bidirectional
flabel metal4 s 23776 0 24096 57456 0 FreeSans 1472 90 0 0 VDD
port 160 nsew power bidirectional
flabel metal4 s 23776 0 24096 56 0 FreeSans 368 0 0 0 VDD
port 160 nsew power bidirectional
flabel metal4 s 23776 57400 24096 57456 0 FreeSans 368 0 0 0 VDD
port 160 nsew power bidirectional
flabel metal4 s 4436 0 4756 57456 0 FreeSans 1472 90 0 0 VSS
port 161 nsew ground bidirectional
flabel metal4 s 4436 0 4756 56 0 FreeSans 368 0 0 0 VSS
port 161 nsew ground bidirectional
flabel metal4 s 4436 57400 4756 57456 0 FreeSans 368 0 0 0 VSS
port 161 nsew ground bidirectional
flabel metal4 s 24436 0 24756 57456 0 FreeSans 1472 90 0 0 VSS
port 161 nsew ground bidirectional
flabel metal4 s 24436 0 24756 56 0 FreeSans 368 0 0 0 VSS
port 161 nsew ground bidirectional
flabel metal4 s 24436 57400 24756 57456 0 FreeSans 368 0 0 0 VSS
port 161 nsew ground bidirectional
flabel metal3 s 28448 224 28560 336 0 FreeSans 448 0 0 0 W1END[0]
port 162 nsew signal input
flabel metal3 s 28448 672 28560 784 0 FreeSans 448 0 0 0 W1END[1]
port 163 nsew signal input
flabel metal3 s 28448 1120 28560 1232 0 FreeSans 448 0 0 0 W1END[2]
port 164 nsew signal input
flabel metal3 s 28448 1568 28560 1680 0 FreeSans 448 0 0 0 W1END[3]
port 165 nsew signal input
flabel metal3 s 28448 5600 28560 5712 0 FreeSans 448 0 0 0 W2END[0]
port 166 nsew signal input
flabel metal3 s 28448 6048 28560 6160 0 FreeSans 448 0 0 0 W2END[1]
port 167 nsew signal input
flabel metal3 s 28448 6496 28560 6608 0 FreeSans 448 0 0 0 W2END[2]
port 168 nsew signal input
flabel metal3 s 28448 6944 28560 7056 0 FreeSans 448 0 0 0 W2END[3]
port 169 nsew signal input
flabel metal3 s 28448 7392 28560 7504 0 FreeSans 448 0 0 0 W2END[4]
port 170 nsew signal input
flabel metal3 s 28448 7840 28560 7952 0 FreeSans 448 0 0 0 W2END[5]
port 171 nsew signal input
flabel metal3 s 28448 8288 28560 8400 0 FreeSans 448 0 0 0 W2END[6]
port 172 nsew signal input
flabel metal3 s 28448 8736 28560 8848 0 FreeSans 448 0 0 0 W2END[7]
port 173 nsew signal input
flabel metal3 s 28448 2016 28560 2128 0 FreeSans 448 0 0 0 W2MID[0]
port 174 nsew signal input
flabel metal3 s 28448 2464 28560 2576 0 FreeSans 448 0 0 0 W2MID[1]
port 175 nsew signal input
flabel metal3 s 28448 2912 28560 3024 0 FreeSans 448 0 0 0 W2MID[2]
port 176 nsew signal input
flabel metal3 s 28448 3360 28560 3472 0 FreeSans 448 0 0 0 W2MID[3]
port 177 nsew signal input
flabel metal3 s 28448 3808 28560 3920 0 FreeSans 448 0 0 0 W2MID[4]
port 178 nsew signal input
flabel metal3 s 28448 4256 28560 4368 0 FreeSans 448 0 0 0 W2MID[5]
port 179 nsew signal input
flabel metal3 s 28448 4704 28560 4816 0 FreeSans 448 0 0 0 W2MID[6]
port 180 nsew signal input
flabel metal3 s 28448 5152 28560 5264 0 FreeSans 448 0 0 0 W2MID[7]
port 181 nsew signal input
flabel metal3 s 28448 16352 28560 16464 0 FreeSans 448 0 0 0 W6END[0]
port 182 nsew signal input
flabel metal3 s 28448 20832 28560 20944 0 FreeSans 448 0 0 0 W6END[10]
port 183 nsew signal input
flabel metal3 s 28448 21280 28560 21392 0 FreeSans 448 0 0 0 W6END[11]
port 184 nsew signal input
flabel metal3 s 28448 16800 28560 16912 0 FreeSans 448 0 0 0 W6END[1]
port 185 nsew signal input
flabel metal3 s 28448 17248 28560 17360 0 FreeSans 448 0 0 0 W6END[2]
port 186 nsew signal input
flabel metal3 s 28448 17696 28560 17808 0 FreeSans 448 0 0 0 W6END[3]
port 187 nsew signal input
flabel metal3 s 28448 18144 28560 18256 0 FreeSans 448 0 0 0 W6END[4]
port 188 nsew signal input
flabel metal3 s 28448 18592 28560 18704 0 FreeSans 448 0 0 0 W6END[5]
port 189 nsew signal input
flabel metal3 s 28448 19040 28560 19152 0 FreeSans 448 0 0 0 W6END[6]
port 190 nsew signal input
flabel metal3 s 28448 19488 28560 19600 0 FreeSans 448 0 0 0 W6END[7]
port 191 nsew signal input
flabel metal3 s 28448 19936 28560 20048 0 FreeSans 448 0 0 0 W6END[8]
port 192 nsew signal input
flabel metal3 s 28448 20384 28560 20496 0 FreeSans 448 0 0 0 W6END[9]
port 193 nsew signal input
flabel metal3 s 28448 9184 28560 9296 0 FreeSans 448 0 0 0 WW4END[0]
port 194 nsew signal input
flabel metal3 s 28448 13664 28560 13776 0 FreeSans 448 0 0 0 WW4END[10]
port 195 nsew signal input
flabel metal3 s 28448 14112 28560 14224 0 FreeSans 448 0 0 0 WW4END[11]
port 196 nsew signal input
flabel metal3 s 28448 14560 28560 14672 0 FreeSans 448 0 0 0 WW4END[12]
port 197 nsew signal input
flabel metal3 s 28448 15008 28560 15120 0 FreeSans 448 0 0 0 WW4END[13]
port 198 nsew signal input
flabel metal3 s 28448 15456 28560 15568 0 FreeSans 448 0 0 0 WW4END[14]
port 199 nsew signal input
flabel metal3 s 28448 15904 28560 16016 0 FreeSans 448 0 0 0 WW4END[15]
port 200 nsew signal input
flabel metal3 s 28448 9632 28560 9744 0 FreeSans 448 0 0 0 WW4END[1]
port 201 nsew signal input
flabel metal3 s 28448 10080 28560 10192 0 FreeSans 448 0 0 0 WW4END[2]
port 202 nsew signal input
flabel metal3 s 28448 10528 28560 10640 0 FreeSans 448 0 0 0 WW4END[3]
port 203 nsew signal input
flabel metal3 s 28448 10976 28560 11088 0 FreeSans 448 0 0 0 WW4END[4]
port 204 nsew signal input
flabel metal3 s 28448 11424 28560 11536 0 FreeSans 448 0 0 0 WW4END[5]
port 205 nsew signal input
flabel metal3 s 28448 11872 28560 11984 0 FreeSans 448 0 0 0 WW4END[6]
port 206 nsew signal input
flabel metal3 s 28448 12320 28560 12432 0 FreeSans 448 0 0 0 WW4END[7]
port 207 nsew signal input
flabel metal3 s 28448 12768 28560 12880 0 FreeSans 448 0 0 0 WW4END[8]
port 208 nsew signal input
flabel metal3 s 28448 13216 28560 13328 0 FreeSans 448 0 0 0 WW4END[9]
port 209 nsew signal input
rlabel metal1 14280 56448 14280 56448 0 VDD
rlabel metal1 14280 55664 14280 55664 0 VSS
rlabel metal3 686 5208 686 5208 0 A_I_top
rlabel metal3 1582 3864 1582 3864 0 A_O_top
rlabel metal3 686 6552 686 6552 0 A_T_top
rlabel metal3 686 9240 686 9240 0 B_I_top
rlabel metal3 16576 40376 16576 40376 0 B_O_top
rlabel metal3 686 10584 686 10584 0 B_T_top
rlabel metal2 25704 21952 25704 21952 0 E1BEG[0]
rlabel metal2 27328 21784 27328 21784 0 E1BEG[1]
rlabel metal3 27874 22680 27874 22680 0 E1BEG[2]
rlabel metal2 25704 23408 25704 23408 0 E1BEG[3]
rlabel metal2 27328 23352 27328 23352 0 E2BEG[0]
rlabel metal2 25480 24304 25480 24304 0 E2BEG[1]
rlabel metal3 27874 24472 27874 24472 0 E2BEG[2]
rlabel metal2 25704 25088 25704 25088 0 E2BEG[3]
rlabel metal2 27328 24920 27328 24920 0 E2BEG[4]
rlabel metal3 27874 25816 27874 25816 0 E2BEG[5]
rlabel metal2 25704 26544 25704 26544 0 E2BEG[6]
rlabel metal2 27272 26600 27272 26600 0 E2BEG[7]
rlabel metal2 25704 27552 25704 27552 0 E2BEGb[0]
rlabel metal2 27272 27272 27272 27272 0 E2BEGb[1]
rlabel metal3 27874 28056 27874 28056 0 E2BEGb[2]
rlabel metal3 27874 28504 27874 28504 0 E2BEGb[3]
rlabel metal3 27874 28952 27874 28952 0 E2BEGb[4]
rlabel metal3 27706 29400 27706 29400 0 E2BEGb[5]
rlabel metal3 27874 29848 27874 29848 0 E2BEGb[6]
rlabel metal3 27706 30296 27706 30296 0 E2BEGb[7]
rlabel metal3 27090 37912 27090 37912 0 E6BEG[0]
rlabel metal2 25704 42448 25704 42448 0 E6BEG[10]
rlabel metal3 27874 42840 27874 42840 0 E6BEG[11]
rlabel metal3 27874 38360 27874 38360 0 E6BEG[1]
rlabel metal3 27706 38808 27706 38808 0 E6BEG[2]
rlabel metal2 25704 39312 25704 39312 0 E6BEG[3]
rlabel metal3 27874 39704 27874 39704 0 E6BEG[4]
rlabel metal2 25704 40320 25704 40320 0 E6BEG[5]
rlabel metal3 27706 40600 27706 40600 0 E6BEG[6]
rlabel metal3 27090 41048 27090 41048 0 E6BEG[7]
rlabel metal3 27874 41496 27874 41496 0 E6BEG[8]
rlabel metal3 27706 41944 27706 41944 0 E6BEG[9]
rlabel metal2 25480 30800 25480 30800 0 EE4BEG[0]
rlabel metal3 27874 35224 27874 35224 0 EE4BEG[10]
rlabel metal3 27706 35672 27706 35672 0 EE4BEG[11]
rlabel metal2 25704 36176 25704 36176 0 EE4BEG[12]
rlabel metal3 27874 36568 27874 36568 0 EE4BEG[13]
rlabel metal2 25480 37072 25480 37072 0 EE4BEG[14]
rlabel metal3 27706 37464 27706 37464 0 EE4BEG[15]
rlabel metal3 28266 31192 28266 31192 0 EE4BEG[1]
rlabel metal3 27090 31640 27090 31640 0 EE4BEG[2]
rlabel metal3 27874 32088 27874 32088 0 EE4BEG[3]
rlabel metal3 27706 32536 27706 32536 0 EE4BEG[4]
rlabel metal2 25704 33040 25704 33040 0 EE4BEG[5]
rlabel metal3 27874 33432 27874 33432 0 EE4BEG[6]
rlabel metal2 25704 34048 25704 34048 0 EE4BEG[7]
rlabel metal3 27706 34328 27706 34328 0 EE4BEG[8]
rlabel metal3 27090 34776 27090 34776 0 EE4BEG[9]
rlabel metal2 1960 22344 1960 22344 0 FrameData[0]
rlabel metal2 2800 23016 2800 23016 0 FrameData[10]
rlabel metal2 3528 24024 3528 24024 0 FrameData[11]
rlabel metal3 784 37016 784 37016 0 FrameData[12]
rlabel metal2 3080 39480 3080 39480 0 FrameData[13]
rlabel metal2 3192 35056 3192 35056 0 FrameData[14]
rlabel metal2 2072 34328 2072 34328 0 FrameData[15]
rlabel metal3 1722 33432 1722 33432 0 FrameData[16]
rlabel metal2 15624 32984 15624 32984 0 FrameData[17]
rlabel metal3 1176 26152 1176 26152 0 FrameData[18]
rlabel metal3 1232 27720 1232 27720 0 FrameData[19]
rlabel metal3 126 13272 126 13272 0 FrameData[1]
rlabel metal3 350 38808 350 38808 0 FrameData[20]
rlabel metal2 2072 12600 2072 12600 0 FrameData[21]
rlabel metal2 13160 25424 13160 25424 0 FrameData[22]
rlabel metal2 17752 24416 17752 24416 0 FrameData[23]
rlabel metal3 18088 21448 18088 21448 0 FrameData[24]
rlabel metal2 18648 21728 18648 21728 0 FrameData[25]
rlabel metal3 2576 20776 2576 20776 0 FrameData[26]
rlabel metal2 6104 44800 6104 44800 0 FrameData[27]
rlabel metal3 2926 49560 2926 49560 0 FrameData[28]
rlabel metal3 1022 50904 1022 50904 0 FrameData[29]
rlabel metal3 1736 14784 1736 14784 0 FrameData[2]
rlabel metal3 2352 22568 2352 22568 0 FrameData[30]
rlabel metal3 238 53592 238 53592 0 FrameData[31]
rlabel metal2 5656 19488 5656 19488 0 FrameData[3]
rlabel metal3 1722 17304 1722 17304 0 FrameData[4]
rlabel metal3 4774 18648 4774 18648 0 FrameData[5]
rlabel metal3 8008 19880 8008 19880 0 FrameData[6]
rlabel metal3 1722 21336 1722 21336 0 FrameData[7]
rlabel metal2 17976 23352 17976 23352 0 FrameData[8]
rlabel metal2 18536 23408 18536 23408 0 FrameData[9]
rlabel metal2 25704 43456 25704 43456 0 FrameData_O[0]
rlabel metal3 27874 47768 27874 47768 0 FrameData_O[10]
rlabel metal3 27818 48216 27818 48216 0 FrameData_O[11]
rlabel metal2 25704 48720 25704 48720 0 FrameData_O[12]
rlabel metal3 27874 49112 27874 49112 0 FrameData_O[13]
rlabel metal2 25704 49728 25704 49728 0 FrameData_O[14]
rlabel metal3 27762 50008 27762 50008 0 FrameData_O[15]
rlabel metal3 27034 50456 27034 50456 0 FrameData_O[16]
rlabel metal3 27874 50904 27874 50904 0 FrameData_O[17]
rlabel metal3 27818 51352 27818 51352 0 FrameData_O[18]
rlabel metal3 27034 51800 27034 51800 0 FrameData_O[19]
rlabel metal3 27762 43736 27762 43736 0 FrameData_O[1]
rlabel metal3 27874 52248 27874 52248 0 FrameData_O[20]
rlabel metal3 26978 52696 26978 52696 0 FrameData_O[21]
rlabel metal3 27762 53144 27762 53144 0 FrameData_O[22]
rlabel metal3 27034 53592 27034 53592 0 FrameData_O[23]
rlabel metal3 27874 54040 27874 54040 0 FrameData_O[24]
rlabel metal3 27034 54488 27034 54488 0 FrameData_O[25]
rlabel metal2 24192 54712 24192 54712 0 FrameData_O[26]
rlabel metal2 23800 53872 23800 53872 0 FrameData_O[27]
rlabel metal3 25074 55832 25074 55832 0 FrameData_O[28]
rlabel metal3 27370 56280 27370 56280 0 FrameData_O[29]
rlabel metal3 27090 44184 27090 44184 0 FrameData_O[2]
rlabel metal3 26922 56728 26922 56728 0 FrameData_O[30]
rlabel metal3 24640 53144 24640 53144 0 FrameData_O[31]
rlabel metal3 27874 44632 27874 44632 0 FrameData_O[3]
rlabel metal3 27818 45080 27818 45080 0 FrameData_O[4]
rlabel metal2 25704 45584 25704 45584 0 FrameData_O[5]
rlabel metal3 27874 45976 27874 45976 0 FrameData_O[6]
rlabel metal2 25704 46592 25704 46592 0 FrameData_O[7]
rlabel metal3 27762 46872 27762 46872 0 FrameData_O[8]
rlabel metal3 27090 47320 27090 47320 0 FrameData_O[9]
rlabel metal2 2072 742 2072 742 0 FrameStrobe[0]
rlabel metal2 20888 52080 20888 52080 0 FrameStrobe[10]
rlabel metal3 24192 52920 24192 52920 0 FrameStrobe[11]
rlabel metal3 20384 52696 20384 52696 0 FrameStrobe[12]
rlabel metal2 19544 126 19544 126 0 FrameStrobe[13]
rlabel metal2 20888 1694 20888 1694 0 FrameStrobe[14]
rlabel metal3 18312 47040 18312 47040 0 FrameStrobe[15]
rlabel metal2 23576 686 23576 686 0 FrameStrobe[16]
rlabel metal2 24920 854 24920 854 0 FrameStrobe[17]
rlabel metal2 23744 50568 23744 50568 0 FrameStrobe[18]
rlabel metal2 27608 798 27608 798 0 FrameStrobe[19]
rlabel metal2 3416 1246 3416 1246 0 FrameStrobe[1]
rlabel metal2 4760 126 4760 126 0 FrameStrobe[2]
rlabel metal2 17864 34888 17864 34888 0 FrameStrobe[3]
rlabel metal2 7448 1582 7448 1582 0 FrameStrobe[4]
rlabel metal2 8792 854 8792 854 0 FrameStrobe[5]
rlabel metal2 20104 52836 20104 52836 0 FrameStrobe[6]
rlabel metal3 22456 51128 22456 51128 0 FrameStrobe[7]
rlabel metal2 21896 53592 21896 53592 0 FrameStrobe[8]
rlabel metal2 22792 27384 22792 27384 0 FrameStrobe[9]
rlabel metal2 2520 55300 2520 55300 0 FrameStrobe_O[0]
rlabel metal3 16016 56280 16016 56280 0 FrameStrobe_O[10]
rlabel metal2 17304 55300 17304 55300 0 FrameStrobe_O[11]
rlabel metal2 18368 56280 18368 56280 0 FrameStrobe_O[12]
rlabel metal2 19544 56826 19544 56826 0 FrameStrobe_O[13]
rlabel metal3 21392 56280 21392 56280 0 FrameStrobe_O[14]
rlabel metal2 22232 57274 22232 57274 0 FrameStrobe_O[15]
rlabel metal2 23576 56826 23576 56826 0 FrameStrobe_O[16]
rlabel metal2 24920 56826 24920 56826 0 FrameStrobe_O[17]
rlabel metal2 26264 57330 26264 57330 0 FrameStrobe_O[18]
rlabel metal2 27608 56714 27608 56714 0 FrameStrobe_O[19]
rlabel metal2 3416 56826 3416 56826 0 FrameStrobe_O[1]
rlabel metal2 4760 57330 4760 57330 0 FrameStrobe_O[2]
rlabel metal2 6104 57274 6104 57274 0 FrameStrobe_O[3]
rlabel metal2 7448 56770 7448 56770 0 FrameStrobe_O[4]
rlabel metal2 9016 56448 9016 56448 0 FrameStrobe_O[5]
rlabel metal2 10584 56504 10584 56504 0 FrameStrobe_O[6]
rlabel metal2 11704 55160 11704 55160 0 FrameStrobe_O[7]
rlabel metal2 13048 56448 13048 56448 0 FrameStrobe_O[8]
rlabel metal2 14616 56504 14616 56504 0 FrameStrobe_O[9]
rlabel metal2 2856 25816 2856 25816 0 Inst_A_IO_1_bidirectional_frame_config_pass.Q
rlabel metal2 15512 39564 15512 39564 0 Inst_B_IO_1_bidirectional_frame_config_pass.Q
rlabel metal2 5544 40264 5544 40264 0 Inst_W_IO_ConfigMem.Inst_frame0_bit0.Q
rlabel metal3 7000 39032 7000 39032 0 Inst_W_IO_ConfigMem.Inst_frame0_bit1.Q
rlabel metal2 4032 23352 4032 23352 0 Inst_W_IO_ConfigMem.Inst_frame0_bit10.Q
rlabel metal2 2520 24416 2520 24416 0 Inst_W_IO_ConfigMem.Inst_frame0_bit11.Q
rlabel metal2 7840 37240 7840 37240 0 Inst_W_IO_ConfigMem.Inst_frame0_bit12.Q
rlabel metal3 6664 38808 6664 38808 0 Inst_W_IO_ConfigMem.Inst_frame0_bit13.Q
rlabel metal3 12544 34888 12544 34888 0 Inst_W_IO_ConfigMem.Inst_frame0_bit14.Q
rlabel metal3 13664 35000 13664 35000 0 Inst_W_IO_ConfigMem.Inst_frame0_bit15.Q
rlabel metal3 16464 31192 16464 31192 0 Inst_W_IO_ConfigMem.Inst_frame0_bit16.Q
rlabel metal3 17528 31864 17528 31864 0 Inst_W_IO_ConfigMem.Inst_frame0_bit17.Q
rlabel metal2 13160 22456 13160 22456 0 Inst_W_IO_ConfigMem.Inst_frame0_bit18.Q
rlabel metal2 11928 19712 11928 19712 0 Inst_W_IO_ConfigMem.Inst_frame0_bit19.Q
rlabel metal2 7224 19096 7224 19096 0 Inst_W_IO_ConfigMem.Inst_frame0_bit2.Q
rlabel metal3 12264 24472 12264 24472 0 Inst_W_IO_ConfigMem.Inst_frame0_bit20.Q
rlabel metal2 10584 20216 10584 20216 0 Inst_W_IO_ConfigMem.Inst_frame0_bit21.Q
rlabel metal2 15512 14840 15512 14840 0 Inst_W_IO_ConfigMem.Inst_frame0_bit22.Q
rlabel metal2 15400 15120 15400 15120 0 Inst_W_IO_ConfigMem.Inst_frame0_bit23.Q
rlabel metal3 15680 15288 15680 15288 0 Inst_W_IO_ConfigMem.Inst_frame0_bit24.Q
rlabel metal3 17080 20776 17080 20776 0 Inst_W_IO_ConfigMem.Inst_frame0_bit25.Q
rlabel metal2 16352 19992 16352 19992 0 Inst_W_IO_ConfigMem.Inst_frame0_bit26.Q
rlabel metal2 11256 17976 11256 17976 0 Inst_W_IO_ConfigMem.Inst_frame0_bit27.Q
rlabel metal2 16016 18536 16016 18536 0 Inst_W_IO_ConfigMem.Inst_frame0_bit28.Q
rlabel metal3 10304 15400 10304 15400 0 Inst_W_IO_ConfigMem.Inst_frame0_bit29.Q
rlabel metal2 7896 21280 7896 21280 0 Inst_W_IO_ConfigMem.Inst_frame0_bit3.Q
rlabel metal3 11788 15288 11788 15288 0 Inst_W_IO_ConfigMem.Inst_frame0_bit30.Q
rlabel metal2 10248 14728 10248 14728 0 Inst_W_IO_ConfigMem.Inst_frame0_bit31.Q
rlabel metal3 9688 9240 9688 9240 0 Inst_W_IO_ConfigMem.Inst_frame0_bit4.Q
rlabel metal2 11592 9128 11592 9128 0 Inst_W_IO_ConfigMem.Inst_frame0_bit5.Q
rlabel metal2 12376 31976 12376 31976 0 Inst_W_IO_ConfigMem.Inst_frame0_bit6.Q
rlabel metal2 13608 32424 13608 32424 0 Inst_W_IO_ConfigMem.Inst_frame0_bit7.Q
rlabel metal2 17472 29624 17472 29624 0 Inst_W_IO_ConfigMem.Inst_frame0_bit8.Q
rlabel metal2 18480 30072 18480 30072 0 Inst_W_IO_ConfigMem.Inst_frame0_bit9.Q
rlabel metal2 3304 32088 3304 32088 0 Inst_W_IO_ConfigMem.Inst_frame1_bit0.Q
rlabel metal2 2296 31920 2296 31920 0 Inst_W_IO_ConfigMem.Inst_frame1_bit1.Q
rlabel metal2 6776 29904 6776 29904 0 Inst_W_IO_ConfigMem.Inst_frame1_bit10.Q
rlabel metal2 5096 29008 5096 29008 0 Inst_W_IO_ConfigMem.Inst_frame1_bit11.Q
rlabel metal2 2856 35168 2856 35168 0 Inst_W_IO_ConfigMem.Inst_frame1_bit12.Q
rlabel metal2 1456 34104 1456 34104 0 Inst_W_IO_ConfigMem.Inst_frame1_bit13.Q
rlabel metal3 12656 38024 12656 38024 0 Inst_W_IO_ConfigMem.Inst_frame1_bit14.Q
rlabel metal3 11536 38024 11536 38024 0 Inst_W_IO_ConfigMem.Inst_frame1_bit15.Q
rlabel metal2 7784 33208 7784 33208 0 Inst_W_IO_ConfigMem.Inst_frame1_bit16.Q
rlabel metal3 7000 32536 7000 32536 0 Inst_W_IO_ConfigMem.Inst_frame1_bit17.Q
rlabel metal2 3304 25928 3304 25928 0 Inst_W_IO_ConfigMem.Inst_frame1_bit18.Q
rlabel metal2 2520 26152 2520 26152 0 Inst_W_IO_ConfigMem.Inst_frame1_bit19.Q
rlabel metal2 11144 16184 11144 16184 0 Inst_W_IO_ConfigMem.Inst_frame1_bit2.Q
rlabel metal2 2912 28840 2912 28840 0 Inst_W_IO_ConfigMem.Inst_frame1_bit20.Q
rlabel metal2 2856 29848 2856 29848 0 Inst_W_IO_ConfigMem.Inst_frame1_bit21.Q
rlabel metal2 14336 24696 14336 24696 0 Inst_W_IO_ConfigMem.Inst_frame1_bit22.Q
rlabel metal2 13384 24584 13384 24584 0 Inst_W_IO_ConfigMem.Inst_frame1_bit23.Q
rlabel metal3 16240 21448 16240 21448 0 Inst_W_IO_ConfigMem.Inst_frame1_bit24.Q
rlabel metal2 17640 21280 17640 21280 0 Inst_W_IO_ConfigMem.Inst_frame1_bit25.Q
rlabel metal3 4816 27832 4816 27832 0 Inst_W_IO_ConfigMem.Inst_frame1_bit26.Q
rlabel metal2 6552 27552 6552 27552 0 Inst_W_IO_ConfigMem.Inst_frame1_bit27.Q
rlabel metal3 6552 10584 6552 10584 0 Inst_W_IO_ConfigMem.Inst_frame1_bit28.Q
rlabel metal3 7112 13720 7112 13720 0 Inst_W_IO_ConfigMem.Inst_frame1_bit29.Q
rlabel metal3 11032 16184 11032 16184 0 Inst_W_IO_ConfigMem.Inst_frame1_bit3.Q
rlabel metal2 1624 14392 1624 14392 0 Inst_W_IO_ConfigMem.Inst_frame1_bit30.Q
rlabel metal2 2632 14784 2632 14784 0 Inst_W_IO_ConfigMem.Inst_frame1_bit31.Q
rlabel metal2 11200 9240 11200 9240 0 Inst_W_IO_ConfigMem.Inst_frame1_bit4.Q
rlabel metal2 12152 11312 12152 11312 0 Inst_W_IO_ConfigMem.Inst_frame1_bit5.Q
rlabel metal3 13328 23912 13328 23912 0 Inst_W_IO_ConfigMem.Inst_frame1_bit6.Q
rlabel metal2 13160 24136 13160 24136 0 Inst_W_IO_ConfigMem.Inst_frame1_bit7.Q
rlabel metal2 14728 23072 14728 23072 0 Inst_W_IO_ConfigMem.Inst_frame1_bit8.Q
rlabel metal3 16632 22344 16632 22344 0 Inst_W_IO_ConfigMem.Inst_frame1_bit9.Q
rlabel metal3 8792 27832 8792 27832 0 Inst_W_IO_ConfigMem.Inst_frame2_bit0.Q
rlabel metal2 10472 28504 10472 28504 0 Inst_W_IO_ConfigMem.Inst_frame2_bit1.Q
rlabel metal2 4032 13048 4032 13048 0 Inst_W_IO_ConfigMem.Inst_frame2_bit10.Q
rlabel metal2 5880 13216 5880 13216 0 Inst_W_IO_ConfigMem.Inst_frame2_bit11.Q
rlabel metal3 6944 38920 6944 38920 0 Inst_W_IO_ConfigMem.Inst_frame2_bit12.Q
rlabel metal3 6552 40376 6552 40376 0 Inst_W_IO_ConfigMem.Inst_frame2_bit13.Q
rlabel metal2 5152 23912 5152 23912 0 Inst_W_IO_ConfigMem.Inst_frame2_bit14.Q
rlabel metal2 6048 30184 6048 30184 0 Inst_W_IO_ConfigMem.Inst_frame2_bit15.Q
rlabel metal2 9800 30464 9800 30464 0 Inst_W_IO_ConfigMem.Inst_frame2_bit16.Q
rlabel metal2 11144 31640 11144 31640 0 Inst_W_IO_ConfigMem.Inst_frame2_bit17.Q
rlabel metal2 7896 24976 7896 24976 0 Inst_W_IO_ConfigMem.Inst_frame2_bit18.Q
rlabel metal2 9240 25368 9240 25368 0 Inst_W_IO_ConfigMem.Inst_frame2_bit19.Q
rlabel metal2 8232 20888 8232 20888 0 Inst_W_IO_ConfigMem.Inst_frame2_bit2.Q
rlabel metal3 8960 12152 8960 12152 0 Inst_W_IO_ConfigMem.Inst_frame2_bit20.Q
rlabel metal2 10696 12432 10696 12432 0 Inst_W_IO_ConfigMem.Inst_frame2_bit21.Q
rlabel metal2 15176 27552 15176 27552 0 Inst_W_IO_ConfigMem.Inst_frame2_bit22.Q
rlabel metal2 15288 28504 15288 28504 0 Inst_W_IO_ConfigMem.Inst_frame2_bit23.Q
rlabel metal2 19096 28336 19096 28336 0 Inst_W_IO_ConfigMem.Inst_frame2_bit24.Q
rlabel metal3 19936 28616 19936 28616 0 Inst_W_IO_ConfigMem.Inst_frame2_bit25.Q
rlabel metal3 12432 39704 12432 39704 0 Inst_W_IO_ConfigMem.Inst_frame2_bit26.Q
rlabel metal3 11424 39480 11424 39480 0 Inst_W_IO_ConfigMem.Inst_frame2_bit27.Q
rlabel metal2 6776 34608 6776 34608 0 Inst_W_IO_ConfigMem.Inst_frame2_bit28.Q
rlabel metal3 4872 34888 4872 34888 0 Inst_W_IO_ConfigMem.Inst_frame2_bit29.Q
rlabel metal2 10360 22680 10360 22680 0 Inst_W_IO_ConfigMem.Inst_frame2_bit3.Q
rlabel metal2 3696 20888 3696 20888 0 Inst_W_IO_ConfigMem.Inst_frame2_bit30.Q
rlabel metal3 2128 19432 2128 19432 0 Inst_W_IO_ConfigMem.Inst_frame2_bit31.Q
rlabel metal3 9240 11368 9240 11368 0 Inst_W_IO_ConfigMem.Inst_frame2_bit4.Q
rlabel metal2 11480 12432 11480 12432 0 Inst_W_IO_ConfigMem.Inst_frame2_bit5.Q
rlabel metal2 12992 27272 12992 27272 0 Inst_W_IO_ConfigMem.Inst_frame2_bit6.Q
rlabel metal3 13440 28616 13440 28616 0 Inst_W_IO_ConfigMem.Inst_frame2_bit7.Q
rlabel metal2 18032 25480 18032 25480 0 Inst_W_IO_ConfigMem.Inst_frame2_bit8.Q
rlabel metal2 19432 26152 19432 26152 0 Inst_W_IO_ConfigMem.Inst_frame2_bit9.Q
rlabel metal2 14728 12488 14728 12488 0 Inst_W_IO_ConfigMem.Inst_frame3_bit22.Q
rlabel metal2 19768 20496 19768 20496 0 Inst_W_IO_ConfigMem.Inst_frame3_bit23.Q
rlabel metal2 16856 35168 16856 35168 0 Inst_W_IO_ConfigMem.Inst_frame3_bit24.Q
rlabel metal3 19320 32536 19320 32536 0 Inst_W_IO_ConfigMem.Inst_frame3_bit25.Q
rlabel metal3 4312 17640 4312 17640 0 Inst_W_IO_ConfigMem.Inst_frame3_bit26.Q
rlabel metal2 5992 16016 5992 16016 0 Inst_W_IO_ConfigMem.Inst_frame3_bit27.Q
rlabel metal3 8008 35672 8008 35672 0 Inst_W_IO_ConfigMem.Inst_frame3_bit28.Q
rlabel metal2 9352 35952 9352 35952 0 Inst_W_IO_ConfigMem.Inst_frame3_bit29.Q
rlabel metal2 4312 22064 4312 22064 0 Inst_W_IO_ConfigMem.Inst_frame3_bit30.Q
rlabel metal2 6440 21560 6440 21560 0 Inst_W_IO_ConfigMem.Inst_frame3_bit31.Q
rlabel metal2 14392 10864 14392 10864 0 Inst_W_IO_switch_matrix.E1BEG0
rlabel metal2 19880 21168 19880 21168 0 Inst_W_IO_switch_matrix.E1BEG1
rlabel metal3 14616 36456 14616 36456 0 Inst_W_IO_switch_matrix.E1BEG2
rlabel metal3 18648 32760 18648 32760 0 Inst_W_IO_switch_matrix.E1BEG3
rlabel metal2 5544 13384 5544 13384 0 Inst_W_IO_switch_matrix.E2BEG0
rlabel metal3 9016 35448 9016 35448 0 Inst_W_IO_switch_matrix.E2BEG1
rlabel metal2 5992 22680 5992 22680 0 Inst_W_IO_switch_matrix.E2BEG2
rlabel metal2 10080 27608 10080 27608 0 Inst_W_IO_switch_matrix.E2BEG3
rlabel metal2 9912 23240 9912 23240 0 Inst_W_IO_switch_matrix.E2BEG4
rlabel metal2 10920 12264 10920 12264 0 Inst_W_IO_switch_matrix.E2BEG5
rlabel metal2 13944 29512 13944 29512 0 Inst_W_IO_switch_matrix.E2BEG6
rlabel metal2 18984 25144 18984 25144 0 Inst_W_IO_switch_matrix.E2BEG7
rlabel metal2 5208 11424 5208 11424 0 Inst_W_IO_switch_matrix.E2BEGb0
rlabel metal2 8400 40264 8400 40264 0 Inst_W_IO_switch_matrix.E2BEGb1
rlabel metal2 5656 24304 5656 24304 0 Inst_W_IO_switch_matrix.E2BEGb2
rlabel metal2 10472 30688 10472 30688 0 Inst_W_IO_switch_matrix.E2BEGb3
rlabel metal2 8568 24640 8568 24640 0 Inst_W_IO_switch_matrix.E2BEGb4
rlabel metal2 10080 12040 10080 12040 0 Inst_W_IO_switch_matrix.E2BEGb5
rlabel metal2 15624 27440 15624 27440 0 Inst_W_IO_switch_matrix.E2BEGb6
rlabel metal2 19488 27720 19488 27720 0 Inst_W_IO_switch_matrix.E2BEGb7
rlabel metal2 5992 28168 5992 28168 0 Inst_W_IO_switch_matrix.E6BEG0
rlabel metal2 7784 10192 7784 10192 0 Inst_W_IO_switch_matrix.E6BEG1
rlabel metal2 13496 35112 13496 35112 0 Inst_W_IO_switch_matrix.E6BEG10
rlabel metal2 17752 32648 17752 32648 0 Inst_W_IO_switch_matrix.E6BEG11
rlabel metal2 2856 12432 2856 12432 0 Inst_W_IO_switch_matrix.E6BEG2
rlabel metal2 6104 39984 6104 39984 0 Inst_W_IO_switch_matrix.E6BEG3
rlabel metal3 6664 21336 6664 21336 0 Inst_W_IO_switch_matrix.E6BEG4
rlabel metal2 11032 8680 11032 8680 0 Inst_W_IO_switch_matrix.E6BEG5
rlabel metal2 13048 32256 13048 32256 0 Inst_W_IO_switch_matrix.E6BEG6
rlabel metal2 17808 30856 17808 30856 0 Inst_W_IO_switch_matrix.E6BEG7
rlabel metal3 2464 23128 2464 23128 0 Inst_W_IO_switch_matrix.E6BEG8
rlabel metal2 8568 37576 8568 37576 0 Inst_W_IO_switch_matrix.E6BEG9
rlabel metal2 12488 39984 12488 39984 0 Inst_W_IO_switch_matrix.EE4BEG0
rlabel metal2 6160 35112 6160 35112 0 Inst_W_IO_switch_matrix.EE4BEG1
rlabel metal3 12768 38248 12768 38248 0 Inst_W_IO_switch_matrix.EE4BEG10
rlabel metal2 7336 32872 7336 32872 0 Inst_W_IO_switch_matrix.EE4BEG11
rlabel metal2 3752 25872 3752 25872 0 Inst_W_IO_switch_matrix.EE4BEG12
rlabel metal2 3192 30576 3192 30576 0 Inst_W_IO_switch_matrix.EE4BEG13
rlabel metal3 14336 24584 14336 24584 0 Inst_W_IO_switch_matrix.EE4BEG14
rlabel metal2 14728 20664 14728 20664 0 Inst_W_IO_switch_matrix.EE4BEG15
rlabel metal3 2744 21000 2744 21000 0 Inst_W_IO_switch_matrix.EE4BEG2
rlabel metal2 3752 32088 3752 32088 0 Inst_W_IO_switch_matrix.EE4BEG3
rlabel metal2 11816 16576 11816 16576 0 Inst_W_IO_switch_matrix.EE4BEG4
rlabel metal2 13608 11256 13608 11256 0 Inst_W_IO_switch_matrix.EE4BEG5
rlabel metal2 13944 24136 13944 24136 0 Inst_W_IO_switch_matrix.EE4BEG6
rlabel metal3 15792 22568 15792 22568 0 Inst_W_IO_switch_matrix.EE4BEG7
rlabel metal2 6160 30408 6160 30408 0 Inst_W_IO_switch_matrix.EE4BEG8
rlabel metal2 2184 34440 2184 34440 0 Inst_W_IO_switch_matrix.EE4BEG9
rlabel metal2 728 854 728 854 0 UserCLK
rlabel metal2 18648 37968 18648 37968 0 UserCLK_regs
rlabel metal2 896 55944 896 55944 0 UserCLKo
rlabel metal3 25690 280 25690 280 0 W1END[0]
rlabel metal3 26698 728 26698 728 0 W1END[1]
rlabel metal3 24626 1176 24626 1176 0 W1END[2]
rlabel metal3 28378 1624 28378 1624 0 W1END[3]
rlabel metal3 19712 16856 19712 16856 0 W2END[0]
rlabel metal2 16968 17248 16968 17248 0 W2END[1]
rlabel metal2 16632 9352 16632 9352 0 W2END[2]
rlabel metal2 15736 18032 15736 18032 0 W2END[3]
rlabel metal2 15176 15456 15176 15456 0 W2END[4]
rlabel metal3 27678 7896 27678 7896 0 W2END[5]
rlabel metal3 28434 8344 28434 8344 0 W2END[6]
rlabel metal2 14728 18424 14728 18424 0 W2END[7]
rlabel metal3 24850 2072 24850 2072 0 W2MID[0]
rlabel metal3 21042 2520 21042 2520 0 W2MID[1]
rlabel metal3 20762 2968 20762 2968 0 W2MID[2]
rlabel metal2 16744 21392 16744 21392 0 W2MID[3]
rlabel metal3 17472 20552 17472 20552 0 W2MID[4]
rlabel metal2 16856 21112 16856 21112 0 W2MID[5]
rlabel metal3 27678 4760 27678 4760 0 W2MID[6]
rlabel via3 15176 18639 15176 18639 0 W2MID[7]
rlabel metal2 18424 25424 18424 25424 0 W6END[0]
rlabel metal3 7896 15400 7896 15400 0 W6END[10]
rlabel metal2 2408 30856 2408 30856 0 W6END[11]
rlabel metal2 5096 24808 5096 24808 0 W6END[1]
rlabel metal3 11312 24360 11312 24360 0 W6END[2]
rlabel metal2 2128 25368 2128 25368 0 W6END[3]
rlabel metal3 28434 18200 28434 18200 0 W6END[4]
rlabel metal2 3304 33824 3304 33824 0 W6END[5]
rlabel metal2 23128 24528 23128 24528 0 W6END[6]
rlabel metal3 952 13832 952 13832 0 W6END[7]
rlabel metal3 15960 23464 15960 23464 0 W6END[8]
rlabel metal2 1848 31416 1848 31416 0 W6END[9]
rlabel metal3 20552 25480 20552 25480 0 WW4END[0]
rlabel metal2 9856 11480 9856 11480 0 WW4END[10]
rlabel metal3 28266 14168 28266 14168 0 WW4END[11]
rlabel metal3 28154 14616 28154 14616 0 WW4END[12]
rlabel metal2 2296 24248 2296 24248 0 WW4END[13]
rlabel metal2 21560 28504 21560 28504 0 WW4END[14]
rlabel metal3 8568 15736 8568 15736 0 WW4END[15]
rlabel metal3 16016 19432 16016 19432 0 WW4END[1]
rlabel metal4 24920 10752 24920 10752 0 WW4END[2]
rlabel metal2 25032 16408 25032 16408 0 WW4END[3]
rlabel metal3 27678 11032 27678 11032 0 WW4END[4]
rlabel metal3 28434 11480 28434 11480 0 WW4END[5]
rlabel metal3 28322 11928 28322 11928 0 WW4END[6]
rlabel metal3 27678 12376 27678 12376 0 WW4END[7]
rlabel metal2 17640 23240 17640 23240 0 WW4END[8]
rlabel metal3 27678 13272 27678 13272 0 WW4END[9]
rlabel metal3 16072 19992 16072 19992 0 _000_
rlabel metal2 15176 18088 15176 18088 0 _001_
rlabel metal2 15400 15792 15400 15792 0 _002_
rlabel metal2 16184 13664 16184 13664 0 _003_
rlabel metal3 10976 21336 10976 21336 0 _004_
rlabel metal2 15960 15148 15960 15148 0 _005_
rlabel metal3 9856 14616 9856 14616 0 _006_
rlabel metal2 15960 17080 15960 17080 0 _007_
rlabel metal2 16240 17528 16240 17528 0 _008_
rlabel metal2 16968 18032 16968 18032 0 _009_
rlabel metal3 16800 18200 16800 18200 0 _010_
rlabel metal2 16744 19432 16744 19432 0 _011_
rlabel metal3 16352 18648 16352 18648 0 _012_
rlabel metal2 13776 16856 13776 16856 0 _013_
rlabel metal2 16072 20384 16072 20384 0 _014_
rlabel metal2 14280 18424 14280 18424 0 _015_
rlabel metal2 15624 17752 15624 17752 0 _016_
rlabel metal3 13552 17080 13552 17080 0 _017_
rlabel metal2 12824 17920 12824 17920 0 _018_
rlabel metal3 10808 19432 10808 19432 0 _019_
rlabel metal3 10192 20776 10192 20776 0 _020_
rlabel metal2 13832 23184 13832 23184 0 _021_
rlabel metal2 11536 20776 11536 20776 0 _022_
rlabel metal2 12936 20328 12936 20328 0 _023_
rlabel metal2 12376 19992 12376 19992 0 _024_
rlabel metal2 11648 23352 11648 23352 0 _025_
rlabel metal2 11816 21784 11816 21784 0 _026_
rlabel metal2 15400 13216 15400 13216 0 _027_
rlabel metal2 16968 14224 16968 14224 0 _028_
rlabel metal3 16632 14504 16632 14504 0 _029_
rlabel metal2 17416 14224 17416 14224 0 _030_
rlabel metal3 15624 15400 15624 15400 0 _031_
rlabel metal2 16296 15400 16296 15400 0 _032_
rlabel metal3 16856 15848 16856 15848 0 _033_
rlabel metal2 10248 16912 10248 16912 0 _034_
rlabel metal2 11256 16072 11256 16072 0 _035_
rlabel metal2 11480 15204 11480 15204 0 _036_
rlabel metal3 10248 14280 10248 14280 0 _037_
rlabel metal2 11144 14952 11144 14952 0 _038_
rlabel metal3 9688 16072 9688 16072 0 _039_
rlabel metal3 10528 15512 10528 15512 0 _040_
rlabel metal2 10584 15456 10584 15456 0 _041_
rlabel metal2 18648 39480 18648 39480 0 clknet_0_UserCLK
rlabel metal2 16408 41944 16408 41944 0 clknet_0_UserCLK_regs
rlabel metal2 15512 36904 15512 36904 0 clknet_1_0__leaf_UserCLK
rlabel metal2 16744 36120 16744 36120 0 clknet_1_0__leaf_UserCLK_regs
rlabel metal2 18424 41104 18424 41104 0 clknet_1_1__leaf_UserCLK_regs
rlabel metal2 2520 5880 2520 5880 0 net1
rlabel metal2 23688 33432 23688 33432 0 net10
rlabel metal3 7448 43624 7448 43624 0 net100
rlabel metal3 19432 53592 19432 53592 0 net101
rlabel metal2 21784 53088 21784 53088 0 net102
rlabel metal2 22680 53144 22680 53144 0 net103
rlabel metal2 20216 55720 20216 55720 0 net104
rlabel metal2 22960 55440 22960 55440 0 net105
rlabel metal3 24360 55272 24360 55272 0 net106
rlabel metal2 21952 52248 21952 52248 0 net107
rlabel metal2 25704 53228 25704 53228 0 net108
rlabel metal2 23576 50680 23576 50680 0 net109
rlabel metal3 20692 23912 20692 23912 0 net11
rlabel metal2 19992 52920 19992 52920 0 net110
rlabel metal3 1848 20888 1848 20888 0 net111
rlabel metal2 5824 55440 5824 55440 0 net112
rlabel metal2 18872 37184 18872 37184 0 net113
rlabel metal2 21112 55272 21112 55272 0 net114
rlabel metal3 14728 54600 14728 54600 0 net115
rlabel metal3 11592 55328 11592 55328 0 net116
rlabel metal2 24360 53256 24360 53256 0 net117
rlabel metal2 22344 53816 22344 53816 0 net118
rlabel metal2 23408 51464 23408 51464 0 net119
rlabel metal2 24528 25592 24528 25592 0 net12
rlabel metal2 1400 54376 1400 54376 0 net120
rlabel metal2 2184 11088 2184 11088 0 net121
rlabel metal2 2296 7588 2296 7588 0 net122
rlabel metal2 9352 24360 9352 24360 0 net13
rlabel metal3 25928 25480 25928 25480 0 net14
rlabel metal2 24696 27216 24696 27216 0 net15
rlabel metal2 19600 24808 19600 24808 0 net16
rlabel metal2 17472 23128 17472 23128 0 net17
rlabel metal2 26264 26992 26264 26992 0 net18
rlabel metal2 26376 27104 26376 27104 0 net19
rlabel metal2 17528 13944 17528 13944 0 net2
rlabel metal2 25816 29568 25816 29568 0 net20
rlabel metal2 9520 25592 9520 25592 0 net21
rlabel metal3 26096 30184 26096 30184 0 net22
rlabel metal2 16184 27776 16184 27776 0 net23
rlabel metal2 20104 28000 20104 28000 0 net24
rlabel metal2 25144 33600 25144 33600 0 net25
rlabel metal2 24696 42672 24696 42672 0 net26
rlabel metal2 2072 17752 2072 17752 0 net27
rlabel metal3 17864 27944 17864 27944 0 net28
rlabel metal2 6888 12096 6888 12096 0 net29
rlabel metal2 13720 15960 13720 15960 0 net3
rlabel metal2 1736 24472 1736 24472 0 net30
rlabel metal2 2352 22344 2352 22344 0 net31
rlabel metal2 1736 19824 1736 19824 0 net32
rlabel metal2 1624 17304 1624 17304 0 net33
rlabel metal2 2072 29736 2072 29736 0 net34
rlabel metal3 1456 32536 1456 32536 0 net35
rlabel metal2 1400 23072 1400 23072 0 net36
rlabel metal2 9688 17192 9688 17192 0 net37
rlabel metal3 4424 16856 4424 16856 0 net38
rlabel metal3 6552 23576 6552 23576 0 net39
rlabel metal2 2296 11536 2296 11536 0 net4
rlabel metal2 2184 23408 2184 23408 0 net40
rlabel metal3 9856 32536 9856 32536 0 net41
rlabel metal3 21672 44296 21672 44296 0 net42
rlabel metal2 26264 39312 26264 39312 0 net43
rlabel metal2 3304 13216 3304 13216 0 net44
rlabel metal3 19908 39704 19908 39704 0 net45
rlabel metal3 21168 41160 21168 41160 0 net46
rlabel metal3 23688 40376 23688 40376 0 net47
rlabel metal3 19264 41832 19264 41832 0 net48
rlabel metal3 21056 40152 21056 40152 0 net49
rlabel metal2 24920 18536 24920 18536 0 net5
rlabel metal2 1176 24080 1176 24080 0 net50
rlabel metal3 17024 43400 17024 43400 0 net51
rlabel metal2 24920 32872 24920 32872 0 net52
rlabel metal2 26376 37352 26376 37352 0 net53
rlabel metal2 26264 37352 26264 37352 0 net54
rlabel metal2 25032 32984 25032 32984 0 net55
rlabel metal2 2744 29400 2744 29400 0 net56
rlabel metal2 15288 26236 15288 26236 0 net57
rlabel metal2 15176 33208 15176 33208 0 net58
rlabel metal2 26376 34832 26376 34832 0 net59
rlabel metal3 22792 21448 22792 21448 0 net6
rlabel metal2 1736 22456 1736 22456 0 net60
rlabel metal2 26376 32872 26376 32872 0 net61
rlabel metal2 12096 16968 12096 16968 0 net62
rlabel metal2 17360 17976 17360 17976 0 net63
rlabel metal2 14616 26432 14616 26432 0 net64
rlabel metal2 16968 24248 16968 24248 0 net65
rlabel metal3 23128 30912 23128 30912 0 net66
rlabel metal2 1736 34552 1736 34552 0 net67
rlabel metal2 2184 40544 2184 40544 0 net68
rlabel metal3 1288 12264 1288 12264 0 net69
rlabel metal2 26376 24248 26376 24248 0 net7
rlabel metal2 26376 49280 26376 49280 0 net70
rlabel metal2 24696 48944 24696 48944 0 net71
rlabel metal2 26376 51240 26376 51240 0 net72
rlabel metal2 24696 49616 24696 49616 0 net73
rlabel metal2 26264 51016 26264 51016 0 net74
rlabel metal2 24920 49392 24920 49392 0 net75
rlabel metal3 21952 52136 21952 52136 0 net76
rlabel metal2 1624 22344 1624 22344 0 net77
rlabel metal2 2240 25256 2240 25256 0 net78
rlabel metal2 2296 42336 2296 42336 0 net79
rlabel metal2 19488 25368 19488 25368 0 net8
rlabel metal2 26208 53704 26208 53704 0 net80
rlabel metal2 24696 52976 24696 52976 0 net81
rlabel metal3 20496 54376 20496 54376 0 net82
rlabel metal3 25872 53704 25872 53704 0 net83
rlabel metal2 26096 55272 26096 55272 0 net84
rlabel metal2 24696 55216 24696 55216 0 net85
rlabel metal2 23128 52864 23128 52864 0 net86
rlabel metal2 22904 52584 22904 52584 0 net87
rlabel metal2 20832 55272 20832 55272 0 net88
rlabel metal2 21560 45864 21560 45864 0 net89
rlabel metal3 20776 12376 20776 12376 0 net9
rlabel metal2 24696 44184 24696 44184 0 net90
rlabel metal2 2520 17696 2520 17696 0 net91
rlabel metal3 27272 31248 27272 31248 0 net92
rlabel metal3 20552 19712 20552 19712 0 net93
rlabel metal3 17248 8120 17248 8120 0 net94
rlabel metal3 22848 45864 22848 45864 0 net95
rlabel metal3 26712 44632 26712 44632 0 net96
rlabel metal2 24920 45584 24920 45584 0 net97
rlabel metal3 21336 48104 21336 48104 0 net98
rlabel metal3 22400 46424 22400 46424 0 net99
<< properties >>
string FIXED_BBOX 0 0 28560 57456
<< end >>
