magic
tech gf180mcuD
magscale 1 10
timestamp 1764970338
<< metal1 >>
rect 672 13354 56784 13388
rect 672 13302 4466 13354
rect 4518 13302 4570 13354
rect 4622 13302 4674 13354
rect 4726 13302 24466 13354
rect 24518 13302 24570 13354
rect 24622 13302 24674 13354
rect 24726 13302 44466 13354
rect 44518 13302 44570 13354
rect 44622 13302 44674 13354
rect 44726 13302 56784 13354
rect 672 13268 56784 13302
rect 2158 13186 2210 13198
rect 2158 13122 2210 13134
rect 3726 13186 3778 13198
rect 3726 13122 3778 13134
rect 5966 13186 6018 13198
rect 5966 13122 6018 13134
rect 7534 13186 7586 13198
rect 7534 13122 7586 13134
rect 9774 13186 9826 13198
rect 9774 13122 9826 13134
rect 11342 13186 11394 13198
rect 11342 13122 11394 13134
rect 21198 13186 21250 13198
rect 21198 13122 21250 13134
rect 22654 13186 22706 13198
rect 22654 13122 22706 13134
rect 48974 13186 49026 13198
rect 48974 13122 49026 13134
rect 51102 13186 51154 13198
rect 51102 13122 51154 13134
rect 54910 13186 54962 13198
rect 54910 13122 54962 13134
rect 25454 13074 25506 13086
rect 8082 13022 8094 13074
rect 8146 13022 8158 13074
rect 10322 13022 10334 13074
rect 10386 13022 10398 13074
rect 13682 13022 13694 13074
rect 13746 13022 13758 13074
rect 14914 13022 14926 13074
rect 14978 13022 14990 13074
rect 17490 13022 17502 13074
rect 17554 13022 17566 13074
rect 18274 13022 18286 13074
rect 18338 13022 18350 13074
rect 52882 13022 52894 13074
rect 52946 13022 52958 13074
rect 25454 13010 25506 13022
rect 2706 12910 2718 12962
rect 2770 12910 2782 12962
rect 4274 12910 4286 12962
rect 4338 12910 4350 12962
rect 6514 12910 6526 12962
rect 6578 12910 6590 12962
rect 11890 12910 11902 12962
rect 11954 12910 11966 12962
rect 12898 12910 12910 12962
rect 12962 12910 12974 12962
rect 15698 12910 15710 12962
rect 15762 12910 15774 12962
rect 16930 12910 16942 12962
rect 16994 12910 17006 12962
rect 21746 12910 21758 12962
rect 21810 12910 21822 12962
rect 22082 12910 22094 12962
rect 22146 12910 22158 12962
rect 25106 12910 25118 12962
rect 25170 12910 25182 12962
rect 44930 12910 44942 12962
rect 44994 12910 45006 12962
rect 46834 12910 46846 12962
rect 46898 12910 46910 12962
rect 48402 12910 48414 12962
rect 48466 12910 48478 12962
rect 50754 12910 50766 12962
rect 50818 12910 50830 12962
rect 52098 12910 52110 12962
rect 52162 12910 52174 12962
rect 54338 12910 54350 12962
rect 54402 12910 54414 12962
rect 19294 12850 19346 12862
rect 19294 12786 19346 12798
rect 20302 12850 20354 12862
rect 20302 12786 20354 12798
rect 24110 12850 24162 12862
rect 24110 12786 24162 12798
rect 47854 12850 47906 12862
rect 47854 12786 47906 12798
rect 49982 12850 50034 12862
rect 49982 12786 50034 12798
rect 45950 12738 46002 12750
rect 45950 12674 46002 12686
rect 672 12570 56784 12604
rect 672 12518 3806 12570
rect 3858 12518 3910 12570
rect 3962 12518 4014 12570
rect 4066 12518 23806 12570
rect 23858 12518 23910 12570
rect 23962 12518 24014 12570
rect 24066 12518 43806 12570
rect 43858 12518 43910 12570
rect 43962 12518 44014 12570
rect 44066 12518 56784 12570
rect 672 12484 56784 12518
rect 2270 12402 2322 12414
rect 2270 12338 2322 12350
rect 6974 12402 7026 12414
rect 6974 12338 7026 12350
rect 8542 12402 8594 12414
rect 8542 12338 8594 12350
rect 10110 12402 10162 12414
rect 10110 12338 10162 12350
rect 11678 12402 11730 12414
rect 11678 12338 11730 12350
rect 14814 12402 14866 12414
rect 14814 12338 14866 12350
rect 16718 12402 16770 12414
rect 16718 12338 16770 12350
rect 22318 12402 22370 12414
rect 22318 12338 22370 12350
rect 23886 12402 23938 12414
rect 23886 12338 23938 12350
rect 47966 12402 48018 12414
rect 47966 12338 48018 12350
rect 49422 12402 49474 12414
rect 49422 12338 49474 12350
rect 52558 12402 52610 12414
rect 52558 12338 52610 12350
rect 54126 12402 54178 12414
rect 54126 12338 54178 12350
rect 55694 12402 55746 12414
rect 55694 12338 55746 12350
rect 5966 12290 6018 12302
rect 3602 12238 3614 12290
rect 3666 12238 3678 12290
rect 5966 12226 6018 12238
rect 13694 12290 13746 12302
rect 27134 12290 27186 12302
rect 18162 12238 18174 12290
rect 18226 12238 18238 12290
rect 19506 12238 19518 12290
rect 19570 12238 19582 12290
rect 13694 12226 13746 12238
rect 27134 12226 27186 12238
rect 27918 12290 27970 12302
rect 29262 12290 29314 12302
rect 28578 12238 28590 12290
rect 28642 12238 28654 12290
rect 27918 12226 27970 12238
rect 29262 12226 29314 12238
rect 37102 12290 37154 12302
rect 37102 12226 37154 12238
rect 37326 12290 37378 12302
rect 37326 12226 37378 12238
rect 44494 12290 44546 12302
rect 44494 12226 44546 12238
rect 45278 12290 45330 12302
rect 45278 12226 45330 12238
rect 13358 12178 13410 12190
rect 20638 12178 20690 12190
rect 27358 12178 27410 12190
rect 5506 12126 5518 12178
rect 5570 12126 5582 12178
rect 7522 12126 7534 12178
rect 7586 12126 7598 12178
rect 10658 12126 10670 12178
rect 10722 12126 10734 12178
rect 12226 12126 12238 12178
rect 12290 12126 12302 12178
rect 15810 12126 15822 12178
rect 15874 12126 15886 12178
rect 17266 12126 17278 12178
rect 17330 12126 17342 12178
rect 18834 12126 18846 12178
rect 18898 12126 18910 12178
rect 21970 12126 21982 12178
rect 22034 12126 22046 12178
rect 13358 12114 13410 12126
rect 20638 12114 20690 12126
rect 27358 12114 27410 12126
rect 29038 12178 29090 12190
rect 29038 12114 29090 12126
rect 36878 12178 36930 12190
rect 36878 12114 36930 12126
rect 37662 12178 37714 12190
rect 37662 12114 37714 12126
rect 44718 12178 44770 12190
rect 46958 12178 47010 12190
rect 46498 12126 46510 12178
rect 46562 12126 46574 12178
rect 52210 12126 52222 12178
rect 52274 12126 52286 12178
rect 44718 12114 44770 12126
rect 46958 12114 47010 12126
rect 12798 12066 12850 12078
rect 21198 12066 21250 12078
rect 36318 12066 36370 12078
rect 2818 12014 2830 12066
rect 2882 12014 2894 12066
rect 4386 12014 4398 12066
rect 4450 12014 4462 12066
rect 9090 12014 9102 12066
rect 9154 12014 9166 12066
rect 15362 12014 15374 12066
rect 15426 12014 15438 12066
rect 23314 12014 23326 12066
rect 23378 12014 23390 12066
rect 12798 12002 12850 12014
rect 21198 12002 21250 12014
rect 36318 12002 36370 12014
rect 38222 12066 38274 12078
rect 38222 12002 38274 12014
rect 46062 12066 46114 12078
rect 50990 12066 51042 12078
rect 48514 12014 48526 12066
rect 48578 12014 48590 12066
rect 48850 12014 48862 12066
rect 48914 12014 48926 12066
rect 53554 12014 53566 12066
rect 53618 12014 53630 12066
rect 55122 12014 55134 12066
rect 55186 12014 55198 12066
rect 46062 12002 46114 12014
rect 50990 12002 51042 12014
rect 5182 11954 5234 11966
rect 5182 11890 5234 11902
rect 5406 11954 5458 11966
rect 5406 11890 5458 11902
rect 50430 11954 50482 11966
rect 50430 11890 50482 11902
rect 672 11786 56784 11820
rect 672 11734 4466 11786
rect 4518 11734 4570 11786
rect 4622 11734 4674 11786
rect 4726 11734 24466 11786
rect 24518 11734 24570 11786
rect 24622 11734 24674 11786
rect 24726 11734 44466 11786
rect 44518 11734 44570 11786
rect 44622 11734 44674 11786
rect 44726 11734 56784 11786
rect 672 11700 56784 11734
rect 4622 11618 4674 11630
rect 4622 11554 4674 11566
rect 6190 11618 6242 11630
rect 6190 11554 6242 11566
rect 7758 11618 7810 11630
rect 7758 11554 7810 11566
rect 10894 11618 10946 11630
rect 10894 11554 10946 11566
rect 13918 11618 13970 11630
rect 13918 11554 13970 11566
rect 15486 11618 15538 11630
rect 15486 11554 15538 11566
rect 17390 11618 17442 11630
rect 17390 11554 17442 11566
rect 20526 11618 20578 11630
rect 20526 11554 20578 11566
rect 30718 11618 30770 11630
rect 30718 11554 30770 11566
rect 30942 11618 30994 11630
rect 50318 11618 50370 11630
rect 47506 11566 47518 11618
rect 47570 11566 47582 11618
rect 30942 11554 30994 11566
rect 50318 11554 50370 11566
rect 51886 11618 51938 11630
rect 51886 11554 51938 11566
rect 53454 11618 53506 11630
rect 53454 11554 53506 11566
rect 2046 11506 2098 11518
rect 31502 11506 31554 11518
rect 13010 11454 13022 11506
rect 13074 11454 13086 11506
rect 16818 11454 16830 11506
rect 16882 11454 16894 11506
rect 2046 11442 2098 11454
rect 31502 11442 31554 11454
rect 34190 11506 34242 11518
rect 34190 11442 34242 11454
rect 34414 11506 34466 11518
rect 49746 11454 49758 11506
rect 49810 11454 49822 11506
rect 34414 11442 34466 11454
rect 1486 11394 1538 11406
rect 24558 11394 24610 11406
rect 3602 11342 3614 11394
rect 3666 11342 3678 11394
rect 5170 11342 5182 11394
rect 5234 11342 5246 11394
rect 6626 11342 6638 11394
rect 6690 11342 6702 11394
rect 8082 11342 8094 11394
rect 8146 11342 8158 11394
rect 11442 11342 11454 11394
rect 11506 11342 11518 11394
rect 13570 11342 13582 11394
rect 13634 11342 13646 11394
rect 14914 11342 14926 11394
rect 14978 11342 14990 11394
rect 18498 11342 18510 11394
rect 18562 11342 18574 11394
rect 19954 11342 19966 11394
rect 20018 11342 20030 11394
rect 22754 11342 22766 11394
rect 22818 11342 22830 11394
rect 1486 11330 1538 11342
rect 24558 11330 24610 11342
rect 34974 11394 35026 11406
rect 34974 11330 35026 11342
rect 47182 11394 47234 11406
rect 48178 11342 48190 11394
rect 48242 11342 48254 11394
rect 51314 11342 51326 11394
rect 51378 11342 51390 11394
rect 52882 11342 52894 11394
rect 52946 11342 52958 11394
rect 54898 11342 54910 11394
rect 54962 11342 54974 11394
rect 47182 11330 47234 11342
rect 1262 11282 1314 11294
rect 1262 11218 1314 11230
rect 2606 11282 2658 11294
rect 21758 11282 21810 11294
rect 12338 11230 12350 11282
rect 12402 11230 12414 11282
rect 19058 11230 19070 11282
rect 19122 11230 19134 11282
rect 2606 11218 2658 11230
rect 21758 11218 21810 11230
rect 23998 11282 24050 11294
rect 23998 11218 24050 11230
rect 25118 11282 25170 11294
rect 25118 11218 25170 11230
rect 42030 11282 42082 11294
rect 42030 11218 42082 11230
rect 46846 11282 46898 11294
rect 46846 11218 46898 11230
rect 49198 11282 49250 11294
rect 49198 11218 49250 11230
rect 54462 11282 54514 11294
rect 54462 11218 54514 11230
rect 55246 11282 55298 11294
rect 55246 11218 55298 11230
rect 672 11002 56784 11036
rect 672 10950 3806 11002
rect 3858 10950 3910 11002
rect 3962 10950 4014 11002
rect 4066 10950 23806 11002
rect 23858 10950 23910 11002
rect 23962 10950 24014 11002
rect 24066 10950 43806 11002
rect 43858 10950 43910 11002
rect 43962 10950 44014 11002
rect 44066 10950 56784 11002
rect 672 10916 56784 10950
rect 3390 10834 3442 10846
rect 3390 10770 3442 10782
rect 7422 10834 7474 10846
rect 7422 10770 7474 10782
rect 8990 10834 9042 10846
rect 8990 10770 9042 10782
rect 10558 10834 10610 10846
rect 10558 10770 10610 10782
rect 13022 10834 13074 10846
rect 13022 10770 13074 10782
rect 14590 10834 14642 10846
rect 14590 10770 14642 10782
rect 16718 10834 16770 10846
rect 16718 10770 16770 10782
rect 21646 10834 21698 10846
rect 21646 10770 21698 10782
rect 49646 10834 49698 10846
rect 49646 10770 49698 10782
rect 51214 10834 51266 10846
rect 51214 10770 51266 10782
rect 52558 10834 52610 10846
rect 52558 10770 52610 10782
rect 54574 10722 54626 10734
rect 2146 10670 2158 10722
rect 2210 10670 2222 10722
rect 6066 10670 6078 10722
rect 6130 10670 6142 10722
rect 18610 10670 18622 10722
rect 18674 10670 18686 10722
rect 19618 10670 19630 10722
rect 19682 10670 19694 10722
rect 37090 10670 37102 10722
rect 37154 10670 37166 10722
rect 54574 10658 54626 10670
rect 56142 10722 56194 10734
rect 56142 10658 56194 10670
rect 42254 10610 42306 10622
rect 4162 10558 4174 10610
rect 4226 10558 4238 10610
rect 8194 10558 8206 10610
rect 8258 10558 8270 10610
rect 16146 10558 16158 10610
rect 16210 10558 16222 10610
rect 17938 10558 17950 10610
rect 18002 10558 18014 10610
rect 21074 10558 21086 10610
rect 21138 10558 21150 10610
rect 48738 10558 48750 10610
rect 48802 10558 48814 10610
rect 50194 10558 50206 10610
rect 50258 10558 50270 10610
rect 52098 10558 52110 10610
rect 52162 10558 52174 10610
rect 42254 10546 42306 10558
rect 41134 10498 41186 10510
rect 2818 10446 2830 10498
rect 2882 10446 2894 10498
rect 6850 10446 6862 10498
rect 6914 10446 6926 10498
rect 9986 10446 9998 10498
rect 10050 10446 10062 10498
rect 11554 10446 11566 10498
rect 11618 10446 11630 10498
rect 14018 10446 14030 10498
rect 14082 10446 14094 10498
rect 15586 10446 15598 10498
rect 15650 10446 15662 10498
rect 41134 10434 41186 10446
rect 41358 10498 41410 10510
rect 41358 10434 41410 10446
rect 41918 10498 41970 10510
rect 41918 10434 41970 10446
rect 42814 10498 42866 10510
rect 42814 10434 42866 10446
rect 48190 10498 48242 10510
rect 53554 10446 53566 10498
rect 53618 10446 53630 10498
rect 55122 10446 55134 10498
rect 55186 10446 55198 10498
rect 48190 10434 48242 10446
rect 1374 10386 1426 10398
rect 1374 10322 1426 10334
rect 20078 10386 20130 10398
rect 20078 10322 20130 10334
rect 20638 10386 20690 10398
rect 20638 10322 20690 10334
rect 37550 10386 37602 10398
rect 37550 10322 37602 10334
rect 37886 10386 37938 10398
rect 37886 10322 37938 10334
rect 47406 10386 47458 10398
rect 47406 10322 47458 10334
rect 47630 10386 47682 10398
rect 47630 10322 47682 10334
rect 672 10218 56784 10252
rect 672 10166 4466 10218
rect 4518 10166 4570 10218
rect 4622 10166 4674 10218
rect 4726 10166 24466 10218
rect 24518 10166 24570 10218
rect 24622 10166 24674 10218
rect 24726 10166 44466 10218
rect 44518 10166 44570 10218
rect 44622 10166 44674 10218
rect 44726 10166 56784 10218
rect 672 10132 56784 10166
rect 17390 10050 17442 10062
rect 17390 9986 17442 9998
rect 17726 10050 17778 10062
rect 17726 9986 17778 9998
rect 26126 10050 26178 10062
rect 26126 9986 26178 9998
rect 26462 10050 26514 10062
rect 26462 9986 26514 9998
rect 35870 10050 35922 10062
rect 35870 9986 35922 9998
rect 36094 10050 36146 10062
rect 36094 9986 36146 9998
rect 41134 10050 41186 10062
rect 41134 9986 41186 9998
rect 41470 10050 41522 10062
rect 41470 9986 41522 9998
rect 5742 9938 5794 9950
rect 1474 9886 1486 9938
rect 1538 9886 1550 9938
rect 5742 9874 5794 9886
rect 9438 9938 9490 9950
rect 9438 9874 9490 9886
rect 20302 9938 20354 9950
rect 20302 9874 20354 9886
rect 25566 9938 25618 9950
rect 49410 9886 49422 9938
rect 49474 9886 49486 9938
rect 50194 9886 50206 9938
rect 50258 9886 50270 9938
rect 50978 9886 50990 9938
rect 51042 9886 51054 9938
rect 51762 9886 51774 9938
rect 51826 9886 51838 9938
rect 25566 9874 25618 9886
rect 6302 9826 6354 9838
rect 1250 9774 1262 9826
rect 1314 9774 1326 9826
rect 3042 9774 3054 9826
rect 3106 9774 3118 9826
rect 5282 9774 5294 9826
rect 5346 9774 5358 9826
rect 6302 9762 6354 9774
rect 9998 9826 10050 9838
rect 9998 9762 10050 9774
rect 10334 9826 10386 9838
rect 20862 9826 20914 9838
rect 10770 9774 10782 9826
rect 10834 9774 10846 9826
rect 10334 9762 10386 9774
rect 20862 9762 20914 9774
rect 23438 9826 23490 9838
rect 23438 9762 23490 9774
rect 36654 9826 36706 9838
rect 36654 9762 36706 9774
rect 42590 9826 42642 9838
rect 42590 9762 42642 9774
rect 44606 9826 44658 9838
rect 44606 9762 44658 9774
rect 48526 9826 48578 9838
rect 52546 9774 52558 9826
rect 52610 9774 52622 9826
rect 54226 9774 54238 9826
rect 54290 9774 54302 9826
rect 48526 9762 48578 9774
rect 2046 9714 2098 9726
rect 2046 9650 2098 9662
rect 4286 9714 4338 9726
rect 4286 9650 4338 9662
rect 6638 9714 6690 9726
rect 6638 9650 6690 9662
rect 11118 9714 11170 9726
rect 21198 9714 21250 9726
rect 16930 9662 16942 9714
rect 16994 9662 17006 9714
rect 11118 9650 11170 9662
rect 21198 9650 21250 9662
rect 23102 9714 23154 9726
rect 23102 9650 23154 9662
rect 23998 9714 24050 9726
rect 42254 9714 42306 9726
rect 41906 9662 41918 9714
rect 41970 9662 41982 9714
rect 23998 9650 24050 9662
rect 42254 9650 42306 9662
rect 43150 9714 43202 9726
rect 43150 9650 43202 9662
rect 44270 9714 44322 9726
rect 44270 9650 44322 9662
rect 45166 9714 45218 9726
rect 45166 9650 45218 9662
rect 48302 9714 48354 9726
rect 53566 9714 53618 9726
rect 48962 9662 48974 9714
rect 49026 9662 49038 9714
rect 48302 9650 48354 9662
rect 53566 9650 53618 9662
rect 55134 9602 55186 9614
rect 55134 9538 55186 9550
rect 672 9434 56784 9468
rect 672 9382 3806 9434
rect 3858 9382 3910 9434
rect 3962 9382 4014 9434
rect 4066 9382 23806 9434
rect 23858 9382 23910 9434
rect 23962 9382 24014 9434
rect 24066 9382 43806 9434
rect 43858 9382 43910 9434
rect 43962 9382 44014 9434
rect 44066 9382 56784 9434
rect 672 9348 56784 9382
rect 2046 9266 2098 9278
rect 2046 9202 2098 9214
rect 51214 9266 51266 9278
rect 51214 9202 51266 9214
rect 53006 9266 53058 9278
rect 53006 9202 53058 9214
rect 10110 9154 10162 9166
rect 3042 9102 3054 9154
rect 3106 9102 3118 9154
rect 6066 9102 6078 9154
rect 6130 9102 6142 9154
rect 10110 9090 10162 9102
rect 52210 8990 52222 9042
rect 52274 8990 52286 9042
rect 10334 8930 10386 8942
rect 2594 8878 2606 8930
rect 2658 8878 2670 8930
rect 10334 8866 10386 8878
rect 22430 8930 22482 8942
rect 22430 8866 22482 8878
rect 47630 8930 47682 8942
rect 47630 8866 47682 8878
rect 49870 8930 49922 8942
rect 50194 8878 50206 8930
rect 50258 8878 50270 8930
rect 53554 8878 53566 8930
rect 53618 8878 53630 8930
rect 54338 8878 54350 8930
rect 54402 8878 54414 8930
rect 55122 8878 55134 8930
rect 55186 8878 55198 8930
rect 55906 8878 55918 8930
rect 55970 8878 55982 8930
rect 49870 8866 49922 8878
rect 3502 8818 3554 8830
rect 3502 8754 3554 8766
rect 3726 8818 3778 8830
rect 3726 8754 3778 8766
rect 6526 8818 6578 8830
rect 6526 8754 6578 8766
rect 6750 8818 6802 8830
rect 6750 8754 6802 8766
rect 10894 8818 10946 8830
rect 10894 8754 10946 8766
rect 11230 8818 11282 8830
rect 11230 8754 11282 8766
rect 22990 8818 23042 8830
rect 22990 8754 23042 8766
rect 23214 8818 23266 8830
rect 23214 8754 23266 8766
rect 46846 8818 46898 8830
rect 46846 8754 46898 8766
rect 47070 8818 47122 8830
rect 47070 8754 47122 8766
rect 49086 8818 49138 8830
rect 49086 8754 49138 8766
rect 49310 8818 49362 8830
rect 49310 8754 49362 8766
rect 672 8650 56784 8684
rect 672 8598 4466 8650
rect 4518 8598 4570 8650
rect 4622 8598 4674 8650
rect 4726 8598 24466 8650
rect 24518 8598 24570 8650
rect 24622 8598 24674 8650
rect 24726 8598 44466 8650
rect 44518 8598 44570 8650
rect 44622 8598 44674 8650
rect 44726 8598 56784 8650
rect 672 8564 56784 8598
rect 8878 8370 8930 8382
rect 1474 8318 1486 8370
rect 1538 8318 1550 8370
rect 8878 8306 8930 8318
rect 34414 8370 34466 8382
rect 34414 8306 34466 8318
rect 34638 8370 34690 8382
rect 34638 8306 34690 8318
rect 35198 8370 35250 8382
rect 35198 8306 35250 8318
rect 39790 8370 39842 8382
rect 39790 8306 39842 8318
rect 40238 8370 40290 8382
rect 40238 8306 40290 8318
rect 48414 8370 48466 8382
rect 48414 8306 48466 8318
rect 48974 8370 49026 8382
rect 48974 8306 49026 8318
rect 49870 8370 49922 8382
rect 50978 8318 50990 8370
rect 51042 8318 51054 8370
rect 53330 8318 53342 8370
rect 53394 8318 53406 8370
rect 49870 8306 49922 8318
rect 5742 8258 5794 8270
rect 2258 8206 2270 8258
rect 2322 8206 2334 8258
rect 5742 8194 5794 8206
rect 9438 8258 9490 8270
rect 9438 8194 9490 8206
rect 20526 8258 20578 8270
rect 20526 8194 20578 8206
rect 21534 8258 21586 8270
rect 21534 8194 21586 8206
rect 22094 8258 22146 8270
rect 22094 8194 22146 8206
rect 50094 8258 50146 8270
rect 52546 8206 52558 8258
rect 52610 8206 52622 8258
rect 54114 8206 54126 8258
rect 54178 8206 54190 8258
rect 50094 8194 50146 8206
rect 5406 8146 5458 8158
rect 5406 8082 5458 8094
rect 6302 8146 6354 8158
rect 6302 8082 6354 8094
rect 9774 8146 9826 8158
rect 9774 8082 9826 8094
rect 19966 8146 20018 8158
rect 19966 8082 20018 8094
rect 20862 8146 20914 8158
rect 20862 8082 20914 8094
rect 22430 8146 22482 8158
rect 48190 8146 48242 8158
rect 40674 8094 40686 8146
rect 40738 8094 40750 8146
rect 22430 8082 22482 8094
rect 48190 8082 48242 8094
rect 50654 8146 50706 8158
rect 50654 8082 50706 8094
rect 51998 8146 52050 8158
rect 51998 8082 52050 8094
rect 55134 8146 55186 8158
rect 55134 8082 55186 8094
rect 672 7866 56784 7900
rect 672 7814 3806 7866
rect 3858 7814 3910 7866
rect 3962 7814 4014 7866
rect 4066 7814 23806 7866
rect 23858 7814 23910 7866
rect 23962 7814 24014 7866
rect 24066 7814 43806 7866
rect 43858 7814 43910 7866
rect 43962 7814 44014 7866
rect 44066 7814 56784 7866
rect 672 7780 56784 7814
rect 53006 7698 53058 7710
rect 53006 7634 53058 7646
rect 56142 7698 56194 7710
rect 56142 7634 56194 7646
rect 9662 7586 9714 7598
rect 9662 7522 9714 7534
rect 18958 7586 19010 7598
rect 18958 7522 19010 7534
rect 19742 7586 19794 7598
rect 19742 7522 19794 7534
rect 50542 7586 50594 7598
rect 50542 7522 50594 7534
rect 54574 7586 54626 7598
rect 54574 7522 54626 7534
rect 9998 7474 10050 7486
rect 9998 7410 10050 7422
rect 19518 7474 19570 7486
rect 19518 7410 19570 7422
rect 50878 7474 50930 7486
rect 52098 7422 52110 7474
rect 52162 7422 52174 7474
rect 53666 7422 53678 7474
rect 53730 7422 53742 7474
rect 50878 7410 50930 7422
rect 10558 7362 10610 7374
rect 10558 7298 10610 7310
rect 31166 7362 31218 7374
rect 31166 7298 31218 7310
rect 51438 7362 51490 7374
rect 55122 7310 55134 7362
rect 55186 7310 55198 7362
rect 51438 7298 51490 7310
rect 30270 7250 30322 7262
rect 30270 7186 30322 7198
rect 30606 7250 30658 7262
rect 30606 7186 30658 7198
rect 672 7082 56784 7116
rect 672 7030 4466 7082
rect 4518 7030 4570 7082
rect 4622 7030 4674 7082
rect 4726 7030 24466 7082
rect 24518 7030 24570 7082
rect 24622 7030 24674 7082
rect 24726 7030 44466 7082
rect 44518 7030 44570 7082
rect 44622 7030 44674 7082
rect 44726 7030 56784 7082
rect 672 6996 56784 7030
rect 4062 6690 4114 6702
rect 4062 6626 4114 6638
rect 14142 6690 14194 6702
rect 14142 6626 14194 6638
rect 20638 6690 20690 6702
rect 20638 6626 20690 6638
rect 21198 6690 21250 6702
rect 21198 6626 21250 6638
rect 23214 6690 23266 6702
rect 23214 6626 23266 6638
rect 23438 6690 23490 6702
rect 23438 6626 23490 6638
rect 37550 6690 37602 6702
rect 37550 6626 37602 6638
rect 38670 6690 38722 6702
rect 38670 6626 38722 6638
rect 41582 6690 41634 6702
rect 52658 6638 52670 6690
rect 52722 6638 52734 6690
rect 54114 6638 54126 6690
rect 54178 6638 54190 6690
rect 41582 6626 41634 6638
rect 4398 6578 4450 6590
rect 3602 6526 3614 6578
rect 3666 6526 3678 6578
rect 4398 6514 4450 6526
rect 21422 6578 21474 6590
rect 21422 6514 21474 6526
rect 23998 6578 24050 6590
rect 23998 6514 24050 6526
rect 37326 6578 37378 6590
rect 38334 6578 38386 6590
rect 37986 6526 37998 6578
rect 38050 6526 38062 6578
rect 37326 6514 37378 6526
rect 38334 6514 38386 6526
rect 39230 6578 39282 6590
rect 39230 6514 39282 6526
rect 41358 6578 41410 6590
rect 53566 6578 53618 6590
rect 42018 6526 42030 6578
rect 42082 6526 42094 6578
rect 41358 6514 41410 6526
rect 53566 6514 53618 6526
rect 55134 6466 55186 6478
rect 55134 6402 55186 6414
rect 672 6298 56784 6332
rect 672 6246 3806 6298
rect 3858 6246 3910 6298
rect 3962 6246 4014 6298
rect 4066 6246 23806 6298
rect 23858 6246 23910 6298
rect 23962 6246 24014 6298
rect 24066 6246 43806 6298
rect 43858 6246 43910 6298
rect 43962 6246 44014 6298
rect 44066 6246 56784 6298
rect 672 6212 56784 6246
rect 53006 6130 53058 6142
rect 53006 6066 53058 6078
rect 56142 6130 56194 6142
rect 56142 6066 56194 6078
rect 20526 6018 20578 6030
rect 54574 6018 54626 6030
rect 13458 5966 13470 6018
rect 13522 5966 13534 6018
rect 14354 5966 14366 6018
rect 14418 5966 14430 6018
rect 15586 5966 15598 6018
rect 15650 5966 15662 6018
rect 19618 5966 19630 6018
rect 19682 5966 19694 6018
rect 31826 5966 31838 6018
rect 31890 5966 31902 6018
rect 20526 5954 20578 5966
rect 54574 5954 54626 5966
rect 13918 5906 13970 5918
rect 13918 5842 13970 5854
rect 14814 5906 14866 5918
rect 14814 5842 14866 5854
rect 20078 5906 20130 5918
rect 52098 5854 52110 5906
rect 52162 5854 52174 5906
rect 53554 5854 53566 5906
rect 53618 5854 53630 5906
rect 55234 5854 55246 5906
rect 55298 5854 55310 5906
rect 20078 5842 20130 5854
rect 30382 5794 30434 5806
rect 30382 5730 30434 5742
rect 30942 5794 30994 5806
rect 30942 5730 30994 5742
rect 32286 5794 32338 5806
rect 32286 5730 32338 5742
rect 15150 5682 15202 5694
rect 15150 5618 15202 5630
rect 30046 5682 30098 5694
rect 30046 5618 30098 5630
rect 32622 5682 32674 5694
rect 32622 5618 32674 5630
rect 672 5514 56784 5548
rect 672 5462 4466 5514
rect 4518 5462 4570 5514
rect 4622 5462 4674 5514
rect 4726 5462 24466 5514
rect 24518 5462 24570 5514
rect 24622 5462 24674 5514
rect 24726 5462 44466 5514
rect 44518 5462 44570 5514
rect 44622 5462 44674 5514
rect 44726 5462 56784 5514
rect 672 5428 56784 5462
rect 2606 5346 2658 5358
rect 2606 5282 2658 5294
rect 2942 5346 2994 5358
rect 2942 5282 2994 5294
rect 15150 5346 15202 5358
rect 15150 5282 15202 5294
rect 28814 5346 28866 5358
rect 28814 5282 28866 5294
rect 52334 5346 52386 5358
rect 52334 5282 52386 5294
rect 2046 5234 2098 5246
rect 2046 5170 2098 5182
rect 3950 5234 4002 5246
rect 3950 5170 4002 5182
rect 6750 5234 6802 5246
rect 6750 5170 6802 5182
rect 12574 5234 12626 5246
rect 12574 5170 12626 5182
rect 13582 5234 13634 5246
rect 13582 5170 13634 5182
rect 27918 5234 27970 5246
rect 27918 5170 27970 5182
rect 28478 5234 28530 5246
rect 28478 5170 28530 5182
rect 47518 5234 47570 5246
rect 47518 5170 47570 5182
rect 51998 5234 52050 5246
rect 51998 5170 52050 5182
rect 52894 5234 52946 5246
rect 54114 5182 54126 5234
rect 54178 5182 54190 5234
rect 52894 5170 52946 5182
rect 4510 5122 4562 5134
rect 4510 5058 4562 5070
rect 4846 5122 4898 5134
rect 4846 5058 4898 5070
rect 7310 5122 7362 5134
rect 7310 5058 7362 5070
rect 7646 5122 7698 5134
rect 7646 5058 7698 5070
rect 13134 5122 13186 5134
rect 13134 5058 13186 5070
rect 14142 5122 14194 5134
rect 14142 5058 14194 5070
rect 14366 5122 14418 5134
rect 14366 5058 14418 5070
rect 14814 5122 14866 5134
rect 14814 5058 14866 5070
rect 46622 5122 46674 5134
rect 46622 5058 46674 5070
rect 46958 5122 47010 5134
rect 46958 5058 47010 5070
rect 51102 5122 51154 5134
rect 51102 5058 51154 5070
rect 51438 5122 51490 5134
rect 51438 5058 51490 5070
rect 53230 5122 53282 5134
rect 54898 5070 54910 5122
rect 54962 5070 54974 5122
rect 53230 5058 53282 5070
rect 53666 4958 53678 5010
rect 53730 4958 53742 5010
rect 672 4730 56784 4764
rect 672 4678 3806 4730
rect 3858 4678 3910 4730
rect 3962 4678 4014 4730
rect 4066 4678 23806 4730
rect 23858 4678 23910 4730
rect 23962 4678 24014 4730
rect 24066 4678 43806 4730
rect 43858 4678 43910 4730
rect 43962 4678 44014 4730
rect 44066 4678 56784 4730
rect 672 4644 56784 4678
rect 54574 4562 54626 4574
rect 54574 4498 54626 4510
rect 56142 4562 56194 4574
rect 56142 4498 56194 4510
rect 4846 4450 4898 4462
rect 4846 4386 4898 4398
rect 13470 4450 13522 4462
rect 13470 4386 13522 4398
rect 36206 4450 36258 4462
rect 39902 4450 39954 4462
rect 36978 4398 36990 4450
rect 37042 4398 37054 4450
rect 36206 4386 36258 4398
rect 39902 4386 39954 4398
rect 41358 4450 41410 4462
rect 41358 4386 41410 4398
rect 49870 4450 49922 4462
rect 49870 4386 49922 4398
rect 51438 4450 51490 4462
rect 51438 4386 51490 4398
rect 51998 4450 52050 4462
rect 53118 4450 53170 4462
rect 52658 4398 52670 4450
rect 52722 4398 52734 4450
rect 51998 4386 52050 4398
rect 53118 4386 53170 4398
rect 5182 4338 5234 4350
rect 5182 4274 5234 4286
rect 36542 4338 36594 4350
rect 36542 4274 36594 4286
rect 41694 4338 41746 4350
rect 41694 4274 41746 4286
rect 52222 4338 52274 4350
rect 52222 4274 52274 4286
rect 5742 4226 5794 4238
rect 5742 4162 5794 4174
rect 42254 4226 42306 4238
rect 53554 4174 53566 4226
rect 53618 4174 53630 4226
rect 55122 4174 55134 4226
rect 55186 4174 55198 4226
rect 42254 4162 42306 4174
rect 39006 4114 39058 4126
rect 39006 4050 39058 4062
rect 39342 4114 39394 4126
rect 39342 4050 39394 4062
rect 48974 4114 49026 4126
rect 48974 4050 49026 4062
rect 49310 4114 49362 4126
rect 49310 4050 49362 4062
rect 672 3946 56784 3980
rect 672 3894 4466 3946
rect 4518 3894 4570 3946
rect 4622 3894 4674 3946
rect 4726 3894 24466 3946
rect 24518 3894 24570 3946
rect 24622 3894 24674 3946
rect 24726 3894 44466 3946
rect 44518 3894 44570 3946
rect 44622 3894 44674 3946
rect 44726 3894 56784 3946
rect 672 3860 56784 3894
rect 9438 3778 9490 3790
rect 9438 3714 9490 3726
rect 9662 3778 9714 3790
rect 9662 3714 9714 3726
rect 18398 3778 18450 3790
rect 18398 3714 18450 3726
rect 18622 3778 18674 3790
rect 18622 3714 18674 3726
rect 33294 3778 33346 3790
rect 33294 3714 33346 3726
rect 35646 3778 35698 3790
rect 35646 3714 35698 3726
rect 36318 3778 36370 3790
rect 36318 3714 36370 3726
rect 36542 3778 36594 3790
rect 36542 3714 36594 3726
rect 43710 3778 43762 3790
rect 43710 3714 43762 3726
rect 43934 3778 43986 3790
rect 43934 3714 43986 3726
rect 51438 3778 51490 3790
rect 51438 3714 51490 3726
rect 51662 3778 51714 3790
rect 51662 3714 51714 3726
rect 8878 3666 8930 3678
rect 8878 3602 8930 3614
rect 15822 3666 15874 3678
rect 15822 3602 15874 3614
rect 32398 3666 32450 3678
rect 32398 3602 32450 3614
rect 32958 3666 33010 3678
rect 32958 3602 33010 3614
rect 35310 3666 35362 3678
rect 35310 3602 35362 3614
rect 37102 3666 37154 3678
rect 37102 3602 37154 3614
rect 50542 3666 50594 3678
rect 52546 3614 52558 3666
rect 52610 3614 52622 3666
rect 54898 3614 54910 3666
rect 54962 3614 54974 3666
rect 50542 3602 50594 3614
rect 10110 3554 10162 3566
rect 10110 3490 10162 3502
rect 10446 3554 10498 3566
rect 49758 3554 49810 3566
rect 15138 3502 15150 3554
rect 15202 3502 15214 3554
rect 10446 3490 10498 3502
rect 49758 3490 49810 3502
rect 49982 3554 50034 3566
rect 54338 3502 54350 3554
rect 54402 3502 54414 3554
rect 49982 3490 50034 3502
rect 11006 3442 11058 3454
rect 11006 3378 11058 3390
rect 15598 3442 15650 3454
rect 15598 3378 15650 3390
rect 19182 3442 19234 3454
rect 19182 3378 19234 3390
rect 34750 3442 34802 3454
rect 52222 3442 52274 3454
rect 44370 3390 44382 3442
rect 44434 3390 44446 3442
rect 34750 3378 34802 3390
rect 52222 3378 52274 3390
rect 53566 3442 53618 3454
rect 53566 3378 53618 3390
rect 672 3162 56784 3196
rect 672 3110 3806 3162
rect 3858 3110 3910 3162
rect 3962 3110 4014 3162
rect 4066 3110 23806 3162
rect 23858 3110 23910 3162
rect 23962 3110 24014 3162
rect 24066 3110 43806 3162
rect 43858 3110 43910 3162
rect 43962 3110 44014 3162
rect 44066 3110 56784 3162
rect 672 3076 56784 3110
rect 54574 2994 54626 3006
rect 54574 2930 54626 2942
rect 56142 2994 56194 3006
rect 56142 2930 56194 2942
rect 21198 2882 21250 2894
rect 21198 2818 21250 2830
rect 22094 2882 22146 2894
rect 29262 2882 29314 2894
rect 28578 2830 28590 2882
rect 28642 2830 28654 2882
rect 22094 2818 22146 2830
rect 29262 2818 29314 2830
rect 32846 2882 32898 2894
rect 32846 2818 32898 2830
rect 37662 2882 37714 2894
rect 37662 2818 37714 2830
rect 21534 2770 21586 2782
rect 21534 2706 21586 2718
rect 24894 2770 24946 2782
rect 24894 2706 24946 2718
rect 25454 2770 25506 2782
rect 25454 2706 25506 2718
rect 25678 2770 25730 2782
rect 25678 2706 25730 2718
rect 29038 2770 29090 2782
rect 29038 2706 29090 2718
rect 31950 2770 32002 2782
rect 37886 2770 37938 2782
rect 32386 2718 32398 2770
rect 32450 2718 32462 2770
rect 52210 2718 52222 2770
rect 52274 2718 52286 2770
rect 53554 2718 53566 2770
rect 53618 2718 53630 2770
rect 31950 2706 32002 2718
rect 37886 2706 37938 2718
rect 3838 2658 3890 2670
rect 3838 2594 3890 2606
rect 38446 2658 38498 2670
rect 52770 2606 52782 2658
rect 52834 2606 52846 2658
rect 55122 2606 55134 2658
rect 55186 2606 55198 2658
rect 38446 2594 38498 2606
rect 4398 2546 4450 2558
rect 4398 2482 4450 2494
rect 4958 2546 5010 2558
rect 4958 2482 5010 2494
rect 672 2378 56784 2412
rect 672 2326 4466 2378
rect 4518 2326 4570 2378
rect 4622 2326 4674 2378
rect 4726 2326 24466 2378
rect 24518 2326 24570 2378
rect 24622 2326 24674 2378
rect 24726 2326 44466 2378
rect 44518 2326 44570 2378
rect 44622 2326 44674 2378
rect 44726 2326 56784 2378
rect 672 2292 56784 2326
rect 6974 2210 7026 2222
rect 6974 2146 7026 2158
rect 7310 2210 7362 2222
rect 7310 2146 7362 2158
rect 14254 2210 14306 2222
rect 14254 2146 14306 2158
rect 14590 2210 14642 2222
rect 14590 2146 14642 2158
rect 17838 2210 17890 2222
rect 17838 2146 17890 2158
rect 18062 2210 18114 2222
rect 18062 2146 18114 2158
rect 21310 2210 21362 2222
rect 21310 2146 21362 2158
rect 21646 2210 21698 2222
rect 21646 2146 21698 2158
rect 28702 2210 28754 2222
rect 28702 2146 28754 2158
rect 28926 2210 28978 2222
rect 28926 2146 28978 2158
rect 2830 2098 2882 2110
rect 2830 2034 2882 2046
rect 20750 2098 20802 2110
rect 20750 2034 20802 2046
rect 25118 2098 25170 2110
rect 25118 2034 25170 2046
rect 29486 2098 29538 2110
rect 52546 2046 52558 2098
rect 52610 2046 52622 2098
rect 54114 2046 54126 2098
rect 54178 2046 54190 2098
rect 54898 2046 54910 2098
rect 54962 2046 54974 2098
rect 29486 2034 29538 2046
rect 2494 1986 2546 1998
rect 2494 1922 2546 1934
rect 3390 1986 3442 1998
rect 3390 1922 3442 1934
rect 3726 1986 3778 1998
rect 3726 1922 3778 1934
rect 24558 1986 24610 1998
rect 24558 1922 24610 1934
rect 30382 1986 30434 1998
rect 30382 1922 30434 1934
rect 30942 1986 30994 1998
rect 30942 1922 30994 1934
rect 51662 1986 51714 1998
rect 51662 1922 51714 1934
rect 24110 1874 24162 1886
rect 2034 1822 2046 1874
rect 2098 1822 2110 1874
rect 6514 1822 6526 1874
rect 6578 1822 6590 1874
rect 13794 1822 13806 1874
rect 13858 1822 13870 1874
rect 17378 1822 17390 1874
rect 17442 1822 17454 1874
rect 24110 1810 24162 1822
rect 31166 1874 31218 1886
rect 31166 1810 31218 1822
rect 51438 1874 51490 1886
rect 53566 1874 53618 1886
rect 52098 1822 52110 1874
rect 52162 1822 52174 1874
rect 51438 1810 51490 1822
rect 53566 1810 53618 1822
rect 672 1594 56784 1628
rect 672 1542 3806 1594
rect 3858 1542 3910 1594
rect 3962 1542 4014 1594
rect 4066 1542 23806 1594
rect 23858 1542 23910 1594
rect 23962 1542 24014 1594
rect 24066 1542 43806 1594
rect 43858 1542 43910 1594
rect 43962 1542 44014 1594
rect 44066 1542 56784 1594
rect 672 1508 56784 1542
rect 53566 1426 53618 1438
rect 53566 1362 53618 1374
rect 56142 1426 56194 1438
rect 56142 1362 56194 1374
rect 2830 1314 2882 1326
rect 2830 1250 2882 1262
rect 51998 1314 52050 1326
rect 51998 1250 52050 1262
rect 50978 1150 50990 1202
rect 51042 1150 51054 1202
rect 52546 1150 52558 1202
rect 52610 1150 52622 1202
rect 55346 1150 55358 1202
rect 55410 1150 55422 1202
rect 672 810 56784 844
rect 672 758 4466 810
rect 4518 758 4570 810
rect 4622 758 4674 810
rect 4726 758 24466 810
rect 24518 758 24570 810
rect 24622 758 24674 810
rect 24726 758 44466 810
rect 44518 758 44570 810
rect 44622 758 44674 810
rect 44726 758 56784 810
rect 672 724 56784 758
<< via1 >>
rect 4466 13302 4518 13354
rect 4570 13302 4622 13354
rect 4674 13302 4726 13354
rect 24466 13302 24518 13354
rect 24570 13302 24622 13354
rect 24674 13302 24726 13354
rect 44466 13302 44518 13354
rect 44570 13302 44622 13354
rect 44674 13302 44726 13354
rect 2158 13134 2210 13186
rect 3726 13134 3778 13186
rect 5966 13134 6018 13186
rect 7534 13134 7586 13186
rect 9774 13134 9826 13186
rect 11342 13134 11394 13186
rect 21198 13134 21250 13186
rect 22654 13134 22706 13186
rect 48974 13134 49026 13186
rect 51102 13134 51154 13186
rect 54910 13134 54962 13186
rect 8094 13022 8146 13074
rect 10334 13022 10386 13074
rect 13694 13022 13746 13074
rect 14926 13022 14978 13074
rect 17502 13022 17554 13074
rect 18286 13022 18338 13074
rect 25454 13022 25506 13074
rect 52894 13022 52946 13074
rect 2718 12910 2770 12962
rect 4286 12910 4338 12962
rect 6526 12910 6578 12962
rect 11902 12910 11954 12962
rect 12910 12910 12962 12962
rect 15710 12910 15762 12962
rect 16942 12910 16994 12962
rect 21758 12910 21810 12962
rect 22094 12910 22146 12962
rect 25118 12910 25170 12962
rect 44942 12910 44994 12962
rect 46846 12910 46898 12962
rect 48414 12910 48466 12962
rect 50766 12910 50818 12962
rect 52110 12910 52162 12962
rect 54350 12910 54402 12962
rect 19294 12798 19346 12850
rect 20302 12798 20354 12850
rect 24110 12798 24162 12850
rect 47854 12798 47906 12850
rect 49982 12798 50034 12850
rect 45950 12686 46002 12738
rect 3806 12518 3858 12570
rect 3910 12518 3962 12570
rect 4014 12518 4066 12570
rect 23806 12518 23858 12570
rect 23910 12518 23962 12570
rect 24014 12518 24066 12570
rect 43806 12518 43858 12570
rect 43910 12518 43962 12570
rect 44014 12518 44066 12570
rect 2270 12350 2322 12402
rect 6974 12350 7026 12402
rect 8542 12350 8594 12402
rect 10110 12350 10162 12402
rect 11678 12350 11730 12402
rect 14814 12350 14866 12402
rect 16718 12350 16770 12402
rect 22318 12350 22370 12402
rect 23886 12350 23938 12402
rect 47966 12350 48018 12402
rect 49422 12350 49474 12402
rect 52558 12350 52610 12402
rect 54126 12350 54178 12402
rect 55694 12350 55746 12402
rect 3614 12238 3666 12290
rect 5966 12238 6018 12290
rect 13694 12238 13746 12290
rect 18174 12238 18226 12290
rect 19518 12238 19570 12290
rect 27134 12238 27186 12290
rect 27918 12238 27970 12290
rect 28590 12238 28642 12290
rect 29262 12238 29314 12290
rect 37102 12238 37154 12290
rect 37326 12238 37378 12290
rect 44494 12238 44546 12290
rect 45278 12238 45330 12290
rect 5518 12126 5570 12178
rect 7534 12126 7586 12178
rect 10670 12126 10722 12178
rect 12238 12126 12290 12178
rect 13358 12126 13410 12178
rect 15822 12126 15874 12178
rect 17278 12126 17330 12178
rect 18846 12126 18898 12178
rect 20638 12126 20690 12178
rect 21982 12126 22034 12178
rect 27358 12126 27410 12178
rect 29038 12126 29090 12178
rect 36878 12126 36930 12178
rect 37662 12126 37714 12178
rect 44718 12126 44770 12178
rect 46510 12126 46562 12178
rect 46958 12126 47010 12178
rect 52222 12126 52274 12178
rect 2830 12014 2882 12066
rect 4398 12014 4450 12066
rect 9102 12014 9154 12066
rect 12798 12014 12850 12066
rect 15374 12014 15426 12066
rect 21198 12014 21250 12066
rect 23326 12014 23378 12066
rect 36318 12014 36370 12066
rect 38222 12014 38274 12066
rect 46062 12014 46114 12066
rect 48526 12014 48578 12066
rect 48862 12014 48914 12066
rect 50990 12014 51042 12066
rect 53566 12014 53618 12066
rect 55134 12014 55186 12066
rect 5182 11902 5234 11954
rect 5406 11902 5458 11954
rect 50430 11902 50482 11954
rect 4466 11734 4518 11786
rect 4570 11734 4622 11786
rect 4674 11734 4726 11786
rect 24466 11734 24518 11786
rect 24570 11734 24622 11786
rect 24674 11734 24726 11786
rect 44466 11734 44518 11786
rect 44570 11734 44622 11786
rect 44674 11734 44726 11786
rect 4622 11566 4674 11618
rect 6190 11566 6242 11618
rect 7758 11566 7810 11618
rect 10894 11566 10946 11618
rect 13918 11566 13970 11618
rect 15486 11566 15538 11618
rect 17390 11566 17442 11618
rect 20526 11566 20578 11618
rect 30718 11566 30770 11618
rect 30942 11566 30994 11618
rect 47518 11566 47570 11618
rect 50318 11566 50370 11618
rect 51886 11566 51938 11618
rect 53454 11566 53506 11618
rect 2046 11454 2098 11506
rect 13022 11454 13074 11506
rect 16830 11454 16882 11506
rect 31502 11454 31554 11506
rect 34190 11454 34242 11506
rect 34414 11454 34466 11506
rect 49758 11454 49810 11506
rect 1486 11342 1538 11394
rect 3614 11342 3666 11394
rect 5182 11342 5234 11394
rect 6638 11342 6690 11394
rect 8094 11342 8146 11394
rect 11454 11342 11506 11394
rect 13582 11342 13634 11394
rect 14926 11342 14978 11394
rect 18510 11342 18562 11394
rect 19966 11342 20018 11394
rect 22766 11342 22818 11394
rect 24558 11342 24610 11394
rect 34974 11342 35026 11394
rect 47182 11342 47234 11394
rect 48190 11342 48242 11394
rect 51326 11342 51378 11394
rect 52894 11342 52946 11394
rect 54910 11342 54962 11394
rect 1262 11230 1314 11282
rect 2606 11230 2658 11282
rect 12350 11230 12402 11282
rect 19070 11230 19122 11282
rect 21758 11230 21810 11282
rect 23998 11230 24050 11282
rect 25118 11230 25170 11282
rect 42030 11230 42082 11282
rect 46846 11230 46898 11282
rect 49198 11230 49250 11282
rect 54462 11230 54514 11282
rect 55246 11230 55298 11282
rect 3806 10950 3858 11002
rect 3910 10950 3962 11002
rect 4014 10950 4066 11002
rect 23806 10950 23858 11002
rect 23910 10950 23962 11002
rect 24014 10950 24066 11002
rect 43806 10950 43858 11002
rect 43910 10950 43962 11002
rect 44014 10950 44066 11002
rect 3390 10782 3442 10834
rect 7422 10782 7474 10834
rect 8990 10782 9042 10834
rect 10558 10782 10610 10834
rect 13022 10782 13074 10834
rect 14590 10782 14642 10834
rect 16718 10782 16770 10834
rect 21646 10782 21698 10834
rect 49646 10782 49698 10834
rect 51214 10782 51266 10834
rect 52558 10782 52610 10834
rect 2158 10670 2210 10722
rect 6078 10670 6130 10722
rect 18622 10670 18674 10722
rect 19630 10670 19682 10722
rect 37102 10670 37154 10722
rect 54574 10670 54626 10722
rect 56142 10670 56194 10722
rect 4174 10558 4226 10610
rect 8206 10558 8258 10610
rect 16158 10558 16210 10610
rect 17950 10558 18002 10610
rect 21086 10558 21138 10610
rect 42254 10558 42306 10610
rect 48750 10558 48802 10610
rect 50206 10558 50258 10610
rect 52110 10558 52162 10610
rect 2830 10446 2882 10498
rect 6862 10446 6914 10498
rect 9998 10446 10050 10498
rect 11566 10446 11618 10498
rect 14030 10446 14082 10498
rect 15598 10446 15650 10498
rect 41134 10446 41186 10498
rect 41358 10446 41410 10498
rect 41918 10446 41970 10498
rect 42814 10446 42866 10498
rect 48190 10446 48242 10498
rect 53566 10446 53618 10498
rect 55134 10446 55186 10498
rect 1374 10334 1426 10386
rect 20078 10334 20130 10386
rect 20638 10334 20690 10386
rect 37550 10334 37602 10386
rect 37886 10334 37938 10386
rect 47406 10334 47458 10386
rect 47630 10334 47682 10386
rect 4466 10166 4518 10218
rect 4570 10166 4622 10218
rect 4674 10166 4726 10218
rect 24466 10166 24518 10218
rect 24570 10166 24622 10218
rect 24674 10166 24726 10218
rect 44466 10166 44518 10218
rect 44570 10166 44622 10218
rect 44674 10166 44726 10218
rect 17390 9998 17442 10050
rect 17726 9998 17778 10050
rect 26126 9998 26178 10050
rect 26462 9998 26514 10050
rect 35870 9998 35922 10050
rect 36094 9998 36146 10050
rect 41134 9998 41186 10050
rect 41470 9998 41522 10050
rect 1486 9886 1538 9938
rect 5742 9886 5794 9938
rect 9438 9886 9490 9938
rect 20302 9886 20354 9938
rect 25566 9886 25618 9938
rect 49422 9886 49474 9938
rect 50206 9886 50258 9938
rect 50990 9886 51042 9938
rect 51774 9886 51826 9938
rect 1262 9774 1314 9826
rect 3054 9774 3106 9826
rect 5294 9774 5346 9826
rect 6302 9774 6354 9826
rect 9998 9774 10050 9826
rect 10334 9774 10386 9826
rect 10782 9774 10834 9826
rect 20862 9774 20914 9826
rect 23438 9774 23490 9826
rect 36654 9774 36706 9826
rect 42590 9774 42642 9826
rect 44606 9774 44658 9826
rect 48526 9774 48578 9826
rect 52558 9774 52610 9826
rect 54238 9774 54290 9826
rect 2046 9662 2098 9714
rect 4286 9662 4338 9714
rect 6638 9662 6690 9714
rect 11118 9662 11170 9714
rect 16942 9662 16994 9714
rect 21198 9662 21250 9714
rect 23102 9662 23154 9714
rect 23998 9662 24050 9714
rect 41918 9662 41970 9714
rect 42254 9662 42306 9714
rect 43150 9662 43202 9714
rect 44270 9662 44322 9714
rect 45166 9662 45218 9714
rect 48302 9662 48354 9714
rect 48974 9662 49026 9714
rect 53566 9662 53618 9714
rect 55134 9550 55186 9602
rect 3806 9382 3858 9434
rect 3910 9382 3962 9434
rect 4014 9382 4066 9434
rect 23806 9382 23858 9434
rect 23910 9382 23962 9434
rect 24014 9382 24066 9434
rect 43806 9382 43858 9434
rect 43910 9382 43962 9434
rect 44014 9382 44066 9434
rect 2046 9214 2098 9266
rect 51214 9214 51266 9266
rect 53006 9214 53058 9266
rect 3054 9102 3106 9154
rect 6078 9102 6130 9154
rect 10110 9102 10162 9154
rect 52222 8990 52274 9042
rect 2606 8878 2658 8930
rect 10334 8878 10386 8930
rect 22430 8878 22482 8930
rect 47630 8878 47682 8930
rect 49870 8878 49922 8930
rect 50206 8878 50258 8930
rect 53566 8878 53618 8930
rect 54350 8878 54402 8930
rect 55134 8878 55186 8930
rect 55918 8878 55970 8930
rect 3502 8766 3554 8818
rect 3726 8766 3778 8818
rect 6526 8766 6578 8818
rect 6750 8766 6802 8818
rect 10894 8766 10946 8818
rect 11230 8766 11282 8818
rect 22990 8766 23042 8818
rect 23214 8766 23266 8818
rect 46846 8766 46898 8818
rect 47070 8766 47122 8818
rect 49086 8766 49138 8818
rect 49310 8766 49362 8818
rect 4466 8598 4518 8650
rect 4570 8598 4622 8650
rect 4674 8598 4726 8650
rect 24466 8598 24518 8650
rect 24570 8598 24622 8650
rect 24674 8598 24726 8650
rect 44466 8598 44518 8650
rect 44570 8598 44622 8650
rect 44674 8598 44726 8650
rect 1486 8318 1538 8370
rect 8878 8318 8930 8370
rect 34414 8318 34466 8370
rect 34638 8318 34690 8370
rect 35198 8318 35250 8370
rect 39790 8318 39842 8370
rect 40238 8318 40290 8370
rect 48414 8318 48466 8370
rect 48974 8318 49026 8370
rect 49870 8318 49922 8370
rect 50990 8318 51042 8370
rect 53342 8318 53394 8370
rect 2270 8206 2322 8258
rect 5742 8206 5794 8258
rect 9438 8206 9490 8258
rect 20526 8206 20578 8258
rect 21534 8206 21586 8258
rect 22094 8206 22146 8258
rect 50094 8206 50146 8258
rect 52558 8206 52610 8258
rect 54126 8206 54178 8258
rect 5406 8094 5458 8146
rect 6302 8094 6354 8146
rect 9774 8094 9826 8146
rect 19966 8094 20018 8146
rect 20862 8094 20914 8146
rect 22430 8094 22482 8146
rect 40686 8094 40738 8146
rect 48190 8094 48242 8146
rect 50654 8094 50706 8146
rect 51998 8094 52050 8146
rect 55134 8094 55186 8146
rect 3806 7814 3858 7866
rect 3910 7814 3962 7866
rect 4014 7814 4066 7866
rect 23806 7814 23858 7866
rect 23910 7814 23962 7866
rect 24014 7814 24066 7866
rect 43806 7814 43858 7866
rect 43910 7814 43962 7866
rect 44014 7814 44066 7866
rect 53006 7646 53058 7698
rect 56142 7646 56194 7698
rect 9662 7534 9714 7586
rect 18958 7534 19010 7586
rect 19742 7534 19794 7586
rect 50542 7534 50594 7586
rect 54574 7534 54626 7586
rect 9998 7422 10050 7474
rect 19518 7422 19570 7474
rect 50878 7422 50930 7474
rect 52110 7422 52162 7474
rect 53678 7422 53730 7474
rect 10558 7310 10610 7362
rect 31166 7310 31218 7362
rect 51438 7310 51490 7362
rect 55134 7310 55186 7362
rect 30270 7198 30322 7250
rect 30606 7198 30658 7250
rect 4466 7030 4518 7082
rect 4570 7030 4622 7082
rect 4674 7030 4726 7082
rect 24466 7030 24518 7082
rect 24570 7030 24622 7082
rect 24674 7030 24726 7082
rect 44466 7030 44518 7082
rect 44570 7030 44622 7082
rect 44674 7030 44726 7082
rect 4062 6638 4114 6690
rect 14142 6638 14194 6690
rect 20638 6638 20690 6690
rect 21198 6638 21250 6690
rect 23214 6638 23266 6690
rect 23438 6638 23490 6690
rect 37550 6638 37602 6690
rect 38670 6638 38722 6690
rect 41582 6638 41634 6690
rect 52670 6638 52722 6690
rect 54126 6638 54178 6690
rect 3614 6526 3666 6578
rect 4398 6526 4450 6578
rect 21422 6526 21474 6578
rect 23998 6526 24050 6578
rect 37326 6526 37378 6578
rect 37998 6526 38050 6578
rect 38334 6526 38386 6578
rect 39230 6526 39282 6578
rect 41358 6526 41410 6578
rect 42030 6526 42082 6578
rect 53566 6526 53618 6578
rect 55134 6414 55186 6466
rect 3806 6246 3858 6298
rect 3910 6246 3962 6298
rect 4014 6246 4066 6298
rect 23806 6246 23858 6298
rect 23910 6246 23962 6298
rect 24014 6246 24066 6298
rect 43806 6246 43858 6298
rect 43910 6246 43962 6298
rect 44014 6246 44066 6298
rect 53006 6078 53058 6130
rect 56142 6078 56194 6130
rect 13470 5966 13522 6018
rect 14366 5966 14418 6018
rect 15598 5966 15650 6018
rect 19630 5966 19682 6018
rect 20526 5966 20578 6018
rect 31838 5966 31890 6018
rect 54574 5966 54626 6018
rect 13918 5854 13970 5906
rect 14814 5854 14866 5906
rect 20078 5854 20130 5906
rect 52110 5854 52162 5906
rect 53566 5854 53618 5906
rect 55246 5854 55298 5906
rect 30382 5742 30434 5794
rect 30942 5742 30994 5794
rect 32286 5742 32338 5794
rect 15150 5630 15202 5682
rect 30046 5630 30098 5682
rect 32622 5630 32674 5682
rect 4466 5462 4518 5514
rect 4570 5462 4622 5514
rect 4674 5462 4726 5514
rect 24466 5462 24518 5514
rect 24570 5462 24622 5514
rect 24674 5462 24726 5514
rect 44466 5462 44518 5514
rect 44570 5462 44622 5514
rect 44674 5462 44726 5514
rect 2606 5294 2658 5346
rect 2942 5294 2994 5346
rect 15150 5294 15202 5346
rect 28814 5294 28866 5346
rect 52334 5294 52386 5346
rect 2046 5182 2098 5234
rect 3950 5182 4002 5234
rect 6750 5182 6802 5234
rect 12574 5182 12626 5234
rect 13582 5182 13634 5234
rect 27918 5182 27970 5234
rect 28478 5182 28530 5234
rect 47518 5182 47570 5234
rect 51998 5182 52050 5234
rect 52894 5182 52946 5234
rect 54126 5182 54178 5234
rect 4510 5070 4562 5122
rect 4846 5070 4898 5122
rect 7310 5070 7362 5122
rect 7646 5070 7698 5122
rect 13134 5070 13186 5122
rect 14142 5070 14194 5122
rect 14366 5070 14418 5122
rect 14814 5070 14866 5122
rect 46622 5070 46674 5122
rect 46958 5070 47010 5122
rect 51102 5070 51154 5122
rect 51438 5070 51490 5122
rect 53230 5070 53282 5122
rect 54910 5070 54962 5122
rect 53678 4958 53730 5010
rect 3806 4678 3858 4730
rect 3910 4678 3962 4730
rect 4014 4678 4066 4730
rect 23806 4678 23858 4730
rect 23910 4678 23962 4730
rect 24014 4678 24066 4730
rect 43806 4678 43858 4730
rect 43910 4678 43962 4730
rect 44014 4678 44066 4730
rect 54574 4510 54626 4562
rect 56142 4510 56194 4562
rect 4846 4398 4898 4450
rect 13470 4398 13522 4450
rect 36206 4398 36258 4450
rect 36990 4398 37042 4450
rect 39902 4398 39954 4450
rect 41358 4398 41410 4450
rect 49870 4398 49922 4450
rect 51438 4398 51490 4450
rect 51998 4398 52050 4450
rect 52670 4398 52722 4450
rect 53118 4398 53170 4450
rect 5182 4286 5234 4338
rect 36542 4286 36594 4338
rect 41694 4286 41746 4338
rect 52222 4286 52274 4338
rect 5742 4174 5794 4226
rect 42254 4174 42306 4226
rect 53566 4174 53618 4226
rect 55134 4174 55186 4226
rect 39006 4062 39058 4114
rect 39342 4062 39394 4114
rect 48974 4062 49026 4114
rect 49310 4062 49362 4114
rect 4466 3894 4518 3946
rect 4570 3894 4622 3946
rect 4674 3894 4726 3946
rect 24466 3894 24518 3946
rect 24570 3894 24622 3946
rect 24674 3894 24726 3946
rect 44466 3894 44518 3946
rect 44570 3894 44622 3946
rect 44674 3894 44726 3946
rect 9438 3726 9490 3778
rect 9662 3726 9714 3778
rect 18398 3726 18450 3778
rect 18622 3726 18674 3778
rect 33294 3726 33346 3778
rect 35646 3726 35698 3778
rect 36318 3726 36370 3778
rect 36542 3726 36594 3778
rect 43710 3726 43762 3778
rect 43934 3726 43986 3778
rect 51438 3726 51490 3778
rect 51662 3726 51714 3778
rect 8878 3614 8930 3666
rect 15822 3614 15874 3666
rect 32398 3614 32450 3666
rect 32958 3614 33010 3666
rect 35310 3614 35362 3666
rect 37102 3614 37154 3666
rect 50542 3614 50594 3666
rect 52558 3614 52610 3666
rect 54910 3614 54962 3666
rect 10110 3502 10162 3554
rect 10446 3502 10498 3554
rect 15150 3502 15202 3554
rect 49758 3502 49810 3554
rect 49982 3502 50034 3554
rect 54350 3502 54402 3554
rect 11006 3390 11058 3442
rect 15598 3390 15650 3442
rect 19182 3390 19234 3442
rect 34750 3390 34802 3442
rect 44382 3390 44434 3442
rect 52222 3390 52274 3442
rect 53566 3390 53618 3442
rect 3806 3110 3858 3162
rect 3910 3110 3962 3162
rect 4014 3110 4066 3162
rect 23806 3110 23858 3162
rect 23910 3110 23962 3162
rect 24014 3110 24066 3162
rect 43806 3110 43858 3162
rect 43910 3110 43962 3162
rect 44014 3110 44066 3162
rect 54574 2942 54626 2994
rect 56142 2942 56194 2994
rect 21198 2830 21250 2882
rect 22094 2830 22146 2882
rect 28590 2830 28642 2882
rect 29262 2830 29314 2882
rect 32846 2830 32898 2882
rect 37662 2830 37714 2882
rect 21534 2718 21586 2770
rect 24894 2718 24946 2770
rect 25454 2718 25506 2770
rect 25678 2718 25730 2770
rect 29038 2718 29090 2770
rect 31950 2718 32002 2770
rect 32398 2718 32450 2770
rect 37886 2718 37938 2770
rect 52222 2718 52274 2770
rect 53566 2718 53618 2770
rect 3838 2606 3890 2658
rect 38446 2606 38498 2658
rect 52782 2606 52834 2658
rect 55134 2606 55186 2658
rect 4398 2494 4450 2546
rect 4958 2494 5010 2546
rect 4466 2326 4518 2378
rect 4570 2326 4622 2378
rect 4674 2326 4726 2378
rect 24466 2326 24518 2378
rect 24570 2326 24622 2378
rect 24674 2326 24726 2378
rect 44466 2326 44518 2378
rect 44570 2326 44622 2378
rect 44674 2326 44726 2378
rect 6974 2158 7026 2210
rect 7310 2158 7362 2210
rect 14254 2158 14306 2210
rect 14590 2158 14642 2210
rect 17838 2158 17890 2210
rect 18062 2158 18114 2210
rect 21310 2158 21362 2210
rect 21646 2158 21698 2210
rect 28702 2158 28754 2210
rect 28926 2158 28978 2210
rect 2830 2046 2882 2098
rect 20750 2046 20802 2098
rect 25118 2046 25170 2098
rect 29486 2046 29538 2098
rect 52558 2046 52610 2098
rect 54126 2046 54178 2098
rect 54910 2046 54962 2098
rect 2494 1934 2546 1986
rect 3390 1934 3442 1986
rect 3726 1934 3778 1986
rect 24558 1934 24610 1986
rect 30382 1934 30434 1986
rect 30942 1934 30994 1986
rect 51662 1934 51714 1986
rect 2046 1822 2098 1874
rect 6526 1822 6578 1874
rect 13806 1822 13858 1874
rect 17390 1822 17442 1874
rect 24110 1822 24162 1874
rect 31166 1822 31218 1874
rect 51438 1822 51490 1874
rect 52110 1822 52162 1874
rect 53566 1822 53618 1874
rect 3806 1542 3858 1594
rect 3910 1542 3962 1594
rect 4014 1542 4066 1594
rect 23806 1542 23858 1594
rect 23910 1542 23962 1594
rect 24014 1542 24066 1594
rect 43806 1542 43858 1594
rect 43910 1542 43962 1594
rect 44014 1542 44066 1594
rect 53566 1374 53618 1426
rect 56142 1374 56194 1426
rect 2830 1262 2882 1314
rect 51998 1262 52050 1314
rect 50990 1150 51042 1202
rect 52558 1150 52610 1202
rect 55358 1150 55410 1202
rect 4466 758 4518 810
rect 4570 758 4622 810
rect 4674 758 4726 810
rect 24466 758 24518 810
rect 24570 758 24622 810
rect 24674 758 24726 810
rect 44466 758 44518 810
rect 44570 758 44622 810
rect 44674 758 44726 810
<< metal2 >>
rect 672 14112 784 14224
rect 1120 14112 1232 14224
rect 1568 14112 1680 14224
rect 2016 14112 2128 14224
rect 2464 14112 2576 14224
rect 2912 14112 3024 14224
rect 3360 14112 3472 14224
rect 3808 14112 3920 14224
rect 4256 14112 4368 14224
rect 4704 14112 4816 14224
rect 5152 14112 5264 14224
rect 5600 14112 5712 14224
rect 6048 14112 6160 14224
rect 6496 14112 6608 14224
rect 6944 14112 7056 14224
rect 7392 14112 7504 14224
rect 7840 14112 7952 14224
rect 8288 14112 8400 14224
rect 8736 14112 8848 14224
rect 9184 14112 9296 14224
rect 9632 14112 9744 14224
rect 10080 14112 10192 14224
rect 10528 14112 10640 14224
rect 10976 14112 11088 14224
rect 11424 14112 11536 14224
rect 11872 14112 11984 14224
rect 12320 14112 12432 14224
rect 12768 14112 12880 14224
rect 13216 14112 13328 14224
rect 13664 14112 13776 14224
rect 14112 14112 14224 14224
rect 14560 14112 14672 14224
rect 15008 14112 15120 14224
rect 15456 14112 15568 14224
rect 15904 14112 16016 14224
rect 16352 14112 16464 14224
rect 16800 14112 16912 14224
rect 17248 14112 17360 14224
rect 17696 14112 17808 14224
rect 18144 14112 18256 14224
rect 18592 14112 18704 14224
rect 19040 14112 19152 14224
rect 19488 14112 19600 14224
rect 19936 14112 20048 14224
rect 20384 14112 20496 14224
rect 20832 14112 20944 14224
rect 21280 14112 21392 14224
rect 21728 14112 21840 14224
rect 22176 14112 22288 14224
rect 22624 14112 22736 14224
rect 23072 14112 23184 14224
rect 23520 14112 23632 14224
rect 23968 14112 24080 14224
rect 24416 14112 24528 14224
rect 24864 14112 24976 14224
rect 25312 14112 25424 14224
rect 25760 14112 25872 14224
rect 26208 14112 26320 14224
rect 26656 14112 26768 14224
rect 27104 14112 27216 14224
rect 27552 14112 27664 14224
rect 28000 14112 28112 14224
rect 28448 14112 28560 14224
rect 28896 14112 29008 14224
rect 29344 14112 29456 14224
rect 29792 14112 29904 14224
rect 30240 14112 30352 14224
rect 30688 14112 30800 14224
rect 31136 14112 31248 14224
rect 31584 14112 31696 14224
rect 31836 14196 31892 14206
rect 364 13076 420 13086
rect 252 12068 308 12078
rect 140 12012 252 12068
rect 140 5460 196 12012
rect 252 12002 308 12012
rect 364 8372 420 13020
rect 700 9716 756 14112
rect 924 12628 980 12638
rect 700 9650 756 9660
rect 812 10836 868 10846
rect 812 9492 868 10780
rect 924 9828 980 12572
rect 1036 12180 1092 12190
rect 1036 10836 1092 12124
rect 1148 11844 1204 14112
rect 1148 11778 1204 11788
rect 1484 13972 1540 13982
rect 1484 11732 1540 13916
rect 1596 11844 1652 14112
rect 2044 12068 2100 14112
rect 2156 13412 2212 13422
rect 2156 13186 2212 13356
rect 2156 13134 2158 13186
rect 2210 13134 2212 13186
rect 2156 13122 2212 13134
rect 2268 12404 2324 12414
rect 2268 12310 2324 12348
rect 2044 12012 2212 12068
rect 1596 11788 1876 11844
rect 1484 11676 1652 11732
rect 1484 11394 1540 11406
rect 1484 11342 1486 11394
rect 1538 11342 1540 11394
rect 1260 11284 1316 11294
rect 1484 11284 1540 11342
rect 1036 10770 1092 10780
rect 1148 11282 1540 11284
rect 1148 11230 1262 11282
rect 1314 11230 1540 11282
rect 1148 11228 1540 11230
rect 924 9762 980 9772
rect 1036 10388 1092 10398
rect 812 9426 868 9436
rect 364 8306 420 8316
rect 140 5394 196 5404
rect 588 6916 644 6926
rect 588 3668 644 6860
rect 1036 5236 1092 10332
rect 1036 5170 1092 5180
rect 1148 4564 1204 11228
rect 1260 11218 1316 11228
rect 1372 10386 1428 10398
rect 1372 10334 1374 10386
rect 1426 10334 1428 10386
rect 1260 9828 1316 9838
rect 1372 9828 1428 10334
rect 1596 10388 1652 11676
rect 1596 10322 1652 10332
rect 1484 9940 1540 9950
rect 1484 9938 1764 9940
rect 1484 9886 1486 9938
rect 1538 9886 1764 9938
rect 1484 9884 1764 9886
rect 1484 9874 1540 9884
rect 1260 9826 1428 9828
rect 1260 9774 1262 9826
rect 1314 9774 1428 9826
rect 1260 9772 1428 9774
rect 1260 4676 1316 9772
rect 1484 9716 1540 9726
rect 1484 8370 1540 9660
rect 1484 8318 1486 8370
rect 1538 8318 1540 8370
rect 1484 8306 1540 8318
rect 1484 8148 1540 8158
rect 1484 4900 1540 8092
rect 1708 5124 1764 9884
rect 1820 9716 1876 11788
rect 2044 11508 2100 11518
rect 2044 11414 2100 11452
rect 2156 10722 2212 12012
rect 2156 10670 2158 10722
rect 2210 10670 2212 10722
rect 2156 10658 2212 10670
rect 2268 11844 2324 11854
rect 2044 9716 2100 9726
rect 1820 9714 2100 9716
rect 1820 9662 2046 9714
rect 2098 9662 2100 9714
rect 1820 9660 2100 9662
rect 2044 9650 2100 9660
rect 1820 9492 1876 9502
rect 2268 9492 2324 11788
rect 2492 11284 2548 14112
rect 2716 12962 2772 12974
rect 2716 12910 2718 12962
rect 2770 12910 2772 12962
rect 2604 11284 2660 11294
rect 2492 11282 2660 11284
rect 2492 11230 2606 11282
rect 2658 11230 2660 11282
rect 2492 11228 2660 11230
rect 2604 11218 2660 11228
rect 1820 7588 1876 9436
rect 2044 9436 2324 9492
rect 2380 10724 2436 10734
rect 2044 9266 2100 9436
rect 2044 9214 2046 9266
rect 2098 9214 2100 9266
rect 2044 9202 2100 9214
rect 2380 9044 2436 10668
rect 2380 8978 2436 8988
rect 2492 10612 2548 10622
rect 1820 7522 1876 7532
rect 2044 8932 2100 8942
rect 1708 5058 1764 5068
rect 1820 5236 1876 5246
rect 1484 4834 1540 4844
rect 1596 5012 1652 5022
rect 1260 4620 1428 4676
rect 1148 4508 1316 4564
rect 588 3602 644 3612
rect 1148 3780 1204 3790
rect 1036 3444 1092 3454
rect 1036 980 1092 3388
rect 1036 914 1092 924
rect 1148 84 1204 3724
rect 1260 980 1316 4508
rect 1260 914 1316 924
rect 1372 196 1428 4620
rect 1596 2996 1652 4956
rect 1596 2930 1652 2940
rect 1708 4340 1764 4350
rect 1708 1764 1764 4284
rect 1596 1708 1764 1764
rect 1596 532 1652 1708
rect 1820 1092 1876 5180
rect 2044 5234 2100 8876
rect 2492 8820 2548 10556
rect 2044 5182 2046 5234
rect 2098 5182 2100 5234
rect 2044 5170 2100 5182
rect 2156 8764 2548 8820
rect 2604 8930 2660 8942
rect 2604 8878 2606 8930
rect 2658 8878 2660 8930
rect 2044 1876 2100 1886
rect 2156 1876 2212 8764
rect 2604 8596 2660 8878
rect 2604 8530 2660 8540
rect 2716 8428 2772 12910
rect 2940 12180 2996 14112
rect 2940 12114 2996 12124
rect 3164 13972 3220 13982
rect 2828 12066 2884 12078
rect 2828 12014 2830 12066
rect 2882 12014 2884 12066
rect 2828 11284 2884 12014
rect 2828 11228 2996 11284
rect 2492 8372 2772 8428
rect 2828 10498 2884 10510
rect 2828 10446 2830 10498
rect 2882 10446 2884 10498
rect 2268 8260 2324 8270
rect 2268 8166 2324 8204
rect 2492 2548 2548 8372
rect 2828 6132 2884 10446
rect 2940 10500 2996 11228
rect 2940 10434 2996 10444
rect 3052 9828 3108 9838
rect 3052 9734 3108 9772
rect 3052 9156 3108 9166
rect 3164 9156 3220 13916
rect 3388 12404 3444 14112
rect 3388 12338 3444 12348
rect 3612 13524 3668 13534
rect 3612 12290 3668 13468
rect 3724 13188 3780 13198
rect 3724 13094 3780 13132
rect 3836 12740 3892 14112
rect 4284 13412 4340 14112
rect 4732 13524 4788 14112
rect 4732 13458 4788 13468
rect 4284 13346 4340 13356
rect 4464 13356 4728 13366
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4464 13290 4728 13300
rect 4284 12964 4340 12974
rect 4284 12870 4340 12908
rect 4956 12964 5012 12974
rect 3836 12684 4340 12740
rect 3804 12572 4068 12582
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 3804 12506 4068 12516
rect 3612 12238 3614 12290
rect 3666 12238 3668 12290
rect 3612 12226 3668 12238
rect 3388 12180 3444 12190
rect 3388 10834 3444 12124
rect 3612 11394 3668 11406
rect 3612 11342 3614 11394
rect 3666 11342 3668 11394
rect 3612 11172 3668 11342
rect 3612 11106 3668 11116
rect 3804 11004 4068 11014
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 3804 10938 4068 10948
rect 3388 10782 3390 10834
rect 3442 10782 3444 10834
rect 3388 10770 3444 10782
rect 4172 10610 4228 10622
rect 4172 10558 4174 10610
rect 4226 10558 4228 10610
rect 4172 9492 4228 10558
rect 4284 9714 4340 12684
rect 4396 12068 4452 12078
rect 4396 12066 4900 12068
rect 4396 12014 4398 12066
rect 4450 12014 4900 12066
rect 4396 12012 4900 12014
rect 4396 12002 4452 12012
rect 4464 11788 4728 11798
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4464 11722 4728 11732
rect 4620 11620 4676 11630
rect 4620 11526 4676 11564
rect 4464 10220 4728 10230
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4464 10154 4728 10164
rect 4284 9662 4286 9714
rect 4338 9662 4340 9714
rect 4284 9650 4340 9662
rect 3804 9436 4068 9446
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 4172 9426 4228 9436
rect 3804 9370 4068 9380
rect 3052 9154 3220 9156
rect 3052 9102 3054 9154
rect 3106 9102 3220 9154
rect 3052 9100 3220 9102
rect 3052 9090 3108 9100
rect 3500 8820 3556 8830
rect 3724 8820 3780 8830
rect 3500 8818 3780 8820
rect 3500 8766 3502 8818
rect 3554 8766 3726 8818
rect 3778 8766 3780 8818
rect 3500 8764 3780 8766
rect 3500 8754 3556 8764
rect 3388 8708 3444 8718
rect 2828 6066 2884 6076
rect 2940 7700 2996 7710
rect 2716 5684 2772 5694
rect 2604 5348 2660 5358
rect 2604 5254 2660 5292
rect 2492 2482 2548 2492
rect 2044 1874 2212 1876
rect 2044 1822 2046 1874
rect 2098 1822 2212 1874
rect 2044 1820 2212 1822
rect 2492 1986 2548 1998
rect 2492 1934 2494 1986
rect 2546 1934 2548 1986
rect 2044 1810 2100 1820
rect 2492 1316 2548 1934
rect 2716 1876 2772 5628
rect 2940 5572 2996 7644
rect 2828 5516 2996 5572
rect 2828 2098 2884 5516
rect 2940 5348 2996 5358
rect 2940 5254 2996 5292
rect 3388 4452 3444 8652
rect 3724 8372 3780 8764
rect 4464 8652 4728 8662
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4464 8586 4728 8596
rect 3724 8306 3780 8316
rect 3804 7868 4068 7878
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 3804 7802 4068 7812
rect 3500 7364 3556 7374
rect 3500 6132 3556 7308
rect 4464 7084 4728 7094
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4464 7018 4728 7028
rect 4060 6692 4116 6702
rect 4060 6690 4228 6692
rect 4060 6638 4062 6690
rect 4114 6638 4228 6690
rect 4060 6636 4228 6638
rect 4060 6626 4116 6636
rect 3612 6580 3668 6590
rect 3612 6486 3668 6524
rect 4172 6580 4228 6636
rect 4396 6580 4452 6590
rect 4172 6578 4452 6580
rect 4172 6526 4398 6578
rect 4450 6526 4452 6578
rect 4172 6524 4452 6526
rect 3804 6300 4068 6310
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 3804 6234 4068 6244
rect 3500 6076 4004 6132
rect 3948 5234 4004 6076
rect 3948 5182 3950 5234
rect 4002 5182 4004 5234
rect 3948 5170 4004 5182
rect 3804 4732 4068 4742
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 3804 4666 4068 4676
rect 4172 4676 4228 6524
rect 4396 6514 4452 6524
rect 4464 5516 4728 5526
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4464 5450 4728 5460
rect 4844 5338 4900 12012
rect 4956 11396 5012 12908
rect 5180 12180 5236 14112
rect 5628 13188 5684 14112
rect 5628 13122 5684 13132
rect 5964 13300 6020 13310
rect 5964 13186 6020 13244
rect 5964 13134 5966 13186
rect 6018 13134 6020 13186
rect 5964 13122 6020 13134
rect 5964 12852 6020 12862
rect 5964 12290 6020 12796
rect 5964 12238 5966 12290
rect 6018 12238 6020 12290
rect 5964 12226 6020 12238
rect 5068 12124 5236 12180
rect 5516 12180 5572 12190
rect 5516 12178 5908 12180
rect 5516 12126 5518 12178
rect 5570 12126 5908 12178
rect 5516 12124 5908 12126
rect 5068 11620 5124 12124
rect 5516 12114 5572 12124
rect 5180 11956 5236 11966
rect 5404 11956 5460 11966
rect 5180 11954 5460 11956
rect 5180 11902 5182 11954
rect 5234 11902 5406 11954
rect 5458 11902 5460 11954
rect 5180 11900 5460 11902
rect 5180 11890 5236 11900
rect 5404 11890 5460 11900
rect 5068 11554 5124 11564
rect 4956 11340 5124 11396
rect 4956 9268 5012 9278
rect 4956 6916 5012 9212
rect 4956 6850 5012 6860
rect 4844 5282 5012 5338
rect 4956 5236 5012 5282
rect 4956 5170 5012 5180
rect 4508 5124 4564 5134
rect 4844 5124 4900 5134
rect 4508 5122 4900 5124
rect 4508 5070 4510 5122
rect 4562 5070 4846 5122
rect 4898 5070 4900 5122
rect 4508 5068 4900 5070
rect 4508 5058 4564 5068
rect 4172 4610 4228 4620
rect 4396 4900 4452 4910
rect 3388 4386 3444 4396
rect 3276 4116 3332 4126
rect 3276 2884 3332 4060
rect 4396 4116 4452 4844
rect 4844 4900 4900 5068
rect 5068 5012 5124 11340
rect 5180 11394 5236 11406
rect 5180 11342 5182 11394
rect 5234 11342 5236 11394
rect 5180 5572 5236 11342
rect 5740 10052 5796 10062
rect 5740 9938 5796 9996
rect 5740 9886 5742 9938
rect 5794 9886 5796 9938
rect 5740 9874 5796 9886
rect 5292 9826 5348 9838
rect 5292 9774 5294 9826
rect 5346 9774 5348 9826
rect 5292 8596 5348 9774
rect 5292 8530 5348 8540
rect 5740 8258 5796 8270
rect 5740 8206 5742 8258
rect 5794 8206 5796 8258
rect 5180 5506 5236 5516
rect 5404 8148 5460 8158
rect 5740 8148 5796 8206
rect 5404 8146 5796 8148
rect 5404 8094 5406 8146
rect 5458 8094 5796 8146
rect 5404 8092 5796 8094
rect 5068 4946 5124 4956
rect 4844 4834 4900 4844
rect 4844 4452 4900 4462
rect 4844 4358 4900 4396
rect 5180 4452 5236 4462
rect 5180 4338 5236 4396
rect 5180 4286 5182 4338
rect 5234 4286 5236 4338
rect 5180 4274 5236 4286
rect 4396 4050 4452 4060
rect 4464 3948 4728 3958
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4464 3882 4728 3892
rect 3804 3164 4068 3174
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 3804 3098 4068 3108
rect 3276 2818 3332 2828
rect 3836 2660 3892 2670
rect 3836 2566 3892 2604
rect 4396 2548 4452 2586
rect 4396 2482 4452 2492
rect 4956 2548 5012 2558
rect 5012 2492 5124 2548
rect 4956 2454 5012 2492
rect 4464 2380 4728 2390
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4464 2314 4728 2324
rect 2828 2046 2830 2098
rect 2882 2046 2884 2098
rect 2828 2034 2884 2046
rect 3388 1988 3444 1998
rect 3388 1894 3444 1932
rect 3724 1988 3780 1998
rect 3724 1894 3780 1932
rect 2716 1810 2772 1820
rect 5068 1652 5124 2492
rect 3804 1596 4068 1606
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 5068 1586 5124 1596
rect 3804 1530 4068 1540
rect 2492 1250 2548 1260
rect 2828 1316 2884 1326
rect 2828 1222 2884 1260
rect 1820 1026 1876 1036
rect 4464 812 4728 822
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4464 746 4728 756
rect 1596 466 1652 476
rect 4508 644 4564 654
rect 1372 130 1428 140
rect 1820 196 1876 206
rect 1820 112 1876 140
rect 4508 112 4564 588
rect 5404 644 5460 8092
rect 5740 4228 5796 4238
rect 5740 4134 5796 4172
rect 5852 1204 5908 12124
rect 5964 11844 6020 11854
rect 5964 7364 6020 11788
rect 6076 10722 6132 14112
rect 6524 13188 6580 14112
rect 6188 13132 6580 13188
rect 6636 13748 6692 13758
rect 6188 11618 6244 13132
rect 6524 12964 6580 12974
rect 6524 12870 6580 12908
rect 6636 12292 6692 13692
rect 6972 12628 7028 14112
rect 7420 13300 7476 14112
rect 7420 13234 7476 13244
rect 7532 13188 7588 13198
rect 7532 13094 7588 13132
rect 6972 12572 7476 12628
rect 6972 12404 7028 12414
rect 6972 12310 7028 12348
rect 6524 12236 6692 12292
rect 6524 11844 6580 12236
rect 6524 11778 6580 11788
rect 6636 12068 6692 12078
rect 6188 11566 6190 11618
rect 6242 11566 6244 11618
rect 6188 11554 6244 11566
rect 6636 11394 6692 12012
rect 6636 11342 6638 11394
rect 6690 11342 6692 11394
rect 6636 11330 6692 11342
rect 7420 10834 7476 12572
rect 7868 12404 7924 14112
rect 8092 13076 8148 13086
rect 8092 12982 8148 13020
rect 8316 12404 8372 14112
rect 8652 12516 8708 12526
rect 7868 12338 7924 12348
rect 7980 12348 8372 12404
rect 8540 12404 8596 12414
rect 7532 12180 7588 12190
rect 7532 12086 7588 12124
rect 7756 11620 7812 11630
rect 7980 11620 8036 12348
rect 8540 12310 8596 12348
rect 7756 11618 8036 11620
rect 7756 11566 7758 11618
rect 7810 11566 8036 11618
rect 7756 11564 8036 11566
rect 7756 11554 7812 11564
rect 7420 10782 7422 10834
rect 7474 10782 7476 10834
rect 7420 10770 7476 10782
rect 8092 11394 8148 11406
rect 8092 11342 8094 11394
rect 8146 11342 8148 11394
rect 6076 10670 6078 10722
rect 6130 10670 6132 10722
rect 6076 10658 6132 10670
rect 6860 10498 6916 10510
rect 6860 10446 6862 10498
rect 6914 10446 6916 10498
rect 6300 9826 6356 9838
rect 6300 9774 6302 9826
rect 6354 9774 6356 9826
rect 6300 9716 6356 9774
rect 6636 9716 6692 9726
rect 6300 9714 6692 9716
rect 6300 9662 6638 9714
rect 6690 9662 6692 9714
rect 6300 9660 6692 9662
rect 6188 9604 6244 9614
rect 6076 9156 6132 9166
rect 6076 9062 6132 9100
rect 6188 7476 6244 9548
rect 6524 8820 6580 8830
rect 6524 8726 6580 8764
rect 6412 8372 6468 8382
rect 6188 7410 6244 7420
rect 6300 8146 6356 8158
rect 6300 8094 6302 8146
rect 6354 8094 6356 8146
rect 5964 7298 6020 7308
rect 6300 6804 6356 8094
rect 6300 6738 6356 6748
rect 6188 6580 6244 6590
rect 6076 5796 6132 5806
rect 6076 3780 6132 5740
rect 6188 4116 6244 6524
rect 6300 6244 6356 6254
rect 6300 4340 6356 6188
rect 6300 4274 6356 4284
rect 6188 4050 6244 4060
rect 6076 3714 6132 3724
rect 5852 1138 5908 1148
rect 6412 868 6468 8316
rect 6524 6916 6580 6926
rect 6524 4564 6580 6860
rect 6524 4498 6580 4508
rect 6636 3444 6692 9660
rect 6748 8820 6804 8830
rect 6748 8726 6804 8764
rect 6860 6468 6916 10446
rect 7532 10388 7588 10398
rect 6860 6402 6916 6412
rect 6972 10276 7028 10286
rect 6972 6244 7028 10220
rect 6748 6188 7028 6244
rect 7196 9716 7252 9726
rect 6748 5234 6804 6188
rect 6748 5182 6750 5234
rect 6802 5182 6804 5234
rect 6748 5170 6804 5182
rect 6860 5908 6916 5918
rect 6860 4564 6916 5852
rect 6860 4498 6916 4508
rect 6636 3378 6692 3388
rect 6748 4452 6804 4462
rect 6748 3332 6804 4396
rect 6748 3266 6804 3276
rect 6972 2212 7028 2222
rect 7196 2212 7252 9660
rect 7532 9268 7588 10332
rect 7532 9202 7588 9212
rect 7980 9380 8036 9390
rect 7868 8820 7924 8830
rect 7308 5124 7364 5134
rect 7644 5124 7700 5134
rect 7308 5122 7700 5124
rect 7308 5070 7310 5122
rect 7362 5070 7646 5122
rect 7698 5070 7700 5122
rect 7308 5068 7700 5070
rect 7308 5058 7364 5068
rect 7644 4340 7700 5068
rect 7644 4274 7700 4284
rect 7420 2660 7476 2670
rect 7308 2212 7364 2222
rect 6972 2210 7364 2212
rect 6972 2158 6974 2210
rect 7026 2158 7310 2210
rect 7362 2158 7364 2210
rect 6972 2156 7364 2158
rect 6972 2146 7028 2156
rect 7308 2146 7364 2156
rect 6524 1876 6580 1886
rect 6524 1782 6580 1820
rect 6412 802 6468 812
rect 7196 1652 7252 1662
rect 5404 578 5460 588
rect 7196 112 7252 1596
rect 7420 1316 7476 2604
rect 7420 1250 7476 1260
rect 7868 644 7924 8764
rect 7980 5796 8036 9324
rect 8092 8708 8148 11342
rect 8540 10724 8596 10734
rect 8092 8642 8148 8652
rect 8204 10610 8260 10622
rect 8204 10558 8206 10610
rect 8258 10558 8260 10610
rect 7980 5730 8036 5740
rect 8204 3388 8260 10558
rect 8316 9492 8372 9502
rect 8316 8260 8372 9436
rect 8316 8194 8372 8204
rect 8428 7476 8484 7486
rect 8428 3892 8484 7420
rect 8540 5908 8596 10668
rect 8652 9156 8708 12460
rect 8764 11818 8820 14112
rect 8988 14084 9044 14094
rect 8988 11956 9044 14028
rect 9212 13188 9268 14112
rect 9212 13122 9268 13132
rect 9212 12964 9268 12974
rect 8988 11890 9044 11900
rect 9100 12066 9156 12078
rect 9100 12014 9102 12066
rect 9154 12014 9156 12066
rect 8764 11762 9044 11818
rect 8988 10834 9044 11762
rect 8988 10782 8990 10834
rect 9042 10782 9044 10834
rect 8988 10770 9044 10782
rect 8652 9090 8708 9100
rect 8876 8820 8932 8830
rect 8876 8370 8932 8764
rect 8876 8318 8878 8370
rect 8930 8318 8932 8370
rect 8876 8306 8932 8318
rect 9100 7924 9156 12014
rect 9212 11508 9268 12908
rect 9436 12964 9492 12974
rect 9212 11442 9268 11452
rect 9324 12628 9380 12638
rect 9212 10500 9268 10510
rect 9212 8036 9268 10444
rect 9324 10164 9380 12572
rect 9324 10098 9380 10108
rect 9436 9938 9492 12908
rect 9436 9886 9438 9938
rect 9490 9886 9492 9938
rect 9436 9874 9492 9886
rect 9548 12740 9604 12750
rect 9548 8820 9604 12684
rect 9660 12404 9716 14112
rect 9772 13188 9828 13198
rect 9772 13094 9828 13132
rect 10108 12628 10164 14112
rect 10332 13300 10388 13310
rect 10332 13074 10388 13244
rect 10332 13022 10334 13074
rect 10386 13022 10388 13074
rect 10332 13010 10388 13022
rect 9660 12338 9716 12348
rect 9996 12572 10164 12628
rect 9996 12180 10052 12572
rect 10108 12404 10164 12414
rect 10556 12404 10612 14112
rect 10780 13524 10836 13534
rect 10108 12402 10612 12404
rect 10108 12350 10110 12402
rect 10162 12350 10612 12402
rect 10108 12348 10612 12350
rect 10668 12404 10724 12414
rect 10108 12338 10164 12348
rect 9996 12124 10612 12180
rect 10108 11956 10164 11966
rect 10108 11396 10164 11900
rect 10108 11330 10164 11340
rect 10332 11396 10388 11406
rect 9996 10498 10052 10510
rect 9996 10446 9998 10498
rect 10050 10446 10052 10498
rect 9996 10164 10052 10446
rect 10332 10276 10388 11340
rect 10556 10834 10612 12124
rect 10668 12178 10724 12348
rect 10668 12126 10670 12178
rect 10722 12126 10724 12178
rect 10668 12114 10724 12126
rect 10556 10782 10558 10834
rect 10610 10782 10612 10834
rect 10556 10770 10612 10782
rect 10780 10388 10836 13468
rect 10892 11620 10948 11630
rect 11004 11620 11060 14112
rect 11340 13412 11396 13422
rect 11340 13186 11396 13356
rect 11340 13134 11342 13186
rect 11394 13134 11396 13186
rect 11340 13122 11396 13134
rect 11452 13188 11508 14112
rect 11900 13188 11956 14112
rect 11452 13122 11508 13132
rect 11788 13132 11956 13188
rect 12236 13860 12292 13870
rect 11564 13076 11620 13086
rect 10892 11618 11060 11620
rect 10892 11566 10894 11618
rect 10946 11566 11060 11618
rect 10892 11564 11060 11566
rect 11116 12292 11172 12302
rect 10892 11554 10948 11564
rect 10332 10210 10388 10220
rect 10668 10332 10836 10388
rect 9996 10098 10052 10108
rect 9996 9828 10052 9838
rect 10332 9828 10388 9838
rect 9996 9826 10164 9828
rect 9996 9774 9998 9826
rect 10050 9774 10164 9826
rect 9996 9772 10164 9774
rect 9996 9762 10052 9772
rect 10108 9268 10164 9772
rect 10332 9734 10388 9772
rect 10108 9154 10164 9212
rect 10108 9102 10110 9154
rect 10162 9102 10164 9154
rect 10108 9090 10164 9102
rect 9548 8754 9604 8764
rect 10108 8932 10164 8942
rect 9436 8258 9492 8270
rect 9436 8206 9438 8258
rect 9490 8206 9492 8258
rect 9436 8148 9492 8206
rect 9772 8148 9828 8158
rect 9436 8146 9828 8148
rect 9436 8094 9774 8146
rect 9826 8094 9828 8146
rect 9436 8092 9828 8094
rect 9212 7970 9268 7980
rect 9100 7858 9156 7868
rect 9660 7588 9716 7598
rect 9660 7494 9716 7532
rect 9660 6916 9716 6926
rect 9324 6804 9380 6814
rect 8764 6692 8820 6702
rect 8764 6132 8820 6636
rect 8764 6066 8820 6076
rect 9212 6356 9268 6366
rect 9212 6020 9268 6300
rect 9212 5954 9268 5964
rect 8540 5852 8820 5908
rect 8428 3826 8484 3836
rect 8652 4564 8708 4574
rect 8092 3332 8260 3388
rect 8092 2100 8148 3332
rect 8092 2034 8148 2044
rect 8652 1428 8708 4508
rect 8764 3332 8820 5852
rect 9212 5460 9268 5470
rect 9212 4788 9268 5404
rect 9212 4722 9268 4732
rect 8876 3780 8932 3790
rect 8876 3666 8932 3724
rect 8876 3614 8878 3666
rect 8930 3614 8932 3666
rect 8876 3602 8932 3614
rect 8764 3266 8820 3276
rect 9324 2884 9380 6748
rect 9660 5796 9716 6860
rect 9772 6356 9828 8092
rect 10108 8148 10164 8876
rect 10332 8932 10388 8942
rect 10332 8838 10388 8876
rect 10108 8082 10164 8092
rect 10668 7812 10724 10332
rect 11116 10276 11172 12236
rect 11116 10210 11172 10220
rect 11452 11394 11508 11406
rect 11452 11342 11454 11394
rect 11506 11342 11508 11394
rect 10668 7746 10724 7756
rect 10780 9826 10836 9838
rect 10780 9774 10782 9826
rect 10834 9774 10836 9826
rect 10780 9716 10836 9774
rect 11116 9716 11172 9726
rect 10780 9714 11172 9716
rect 10780 9662 11118 9714
rect 11170 9662 11172 9714
rect 10780 9660 11172 9662
rect 9996 7588 10052 7598
rect 9996 7474 10052 7532
rect 9996 7422 9998 7474
rect 10050 7422 10052 7474
rect 9996 7410 10052 7422
rect 10556 7364 10612 7374
rect 10556 7270 10612 7308
rect 9772 6290 9828 6300
rect 9660 5730 9716 5740
rect 10220 6132 10276 6142
rect 9884 5236 9940 5246
rect 9884 4564 9940 5180
rect 9884 4498 9940 4508
rect 10108 5236 10164 5246
rect 9996 4004 10052 4014
rect 10108 4004 10164 5180
rect 10220 4228 10276 6076
rect 10220 4162 10276 4172
rect 10668 4228 10724 4238
rect 10052 3948 10164 4004
rect 9996 3938 10052 3948
rect 9436 3780 9492 3790
rect 9660 3780 9716 3790
rect 9436 3778 10612 3780
rect 9436 3726 9438 3778
rect 9490 3726 9662 3778
rect 9714 3726 10612 3778
rect 9436 3724 10612 3726
rect 9436 3714 9492 3724
rect 9660 3714 9716 3724
rect 10108 3556 10164 3566
rect 10444 3556 10500 3566
rect 10108 3554 10500 3556
rect 10108 3502 10110 3554
rect 10162 3502 10446 3554
rect 10498 3502 10500 3554
rect 10108 3500 10500 3502
rect 10108 3388 10164 3500
rect 10444 3490 10500 3500
rect 9996 3332 10164 3388
rect 9324 2818 9380 2828
rect 9884 3276 10052 3332
rect 8652 1362 8708 1372
rect 7868 578 7924 588
rect 9884 112 9940 3276
rect 10556 1652 10612 3724
rect 10668 3444 10724 4172
rect 10668 3378 10724 3388
rect 10556 1586 10612 1596
rect 10780 420 10836 9660
rect 11116 9650 11172 9660
rect 10892 8820 10948 8830
rect 11228 8820 11284 8830
rect 10892 8818 11284 8820
rect 10892 8766 10894 8818
rect 10946 8766 11230 8818
rect 11282 8766 11284 8818
rect 10892 8764 11284 8766
rect 10892 8754 10948 8764
rect 10892 8148 10948 8158
rect 10892 2772 10948 8092
rect 11228 5684 11284 8764
rect 11452 8148 11508 11342
rect 11564 10724 11620 13020
rect 11676 12404 11732 12414
rect 11788 12404 11844 13132
rect 11676 12402 11844 12404
rect 11676 12350 11678 12402
rect 11730 12350 11844 12402
rect 11676 12348 11844 12350
rect 11900 12962 11956 12974
rect 11900 12910 11902 12962
rect 11954 12910 11956 12962
rect 11676 12338 11732 12348
rect 11564 10668 11732 10724
rect 11564 10500 11620 10510
rect 11564 10406 11620 10444
rect 11676 8820 11732 10668
rect 11900 9716 11956 12910
rect 11900 9650 11956 9660
rect 12012 12180 12068 12190
rect 11676 8754 11732 8764
rect 11788 9156 11844 9166
rect 11452 8082 11508 8092
rect 11788 7476 11844 9100
rect 12012 7812 12068 12124
rect 12236 12178 12292 13804
rect 12236 12126 12238 12178
rect 12290 12126 12292 12178
rect 12236 12114 12292 12126
rect 12348 11282 12404 14112
rect 12684 13188 12740 13198
rect 12684 12068 12740 13132
rect 12796 12292 12852 14112
rect 13244 13412 13300 14112
rect 13244 13346 13300 13356
rect 13692 13300 13748 14112
rect 13692 13244 13972 13300
rect 13692 13076 13748 13086
rect 13692 12982 13748 13020
rect 12908 12964 12964 12974
rect 12908 12870 12964 12908
rect 13580 12516 13636 12526
rect 13356 12292 13412 12302
rect 12796 12236 12964 12292
rect 12796 12068 12852 12078
rect 12684 12066 12852 12068
rect 12684 12014 12798 12066
rect 12850 12014 12852 12066
rect 12684 12012 12852 12014
rect 12796 12002 12852 12012
rect 12348 11230 12350 11282
rect 12402 11230 12404 11282
rect 12348 11218 12404 11230
rect 12908 10836 12964 12236
rect 13356 12178 13412 12236
rect 13356 12126 13358 12178
rect 13410 12126 13412 12178
rect 13356 12114 13412 12126
rect 13468 12180 13524 12190
rect 13020 11508 13076 11518
rect 13468 11508 13524 12124
rect 13580 11732 13636 12460
rect 13804 12404 13860 12414
rect 13692 12292 13748 12330
rect 13692 12226 13748 12236
rect 13580 11666 13636 11676
rect 13692 12068 13748 12078
rect 13020 11506 13524 11508
rect 13020 11454 13022 11506
rect 13074 11454 13524 11506
rect 13020 11452 13524 11454
rect 13020 11442 13076 11452
rect 13580 11394 13636 11406
rect 13580 11342 13582 11394
rect 13634 11342 13636 11394
rect 13020 10836 13076 10846
rect 12908 10834 13076 10836
rect 12908 10782 13022 10834
rect 13074 10782 13076 10834
rect 12908 10780 13076 10782
rect 13020 10770 13076 10780
rect 12572 10724 12628 10734
rect 12460 10164 12516 10174
rect 12460 9940 12516 10108
rect 12460 9874 12516 9884
rect 12012 7746 12068 7756
rect 11676 7420 11844 7476
rect 11900 7476 11956 7486
rect 11676 5908 11732 7420
rect 11900 6132 11956 7420
rect 11900 6066 11956 6076
rect 11676 5842 11732 5852
rect 11788 6020 11844 6030
rect 11228 5618 11284 5628
rect 11788 4004 11844 5964
rect 12572 5234 12628 10668
rect 13244 10276 13300 10286
rect 13132 9604 13188 9614
rect 13020 8932 13076 8942
rect 12572 5182 12574 5234
rect 12626 5182 12628 5234
rect 12572 5170 12628 5182
rect 12796 7364 12852 7374
rect 11788 3938 11844 3948
rect 12572 4676 12628 4686
rect 11004 3444 11060 3482
rect 11004 3378 11060 3388
rect 10892 2706 10948 2716
rect 11116 3332 11172 3342
rect 11116 1540 11172 3276
rect 11116 1474 11172 1484
rect 10780 354 10836 364
rect 12572 112 12628 4620
rect 12796 3332 12852 7308
rect 13020 7252 13076 8876
rect 13132 7364 13188 9548
rect 13244 8932 13300 10220
rect 13244 8866 13300 8876
rect 13468 8372 13524 8382
rect 13468 7588 13524 8316
rect 13468 7522 13524 7532
rect 13132 7298 13188 7308
rect 13020 7186 13076 7196
rect 12908 7140 12964 7150
rect 12908 6132 12964 7084
rect 12908 6066 12964 6076
rect 13468 6020 13524 6030
rect 13580 6020 13636 11342
rect 13692 10276 13748 12012
rect 13804 10388 13860 12348
rect 13916 11618 13972 13244
rect 14028 12404 14084 12414
rect 14028 12180 14084 12348
rect 14028 12114 14084 12124
rect 13916 11566 13918 11618
rect 13970 11566 13972 11618
rect 13916 11554 13972 11566
rect 14140 10836 14196 14112
rect 14588 13076 14644 14112
rect 14588 13010 14644 13020
rect 14924 13076 14980 13086
rect 14924 12982 14980 13020
rect 14140 10770 14196 10780
rect 14252 12516 14308 12526
rect 13804 10322 13860 10332
rect 14028 10498 14084 10510
rect 14028 10446 14030 10498
rect 14082 10446 14084 10498
rect 13692 10210 13748 10220
rect 14028 10164 14084 10446
rect 14028 10098 14084 10108
rect 14252 10052 14308 12460
rect 14812 12404 14868 12414
rect 15036 12404 15092 14112
rect 15260 13860 15316 13870
rect 14812 12402 15092 12404
rect 14812 12350 14814 12402
rect 14866 12350 15092 12402
rect 14812 12348 15092 12350
rect 15148 13748 15204 13758
rect 14812 12338 14868 12348
rect 15148 11844 15204 13692
rect 15148 11778 15204 11788
rect 14924 11396 14980 11406
rect 14252 9986 14308 9996
rect 14364 11394 14980 11396
rect 14364 11342 14926 11394
rect 14978 11342 14980 11394
rect 14364 11340 14980 11342
rect 14252 8932 14308 8942
rect 13692 8708 13748 8718
rect 13692 7028 13748 8652
rect 13692 6962 13748 6972
rect 14140 7028 14196 7038
rect 13468 6018 13636 6020
rect 13468 5966 13470 6018
rect 13522 5966 13636 6018
rect 13468 5964 13636 5966
rect 13804 6804 13860 6814
rect 13468 5954 13524 5964
rect 13580 5348 13636 5358
rect 13580 5234 13636 5292
rect 13580 5182 13582 5234
rect 13634 5182 13636 5234
rect 13580 5170 13636 5182
rect 13132 5124 13188 5134
rect 13132 5122 13524 5124
rect 13132 5070 13134 5122
rect 13186 5070 13524 5122
rect 13132 5068 13524 5070
rect 13132 5058 13188 5068
rect 13468 4900 13524 5068
rect 13468 4450 13524 4844
rect 13468 4398 13470 4450
rect 13522 4398 13524 4450
rect 13468 4386 13524 4398
rect 13132 4228 13188 4238
rect 13132 4116 13188 4172
rect 13132 4060 13412 4116
rect 12796 3266 12852 3276
rect 13244 3892 13300 3902
rect 13244 2548 13300 3836
rect 13356 3108 13412 4060
rect 13356 3042 13412 3052
rect 13244 2482 13300 2492
rect 13580 2884 13636 2894
rect 13132 2436 13188 2446
rect 13132 644 13188 2380
rect 13356 2324 13412 2334
rect 13356 1876 13412 2268
rect 13356 1810 13412 1820
rect 13132 578 13188 588
rect 13580 532 13636 2828
rect 13804 1874 13860 6748
rect 14140 6692 14196 6972
rect 13916 6690 14196 6692
rect 13916 6638 14142 6690
rect 14194 6638 14196 6690
rect 13916 6636 14196 6638
rect 13916 5906 13972 6636
rect 14140 6626 14196 6636
rect 13916 5854 13918 5906
rect 13970 5854 13972 5906
rect 13916 5842 13972 5854
rect 13804 1822 13806 1874
rect 13858 1822 13860 1874
rect 13804 1810 13860 1822
rect 13916 5684 13972 5694
rect 13916 980 13972 5628
rect 14252 5460 14308 8876
rect 14364 6018 14420 11340
rect 14924 11330 14980 11340
rect 14924 11172 14980 11182
rect 15148 11172 15204 11182
rect 14980 11116 15092 11172
rect 14924 11106 14980 11116
rect 14588 10836 14644 10846
rect 14588 10742 14644 10780
rect 14924 8820 14980 8830
rect 14812 8484 14868 8494
rect 14364 5966 14366 6018
rect 14418 5966 14420 6018
rect 14364 5954 14420 5966
rect 14476 8428 14812 8484
rect 14476 5908 14532 8428
rect 14812 8418 14868 8428
rect 14924 6468 14980 8764
rect 15036 8036 15092 11116
rect 15148 8372 15204 11116
rect 15260 9118 15316 13804
rect 15372 12068 15428 12078
rect 15372 11974 15428 12012
rect 15484 11618 15540 14112
rect 15820 13524 15876 13534
rect 15484 11566 15486 11618
rect 15538 11566 15540 11618
rect 15484 11554 15540 11566
rect 15708 12962 15764 12974
rect 15708 12910 15710 12962
rect 15762 12910 15764 12962
rect 15708 10612 15764 12910
rect 15820 12178 15876 13468
rect 15820 12126 15822 12178
rect 15874 12126 15876 12178
rect 15820 12114 15876 12126
rect 15932 10836 15988 14112
rect 16380 13076 16436 14112
rect 16380 13010 16436 13020
rect 16716 12404 16772 12414
rect 16828 12404 16884 14112
rect 16940 12962 16996 12974
rect 16940 12910 16942 12962
rect 16994 12910 16996 12962
rect 16940 12516 16996 12910
rect 17276 12964 17332 14112
rect 17500 13076 17556 13086
rect 17500 12982 17556 13020
rect 17276 12908 17444 12964
rect 16940 12450 16996 12460
rect 16716 12402 16884 12404
rect 16716 12350 16718 12402
rect 16770 12350 16884 12402
rect 16716 12348 16884 12350
rect 16716 12338 16772 12348
rect 17164 12292 17220 12302
rect 15932 10770 15988 10780
rect 16268 12180 16324 12190
rect 16156 10724 16212 10734
rect 15708 10556 16100 10612
rect 15596 10500 15652 10510
rect 15596 10498 15988 10500
rect 15596 10446 15598 10498
rect 15650 10446 15988 10498
rect 15596 10444 15988 10446
rect 15596 10434 15652 10444
rect 15820 9940 15876 9950
rect 15260 9062 15428 9118
rect 15148 8306 15204 8316
rect 15260 8932 15316 8942
rect 15036 7970 15092 7980
rect 14924 6402 14980 6412
rect 15260 6356 15316 8876
rect 15260 6290 15316 6300
rect 14476 5842 14532 5852
rect 14812 6188 15092 6244
rect 14812 5906 14868 6188
rect 14812 5854 14814 5906
rect 14866 5854 14868 5906
rect 14812 5842 14868 5854
rect 14924 6020 14980 6030
rect 14252 5394 14308 5404
rect 14812 5684 14868 5694
rect 14140 5124 14196 5134
rect 14364 5124 14420 5134
rect 14140 5122 14420 5124
rect 14140 5070 14142 5122
rect 14194 5070 14366 5122
rect 14418 5070 14420 5122
rect 14140 5068 14420 5070
rect 14140 5058 14196 5068
rect 14028 2884 14084 2894
rect 14028 1428 14084 2828
rect 14028 1362 14084 1372
rect 14140 2436 14196 2446
rect 13916 914 13972 924
rect 14140 868 14196 2380
rect 14252 2212 14308 2222
rect 14252 2118 14308 2156
rect 14252 1764 14308 1774
rect 14252 1428 14308 1708
rect 14252 1362 14308 1372
rect 14140 802 14196 812
rect 13580 466 13636 476
rect 14364 196 14420 5068
rect 14812 5122 14868 5628
rect 14812 5070 14814 5122
rect 14866 5070 14868 5122
rect 14812 4676 14868 5070
rect 14812 4610 14868 4620
rect 14924 4564 14980 5964
rect 15036 5908 15092 6188
rect 15372 6020 15428 9062
rect 15484 8260 15540 8270
rect 15484 6580 15540 8204
rect 15484 6514 15540 6524
rect 15596 8148 15652 8158
rect 15148 5964 15428 6020
rect 15596 6018 15652 8092
rect 15596 5966 15598 6018
rect 15650 5966 15652 6018
rect 15148 5908 15204 5964
rect 15596 5954 15652 5966
rect 15036 5852 15204 5908
rect 15036 5348 15092 5852
rect 15484 5796 15540 5806
rect 15148 5684 15204 5694
rect 15148 5590 15204 5628
rect 15148 5348 15204 5358
rect 15036 5346 15204 5348
rect 15036 5294 15150 5346
rect 15202 5294 15204 5346
rect 15036 5292 15204 5294
rect 15148 5282 15204 5292
rect 14924 4498 14980 4508
rect 15260 4564 15316 4574
rect 15260 4452 15316 4508
rect 15036 4396 15316 4452
rect 15036 4340 15092 4396
rect 14700 4284 15092 4340
rect 14700 3780 14756 4284
rect 15484 4228 15540 5740
rect 15484 4162 15540 4172
rect 15036 4116 15092 4126
rect 15092 4060 15204 4116
rect 15036 4050 15092 4060
rect 15148 3892 15204 4060
rect 15148 3826 15204 3836
rect 15820 3892 15876 9884
rect 15932 8484 15988 10444
rect 15932 8418 15988 8428
rect 16044 8260 16100 10556
rect 16156 10610 16212 10668
rect 16156 10558 16158 10610
rect 16210 10558 16212 10610
rect 16156 10546 16212 10558
rect 16044 8194 16100 8204
rect 16156 9268 16212 9278
rect 16156 6804 16212 9212
rect 16268 7700 16324 12124
rect 16940 12068 16996 12078
rect 16828 11732 16884 11742
rect 16828 11506 16884 11676
rect 16828 11454 16830 11506
rect 16882 11454 16884 11506
rect 16828 11442 16884 11454
rect 16716 10836 16772 10846
rect 16716 10742 16772 10780
rect 16268 7634 16324 7644
rect 16604 10388 16660 10398
rect 16156 6738 16212 6748
rect 16492 7028 16548 7038
rect 16380 6692 16436 6702
rect 16380 6580 16436 6636
rect 15820 3826 15876 3836
rect 15932 6524 16436 6580
rect 14700 3714 14756 3724
rect 15820 3668 15876 3678
rect 15148 3666 15876 3668
rect 15148 3614 15822 3666
rect 15874 3614 15876 3666
rect 15148 3612 15876 3614
rect 15148 3554 15204 3612
rect 15148 3502 15150 3554
rect 15202 3502 15204 3554
rect 15148 3490 15204 3502
rect 14588 2212 14644 2222
rect 14588 2118 14644 2156
rect 14476 1540 14532 1550
rect 14476 868 14532 1484
rect 14476 802 14532 812
rect 14364 130 14420 140
rect 15260 112 15316 3612
rect 15820 3602 15876 3612
rect 15596 3444 15652 3454
rect 15932 3444 15988 6524
rect 16156 5908 16212 5918
rect 15596 3442 15988 3444
rect 15596 3390 15598 3442
rect 15650 3390 15988 3442
rect 15596 3388 15988 3390
rect 16044 5124 16100 5134
rect 15596 3378 15652 3388
rect 16044 2660 16100 5068
rect 16156 4452 16212 5852
rect 16492 5348 16548 6972
rect 16604 5908 16660 10332
rect 16828 10388 16884 10398
rect 16716 10164 16772 10174
rect 16716 7588 16772 10108
rect 16828 9604 16884 10332
rect 16940 9714 16996 12012
rect 17164 10164 17220 12236
rect 17276 12180 17332 12190
rect 17276 12086 17332 12124
rect 17388 11618 17444 12908
rect 17724 12292 17780 14112
rect 17724 12226 17780 12236
rect 17948 12740 18004 12750
rect 17388 11566 17390 11618
rect 17442 11566 17444 11618
rect 17388 11554 17444 11566
rect 17724 11844 17780 11854
rect 17164 10098 17220 10108
rect 17388 10052 17444 10062
rect 17724 10052 17780 11788
rect 17948 11732 18004 12684
rect 18172 12290 18228 14112
rect 18284 13972 18340 13982
rect 18284 13074 18340 13916
rect 18396 13524 18452 13534
rect 18396 13300 18452 13468
rect 18396 13234 18452 13244
rect 18284 13022 18286 13074
rect 18338 13022 18340 13074
rect 18284 13010 18340 13022
rect 18620 13076 18676 14112
rect 18620 13010 18676 13020
rect 18956 13076 19012 13086
rect 18844 12964 18900 12974
rect 18732 12516 18788 12526
rect 18172 12238 18174 12290
rect 18226 12238 18228 12290
rect 18172 12226 18228 12238
rect 18620 12292 18676 12302
rect 17948 11666 18004 11676
rect 18508 11508 18564 11518
rect 18508 11394 18564 11452
rect 18508 11342 18510 11394
rect 18562 11342 18564 11394
rect 18508 11330 18564 11342
rect 17948 10948 18004 10958
rect 17388 10050 17780 10052
rect 17388 9998 17390 10050
rect 17442 9998 17726 10050
rect 17778 9998 17780 10050
rect 17388 9996 17780 9998
rect 17388 9986 17444 9996
rect 17724 9986 17780 9996
rect 17836 10836 17892 10846
rect 16940 9662 16942 9714
rect 16994 9662 16996 9714
rect 16940 9650 16996 9662
rect 16828 9538 16884 9548
rect 16716 7522 16772 7532
rect 16604 5842 16660 5852
rect 16492 5282 16548 5292
rect 16716 5572 16772 5582
rect 16716 4900 16772 5516
rect 16716 4834 16772 4844
rect 16156 4386 16212 4396
rect 16492 3892 16548 3902
rect 16044 2594 16100 2604
rect 16156 3556 16212 3566
rect 16156 308 16212 3500
rect 16380 3556 16436 3566
rect 16380 1316 16436 3500
rect 16492 1988 16548 3836
rect 17836 3444 17892 10780
rect 17948 10610 18004 10892
rect 18172 10948 18228 10958
rect 17948 10558 17950 10610
rect 18002 10558 18004 10610
rect 17948 10546 18004 10558
rect 18060 10724 18116 10734
rect 18060 9044 18116 10668
rect 18060 8978 18116 8988
rect 18172 7140 18228 10892
rect 18620 10722 18676 12236
rect 18620 10670 18622 10722
rect 18674 10670 18676 10722
rect 18620 10658 18676 10670
rect 18396 10052 18452 10062
rect 18284 9492 18340 9502
rect 18284 8484 18340 9436
rect 18396 8708 18452 9996
rect 18732 9940 18788 12460
rect 18844 12178 18900 12908
rect 18844 12126 18846 12178
rect 18898 12126 18900 12178
rect 18844 12114 18900 12126
rect 18732 9874 18788 9884
rect 18396 8642 18452 8652
rect 18508 9716 18564 9726
rect 18284 8428 18452 8484
rect 18172 7074 18228 7084
rect 18284 7700 18340 7710
rect 18172 6804 18228 6814
rect 17836 3378 17892 3388
rect 18060 4788 18116 4798
rect 16940 2660 16996 2670
rect 16492 1922 16548 1932
rect 16828 2548 16884 2558
rect 16828 1428 16884 2492
rect 16940 1652 16996 2604
rect 17836 2212 17892 2222
rect 18060 2212 18116 4732
rect 17836 2210 18116 2212
rect 17836 2158 17838 2210
rect 17890 2158 18062 2210
rect 18114 2158 18116 2210
rect 17836 2156 18116 2158
rect 17836 2146 17892 2156
rect 18060 2146 18116 2156
rect 17388 1876 17444 1886
rect 17388 1782 17444 1820
rect 16940 1586 16996 1596
rect 18172 1540 18228 6748
rect 18284 4676 18340 7644
rect 18396 7140 18452 8428
rect 18508 8148 18564 9660
rect 18508 8082 18564 8092
rect 18956 7812 19012 13020
rect 19068 11282 19124 14112
rect 19292 12852 19348 12862
rect 19292 12758 19348 12796
rect 19516 12290 19572 14112
rect 19964 12852 20020 14112
rect 19964 12786 20020 12796
rect 20300 12850 20356 12862
rect 20300 12798 20302 12850
rect 20354 12798 20356 12850
rect 19516 12238 19518 12290
rect 19570 12238 19572 12290
rect 19516 12226 19572 12238
rect 19740 12740 19796 12750
rect 19068 11230 19070 11282
rect 19122 11230 19124 11282
rect 19068 11218 19124 11230
rect 19292 12068 19348 12078
rect 18396 7074 18452 7084
rect 18844 7756 19012 7812
rect 19180 7812 19236 7822
rect 18284 4610 18340 4620
rect 18396 5460 18452 5470
rect 18396 3780 18452 5404
rect 18732 4452 18788 4462
rect 18620 3780 18676 3790
rect 18396 3778 18676 3780
rect 18396 3726 18398 3778
rect 18450 3726 18622 3778
rect 18674 3726 18676 3778
rect 18396 3724 18676 3726
rect 18396 3714 18452 3724
rect 18620 3714 18676 3724
rect 18732 2548 18788 4396
rect 18844 3108 18900 7756
rect 18956 7588 19012 7598
rect 18956 7494 19012 7532
rect 19180 6244 19236 7756
rect 19180 6178 19236 6188
rect 19180 3444 19236 3482
rect 19180 3378 19236 3388
rect 18844 3042 18900 3052
rect 18732 2482 18788 2492
rect 19292 2324 19348 12012
rect 19628 11284 19684 11294
rect 19628 10722 19684 11228
rect 19628 10670 19630 10722
rect 19682 10670 19684 10722
rect 19628 10658 19684 10670
rect 19740 10388 19796 12684
rect 20300 12628 20356 12798
rect 20300 12562 20356 12572
rect 20188 12292 20244 12302
rect 19964 11396 20020 11406
rect 19740 10322 19796 10332
rect 19852 11394 20020 11396
rect 19852 11342 19966 11394
rect 20018 11342 20020 11394
rect 19852 11340 20020 11342
rect 19404 9492 19460 9502
rect 19404 2884 19460 9436
rect 19852 9268 19908 11340
rect 19964 11330 20020 11340
rect 20188 11396 20244 12236
rect 20412 11620 20468 14112
rect 20636 12628 20692 12638
rect 20636 12178 20692 12572
rect 20636 12126 20638 12178
rect 20690 12126 20692 12178
rect 20636 12114 20692 12126
rect 20524 11620 20580 11630
rect 20412 11618 20580 11620
rect 20412 11566 20526 11618
rect 20578 11566 20580 11618
rect 20412 11564 20580 11566
rect 20524 11554 20580 11564
rect 20188 11330 20244 11340
rect 20412 11396 20468 11406
rect 20412 11172 20468 11340
rect 20412 11106 20468 11116
rect 20636 11172 20692 11182
rect 20636 10836 20692 11116
rect 20636 10770 20692 10780
rect 20860 10836 20916 14112
rect 20860 10770 20916 10780
rect 20972 13636 21028 13646
rect 20300 10500 20356 10510
rect 20076 10388 20132 10398
rect 20076 10294 20132 10332
rect 19852 9202 19908 9212
rect 19964 10276 20020 10286
rect 19964 9044 20020 10220
rect 20076 10164 20132 10174
rect 20076 9268 20132 10108
rect 20300 9938 20356 10444
rect 20636 10388 20692 10398
rect 20636 10294 20692 10332
rect 20300 9886 20302 9938
rect 20354 9886 20356 9938
rect 20300 9874 20356 9886
rect 20860 9826 20916 9838
rect 20860 9774 20862 9826
rect 20914 9774 20916 9826
rect 20860 9716 20916 9774
rect 20860 9650 20916 9660
rect 20076 9202 20132 9212
rect 19964 8978 20020 8988
rect 19628 8484 19684 8494
rect 19516 7476 19572 7486
rect 19516 7382 19572 7420
rect 19628 6018 19684 8428
rect 19740 8372 19796 8382
rect 19740 7586 19796 8316
rect 20524 8258 20580 8270
rect 20524 8206 20526 8258
rect 20578 8206 20580 8258
rect 19964 8146 20020 8158
rect 19964 8094 19966 8146
rect 20018 8094 20020 8146
rect 19964 7924 20020 8094
rect 20524 8148 20580 8206
rect 20860 8148 20916 8158
rect 20524 8146 20916 8148
rect 20524 8094 20862 8146
rect 20914 8094 20916 8146
rect 20524 8092 20916 8094
rect 19964 7858 20020 7868
rect 20524 7924 20580 7934
rect 19740 7534 19742 7586
rect 19794 7534 19796 7586
rect 19740 7476 19796 7534
rect 19740 7410 19796 7420
rect 20412 7700 20468 7710
rect 20412 6916 20468 7644
rect 20412 6850 20468 6860
rect 20524 6020 20580 7868
rect 20860 7476 20916 8092
rect 20860 7410 20916 7420
rect 20860 7252 20916 7262
rect 20860 6916 20916 7196
rect 20860 6850 20916 6860
rect 20636 6692 20692 6702
rect 20972 6692 21028 13580
rect 21196 13188 21252 13198
rect 21196 13094 21252 13132
rect 21196 12066 21252 12078
rect 21196 12014 21198 12066
rect 21250 12014 21252 12066
rect 21084 11732 21140 11742
rect 21084 10610 21140 11676
rect 21084 10558 21086 10610
rect 21138 10558 21140 10610
rect 21084 10546 21140 10558
rect 21196 9940 21252 12014
rect 21308 11284 21364 14112
rect 21756 13188 21812 14112
rect 21756 13122 21812 13132
rect 21756 12964 21812 12974
rect 21756 12870 21812 12908
rect 22092 12962 22148 12974
rect 22092 12910 22094 12962
rect 22146 12910 22148 12962
rect 22092 12516 22148 12910
rect 22092 12450 22148 12460
rect 22204 12404 22260 14112
rect 22652 13186 22708 14112
rect 22652 13134 22654 13186
rect 22706 13134 22708 13186
rect 22652 13122 22708 13134
rect 22428 12740 22484 12750
rect 22316 12404 22372 12414
rect 22204 12402 22372 12404
rect 22204 12350 22318 12402
rect 22370 12350 22372 12402
rect 22204 12348 22372 12350
rect 22316 12338 22372 12348
rect 21980 12180 22036 12190
rect 21980 12178 22148 12180
rect 21980 12126 21982 12178
rect 22034 12126 22148 12178
rect 21980 12124 22148 12126
rect 21980 12114 22036 12124
rect 21756 11844 21812 11854
rect 21812 11788 22036 11844
rect 21756 11778 21812 11788
rect 21980 11620 22036 11788
rect 21980 11554 22036 11564
rect 22092 11396 22148 12124
rect 21868 11340 22148 11396
rect 21756 11284 21812 11294
rect 21308 11282 21812 11284
rect 21308 11230 21758 11282
rect 21810 11230 21812 11282
rect 21308 11228 21812 11230
rect 21756 11218 21812 11228
rect 21644 10836 21700 10846
rect 21644 10742 21700 10780
rect 21868 10724 21924 11340
rect 21868 10658 21924 10668
rect 22092 11172 22148 11182
rect 21756 10388 21812 10398
rect 21756 10276 21812 10332
rect 21756 10220 22036 10276
rect 20636 6598 20692 6636
rect 20748 6636 21028 6692
rect 21084 9884 21252 9940
rect 21644 9940 21700 9950
rect 19628 5966 19630 6018
rect 19682 5966 19684 6018
rect 19628 5954 19684 5966
rect 20076 6018 20580 6020
rect 20076 5966 20526 6018
rect 20578 5966 20580 6018
rect 20076 5964 20580 5966
rect 20076 5906 20132 5964
rect 20524 5954 20580 5964
rect 20076 5854 20078 5906
rect 20130 5854 20132 5906
rect 20076 5842 20132 5854
rect 19964 5572 20020 5582
rect 19964 3780 20020 5516
rect 20412 4228 20468 4238
rect 20076 4004 20132 4014
rect 20076 3892 20132 3948
rect 20076 3836 20356 3892
rect 19964 3724 20244 3780
rect 19404 2818 19460 2828
rect 19292 2258 19348 2268
rect 20188 2324 20244 3724
rect 20188 2258 20244 2268
rect 18172 1474 18228 1484
rect 20300 1540 20356 3836
rect 20412 2884 20468 4172
rect 20748 3388 20804 6636
rect 21084 6580 21140 9884
rect 21196 9716 21252 9726
rect 21196 9622 21252 9660
rect 21532 8260 21588 8270
rect 21532 8166 21588 8204
rect 21532 7140 21588 7150
rect 21196 6690 21252 6702
rect 21196 6638 21198 6690
rect 21250 6638 21252 6690
rect 21196 6580 21252 6638
rect 21420 6580 21476 6590
rect 21196 6578 21476 6580
rect 21196 6526 21422 6578
rect 21474 6526 21476 6578
rect 21196 6524 21476 6526
rect 21084 6514 21140 6524
rect 20860 6356 20916 6366
rect 20860 4452 20916 6300
rect 21420 5908 21476 6524
rect 21532 6356 21588 7084
rect 21532 6290 21588 6300
rect 21420 5842 21476 5852
rect 20860 4386 20916 4396
rect 20972 5236 21028 5246
rect 20972 4116 21028 5180
rect 21196 4676 21252 4686
rect 20972 4050 21028 4060
rect 21084 4228 21140 4238
rect 20748 3332 20916 3388
rect 20412 2818 20468 2828
rect 20748 2100 20804 2110
rect 20748 2006 20804 2044
rect 20860 1764 20916 3332
rect 20860 1698 20916 1708
rect 20972 2212 21028 2222
rect 20300 1474 20356 1484
rect 16828 1362 16884 1372
rect 16380 1250 16436 1260
rect 20748 1316 20804 1326
rect 20636 980 20692 990
rect 20748 980 20804 1260
rect 20972 1316 21028 2156
rect 20972 1250 21028 1260
rect 21084 1092 21140 4172
rect 21196 2884 21252 4620
rect 21196 2882 21588 2884
rect 21196 2830 21198 2882
rect 21250 2830 21588 2882
rect 21196 2828 21588 2830
rect 21196 2818 21252 2828
rect 21532 2770 21588 2828
rect 21532 2718 21534 2770
rect 21586 2718 21588 2770
rect 21532 2706 21588 2718
rect 21196 2324 21252 2334
rect 21196 1988 21252 2268
rect 21308 2212 21364 2222
rect 21644 2212 21700 9884
rect 21868 9156 21924 9166
rect 21868 8372 21924 9100
rect 21868 8306 21924 8316
rect 21868 7812 21924 7822
rect 21868 7140 21924 7756
rect 21980 7252 22036 10220
rect 22092 10052 22148 11116
rect 22092 9986 22148 9996
rect 22428 9492 22484 12684
rect 23100 12404 23156 14112
rect 23100 12338 23156 12348
rect 23436 13412 23492 13422
rect 23324 12068 23380 12078
rect 23324 11974 23380 12012
rect 23436 11732 23492 13356
rect 23548 13076 23604 14112
rect 23548 13010 23604 13020
rect 23660 13188 23716 13198
rect 23660 12404 23716 13132
rect 23996 13188 24052 14112
rect 24444 13524 24500 14112
rect 23996 13122 24052 13132
rect 24220 13468 24500 13524
rect 24108 13076 24164 13086
rect 24108 12850 24164 13020
rect 24108 12798 24110 12850
rect 24162 12798 24164 12850
rect 24108 12786 24164 12798
rect 23804 12572 24068 12582
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 23804 12506 24068 12516
rect 23884 12404 23940 12414
rect 23660 12348 23828 12404
rect 23772 12180 23828 12348
rect 23884 12310 23940 12348
rect 24220 12404 24276 13468
rect 24892 13412 24948 14112
rect 24464 13356 24728 13366
rect 24892 13356 25060 13412
rect 24332 13300 24388 13310
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24464 13290 24728 13300
rect 24332 13188 24388 13244
rect 24332 13132 24500 13188
rect 24444 13076 24500 13132
rect 24556 13076 24612 13086
rect 24444 13020 24556 13076
rect 24556 13010 24612 13020
rect 24220 12338 24276 12348
rect 24892 12964 24948 12974
rect 23772 12114 23828 12124
rect 24332 11844 24388 11854
rect 23436 11676 23604 11732
rect 22764 11394 22820 11406
rect 22764 11342 22766 11394
rect 22818 11342 22820 11394
rect 22764 10052 22820 11342
rect 22764 9986 22820 9996
rect 23436 9826 23492 9838
rect 23436 9774 23438 9826
rect 23490 9774 23492 9826
rect 22428 9426 22484 9436
rect 23100 9716 23156 9726
rect 23436 9716 23492 9774
rect 23100 9714 23492 9716
rect 23100 9662 23102 9714
rect 23154 9662 23492 9714
rect 23100 9660 23492 9662
rect 22428 8930 22484 8942
rect 22428 8878 22430 8930
rect 22482 8878 22484 8930
rect 22428 8820 22484 8878
rect 22428 8754 22484 8764
rect 22988 8818 23044 8830
rect 22988 8766 22990 8818
rect 23042 8766 23044 8818
rect 22988 8372 23044 8766
rect 23100 8596 23156 9660
rect 23436 9380 23492 9390
rect 23100 8530 23156 8540
rect 23212 8818 23268 8830
rect 23212 8766 23214 8818
rect 23266 8766 23268 8818
rect 23212 8372 23268 8766
rect 23436 8596 23492 9324
rect 23548 9156 23604 11676
rect 24332 11620 24388 11788
rect 24464 11788 24728 11798
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24464 11722 24728 11732
rect 24892 11732 24948 12908
rect 25004 12516 25060 13356
rect 25340 13300 25396 14112
rect 25788 13860 25844 14112
rect 25788 13794 25844 13804
rect 25676 13636 25732 13646
rect 25676 13524 25732 13580
rect 25900 13636 25956 13646
rect 25676 13468 25844 13524
rect 25340 13244 25732 13300
rect 25452 13076 25508 13086
rect 25452 12982 25508 13020
rect 25116 12964 25172 12974
rect 25116 12962 25396 12964
rect 25116 12910 25118 12962
rect 25170 12910 25396 12962
rect 25116 12908 25396 12910
rect 25116 12898 25172 12908
rect 25004 12450 25060 12460
rect 24892 11666 24948 11676
rect 24332 11564 24500 11620
rect 23996 11282 24052 11294
rect 23996 11230 23998 11282
rect 24050 11230 24052 11282
rect 23996 11172 24052 11230
rect 23996 11106 24052 11116
rect 23804 11004 24068 11014
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 23804 10938 24068 10948
rect 24444 10948 24500 11564
rect 24556 11394 24612 11406
rect 24556 11342 24558 11394
rect 24610 11342 24612 11394
rect 24556 11172 24612 11342
rect 25116 11284 25172 11294
rect 25116 11282 25284 11284
rect 25116 11230 25118 11282
rect 25170 11230 25284 11282
rect 25116 11228 25284 11230
rect 25116 11218 25172 11228
rect 24556 11106 24612 11116
rect 24444 10882 24500 10892
rect 25004 10836 25060 10846
rect 24464 10220 24728 10230
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24464 10154 24728 10164
rect 25004 9940 25060 10780
rect 25004 9874 25060 9884
rect 25228 9828 25284 11228
rect 25340 9940 25396 12908
rect 25564 9940 25620 9950
rect 25340 9938 25620 9940
rect 25340 9886 25566 9938
rect 25618 9886 25620 9938
rect 25340 9884 25620 9886
rect 25564 9874 25620 9884
rect 25228 9762 25284 9772
rect 23996 9714 24052 9726
rect 23996 9662 23998 9714
rect 24050 9662 24052 9714
rect 23548 9090 23604 9100
rect 23660 9604 23716 9614
rect 23436 8530 23492 8540
rect 22988 8316 23268 8372
rect 22092 8258 22148 8270
rect 22092 8206 22094 8258
rect 22146 8206 22148 8258
rect 22092 8148 22148 8206
rect 22092 8082 22148 8092
rect 22316 8260 22372 8270
rect 21980 7186 22036 7196
rect 21868 7074 21924 7084
rect 21868 6132 21924 6142
rect 21868 5684 21924 6076
rect 21868 5618 21924 5628
rect 22092 5796 22148 5806
rect 22092 5572 22148 5740
rect 22092 5506 22148 5516
rect 22316 3388 22372 8204
rect 23212 8260 23268 8316
rect 23212 8194 23268 8204
rect 22428 8148 22484 8158
rect 22428 8054 22484 8092
rect 23212 8036 23268 8046
rect 23212 6692 23268 7980
rect 23660 7700 23716 9548
rect 23996 9604 24052 9662
rect 23996 9538 24052 9548
rect 23804 9436 24068 9446
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 23804 9370 24068 9380
rect 25228 8932 25284 8942
rect 24464 8652 24728 8662
rect 24332 8596 24388 8606
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24464 8586 24728 8596
rect 23804 7868 24068 7878
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 23804 7802 24068 7812
rect 24332 7700 24388 8540
rect 24556 8036 24612 8046
rect 24444 7700 24500 7710
rect 23660 7644 23828 7700
rect 24332 7644 24444 7700
rect 23436 7476 23492 7486
rect 23436 7252 23492 7420
rect 23660 7476 23716 7486
rect 23436 7196 23604 7252
rect 23436 6692 23492 6702
rect 23212 6690 23492 6692
rect 23212 6638 23214 6690
rect 23266 6638 23438 6690
rect 23490 6638 23492 6690
rect 23212 6636 23492 6638
rect 23212 6626 23268 6636
rect 23436 6626 23492 6636
rect 22764 6580 22820 6590
rect 21756 3332 21812 3342
rect 21756 2996 21812 3276
rect 22092 3332 22148 3342
rect 22316 3332 22484 3388
rect 21756 2930 21812 2940
rect 21868 3108 21924 3118
rect 21868 2436 21924 3052
rect 22092 2882 22148 3276
rect 22092 2830 22094 2882
rect 22146 2830 22148 2882
rect 22092 2818 22148 2830
rect 21868 2370 21924 2380
rect 21308 2210 21700 2212
rect 21308 2158 21310 2210
rect 21362 2158 21646 2210
rect 21698 2158 21700 2210
rect 21308 2156 21700 2158
rect 21308 2146 21364 2156
rect 21644 2146 21700 2156
rect 21532 1988 21588 1998
rect 21196 1932 21532 1988
rect 21532 1922 21588 1932
rect 21644 1764 21700 1774
rect 21084 1026 21140 1036
rect 21308 1204 21364 1214
rect 20860 980 20916 990
rect 20748 924 20860 980
rect 19964 532 20020 542
rect 16156 242 16212 252
rect 17948 420 18004 430
rect 17948 112 18004 364
rect 1148 18 1204 28
rect 1792 0 1904 112
rect 4480 0 4592 112
rect 7168 0 7280 112
rect 9856 0 9968 112
rect 12544 0 12656 112
rect 15232 0 15344 112
rect 17920 0 18032 112
rect 19964 84 20020 476
rect 20636 112 20692 924
rect 20860 914 20916 924
rect 19964 18 20020 28
rect 20608 0 20720 112
rect 21308 84 21364 1148
rect 21532 1204 21588 1214
rect 21532 308 21588 1148
rect 21644 868 21700 1708
rect 21644 802 21700 812
rect 21532 242 21588 252
rect 22428 308 22484 3332
rect 22764 3332 22820 6524
rect 23324 6468 23380 6478
rect 23324 4788 23380 6412
rect 23324 4722 23380 4732
rect 23436 5236 23492 5246
rect 23436 4676 23492 5180
rect 23548 5012 23604 7196
rect 23660 7028 23716 7420
rect 23660 6962 23716 6972
rect 23772 6804 23828 7644
rect 24444 7634 24500 7644
rect 24556 7364 24612 7980
rect 23660 6748 23828 6804
rect 23884 7308 24612 7364
rect 23660 5236 23716 6748
rect 23772 6580 23828 6590
rect 23884 6580 23940 7308
rect 25228 7140 25284 8876
rect 25340 8820 25396 8830
rect 25340 7364 25396 8764
rect 25340 7298 25396 7308
rect 24464 7084 24728 7094
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 25228 7074 25284 7084
rect 24464 7018 24728 7028
rect 25452 7028 25508 7038
rect 25116 6804 25172 6814
rect 23828 6524 23940 6580
rect 23996 6580 24052 6590
rect 25116 6580 25172 6748
rect 25116 6524 25396 6580
rect 23772 6514 23828 6524
rect 23996 6486 24052 6524
rect 24220 6356 24276 6366
rect 23804 6300 24068 6310
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 23804 6234 24068 6244
rect 24108 6020 24164 6030
rect 24220 6020 24276 6300
rect 24164 5964 24276 6020
rect 24332 6076 25060 6132
rect 24108 5954 24164 5964
rect 24332 5908 24388 6076
rect 24220 5852 24388 5908
rect 24556 5908 24612 5918
rect 24220 5572 24276 5852
rect 24556 5684 24612 5852
rect 24220 5506 24276 5516
rect 24332 5628 24612 5684
rect 24332 5460 24388 5628
rect 24892 5572 24948 5582
rect 24464 5516 24728 5526
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24464 5450 24728 5460
rect 24332 5394 24388 5404
rect 23660 5170 23716 5180
rect 23548 4946 23604 4956
rect 24892 4900 24948 5516
rect 25004 5460 25060 6076
rect 25004 5394 25060 5404
rect 24892 4834 24948 4844
rect 25228 4900 25284 4910
rect 23804 4732 24068 4742
rect 23660 4676 23716 4686
rect 23436 4620 23604 4676
rect 22764 3266 22820 3276
rect 23548 3108 23604 4620
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 23804 4666 24068 4676
rect 24220 4676 24276 4686
rect 23660 3388 23716 4620
rect 24220 4004 24276 4620
rect 25228 4228 25284 4844
rect 25228 4162 25284 4172
rect 25340 4004 25396 6524
rect 25452 4676 25508 6972
rect 25452 4610 25508 4620
rect 24220 3938 24276 3948
rect 24464 3948 24728 3958
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 25340 3938 25396 3948
rect 25564 4452 25620 4462
rect 24464 3882 24728 3892
rect 25564 3668 25620 4396
rect 25564 3602 25620 3612
rect 25676 3388 25732 13244
rect 25788 13188 25844 13468
rect 25788 13122 25844 13132
rect 25900 11620 25956 13580
rect 26236 13300 26292 14112
rect 26236 13234 26292 13244
rect 26348 13524 26404 13534
rect 25900 11554 25956 11564
rect 26012 12964 26068 12974
rect 26012 10388 26068 12908
rect 25788 10332 26068 10388
rect 25788 8260 25844 10332
rect 26348 10276 26404 13468
rect 26684 10612 26740 14112
rect 27132 13300 27188 14112
rect 27244 13300 27300 13310
rect 27132 13244 27244 13300
rect 27244 13234 27300 13244
rect 27132 12628 27188 12638
rect 27132 12292 27188 12572
rect 27132 12290 27412 12292
rect 27132 12238 27134 12290
rect 27186 12238 27412 12290
rect 27132 12236 27412 12238
rect 27132 12226 27188 12236
rect 27356 12178 27412 12236
rect 27356 12126 27358 12178
rect 27410 12126 27412 12178
rect 27356 12114 27412 12126
rect 27356 11956 27412 11966
rect 27356 11172 27412 11900
rect 27580 11956 27636 14112
rect 27804 13972 27860 13982
rect 27580 11890 27636 11900
rect 27692 13748 27748 13758
rect 27356 11106 27412 11116
rect 26796 10612 26852 10622
rect 26684 10556 26796 10612
rect 26796 10546 26852 10556
rect 26348 10210 26404 10220
rect 27020 10388 27076 10398
rect 26012 10164 26068 10174
rect 26012 9268 26068 10108
rect 26124 10052 26180 10062
rect 26460 10052 26516 10062
rect 27020 10052 27076 10332
rect 26124 10050 27076 10052
rect 26124 9998 26126 10050
rect 26178 9998 26462 10050
rect 26514 9998 27076 10050
rect 26124 9996 27076 9998
rect 26124 9986 26180 9996
rect 26460 9986 26516 9996
rect 26012 9202 26068 9212
rect 26348 8652 26628 8708
rect 25788 8194 25844 8204
rect 26236 8484 26292 8494
rect 26236 8260 26292 8428
rect 26348 8372 26404 8652
rect 26572 8596 26628 8652
rect 26796 8596 26852 8606
rect 26572 8540 26796 8596
rect 26796 8530 26852 8540
rect 26348 8306 26404 8316
rect 26236 8194 26292 8204
rect 26908 8260 26964 8270
rect 26908 8036 26964 8204
rect 27020 8036 27076 8046
rect 26908 7980 27020 8036
rect 27020 7970 27076 7980
rect 26012 7700 26068 7710
rect 25788 5236 25844 5246
rect 25788 4676 25844 5180
rect 25788 4610 25844 4620
rect 25900 4452 25956 4462
rect 23660 3332 24276 3388
rect 23548 3042 23604 3052
rect 23660 3220 23716 3230
rect 23660 2212 23716 3164
rect 23804 3164 24068 3174
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 23804 3098 24068 3108
rect 24220 3108 24276 3332
rect 25452 3332 25732 3388
rect 25788 3892 25844 3902
rect 25788 3332 25844 3836
rect 24220 3042 24276 3052
rect 25228 3220 25284 3230
rect 24892 2772 24948 2782
rect 24892 2678 24948 2716
rect 25228 2548 25284 3164
rect 25452 2772 25508 3332
rect 25788 3266 25844 3276
rect 25676 2772 25732 2782
rect 25452 2770 25732 2772
rect 25452 2718 25454 2770
rect 25506 2718 25678 2770
rect 25730 2718 25732 2770
rect 25452 2716 25732 2718
rect 25452 2706 25508 2716
rect 25676 2706 25732 2716
rect 24220 2492 25060 2548
rect 24220 2436 24276 2492
rect 24220 2370 24276 2380
rect 24464 2380 24728 2390
rect 24332 2324 24388 2334
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24464 2314 24728 2324
rect 24332 2212 24388 2268
rect 23660 2156 23940 2212
rect 24332 2156 24724 2212
rect 23772 1988 23828 1998
rect 23772 1738 23828 1932
rect 23660 1682 23828 1738
rect 23884 1764 23940 2156
rect 24556 1986 24612 1998
rect 24556 1934 24558 1986
rect 24610 1934 24612 1986
rect 24108 1876 24164 1886
rect 24556 1876 24612 1934
rect 24108 1874 24612 1876
rect 24108 1822 24110 1874
rect 24162 1822 24612 1874
rect 24108 1820 24612 1822
rect 24108 1810 24164 1820
rect 23884 1698 23940 1708
rect 23324 1652 23380 1662
rect 23660 1652 23716 1682
rect 23380 1596 23716 1652
rect 23804 1596 24068 1606
rect 23324 1586 23380 1596
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 23804 1530 24068 1540
rect 23548 1428 23604 1438
rect 24220 1428 24276 1820
rect 24668 1764 24724 2156
rect 24668 1698 24724 1708
rect 24444 1428 24500 1438
rect 23604 1372 24276 1428
rect 24332 1372 24444 1428
rect 23548 1362 23604 1372
rect 23996 1204 24052 1214
rect 24332 1204 24388 1372
rect 24444 1362 24500 1372
rect 24052 1148 24388 1204
rect 23996 1138 24052 1148
rect 23324 980 23380 990
rect 23380 924 23492 980
rect 23324 914 23380 924
rect 22428 242 22484 252
rect 23324 756 23380 766
rect 23324 112 23380 700
rect 23436 532 23492 924
rect 24332 924 24948 980
rect 24332 868 24388 924
rect 24892 868 24948 924
rect 24332 802 24388 812
rect 24464 812 24728 822
rect 23436 466 23492 476
rect 24220 756 24276 766
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24892 802 24948 812
rect 24464 746 24728 756
rect 25004 756 25060 2492
rect 25228 2482 25284 2492
rect 25116 2100 25172 2110
rect 25116 2006 25172 2044
rect 24220 420 24276 700
rect 25004 690 25060 700
rect 25228 1764 25284 1774
rect 25228 644 25284 1708
rect 25676 1428 25732 1438
rect 25676 1092 25732 1372
rect 25676 1026 25732 1036
rect 25228 578 25284 588
rect 25900 420 25956 4396
rect 24220 364 25956 420
rect 26012 112 26068 7644
rect 27468 7252 27524 7262
rect 27468 6692 27524 7196
rect 27468 6626 27524 6636
rect 26908 6580 26964 6590
rect 26964 6524 27076 6580
rect 26908 6514 26964 6524
rect 26796 6244 26852 6254
rect 26572 6188 26796 6244
rect 26572 5460 26628 6188
rect 26796 6178 26852 6188
rect 26908 5796 26964 5806
rect 26572 5394 26628 5404
rect 26796 5460 26852 5470
rect 26796 5012 26852 5404
rect 26796 4946 26852 4956
rect 26124 3332 26180 3342
rect 26124 2996 26180 3276
rect 26124 2930 26180 2940
rect 26908 2996 26964 5740
rect 27020 5012 27076 6524
rect 27020 4946 27076 4956
rect 27132 5460 27188 5470
rect 26908 2930 26964 2940
rect 27020 3556 27076 3566
rect 27020 1204 27076 3500
rect 27132 1652 27188 5404
rect 27244 4228 27300 4238
rect 27244 2884 27300 4172
rect 27244 2818 27300 2828
rect 27692 2660 27748 13692
rect 27804 11284 27860 13916
rect 27916 12628 27972 12638
rect 27916 12290 27972 12572
rect 27916 12238 27918 12290
rect 27970 12238 27972 12290
rect 27916 12226 27972 12238
rect 28028 11844 28084 14112
rect 28028 11778 28084 11788
rect 28140 12516 28196 12526
rect 27804 11218 27860 11228
rect 27916 10276 27972 10286
rect 27916 7252 27972 10220
rect 27916 7186 27972 7196
rect 28028 9828 28084 9838
rect 27916 6132 27972 6142
rect 27916 5234 27972 6076
rect 28028 6020 28084 9772
rect 28140 9156 28196 12460
rect 28252 12404 28308 12414
rect 28252 11060 28308 12348
rect 28252 10994 28308 11004
rect 28364 12292 28420 12302
rect 28140 9090 28196 9100
rect 28252 10724 28308 10734
rect 28252 8148 28308 10668
rect 28364 9828 28420 12236
rect 28476 10164 28532 14112
rect 28924 13972 28980 14112
rect 28924 13906 28980 13916
rect 28700 12852 28756 12862
rect 28588 12290 28644 12302
rect 28588 12238 28590 12290
rect 28642 12238 28644 12290
rect 28588 11732 28644 12238
rect 28588 11666 28644 11676
rect 28476 10108 28644 10164
rect 28364 9762 28420 9772
rect 28588 9156 28644 10108
rect 28700 9380 28756 12796
rect 28924 12628 28980 12638
rect 28924 10164 28980 12572
rect 29260 12628 29316 12638
rect 29260 12292 29316 12572
rect 29036 12290 29316 12292
rect 29036 12238 29262 12290
rect 29314 12238 29316 12290
rect 29036 12236 29316 12238
rect 29036 12178 29092 12236
rect 29260 12226 29316 12236
rect 29036 12126 29038 12178
rect 29090 12126 29092 12178
rect 29036 12114 29092 12126
rect 28924 10098 28980 10108
rect 29148 11172 29204 11182
rect 29148 9716 29204 11116
rect 29372 11172 29428 14112
rect 29372 11106 29428 11116
rect 29484 13412 29540 13422
rect 29148 9650 29204 9660
rect 28700 9314 28756 9324
rect 29260 9268 29316 9278
rect 28588 9100 28868 9156
rect 28252 8082 28308 8092
rect 28476 8484 28532 8494
rect 28364 6804 28420 6814
rect 28364 6244 28420 6748
rect 28364 6178 28420 6188
rect 28028 5954 28084 5964
rect 28476 5684 28532 8428
rect 28812 8260 28868 9100
rect 28812 8194 28868 8204
rect 28924 8372 28980 8382
rect 28476 5618 28532 5628
rect 28700 5908 28756 5918
rect 27916 5182 27918 5234
rect 27970 5182 27972 5234
rect 27916 5170 27972 5182
rect 28476 5236 28532 5246
rect 28476 5142 28532 5180
rect 28476 4676 28532 4686
rect 27804 4564 27860 4574
rect 27804 4228 27860 4508
rect 27804 4162 27860 4172
rect 27692 2594 27748 2604
rect 28140 2884 28196 2894
rect 28028 2100 28084 2110
rect 27244 1652 27300 1662
rect 27132 1596 27244 1652
rect 27244 1586 27300 1596
rect 27132 1204 27188 1214
rect 27020 1148 27132 1204
rect 27132 1138 27188 1148
rect 28028 1204 28084 2044
rect 28028 1138 28084 1148
rect 28140 644 28196 2828
rect 28476 2660 28532 4620
rect 28588 4228 28644 4238
rect 28588 3332 28644 4172
rect 28588 3266 28644 3276
rect 28700 3108 28756 5852
rect 28812 5348 28868 5358
rect 28812 5254 28868 5292
rect 28924 4676 28980 8316
rect 28924 4610 28980 4620
rect 29148 6692 29204 6702
rect 28588 3052 28756 3108
rect 28588 2882 28644 3052
rect 28588 2830 28590 2882
rect 28642 2830 28644 2882
rect 28588 2818 28644 2830
rect 29036 2884 29092 2894
rect 29036 2770 29092 2828
rect 29036 2718 29038 2770
rect 29090 2718 29092 2770
rect 29036 2706 29092 2718
rect 28476 2594 28532 2604
rect 28252 2548 28308 2558
rect 28252 2100 28308 2492
rect 28700 2548 28756 2558
rect 28252 2034 28308 2044
rect 28588 2212 28644 2222
rect 28588 1092 28644 2156
rect 28700 2212 28756 2492
rect 28924 2212 28980 2222
rect 28700 2210 28980 2212
rect 28700 2158 28702 2210
rect 28754 2158 28926 2210
rect 28978 2158 28980 2210
rect 28700 2156 28980 2158
rect 28700 2146 28756 2156
rect 28924 2146 28980 2156
rect 28588 1026 28644 1036
rect 28140 578 28196 588
rect 26796 532 26852 542
rect 26796 308 26852 476
rect 27020 420 27076 430
rect 28140 420 28196 430
rect 27076 364 28140 420
rect 27020 354 27076 364
rect 28140 354 28196 364
rect 29148 298 29204 6636
rect 29260 4564 29316 9212
rect 29484 7588 29540 13356
rect 29820 13412 29876 14112
rect 29820 13346 29876 13356
rect 30268 12516 30324 14112
rect 30716 14084 30772 14112
rect 30716 14018 30772 14028
rect 30268 12450 30324 12460
rect 30380 13748 30436 13758
rect 30156 12068 30212 12078
rect 30156 11732 30212 12012
rect 30156 11666 30212 11676
rect 30268 10500 30324 10510
rect 29484 7522 29540 7532
rect 29596 9604 29652 9614
rect 29260 4498 29316 4508
rect 29372 7476 29428 7486
rect 29260 2884 29316 2894
rect 29260 2790 29316 2828
rect 29372 2548 29428 7420
rect 29372 2482 29428 2492
rect 29484 5236 29540 5246
rect 29484 2098 29540 5180
rect 29484 2046 29486 2098
rect 29538 2046 29540 2098
rect 29484 2034 29540 2046
rect 29596 1540 29652 9548
rect 30268 9380 30324 10444
rect 29820 9324 30324 9380
rect 29708 7476 29764 7486
rect 29708 2772 29764 7420
rect 29820 6468 29876 9324
rect 30044 9156 30100 9166
rect 30044 8148 30100 9100
rect 30156 9044 30212 9054
rect 30156 8372 30212 8988
rect 30156 8306 30212 8316
rect 30044 8082 30100 8092
rect 30268 7250 30324 7262
rect 30268 7198 30270 7250
rect 30322 7198 30324 7250
rect 30044 7140 30100 7150
rect 30044 6580 30100 7084
rect 30044 6514 30100 6524
rect 30156 6804 30212 6814
rect 29820 6402 29876 6412
rect 30044 5796 30100 5806
rect 30044 5682 30100 5740
rect 30044 5630 30046 5682
rect 30098 5630 30100 5682
rect 29708 2706 29764 2716
rect 29820 4564 29876 4574
rect 29820 1988 29876 4508
rect 30044 3332 30100 5630
rect 30156 5124 30212 6748
rect 30156 5058 30212 5068
rect 30268 6468 30324 7198
rect 30380 6692 30436 13692
rect 31052 12068 31108 12078
rect 30716 11844 30772 11854
rect 30716 11620 30772 11788
rect 30940 11620 30996 11630
rect 30716 11618 30996 11620
rect 30716 11566 30718 11618
rect 30770 11566 30942 11618
rect 30994 11566 30996 11618
rect 30716 11564 30996 11566
rect 30716 11554 30772 11564
rect 30940 11554 30996 11564
rect 31052 10724 31108 12012
rect 31052 10658 31108 10668
rect 31164 7588 31220 14112
rect 31388 13524 31444 13534
rect 31388 10724 31444 13468
rect 31500 11620 31556 11630
rect 31500 11506 31556 11564
rect 31500 11454 31502 11506
rect 31554 11454 31556 11506
rect 31500 11442 31556 11454
rect 31388 10658 31444 10668
rect 31612 10052 31668 14112
rect 31836 13076 31892 14140
rect 32032 14112 32144 14224
rect 32480 14112 32592 14224
rect 32928 14112 33040 14224
rect 33376 14112 33488 14224
rect 33824 14112 33936 14224
rect 34272 14112 34384 14224
rect 34720 14112 34832 14224
rect 35168 14112 35280 14224
rect 35616 14112 35728 14224
rect 36064 14112 36176 14224
rect 36512 14112 36624 14224
rect 36960 14112 37072 14224
rect 37408 14112 37520 14224
rect 37856 14112 37968 14224
rect 38304 14112 38416 14224
rect 38752 14112 38864 14224
rect 39200 14112 39312 14224
rect 39648 14112 39760 14224
rect 40096 14112 40208 14224
rect 40544 14112 40656 14224
rect 40992 14112 41104 14224
rect 41440 14112 41552 14224
rect 41888 14112 42000 14224
rect 42336 14112 42448 14224
rect 42784 14112 42896 14224
rect 43232 14112 43344 14224
rect 43680 14112 43792 14224
rect 44128 14112 44240 14224
rect 44576 14112 44688 14224
rect 45024 14112 45136 14224
rect 45472 14112 45584 14224
rect 45920 14112 46032 14224
rect 46368 14112 46480 14224
rect 46816 14112 46928 14224
rect 47264 14112 47376 14224
rect 47712 14112 47824 14224
rect 48160 14112 48272 14224
rect 48608 14112 48720 14224
rect 49056 14112 49168 14224
rect 49504 14112 49616 14224
rect 49952 14112 50064 14224
rect 50400 14112 50512 14224
rect 50848 14112 50960 14224
rect 51296 14112 51408 14224
rect 51744 14112 51856 14224
rect 52192 14112 52304 14224
rect 52640 14112 52752 14224
rect 53088 14112 53200 14224
rect 53536 14112 53648 14224
rect 53984 14112 54096 14224
rect 54432 14112 54544 14224
rect 54880 14112 54992 14224
rect 55328 14112 55440 14224
rect 55776 14112 55888 14224
rect 56224 14112 56336 14224
rect 56672 14112 56784 14224
rect 31836 13010 31892 13020
rect 31836 12180 31892 12190
rect 31612 9986 31668 9996
rect 31724 11956 31780 11966
rect 31052 7532 31220 7588
rect 31500 9268 31556 9278
rect 30380 6626 30436 6636
rect 30604 7250 30660 7262
rect 30604 7198 30606 7250
rect 30658 7198 30660 7250
rect 30604 6468 30660 7198
rect 30268 6412 30660 6468
rect 30716 7252 30772 7262
rect 30268 4900 30324 6412
rect 30380 5796 30436 5806
rect 30380 5702 30436 5740
rect 30268 4834 30324 4844
rect 30716 4900 30772 7196
rect 30716 4834 30772 4844
rect 30828 7140 30884 7150
rect 30044 3266 30100 3276
rect 30492 3444 30548 3454
rect 30828 3388 30884 7084
rect 30940 5796 30996 5806
rect 30940 5702 30996 5740
rect 31052 5348 31108 7532
rect 31164 7362 31220 7374
rect 31164 7310 31166 7362
rect 31218 7310 31220 7362
rect 31164 7252 31220 7310
rect 31164 7186 31220 7196
rect 31052 5282 31108 5292
rect 31164 6468 31220 6478
rect 31052 5124 31108 5134
rect 31052 4340 31108 5068
rect 31052 4274 31108 4284
rect 29820 1922 29876 1932
rect 30380 1988 30436 1998
rect 30380 1894 30436 1932
rect 29596 1474 29652 1484
rect 30492 1428 30548 3388
rect 30716 3332 30884 3388
rect 30940 4116 30996 4126
rect 30716 2884 30772 3332
rect 30716 2818 30772 2828
rect 30604 2772 30660 2782
rect 30604 1764 30660 2716
rect 30940 2212 30996 4060
rect 31164 3444 31220 6412
rect 31500 6356 31556 9212
rect 31724 9044 31780 11900
rect 31836 10724 31892 12124
rect 32060 10836 32116 14112
rect 32060 10770 32116 10780
rect 32284 12180 32340 12190
rect 31836 10658 31892 10668
rect 32284 9604 32340 12124
rect 32508 11956 32564 14112
rect 32956 12852 33012 14112
rect 33292 13188 33348 13198
rect 32956 12786 33012 12796
rect 33180 12852 33236 12862
rect 32508 11890 32564 11900
rect 32844 11844 32900 11854
rect 32284 9538 32340 9548
rect 32508 9604 32564 9614
rect 32508 9044 32564 9548
rect 31724 8988 32004 9044
rect 31836 8820 31892 8830
rect 31612 7700 31668 7710
rect 31612 7140 31668 7644
rect 31612 7074 31668 7084
rect 31724 7588 31780 7598
rect 31500 6290 31556 6300
rect 31724 4340 31780 7532
rect 31836 6356 31892 8764
rect 31948 7140 32004 8988
rect 32508 8978 32564 8988
rect 32844 8484 32900 11788
rect 33068 11844 33124 11854
rect 32956 10612 33012 10622
rect 32956 8708 33012 10556
rect 32956 8642 33012 8652
rect 32844 8428 33012 8484
rect 31948 7074 32004 7084
rect 32844 7700 32900 7710
rect 31836 6290 31892 6300
rect 32060 6468 32116 6478
rect 31836 6020 31892 6030
rect 31836 5926 31892 5964
rect 31724 4274 31780 4284
rect 32060 3538 32116 6412
rect 32172 5908 32228 5918
rect 32172 5572 32228 5852
rect 32284 5794 32340 5806
rect 32284 5742 32286 5794
rect 32338 5742 32340 5794
rect 32284 5684 32340 5742
rect 32620 5684 32676 5694
rect 32284 5682 32676 5684
rect 32284 5630 32622 5682
rect 32674 5630 32676 5682
rect 32284 5628 32676 5630
rect 32172 5516 32564 5572
rect 32396 5124 32452 5134
rect 32396 3666 32452 5068
rect 32396 3614 32398 3666
rect 32450 3614 32452 3666
rect 32396 3602 32452 3614
rect 32060 3482 32228 3538
rect 31164 3378 31220 3388
rect 31052 3332 31108 3342
rect 31052 2884 31108 3276
rect 31052 2818 31108 2828
rect 31276 3332 32116 3388
rect 31276 2772 31332 3332
rect 31276 2706 31332 2716
rect 31948 2772 32004 2782
rect 31948 2678 32004 2716
rect 30940 2146 30996 2156
rect 30940 1986 30996 1998
rect 30940 1934 30942 1986
rect 30994 1934 30996 1986
rect 30940 1876 30996 1934
rect 31164 1876 31220 1886
rect 30940 1874 31220 1876
rect 30940 1822 31166 1874
rect 31218 1822 31220 1874
rect 30940 1820 31220 1822
rect 30604 1698 30660 1708
rect 31164 1652 31220 1820
rect 31164 1586 31220 1596
rect 30492 1362 30548 1372
rect 31836 1540 31892 1550
rect 31836 1092 31892 1484
rect 31836 1026 31892 1036
rect 32060 1092 32116 3332
rect 32060 1026 32116 1036
rect 32172 756 32228 3482
rect 32508 3388 32564 5516
rect 32172 690 32228 700
rect 32284 3332 32564 3388
rect 26796 242 26852 252
rect 28700 242 29204 298
rect 28700 112 28756 242
rect 31388 196 31444 206
rect 31388 112 31444 140
rect 32284 196 32340 3332
rect 32396 2772 32452 2782
rect 32396 2678 32452 2716
rect 32396 2436 32452 2446
rect 32396 2212 32452 2380
rect 32396 2146 32452 2156
rect 32620 1876 32676 5628
rect 32844 4452 32900 7644
rect 32956 5908 33012 8428
rect 32956 5842 33012 5852
rect 32844 4386 32900 4396
rect 32956 5572 33012 5582
rect 32956 4228 33012 5516
rect 33068 5124 33124 11788
rect 33180 9604 33236 12796
rect 33180 9538 33236 9548
rect 33292 7924 33348 13132
rect 33404 12068 33460 14112
rect 33404 12002 33460 12012
rect 33628 13076 33684 13086
rect 33404 11620 33460 11630
rect 33404 8036 33460 11564
rect 33628 11284 33684 13020
rect 33628 11218 33684 11228
rect 33740 12068 33796 12078
rect 33628 10500 33684 10510
rect 33628 9940 33684 10444
rect 33740 10276 33796 12012
rect 33852 11844 33908 14112
rect 33852 11778 33908 11788
rect 33964 13860 34020 13870
rect 33964 11620 34020 13804
rect 33740 10210 33796 10220
rect 33852 11564 34020 11620
rect 34076 13412 34132 13422
rect 33852 10052 33908 11564
rect 33964 10948 34020 10958
rect 33964 10276 34020 10892
rect 33964 10210 34020 10220
rect 33852 9996 34020 10052
rect 33628 9874 33684 9884
rect 33628 9716 33684 9726
rect 33404 7970 33460 7980
rect 33516 8148 33572 8158
rect 33292 7858 33348 7868
rect 33180 7364 33236 7374
rect 33404 7364 33460 7374
rect 33236 7308 33348 7364
rect 33180 7298 33236 7308
rect 33068 5058 33124 5068
rect 33292 5124 33348 7308
rect 33404 5236 33460 7308
rect 33516 5908 33572 8092
rect 33628 7924 33684 9660
rect 33852 9604 33908 9614
rect 33628 7858 33684 7868
rect 33740 9380 33796 9390
rect 33516 5842 33572 5852
rect 33628 7588 33684 7598
rect 33404 5170 33460 5180
rect 33292 5058 33348 5068
rect 33628 5012 33684 7532
rect 33740 6916 33796 9324
rect 33740 6850 33796 6860
rect 33740 6692 33796 6702
rect 33740 5236 33796 6636
rect 33852 5460 33908 9548
rect 33964 8596 34020 9996
rect 34076 9940 34132 13356
rect 34300 12740 34356 14112
rect 34748 13636 34804 14112
rect 34748 13570 34804 13580
rect 35084 13636 35140 13646
rect 34300 12674 34356 12684
rect 34860 12292 34916 12302
rect 34524 11956 34580 11966
rect 34188 11508 34244 11518
rect 34412 11508 34468 11518
rect 34244 11506 34468 11508
rect 34244 11454 34414 11506
rect 34466 11454 34468 11506
rect 34244 11452 34468 11454
rect 34188 11414 34244 11452
rect 34412 11442 34468 11452
rect 34076 9874 34132 9884
rect 34300 11172 34356 11182
rect 33964 8540 34244 8596
rect 33852 5394 33908 5404
rect 34076 5236 34132 5246
rect 33740 5180 34076 5236
rect 34076 5170 34132 5180
rect 33628 4946 33684 4956
rect 32844 4172 33012 4228
rect 33292 4340 33348 4350
rect 32844 2882 32900 4172
rect 33292 3778 33348 4284
rect 33292 3726 33294 3778
rect 33346 3726 33348 3778
rect 32956 3668 33012 3678
rect 33292 3668 33348 3726
rect 32956 3666 33348 3668
rect 32956 3614 32958 3666
rect 33010 3614 33348 3666
rect 32956 3612 33348 3614
rect 32956 3602 33012 3612
rect 33516 3556 33572 3566
rect 33516 3220 33572 3500
rect 33516 3154 33572 3164
rect 32844 2830 32846 2882
rect 32898 2830 32900 2882
rect 32844 2818 32900 2830
rect 34188 2436 34244 8540
rect 34300 3388 34356 11116
rect 34412 8372 34468 8382
rect 34524 8372 34580 11900
rect 34748 11956 34804 11966
rect 34748 9268 34804 11900
rect 34748 9202 34804 9212
rect 34636 8372 34692 8382
rect 34412 8370 34692 8372
rect 34412 8318 34414 8370
rect 34466 8318 34638 8370
rect 34690 8318 34692 8370
rect 34412 8316 34692 8318
rect 34412 8306 34468 8316
rect 34636 8306 34692 8316
rect 34860 8148 34916 12236
rect 34972 11396 35028 11406
rect 34972 11302 35028 11340
rect 35084 9492 35140 13580
rect 35196 10164 35252 14112
rect 35644 12180 35700 14112
rect 36092 12404 36148 14112
rect 36092 12338 36148 12348
rect 36204 12740 36260 12750
rect 35644 12114 35700 12124
rect 35980 12180 36036 12190
rect 35196 10098 35252 10108
rect 35644 11844 35700 11854
rect 34972 9436 35140 9492
rect 34972 8820 35028 9436
rect 34972 8754 35028 8764
rect 35084 9268 35140 9278
rect 34860 8082 34916 8092
rect 35084 6020 35140 9212
rect 35532 8932 35588 8942
rect 35308 8820 35364 8830
rect 35196 8372 35252 8382
rect 35196 8278 35252 8316
rect 35084 5954 35140 5964
rect 35196 7140 35252 7150
rect 34636 4900 34692 4910
rect 34300 3332 34580 3388
rect 34188 2370 34244 2380
rect 32620 1820 32900 1876
rect 32732 1204 32788 1214
rect 32396 1148 32732 1204
rect 32396 532 32452 1148
rect 32732 1138 32788 1148
rect 32396 466 32452 476
rect 32844 420 32900 1820
rect 32844 354 32900 364
rect 34076 1652 34132 1662
rect 32284 130 32340 140
rect 34076 112 34132 1596
rect 34524 756 34580 3332
rect 34636 1540 34692 4844
rect 34972 4788 35028 4798
rect 34972 4452 35028 4732
rect 34972 4386 35028 4396
rect 35196 4452 35252 7084
rect 35308 6132 35364 8764
rect 35420 7476 35476 7486
rect 35420 7140 35476 7420
rect 35420 7074 35476 7084
rect 35532 6804 35588 8876
rect 35532 6738 35588 6748
rect 35308 6066 35364 6076
rect 35196 4386 35252 4396
rect 35308 5348 35364 5358
rect 35196 4004 35252 4014
rect 34636 1474 34692 1484
rect 34748 3442 34804 3454
rect 34748 3390 34750 3442
rect 34802 3390 34804 3442
rect 34524 690 34580 700
rect 34748 308 34804 3390
rect 35196 2884 35252 3948
rect 35308 3892 35364 5292
rect 35308 3826 35364 3836
rect 35644 3780 35700 11788
rect 35868 10052 35924 10062
rect 35868 9958 35924 9996
rect 35756 9716 35812 9726
rect 35756 5572 35812 9660
rect 35868 9604 35924 9614
rect 35868 6468 35924 9548
rect 35868 6402 35924 6412
rect 35756 5506 35812 5516
rect 35868 6020 35924 6030
rect 35420 3778 35700 3780
rect 35420 3726 35646 3778
rect 35698 3726 35700 3778
rect 35420 3724 35700 3726
rect 35308 3668 35364 3678
rect 35420 3668 35476 3724
rect 35644 3714 35700 3724
rect 35756 4900 35812 4910
rect 35308 3666 35476 3668
rect 35308 3614 35310 3666
rect 35362 3614 35476 3666
rect 35308 3612 35476 3614
rect 35308 3602 35364 3612
rect 35196 2818 35252 2828
rect 35308 2996 35364 3006
rect 35308 2324 35364 2940
rect 35308 2258 35364 2268
rect 35756 2324 35812 4844
rect 35868 2660 35924 5964
rect 35980 4340 36036 12124
rect 36092 10052 36148 10062
rect 36092 9958 36148 9996
rect 36204 6916 36260 12684
rect 36316 12068 36372 12078
rect 36316 11974 36372 12012
rect 36540 8932 36596 14112
rect 36988 12718 37044 14112
rect 36652 12662 37044 12718
rect 37324 13300 37380 13310
rect 36652 11620 36708 12662
rect 36652 11554 36708 11564
rect 36764 12516 36820 12526
rect 36764 11172 36820 12460
rect 37100 12292 37156 12302
rect 36876 12236 37100 12292
rect 36876 12178 36932 12236
rect 37100 12198 37156 12236
rect 37324 12292 37380 13244
rect 37436 12404 37492 14112
rect 37436 12348 37828 12404
rect 37324 12290 37716 12292
rect 37324 12238 37326 12290
rect 37378 12238 37716 12290
rect 37324 12236 37716 12238
rect 37324 12226 37380 12236
rect 36876 12126 36878 12178
rect 36930 12126 36932 12178
rect 36876 12114 36932 12126
rect 37660 12178 37716 12236
rect 37660 12126 37662 12178
rect 37714 12126 37716 12178
rect 37660 12114 37716 12126
rect 37772 11620 37828 12348
rect 37884 11844 37940 14112
rect 38220 12066 38276 12078
rect 38220 12014 38222 12066
rect 38274 12014 38276 12066
rect 38220 11956 38276 12014
rect 38332 12068 38388 14112
rect 38780 13300 38836 14112
rect 38780 13234 38836 13244
rect 38556 12740 38612 12750
rect 38556 12516 38612 12684
rect 39228 12516 39284 14112
rect 39676 13524 39732 14112
rect 39676 13458 39732 13468
rect 38556 12460 39284 12516
rect 39340 13300 39396 13310
rect 39340 12180 39396 13244
rect 39340 12114 39396 12124
rect 38332 12002 38388 12012
rect 38220 11890 38276 11900
rect 38780 11956 38836 11966
rect 37884 11778 37940 11788
rect 37772 11564 38052 11620
rect 36764 11106 36820 11116
rect 37100 10724 37156 10734
rect 37100 10630 37156 10668
rect 37548 10388 37604 10398
rect 37884 10388 37940 10398
rect 37548 10386 37940 10388
rect 37548 10334 37550 10386
rect 37602 10334 37886 10386
rect 37938 10334 37940 10386
rect 37548 10332 37940 10334
rect 37548 10322 37604 10332
rect 37212 9940 37268 9950
rect 36652 9828 36708 9838
rect 36652 9734 36708 9772
rect 36540 8866 36596 8876
rect 37100 8484 37156 8494
rect 36204 6850 36260 6860
rect 36876 7028 36932 7038
rect 36540 5460 36596 5470
rect 36316 4788 36372 4798
rect 36204 4452 36260 4462
rect 36204 4358 36260 4396
rect 35980 4274 36036 4284
rect 36204 4004 36260 4014
rect 36204 3388 36260 3948
rect 36316 3780 36372 4732
rect 36540 4788 36596 5404
rect 36540 4722 36596 4732
rect 36540 4452 36596 4462
rect 36876 4452 36932 6972
rect 36988 6916 37044 6926
rect 36988 6580 37044 6860
rect 36988 6514 37044 6524
rect 37100 6468 37156 8428
rect 37212 6580 37268 9884
rect 37772 9492 37828 9502
rect 37772 8596 37828 9436
rect 37772 8530 37828 8540
rect 37884 7028 37940 10332
rect 37996 9492 38052 11564
rect 38332 11284 38388 11294
rect 38108 10164 38164 10174
rect 38108 9604 38164 10108
rect 38108 9538 38164 9548
rect 37996 9426 38052 9436
rect 38332 7252 38388 11228
rect 38780 8148 38836 11900
rect 39676 11284 39732 11294
rect 39340 11060 39396 11070
rect 39340 10836 39396 11004
rect 39340 10770 39396 10780
rect 39676 10612 39732 11228
rect 39676 10546 39732 10556
rect 40124 9156 40180 14112
rect 40236 12964 40292 12974
rect 40236 10948 40292 12908
rect 40236 10882 40292 10892
rect 40348 11620 40404 11630
rect 40236 10388 40292 10398
rect 40236 9828 40292 10332
rect 40236 9762 40292 9772
rect 40012 9100 40180 9156
rect 39788 8372 39844 8382
rect 39788 8278 39844 8316
rect 38780 8082 38836 8092
rect 38612 8036 38668 8046
rect 38444 7980 38612 8036
rect 38444 7476 38500 7980
rect 38612 7970 38668 7980
rect 38780 7924 38836 7934
rect 38612 7476 38668 7486
rect 38444 7410 38500 7420
rect 38556 7420 38612 7476
rect 38556 7410 38668 7420
rect 38556 7252 38612 7410
rect 38332 7196 38612 7252
rect 37884 6962 37940 6972
rect 37548 6690 37604 6702
rect 37548 6638 37550 6690
rect 37602 6638 37604 6690
rect 37212 6514 37268 6524
rect 37324 6580 37380 6590
rect 37548 6580 37604 6638
rect 38668 6690 38724 6702
rect 38668 6638 38670 6690
rect 38722 6638 38724 6690
rect 37324 6578 37604 6580
rect 37324 6526 37326 6578
rect 37378 6526 37604 6578
rect 37324 6524 37604 6526
rect 37996 6578 38052 6590
rect 37996 6526 37998 6578
rect 38050 6526 38052 6578
rect 37100 6402 37156 6412
rect 36988 6132 37044 6142
rect 36988 4676 37044 6076
rect 37324 5908 37380 6524
rect 37996 6356 38052 6526
rect 38332 6580 38388 6590
rect 38668 6580 38724 6638
rect 38332 6578 38724 6580
rect 38332 6526 38334 6578
rect 38386 6526 38724 6578
rect 38332 6524 38724 6526
rect 38332 6514 38388 6524
rect 37996 6290 38052 6300
rect 37324 5842 37380 5852
rect 36988 4610 37044 4620
rect 37548 5236 37604 5246
rect 36988 4452 37044 4462
rect 36876 4450 37044 4452
rect 36876 4398 36990 4450
rect 37042 4398 37044 4450
rect 36876 4396 37044 4398
rect 36540 4338 36596 4396
rect 36988 4386 37044 4396
rect 36540 4286 36542 4338
rect 36594 4286 36596 4338
rect 36540 4274 36596 4286
rect 36652 4340 36708 4350
rect 36540 3780 36596 3790
rect 36316 3778 36596 3780
rect 36316 3726 36318 3778
rect 36370 3726 36542 3778
rect 36594 3726 36596 3778
rect 36316 3724 36596 3726
rect 36316 3714 36372 3724
rect 36540 3714 36596 3724
rect 35868 2594 35924 2604
rect 36092 3332 36260 3388
rect 35756 2258 35812 2268
rect 36092 1764 36148 3332
rect 36652 2996 36708 4284
rect 37100 3780 37156 3790
rect 37100 3666 37156 3724
rect 37100 3614 37102 3666
rect 37154 3614 37156 3666
rect 37100 3602 37156 3614
rect 36652 2930 36708 2940
rect 36876 3444 36932 3454
rect 36876 2100 36932 3388
rect 36876 2034 36932 2044
rect 36092 1698 36148 1708
rect 37548 1652 37604 5180
rect 38220 5236 38276 5246
rect 38220 3332 38276 5180
rect 38444 3388 38500 6524
rect 38556 6244 38612 6254
rect 38556 5460 38612 6188
rect 38556 5404 38724 5460
rect 38668 4228 38724 5404
rect 38780 5124 38836 7868
rect 39004 6580 39060 6590
rect 39004 6356 39060 6524
rect 39228 6580 39284 6590
rect 39228 6486 39284 6524
rect 39004 6290 39060 6300
rect 38780 5058 38836 5068
rect 39900 4564 39956 4574
rect 39900 4450 39956 4508
rect 39900 4398 39902 4450
rect 39954 4398 39956 4450
rect 39900 4386 39956 4398
rect 38668 4162 38724 4172
rect 39004 4116 39060 4126
rect 39340 4116 39396 4126
rect 39004 4114 39396 4116
rect 39004 4062 39006 4114
rect 39058 4062 39342 4114
rect 39394 4062 39396 4114
rect 39004 4060 39396 4062
rect 39004 3444 39060 4060
rect 39340 4050 39396 4060
rect 40012 4004 40068 9100
rect 40236 8372 40292 8382
rect 40236 8278 40292 8316
rect 40348 7140 40404 11564
rect 40572 10836 40628 14112
rect 41020 13076 41076 14112
rect 41468 13188 41524 14112
rect 41468 13122 41524 13132
rect 41020 13010 41076 13020
rect 41916 11956 41972 14112
rect 40572 10770 40628 10780
rect 41020 11900 41972 11956
rect 42140 12740 42196 12750
rect 40124 7084 40404 7140
rect 40684 8146 40740 8158
rect 40684 8094 40686 8146
rect 40738 8094 40740 8146
rect 40684 7140 40740 8094
rect 40124 6916 40180 7084
rect 40684 7074 40740 7084
rect 40460 7028 40516 7038
rect 40124 6850 40180 6860
rect 40348 6916 40404 6926
rect 40236 6804 40292 6814
rect 40236 4452 40292 6748
rect 40348 4564 40404 6860
rect 40460 5348 40516 6972
rect 40460 5282 40516 5292
rect 40572 5908 40628 5918
rect 40348 4498 40404 4508
rect 40236 4386 40292 4396
rect 40012 3938 40068 3948
rect 38220 3266 38276 3276
rect 38332 3332 38500 3388
rect 38556 3388 39060 3444
rect 37660 2884 37716 2894
rect 37716 2828 37940 2884
rect 37660 2790 37716 2828
rect 37884 2770 37940 2828
rect 37884 2718 37886 2770
rect 37938 2718 37940 2770
rect 37884 2706 37940 2718
rect 38332 2660 38388 3332
rect 38332 2594 38388 2604
rect 38444 2658 38500 2670
rect 38444 2606 38446 2658
rect 38498 2606 38500 2658
rect 38444 2548 38500 2606
rect 38444 2482 38500 2492
rect 38556 1764 38612 3388
rect 40572 2772 40628 5852
rect 41020 4116 41076 11900
rect 41692 11732 41748 11742
rect 41132 10500 41188 10510
rect 41132 10406 41188 10444
rect 41356 10500 41412 10510
rect 41356 10406 41412 10444
rect 41132 10164 41188 10174
rect 41132 10050 41188 10108
rect 41132 9998 41134 10050
rect 41186 9998 41188 10050
rect 41132 9986 41188 9998
rect 41468 10164 41524 10174
rect 41468 10050 41524 10108
rect 41468 9998 41470 10050
rect 41522 9998 41524 10050
rect 41468 9986 41524 9998
rect 41244 9716 41300 9726
rect 41244 8036 41300 9660
rect 41244 7970 41300 7980
rect 41580 7700 41636 7710
rect 41580 7028 41636 7644
rect 41580 6962 41636 6972
rect 41580 6690 41636 6702
rect 41580 6638 41582 6690
rect 41634 6638 41636 6690
rect 41020 4050 41076 4060
rect 41244 6580 41300 6590
rect 40572 2706 40628 2716
rect 40348 2660 40404 2670
rect 38556 1698 38612 1708
rect 38668 2100 38724 2110
rect 37548 1586 37604 1596
rect 38668 1540 38724 2044
rect 38668 1474 38724 1484
rect 40236 1764 40292 1774
rect 39452 1316 39508 1326
rect 34748 242 34804 252
rect 36764 420 36820 430
rect 36764 112 36820 364
rect 39452 112 39508 1260
rect 40236 532 40292 1708
rect 40348 1428 40404 2604
rect 40348 1362 40404 1372
rect 41244 1428 41300 6524
rect 41356 6580 41412 6590
rect 41580 6580 41636 6638
rect 41356 6578 41636 6580
rect 41356 6526 41358 6578
rect 41410 6526 41636 6578
rect 41356 6524 41636 6526
rect 41692 6580 41748 11676
rect 42028 11282 42084 11294
rect 42028 11230 42030 11282
rect 42082 11230 42084 11282
rect 41804 11172 41860 11182
rect 41804 9940 41860 11116
rect 42028 10612 42084 11230
rect 42028 10546 42084 10556
rect 41916 10500 41972 10510
rect 41916 10406 41972 10444
rect 42140 10276 42196 12684
rect 42364 12628 42420 14112
rect 42364 12562 42420 12572
rect 42812 12292 42868 14112
rect 42812 12226 42868 12236
rect 43036 12180 43092 12190
rect 42252 10612 42308 10622
rect 42252 10518 42308 10556
rect 42700 10612 42756 10622
rect 42140 10210 42196 10220
rect 41804 9874 41860 9884
rect 42588 9826 42644 9838
rect 42588 9774 42590 9826
rect 42642 9774 42644 9826
rect 41916 9714 41972 9726
rect 41916 9662 41918 9714
rect 41970 9662 41972 9714
rect 41916 9044 41972 9662
rect 42252 9716 42308 9726
rect 42588 9716 42644 9774
rect 42252 9714 42644 9716
rect 42252 9662 42254 9714
rect 42306 9662 42644 9714
rect 42252 9660 42644 9662
rect 42252 9156 42308 9660
rect 42700 9604 42756 10556
rect 42700 9538 42756 9548
rect 42812 10498 42868 10510
rect 42812 10446 42814 10498
rect 42866 10446 42868 10498
rect 42252 9090 42308 9100
rect 42364 9492 42420 9502
rect 41916 8978 41972 8988
rect 41356 6356 41412 6524
rect 41692 6514 41748 6524
rect 41916 7700 41972 7710
rect 41356 6290 41412 6300
rect 41916 6132 41972 7644
rect 42028 6578 42084 6590
rect 42028 6526 42030 6578
rect 42082 6526 42084 6578
rect 42028 6468 42084 6526
rect 42028 6402 42084 6412
rect 41916 6066 41972 6076
rect 42140 5348 42196 5358
rect 41804 5012 41860 5022
rect 41356 4452 41412 4462
rect 41356 4358 41412 4396
rect 41692 4452 41748 4462
rect 41692 4338 41748 4396
rect 41692 4286 41694 4338
rect 41746 4286 41748 4338
rect 41692 4274 41748 4286
rect 41692 4116 41748 4126
rect 41692 3556 41748 4060
rect 41692 3490 41748 3500
rect 41804 2436 41860 4956
rect 41916 3668 41972 3678
rect 41916 3108 41972 3612
rect 41916 3052 42084 3108
rect 42028 2884 42084 3052
rect 42028 2818 42084 2828
rect 41804 2370 41860 2380
rect 41916 2212 41972 2222
rect 41972 2156 42084 2212
rect 41916 2146 41972 2156
rect 41244 1362 41300 1372
rect 42028 1092 42084 2156
rect 42028 1026 42084 1036
rect 40236 466 40292 476
rect 40460 532 40516 542
rect 40460 196 40516 476
rect 40460 130 40516 140
rect 42140 112 42196 5292
rect 42252 4226 42308 4238
rect 42252 4174 42254 4226
rect 42306 4174 42308 4226
rect 42252 3668 42308 4174
rect 42364 3892 42420 9436
rect 42812 5012 42868 10446
rect 42924 9604 42980 9614
rect 42924 8596 42980 9548
rect 42924 8530 42980 8540
rect 42812 4946 42868 4956
rect 42364 3826 42420 3836
rect 42252 3602 42308 3612
rect 42364 3444 42420 3454
rect 42252 2996 42308 3006
rect 42252 1652 42308 2940
rect 42364 2324 42420 3388
rect 42364 2258 42420 2268
rect 43036 2100 43092 12124
rect 43260 11620 43316 14112
rect 43596 13972 43652 13982
rect 43260 11554 43316 11564
rect 43484 12292 43540 12302
rect 43148 9714 43204 9726
rect 43148 9662 43150 9714
rect 43202 9662 43204 9714
rect 43148 9156 43204 9662
rect 43148 9090 43204 9100
rect 43484 6244 43540 12236
rect 43596 10836 43652 13916
rect 43708 13636 43764 14112
rect 43708 13570 43764 13580
rect 44156 13412 44212 14112
rect 44604 13860 44660 14112
rect 44604 13794 44660 13804
rect 44156 13356 44324 13412
rect 44156 13188 44212 13198
rect 43804 12572 44068 12582
rect 43860 12516 43908 12572
rect 43964 12516 44012 12572
rect 43804 12506 44068 12516
rect 44044 11508 44100 11518
rect 44044 11172 44100 11452
rect 44156 11284 44212 13132
rect 44156 11218 44212 11228
rect 44044 11106 44100 11116
rect 44268 11060 44324 13356
rect 44464 13356 44728 13366
rect 44520 13300 44568 13356
rect 44624 13300 44672 13356
rect 44464 13290 44728 13300
rect 44940 12964 44996 12974
rect 44940 12870 44996 12908
rect 44492 12292 44548 12302
rect 44548 12236 44772 12292
rect 44492 12198 44548 12236
rect 44716 12178 44772 12236
rect 44716 12126 44718 12178
rect 44770 12126 44772 12178
rect 44716 12114 44772 12126
rect 44464 11788 44728 11798
rect 44520 11732 44568 11788
rect 44624 11732 44672 11788
rect 44464 11722 44728 11732
rect 43804 11004 44068 11014
rect 43860 10948 43908 11004
rect 43964 10948 44012 11004
rect 43804 10938 44068 10948
rect 44156 11004 44324 11060
rect 43708 10836 43764 10846
rect 43596 10780 43708 10836
rect 43708 10770 43764 10780
rect 44156 9716 44212 11004
rect 44268 10276 44324 10286
rect 44268 10052 44324 10220
rect 44464 10220 44728 10230
rect 44520 10164 44568 10220
rect 44624 10164 44672 10220
rect 44464 10154 44728 10164
rect 44268 9996 44884 10052
rect 44604 9826 44660 9838
rect 44604 9774 44606 9826
rect 44658 9774 44660 9826
rect 44156 9650 44212 9660
rect 44268 9716 44324 9726
rect 44604 9716 44660 9774
rect 44268 9714 44660 9716
rect 44268 9662 44270 9714
rect 44322 9662 44660 9714
rect 44268 9660 44660 9662
rect 43804 9436 44068 9446
rect 43860 9380 43908 9436
rect 43964 9380 44012 9436
rect 43804 9370 44068 9380
rect 44044 8708 44100 8718
rect 43596 8484 43652 8494
rect 43596 8036 43652 8428
rect 44044 8372 44100 8652
rect 44044 8316 44212 8372
rect 43596 7970 43652 7980
rect 44156 7924 44212 8316
rect 44268 8148 44324 9660
rect 44464 8652 44728 8662
rect 44520 8596 44568 8652
rect 44624 8596 44672 8652
rect 44464 8586 44728 8596
rect 44268 8082 44324 8092
rect 43804 7868 44068 7878
rect 43860 7812 43908 7868
rect 43964 7812 44012 7868
rect 44156 7858 44212 7868
rect 43804 7802 44068 7812
rect 43820 7476 43876 7486
rect 43820 7252 43876 7420
rect 43820 7186 43876 7196
rect 44464 7084 44728 7094
rect 44268 7028 44324 7038
rect 44520 7028 44568 7084
rect 44624 7028 44672 7084
rect 44464 7018 44728 7028
rect 43804 6300 44068 6310
rect 43860 6244 43908 6300
rect 43964 6244 44012 6300
rect 43804 6234 44068 6244
rect 43484 6178 43540 6188
rect 43596 6132 43652 6142
rect 43596 5684 43652 6076
rect 43596 5618 43652 5628
rect 44268 5684 44324 6972
rect 44268 5618 44324 5628
rect 44464 5516 44728 5526
rect 44520 5460 44568 5516
rect 44624 5460 44672 5516
rect 44464 5450 44728 5460
rect 43596 4844 44212 4900
rect 43596 4788 43652 4844
rect 43484 4732 43652 4788
rect 44156 4788 44212 4844
rect 43804 4732 44068 4742
rect 43484 4676 43540 4732
rect 43860 4676 43908 4732
rect 43964 4676 44012 4732
rect 44156 4722 44212 4732
rect 43804 4666 44068 4676
rect 43484 4610 43540 4620
rect 43596 4564 43652 4574
rect 43484 4452 43540 4462
rect 43484 3332 43540 4396
rect 43484 3266 43540 3276
rect 43596 3108 43652 4508
rect 44464 3948 44728 3958
rect 43708 3892 43764 3902
rect 44520 3892 44568 3948
rect 44624 3892 44672 3948
rect 44464 3882 44728 3892
rect 43708 3780 43764 3836
rect 43932 3780 43988 3790
rect 43708 3778 43988 3780
rect 43708 3726 43710 3778
rect 43762 3726 43934 3778
rect 43986 3726 43988 3778
rect 43708 3724 43988 3726
rect 43708 3714 43764 3724
rect 43932 3714 43988 3724
rect 44380 3444 44436 3482
rect 44380 3378 44436 3388
rect 44828 3388 44884 9996
rect 45052 9604 45108 14112
rect 45500 13636 45556 14112
rect 45388 13580 45556 13636
rect 45724 14084 45780 14094
rect 45388 12852 45444 13580
rect 45388 12786 45444 12796
rect 45500 12964 45556 12974
rect 45276 12292 45332 12302
rect 45276 12198 45332 12236
rect 45164 9716 45220 9726
rect 45164 9622 45220 9660
rect 45052 9538 45108 9548
rect 45276 8820 45332 8830
rect 45276 7700 45332 8764
rect 45276 7634 45332 7644
rect 45388 7028 45444 7038
rect 45388 6468 45444 6972
rect 45276 6412 45444 6468
rect 45276 5236 45332 6412
rect 45276 5170 45332 5180
rect 45388 6244 45444 6254
rect 45388 4004 45444 6188
rect 45388 3938 45444 3948
rect 44828 3332 44996 3388
rect 43804 3164 44068 3174
rect 43860 3108 43908 3164
rect 43964 3108 44012 3164
rect 43804 3098 44068 3108
rect 43596 3042 43652 3052
rect 44464 2380 44728 2390
rect 44520 2324 44568 2380
rect 44624 2324 44672 2380
rect 44464 2314 44728 2324
rect 43036 2034 43092 2044
rect 44268 1876 44324 1886
rect 42252 1586 42308 1596
rect 43804 1596 44068 1606
rect 43860 1540 43908 1596
rect 43964 1540 44012 1596
rect 43804 1530 44068 1540
rect 44268 868 44324 1820
rect 44828 1092 44884 1102
rect 44268 802 44324 812
rect 44464 812 44728 822
rect 44520 756 44568 812
rect 44624 756 44672 812
rect 44464 746 44728 756
rect 44828 112 44884 1036
rect 44940 868 44996 3332
rect 45500 2996 45556 12908
rect 45612 11844 45668 11854
rect 45612 4452 45668 11788
rect 45724 11732 45780 14028
rect 45948 13188 46004 14112
rect 45948 13132 46228 13188
rect 45948 12738 46004 12750
rect 45948 12686 45950 12738
rect 46002 12686 46004 12738
rect 45948 12516 46004 12686
rect 45948 12450 46004 12460
rect 46060 12068 46116 12078
rect 46060 11974 46116 12012
rect 45724 11666 45780 11676
rect 45948 11620 46004 11630
rect 45612 4386 45668 4396
rect 45724 9044 45780 9054
rect 45724 4116 45780 8988
rect 45948 4340 46004 11564
rect 45948 4284 46116 4340
rect 45724 4060 46004 4116
rect 45500 2930 45556 2940
rect 45836 3220 45892 3230
rect 44940 802 44996 812
rect 45276 1764 45332 1774
rect 45276 308 45332 1708
rect 45836 1204 45892 3164
rect 45948 3108 46004 4060
rect 45948 3042 46004 3052
rect 45836 1138 45892 1148
rect 46060 1204 46116 4284
rect 46060 1138 46116 1148
rect 46172 420 46228 13132
rect 46396 12180 46452 14112
rect 46844 13188 46900 14112
rect 46844 13122 46900 13132
rect 46844 12964 46900 12974
rect 46844 12870 46900 12908
rect 46284 12124 46452 12180
rect 46508 12178 46564 12190
rect 46508 12126 46510 12178
rect 46562 12126 46564 12178
rect 46284 3388 46340 12124
rect 46508 12068 46564 12126
rect 46956 12180 47012 12190
rect 46956 12086 47012 12124
rect 46732 12068 46788 12078
rect 46508 12002 46564 12012
rect 46620 12012 46732 12068
rect 46620 7924 46676 12012
rect 46732 12002 46788 12012
rect 47180 11394 47236 11406
rect 47180 11342 47182 11394
rect 47234 11342 47236 11394
rect 46844 11284 46900 11294
rect 47180 11284 47236 11342
rect 46620 7858 46676 7868
rect 46732 11282 47236 11284
rect 46732 11230 46846 11282
rect 46898 11230 47236 11282
rect 46732 11228 47236 11230
rect 46732 6804 46788 11228
rect 46844 11218 46900 11228
rect 47292 11172 47348 14112
rect 47516 11620 47572 11630
rect 47740 11620 47796 14112
rect 47852 13412 47908 13422
rect 47852 12850 47908 13356
rect 48188 13188 48244 14112
rect 48188 13122 48244 13132
rect 47852 12798 47854 12850
rect 47906 12798 47908 12850
rect 47852 12786 47908 12798
rect 47964 13076 48020 13086
rect 47516 11618 47796 11620
rect 47516 11566 47518 11618
rect 47570 11566 47796 11618
rect 47516 11564 47796 11566
rect 47852 12404 47908 12414
rect 47516 11554 47572 11564
rect 47180 11116 47348 11172
rect 46956 10836 47012 10846
rect 46956 9604 47012 10780
rect 47180 9940 47236 11116
rect 47740 10612 47796 10622
rect 47180 9874 47236 9884
rect 47292 10500 47348 10510
rect 46956 9538 47012 9548
rect 46844 8820 46900 8830
rect 46844 8726 46900 8764
rect 47068 8820 47124 8830
rect 47068 8726 47124 8764
rect 46732 6738 46788 6748
rect 47068 7924 47124 7934
rect 46620 5124 46676 5134
rect 46956 5124 47012 5134
rect 46620 5122 47012 5124
rect 46620 5070 46622 5122
rect 46674 5070 46958 5122
rect 47010 5070 47012 5122
rect 46620 5068 47012 5070
rect 46284 3332 46452 3388
rect 46396 644 46452 3332
rect 46620 1316 46676 5068
rect 46956 5058 47012 5068
rect 47068 4788 47124 7868
rect 47068 4722 47124 4732
rect 46620 1250 46676 1260
rect 47292 1316 47348 10444
rect 47404 10388 47460 10398
rect 47628 10388 47684 10398
rect 47404 10386 47684 10388
rect 47404 10334 47406 10386
rect 47458 10334 47630 10386
rect 47682 10334 47684 10386
rect 47404 10332 47684 10334
rect 47404 10164 47460 10332
rect 47628 10322 47684 10332
rect 47404 10098 47460 10108
rect 47740 9156 47796 10556
rect 47404 9100 47796 9156
rect 47404 6132 47460 9100
rect 47852 9044 47908 12348
rect 47964 12402 48020 13020
rect 47964 12350 47966 12402
rect 48018 12350 48020 12402
rect 47964 12338 48020 12350
rect 48412 12962 48468 12974
rect 48412 12910 48414 12962
rect 48466 12910 48468 12962
rect 48076 12292 48132 12302
rect 47852 8978 47908 8988
rect 47964 10276 48020 10286
rect 47628 8930 47684 8942
rect 47628 8878 47630 8930
rect 47682 8878 47684 8930
rect 47404 6066 47460 6076
rect 47516 6692 47572 6702
rect 47516 5234 47572 6636
rect 47516 5182 47518 5234
rect 47570 5182 47572 5234
rect 47516 5170 47572 5182
rect 47628 2996 47684 8878
rect 47628 2930 47684 2940
rect 47740 8820 47796 8830
rect 47740 2660 47796 8764
rect 47964 7028 48020 10220
rect 48076 10164 48132 12236
rect 48412 11844 48468 12910
rect 48636 12404 48692 14112
rect 49084 13636 49140 14112
rect 49084 13570 49140 13580
rect 48972 13188 49028 13198
rect 48972 13094 49028 13132
rect 48636 12338 48692 12348
rect 49420 12404 49476 12414
rect 49420 12310 49476 12348
rect 48412 11778 48468 11788
rect 48524 12066 48580 12078
rect 48524 12014 48526 12066
rect 48578 12014 48580 12066
rect 48188 11396 48244 11406
rect 48188 11302 48244 11340
rect 48076 10098 48132 10108
rect 48188 10498 48244 10510
rect 48188 10446 48190 10498
rect 48242 10446 48244 10498
rect 48076 8372 48132 8382
rect 48188 8372 48244 10446
rect 48524 10052 48580 12014
rect 48860 12066 48916 12078
rect 48860 12014 48862 12066
rect 48914 12014 48916 12066
rect 48748 10610 48804 10622
rect 48748 10558 48750 10610
rect 48802 10558 48804 10610
rect 48524 9996 48692 10052
rect 48524 9826 48580 9838
rect 48524 9774 48526 9826
rect 48578 9774 48580 9826
rect 48300 9716 48356 9726
rect 48524 9716 48580 9774
rect 48300 9714 48580 9716
rect 48300 9662 48302 9714
rect 48354 9662 48580 9714
rect 48300 9660 48580 9662
rect 48300 9604 48356 9660
rect 48300 9538 48356 9548
rect 48412 8372 48468 8382
rect 48188 8316 48356 8372
rect 48076 8148 48132 8316
rect 48188 8148 48244 8158
rect 48076 8146 48244 8148
rect 48076 8094 48190 8146
rect 48242 8094 48244 8146
rect 48076 8092 48244 8094
rect 48188 8082 48244 8092
rect 47964 6962 48020 6972
rect 48300 5572 48356 8316
rect 48412 8278 48468 8316
rect 48300 5506 48356 5516
rect 48524 6804 48580 6814
rect 47740 2594 47796 2604
rect 48300 4228 48356 4238
rect 47292 1250 47348 1260
rect 47516 1652 47572 1662
rect 46396 578 46452 588
rect 46172 354 46228 364
rect 45276 242 45332 252
rect 47516 112 47572 1596
rect 48300 756 48356 4172
rect 48524 4228 48580 6748
rect 48636 5236 48692 9996
rect 48748 5908 48804 10558
rect 48860 7252 48916 12014
rect 49532 11620 49588 14112
rect 49980 13524 50036 14112
rect 49980 13458 50036 13468
rect 49980 12850 50036 12862
rect 49980 12798 49982 12850
rect 50034 12798 50036 12850
rect 49532 11554 49588 11564
rect 49644 11956 49700 11966
rect 49980 11956 50036 12798
rect 50428 12404 50484 14112
rect 50428 12338 50484 12348
rect 50764 12962 50820 12974
rect 50764 12910 50766 12962
rect 50818 12910 50820 12962
rect 50428 11956 50484 11966
rect 49980 11954 50484 11956
rect 49980 11902 50430 11954
rect 50482 11902 50484 11954
rect 49980 11900 50484 11902
rect 49196 11396 49252 11406
rect 49196 11282 49252 11340
rect 49196 11230 49198 11282
rect 49250 11230 49252 11282
rect 49196 11218 49252 11230
rect 49644 11284 49700 11900
rect 50316 11620 50372 11630
rect 50316 11526 50372 11564
rect 49756 11508 49812 11518
rect 49756 11414 49812 11452
rect 50428 11396 50484 11900
rect 50316 11340 50484 11396
rect 49644 11228 49812 11284
rect 49644 11060 49700 11070
rect 49644 10834 49700 11004
rect 49644 10782 49646 10834
rect 49698 10782 49700 10834
rect 49644 10770 49700 10782
rect 49420 10388 49476 10398
rect 49420 9938 49476 10332
rect 49420 9886 49422 9938
rect 49474 9886 49476 9938
rect 49420 9874 49476 9886
rect 49532 10164 49588 10174
rect 48972 9714 49028 9726
rect 48972 9662 48974 9714
rect 49026 9662 49028 9714
rect 48972 8932 49028 9662
rect 48972 8866 49028 8876
rect 49084 8820 49140 8830
rect 49308 8820 49364 8830
rect 49084 8818 49476 8820
rect 49084 8766 49086 8818
rect 49138 8766 49310 8818
rect 49362 8766 49476 8818
rect 49084 8764 49476 8766
rect 49084 8754 49140 8764
rect 49308 8754 49364 8764
rect 48972 8372 49028 8382
rect 48972 8278 49028 8316
rect 48860 7186 48916 7196
rect 48972 7028 49028 7038
rect 48972 6244 49028 6972
rect 48972 6178 49028 6188
rect 48748 5842 48804 5852
rect 48860 6132 48916 6142
rect 48636 5170 48692 5180
rect 48748 5684 48804 5694
rect 48748 4900 48804 5628
rect 48748 4834 48804 4844
rect 48524 4162 48580 4172
rect 48860 980 48916 6076
rect 48972 4116 49028 4126
rect 48972 4022 49028 4060
rect 49308 4116 49364 4126
rect 49308 4022 49364 4060
rect 48860 914 48916 924
rect 48300 690 48356 700
rect 49420 196 49476 8764
rect 49532 4788 49588 10108
rect 49532 4722 49588 4732
rect 49644 9156 49700 9166
rect 49644 2772 49700 9100
rect 49756 8372 49812 11228
rect 50204 10724 50260 10734
rect 50204 10610 50260 10668
rect 50204 10558 50206 10610
rect 50258 10558 50260 10610
rect 50204 10546 50260 10558
rect 50204 10276 50260 10286
rect 50204 9938 50260 10220
rect 50204 9886 50206 9938
rect 50258 9886 50260 9938
rect 50204 9874 50260 9886
rect 49868 8932 49924 8942
rect 49868 8838 49924 8876
rect 50204 8930 50260 8942
rect 50204 8878 50206 8930
rect 50258 8878 50260 8930
rect 49868 8372 49924 8382
rect 49756 8370 49924 8372
rect 49756 8318 49870 8370
rect 49922 8318 49924 8370
rect 49756 8316 49924 8318
rect 49868 8260 49924 8316
rect 50092 8260 50148 8270
rect 49868 8258 50148 8260
rect 49868 8206 50094 8258
rect 50146 8206 50148 8258
rect 49868 8204 50148 8206
rect 50092 8194 50148 8204
rect 50204 6580 50260 8878
rect 50316 7924 50372 11340
rect 50764 9044 50820 12910
rect 50876 11620 50932 14112
rect 51100 13636 51156 13646
rect 51100 13186 51156 13580
rect 51100 13134 51102 13186
rect 51154 13134 51156 13186
rect 51100 13122 51156 13134
rect 50988 12068 51044 12078
rect 50988 11974 51044 12012
rect 50876 11554 50932 11564
rect 51212 11844 51268 11854
rect 51212 10834 51268 11788
rect 51324 11732 51380 14112
rect 51772 13076 51828 14112
rect 52220 13188 52276 14112
rect 52220 13122 52276 13132
rect 51772 13010 51828 13020
rect 51324 11666 51380 11676
rect 52108 12962 52164 12974
rect 52108 12910 52110 12962
rect 52162 12910 52164 12962
rect 51884 11620 51940 11630
rect 51884 11526 51940 11564
rect 51212 10782 51214 10834
rect 51266 10782 51268 10834
rect 51212 10770 51268 10782
rect 51324 11394 51380 11406
rect 51324 11342 51326 11394
rect 51378 11342 51380 11394
rect 50988 10500 51044 10510
rect 50988 9938 51044 10444
rect 50988 9886 50990 9938
rect 51042 9886 51044 9938
rect 50988 9874 51044 9886
rect 51100 9716 51156 9726
rect 50764 8988 50932 9044
rect 50764 8484 50820 8494
rect 50652 8148 50708 8158
rect 50316 7858 50372 7868
rect 50428 8146 50708 8148
rect 50428 8094 50654 8146
rect 50706 8094 50708 8146
rect 50428 8092 50708 8094
rect 49868 6524 50260 6580
rect 49868 4450 49924 6524
rect 50428 4564 50484 8092
rect 50652 8082 50708 8092
rect 50764 7700 50820 8428
rect 50540 7644 50820 7700
rect 50876 7700 50932 8988
rect 50988 8372 51044 8382
rect 50988 8278 51044 8316
rect 50876 7644 51044 7700
rect 50540 7586 50596 7644
rect 50540 7534 50542 7586
rect 50594 7534 50596 7586
rect 50540 7522 50596 7534
rect 50764 7476 50820 7644
rect 50876 7476 50932 7486
rect 50764 7474 50932 7476
rect 50764 7422 50878 7474
rect 50930 7422 50932 7474
rect 50764 7420 50932 7422
rect 50876 7410 50932 7420
rect 50988 6132 51044 7644
rect 50988 6066 51044 6076
rect 51100 5908 51156 9660
rect 51212 9380 51268 9390
rect 51212 9266 51268 9324
rect 51212 9214 51214 9266
rect 51266 9214 51268 9266
rect 51212 9202 51268 9214
rect 51324 9268 51380 11342
rect 52108 10836 52164 12910
rect 52668 12964 52724 14112
rect 52892 13524 52948 13534
rect 52892 13074 52948 13468
rect 52892 13022 52894 13074
rect 52946 13022 52948 13074
rect 52892 13010 52948 13022
rect 52668 12908 52836 12964
rect 52556 12404 52612 12414
rect 52556 12310 52612 12348
rect 52220 12180 52276 12190
rect 52220 12178 52500 12180
rect 52220 12126 52222 12178
rect 52274 12126 52500 12178
rect 52220 12124 52500 12126
rect 52220 12114 52276 12124
rect 52108 10780 52388 10836
rect 52108 10612 52164 10622
rect 52108 10518 52164 10556
rect 51772 9940 51828 9950
rect 51772 9846 51828 9884
rect 51324 9202 51380 9212
rect 52220 9042 52276 9054
rect 52220 8990 52222 9042
rect 52274 8990 52276 9042
rect 51996 8148 52052 8158
rect 51996 8054 52052 8092
rect 52108 7474 52164 7486
rect 52108 7422 52110 7474
rect 52162 7422 52164 7474
rect 51436 7364 51492 7374
rect 51436 7362 51604 7364
rect 51436 7310 51438 7362
rect 51490 7310 51604 7362
rect 51436 7308 51604 7310
rect 51436 7298 51492 7308
rect 50988 5852 51156 5908
rect 50428 4498 50484 4508
rect 50540 4676 50596 4686
rect 49868 4398 49870 4450
rect 49922 4398 49924 4450
rect 49868 4386 49924 4398
rect 50540 3666 50596 4620
rect 50540 3614 50542 3666
rect 50594 3614 50596 3666
rect 50540 3602 50596 3614
rect 49756 3556 49812 3566
rect 49980 3556 50036 3566
rect 49756 3554 50036 3556
rect 49756 3502 49758 3554
rect 49810 3502 49982 3554
rect 50034 3502 50036 3554
rect 49756 3500 50036 3502
rect 49756 3332 49812 3500
rect 49980 3490 50036 3500
rect 49756 3266 49812 3276
rect 49644 2706 49700 2716
rect 50988 1202 51044 5852
rect 51100 5124 51156 5134
rect 51436 5124 51492 5134
rect 51100 5122 51492 5124
rect 51100 5070 51102 5122
rect 51154 5070 51438 5122
rect 51490 5070 51492 5122
rect 51100 5068 51492 5070
rect 51100 1652 51156 5068
rect 51436 5058 51492 5068
rect 51548 4900 51604 7308
rect 52108 6916 52164 7422
rect 52108 6850 52164 6860
rect 52220 6692 52276 8990
rect 52332 7588 52388 10780
rect 52332 7522 52388 7532
rect 52220 6626 52276 6636
rect 52108 5906 52164 5918
rect 52108 5854 52110 5906
rect 52162 5854 52164 5906
rect 51324 4844 51604 4900
rect 51884 5460 51940 5470
rect 51324 3220 51380 4844
rect 51436 4452 51492 4490
rect 51884 4452 51940 5404
rect 51996 5236 52052 5246
rect 51996 5142 52052 5180
rect 51996 4452 52052 4462
rect 51884 4450 52052 4452
rect 51884 4398 51998 4450
rect 52050 4398 52052 4450
rect 51884 4396 52052 4398
rect 51436 4386 51492 4396
rect 51996 4386 52052 4396
rect 51436 4228 51492 4238
rect 51436 3780 51492 4172
rect 51660 3780 51716 3790
rect 51436 3778 51716 3780
rect 51436 3726 51438 3778
rect 51490 3726 51662 3778
rect 51714 3726 51716 3778
rect 51436 3724 51716 3726
rect 51436 3714 51492 3724
rect 51660 3714 51716 3724
rect 51324 3154 51380 3164
rect 52108 2100 52164 5854
rect 52444 5684 52500 12124
rect 52556 11732 52612 11742
rect 52556 10834 52612 11676
rect 52780 11620 52836 12908
rect 53116 12404 53172 14112
rect 53116 12338 53172 12348
rect 53564 12292 53620 14112
rect 53900 12628 53956 12638
rect 53564 12236 53732 12292
rect 53564 12066 53620 12078
rect 53564 12014 53566 12066
rect 53618 12014 53620 12066
rect 53452 11620 53508 11630
rect 52780 11618 53508 11620
rect 52780 11566 53454 11618
rect 53506 11566 53508 11618
rect 52780 11564 53508 11566
rect 53452 11554 53508 11564
rect 52556 10782 52558 10834
rect 52610 10782 52612 10834
rect 52556 10770 52612 10782
rect 52892 11394 52948 11406
rect 52892 11342 52894 11394
rect 52946 11342 52948 11394
rect 52556 9828 52612 9838
rect 52556 9734 52612 9772
rect 52780 9044 52836 9054
rect 52668 8932 52724 8942
rect 52556 8260 52612 8270
rect 52556 8166 52612 8204
rect 52668 6690 52724 8876
rect 52668 6638 52670 6690
rect 52722 6638 52724 6690
rect 52668 6626 52724 6638
rect 52444 5618 52500 5628
rect 52332 5460 52388 5470
rect 52332 5346 52388 5404
rect 52332 5294 52334 5346
rect 52386 5294 52388 5346
rect 52332 5282 52388 5294
rect 52668 5012 52724 5022
rect 52780 5012 52836 8988
rect 52892 7028 52948 11342
rect 53564 10724 53620 12014
rect 53452 10668 53620 10724
rect 53004 9268 53060 9278
rect 53004 9174 53060 9212
rect 53340 8372 53396 8382
rect 53340 8278 53396 8316
rect 53452 8036 53508 10668
rect 53564 10498 53620 10510
rect 53564 10446 53566 10498
rect 53618 10446 53620 10498
rect 53564 10388 53620 10446
rect 53564 10322 53620 10332
rect 53564 9716 53620 9726
rect 53676 9716 53732 12236
rect 53564 9714 53732 9716
rect 53564 9662 53566 9714
rect 53618 9662 53732 9714
rect 53564 9660 53732 9662
rect 53788 11956 53844 11966
rect 53564 9650 53620 9660
rect 53788 9604 53844 11900
rect 53676 9548 53844 9604
rect 53564 8930 53620 8942
rect 53564 8878 53566 8930
rect 53618 8878 53620 8930
rect 53564 8708 53620 8878
rect 53564 8642 53620 8652
rect 53676 8484 53732 9548
rect 53452 7970 53508 7980
rect 53564 8428 53732 8484
rect 53004 7812 53060 7822
rect 53004 7698 53060 7756
rect 53004 7646 53006 7698
rect 53058 7646 53060 7698
rect 53004 7634 53060 7646
rect 52892 6962 52948 6972
rect 53564 6578 53620 8428
rect 53900 8148 53956 12572
rect 54012 9268 54068 14112
rect 54236 13524 54292 13534
rect 54124 13076 54180 13086
rect 54124 12402 54180 13020
rect 54124 12350 54126 12402
rect 54178 12350 54180 12402
rect 54124 12338 54180 12350
rect 54236 10276 54292 13468
rect 54348 12962 54404 12974
rect 54348 12910 54350 12962
rect 54402 12910 54404 12962
rect 54348 11172 54404 12910
rect 54460 11844 54516 14112
rect 54908 13412 54964 14112
rect 54908 13346 54964 13356
rect 55356 13300 55412 14112
rect 55356 13234 55412 13244
rect 54908 13188 54964 13198
rect 54908 13094 54964 13132
rect 55468 13076 55524 13086
rect 55132 12068 55188 12078
rect 54460 11778 54516 11788
rect 54796 12066 55188 12068
rect 54796 12014 55134 12066
rect 55186 12014 55188 12066
rect 54796 12012 55188 12014
rect 54348 11106 54404 11116
rect 54460 11282 54516 11294
rect 54460 11230 54462 11282
rect 54514 11230 54516 11282
rect 54236 10210 54292 10220
rect 54012 9202 54068 9212
rect 54236 9826 54292 9838
rect 54236 9774 54238 9826
rect 54290 9774 54292 9826
rect 53900 8082 53956 8092
rect 54124 8258 54180 8270
rect 54124 8206 54126 8258
rect 54178 8206 54180 8258
rect 53564 6526 53566 6578
rect 53618 6526 53620 6578
rect 53564 6514 53620 6526
rect 53676 7474 53732 7486
rect 53676 7422 53678 7474
rect 53730 7422 53732 7474
rect 53004 6132 53060 6142
rect 53004 6038 53060 6076
rect 53564 6020 53620 6030
rect 53564 5906 53620 5964
rect 53564 5854 53566 5906
rect 53618 5854 53620 5906
rect 53564 5842 53620 5854
rect 52892 5236 52948 5246
rect 53676 5236 53732 7422
rect 54124 7476 54180 8206
rect 54124 7410 54180 7420
rect 54124 6690 54180 6702
rect 54124 6638 54126 6690
rect 54178 6638 54180 6690
rect 54124 5796 54180 6638
rect 54124 5730 54180 5740
rect 52892 5142 52948 5180
rect 53564 5180 53732 5236
rect 54124 5572 54180 5582
rect 54124 5234 54180 5516
rect 54124 5182 54126 5234
rect 54178 5182 54180 5234
rect 53228 5124 53284 5134
rect 53116 5068 53228 5124
rect 52892 5012 52948 5022
rect 52780 4956 52892 5012
rect 52444 4900 52500 4910
rect 52220 4452 52276 4462
rect 52220 4338 52276 4396
rect 52220 4286 52222 4338
rect 52274 4286 52276 4338
rect 52220 4274 52276 4286
rect 52220 3442 52276 3454
rect 52220 3390 52222 3442
rect 52274 3390 52276 3442
rect 52220 3388 52276 3390
rect 52220 3332 52388 3388
rect 52220 3108 52276 3118
rect 52220 2770 52276 3052
rect 52220 2718 52222 2770
rect 52274 2718 52276 2770
rect 52220 2706 52276 2718
rect 52108 2034 52164 2044
rect 52220 2436 52276 2446
rect 51660 1986 51716 1998
rect 51660 1934 51662 1986
rect 51714 1934 51716 1986
rect 51436 1876 51492 1886
rect 51660 1876 51716 1934
rect 51436 1874 51716 1876
rect 51436 1822 51438 1874
rect 51490 1822 51716 1874
rect 51436 1820 51716 1822
rect 52108 1876 52164 1886
rect 51436 1764 51492 1820
rect 52108 1782 52164 1820
rect 51436 1698 51492 1708
rect 51100 1586 51156 1596
rect 50988 1150 50990 1202
rect 51042 1150 51044 1202
rect 50988 1138 51044 1150
rect 51996 1314 52052 1326
rect 51996 1262 51998 1314
rect 52050 1262 52052 1314
rect 51996 980 52052 1262
rect 51996 914 52052 924
rect 52220 532 52276 2380
rect 52332 1204 52388 3332
rect 52444 2212 52500 4844
rect 52668 4450 52724 4956
rect 52892 4946 52948 4956
rect 52668 4398 52670 4450
rect 52722 4398 52724 4450
rect 52668 4386 52724 4398
rect 53116 4450 53172 5068
rect 53228 5030 53284 5068
rect 53564 4676 53620 5180
rect 54124 5170 54180 5182
rect 53676 5012 53732 5022
rect 53676 4918 53732 4956
rect 53564 4610 53620 4620
rect 53116 4398 53118 4450
rect 53170 4398 53172 4450
rect 53116 4386 53172 4398
rect 54236 4340 54292 9774
rect 54348 8930 54404 8942
rect 54348 8878 54350 8930
rect 54402 8878 54404 8930
rect 54348 8596 54404 8878
rect 54348 8530 54404 8540
rect 54236 4274 54292 4284
rect 53564 4226 53620 4238
rect 53564 4174 53566 4226
rect 53618 4174 53620 4226
rect 52556 3892 52612 3902
rect 52556 3666 52612 3836
rect 52556 3614 52558 3666
rect 52610 3614 52612 3666
rect 52556 3602 52612 3614
rect 53564 3668 53620 4174
rect 53564 3602 53620 3612
rect 54348 3556 54404 3566
rect 54460 3556 54516 11230
rect 54572 10722 54628 10734
rect 54572 10670 54574 10722
rect 54626 10670 54628 10722
rect 54572 10164 54628 10670
rect 54572 10098 54628 10108
rect 54572 7586 54628 7598
rect 54572 7534 54574 7586
rect 54626 7534 54628 7586
rect 54572 7252 54628 7534
rect 54572 7186 54628 7196
rect 54572 6018 54628 6030
rect 54572 5966 54574 6018
rect 54626 5966 54628 6018
rect 54572 5908 54628 5966
rect 54572 5842 54628 5852
rect 54796 4900 54852 12012
rect 55132 12002 55188 12012
rect 54908 11394 54964 11406
rect 54908 11342 54910 11394
rect 54962 11342 54964 11394
rect 54908 11284 54964 11342
rect 55244 11284 55300 11294
rect 54908 11282 55300 11284
rect 54908 11230 55246 11282
rect 55298 11230 55300 11282
rect 54908 11228 55300 11230
rect 54908 6468 54964 11228
rect 55244 11218 55300 11228
rect 55468 11060 55524 13020
rect 55692 12404 55748 12414
rect 55692 12310 55748 12348
rect 55804 11956 55860 14112
rect 55804 11890 55860 11900
rect 55916 13972 55972 13982
rect 55468 10994 55524 11004
rect 55692 11284 55748 11294
rect 55580 10836 55636 10846
rect 55132 10500 55188 10510
rect 54908 6402 54964 6412
rect 55020 10498 55188 10500
rect 55020 10446 55134 10498
rect 55186 10446 55188 10498
rect 55020 10444 55188 10446
rect 55020 5236 55076 10444
rect 55132 10434 55188 10444
rect 55468 10388 55524 10398
rect 55132 9602 55188 9614
rect 55132 9550 55134 9602
rect 55186 9550 55188 9602
rect 55132 9492 55188 9550
rect 55132 9426 55188 9436
rect 55132 8930 55188 8942
rect 55132 8878 55134 8930
rect 55186 8878 55188 8930
rect 55132 8820 55188 8878
rect 55132 8754 55188 8764
rect 55468 8372 55524 10332
rect 55580 9940 55636 10780
rect 55580 9874 55636 9884
rect 55132 8316 55524 8372
rect 55692 8372 55748 11228
rect 55916 9380 55972 13916
rect 56252 12516 56308 14112
rect 56252 12450 56308 12460
rect 55916 9314 55972 9324
rect 56028 12180 56084 12190
rect 55132 8146 55188 8316
rect 55692 8306 55748 8316
rect 55916 8930 55972 8942
rect 55916 8878 55918 8930
rect 55970 8878 55972 8930
rect 55132 8094 55134 8146
rect 55186 8094 55188 8146
rect 55132 8082 55188 8094
rect 55916 8148 55972 8878
rect 55916 8082 55972 8092
rect 56028 7812 56084 12124
rect 56140 10722 56196 10734
rect 56140 10670 56142 10722
rect 56194 10670 56196 10722
rect 56140 9044 56196 10670
rect 56140 8978 56196 8988
rect 56028 7746 56084 7756
rect 56140 7700 56196 7710
rect 56140 7606 56196 7644
rect 55132 7364 55188 7374
rect 55132 7270 55188 7308
rect 56140 6804 56196 6814
rect 55132 6466 55188 6478
rect 55132 6414 55134 6466
rect 55186 6414 55188 6466
rect 55132 6356 55188 6414
rect 55132 6290 55188 6300
rect 56140 6130 56196 6748
rect 56140 6078 56142 6130
rect 56194 6078 56196 6130
rect 56140 6066 56196 6078
rect 56700 6132 56756 14112
rect 56700 6066 56756 6076
rect 55020 5170 55076 5180
rect 55244 5906 55300 5918
rect 55244 5854 55246 5906
rect 55298 5854 55300 5906
rect 54908 5124 54964 5134
rect 54908 5030 54964 5068
rect 54796 4834 54852 4844
rect 54572 4564 54628 4574
rect 54572 4470 54628 4508
rect 55132 4226 55188 4238
rect 55132 4174 55134 4226
rect 55186 4174 55188 4226
rect 55132 3780 55188 4174
rect 55132 3714 55188 3724
rect 54908 3668 54964 3678
rect 54908 3574 54964 3612
rect 54348 3554 54516 3556
rect 54348 3502 54350 3554
rect 54402 3502 54516 3554
rect 54348 3500 54516 3502
rect 54348 3490 54404 3500
rect 53564 3444 53620 3482
rect 53564 3378 53620 3388
rect 54572 3220 54628 3230
rect 52444 2146 52500 2156
rect 52556 2996 52612 3006
rect 52556 2098 52612 2940
rect 54572 2994 54628 3164
rect 54572 2942 54574 2994
rect 54626 2942 54628 2994
rect 54572 2930 54628 2942
rect 53564 2772 53620 2782
rect 53564 2678 53620 2716
rect 52780 2660 52836 2670
rect 52780 2566 52836 2604
rect 55132 2658 55188 2670
rect 55132 2606 55134 2658
rect 55186 2606 55188 2658
rect 52556 2046 52558 2098
rect 52610 2046 52612 2098
rect 52556 2034 52612 2046
rect 54124 2548 54180 2558
rect 54124 2098 54180 2492
rect 54124 2046 54126 2098
rect 54178 2046 54180 2098
rect 54124 2034 54180 2046
rect 54908 2324 54964 2334
rect 54908 2098 54964 2268
rect 54908 2046 54910 2098
rect 54962 2046 54964 2098
rect 54908 2034 54964 2046
rect 53564 1876 53620 1886
rect 53564 1782 53620 1820
rect 55132 1540 55188 2606
rect 55244 2436 55300 5854
rect 56140 5460 56196 5470
rect 55244 2370 55300 2380
rect 55356 4788 55412 4798
rect 55132 1474 55188 1484
rect 53564 1428 53620 1438
rect 53564 1334 53620 1372
rect 52332 1138 52388 1148
rect 52556 1316 52612 1326
rect 52556 1202 52612 1260
rect 52556 1150 52558 1202
rect 52610 1150 52612 1202
rect 52556 1138 52612 1150
rect 55356 1202 55412 4732
rect 56140 4562 56196 5404
rect 56140 4510 56142 4562
rect 56194 4510 56196 4562
rect 56140 4498 56196 4510
rect 56140 4116 56196 4126
rect 56140 2994 56196 4060
rect 56140 2942 56142 2994
rect 56194 2942 56196 2994
rect 56140 2930 56196 2942
rect 56812 3444 56868 3454
rect 56140 2772 56196 2782
rect 56140 1426 56196 2716
rect 56140 1374 56142 1426
rect 56194 1374 56196 1426
rect 56140 1362 56196 1374
rect 56476 2660 56532 2670
rect 55356 1150 55358 1202
rect 55410 1150 55412 1202
rect 55356 1138 55412 1150
rect 52220 466 52276 476
rect 52892 868 52948 878
rect 49420 130 49476 140
rect 50204 196 50260 206
rect 50204 112 50260 140
rect 52892 112 52948 812
rect 55580 756 55636 766
rect 55580 112 55636 700
rect 21308 18 21364 28
rect 23296 0 23408 112
rect 25984 0 26096 112
rect 28672 0 28784 112
rect 31360 0 31472 112
rect 34048 0 34160 112
rect 36736 0 36848 112
rect 39424 0 39536 112
rect 42112 0 42224 112
rect 44800 0 44912 112
rect 47488 0 47600 112
rect 50176 0 50288 112
rect 52864 0 52976 112
rect 55552 0 55664 112
rect 56476 84 56532 2604
rect 56812 532 56868 3388
rect 56812 466 56868 476
rect 56476 18 56532 28
<< via2 >>
rect 31836 14140 31892 14196
rect 364 13020 420 13076
rect 252 12012 308 12068
rect 924 12572 980 12628
rect 700 9660 756 9716
rect 812 10780 868 10836
rect 1036 12124 1092 12180
rect 1148 11788 1204 11844
rect 1484 13916 1540 13972
rect 2156 13356 2212 13412
rect 2268 12402 2324 12404
rect 2268 12350 2270 12402
rect 2270 12350 2322 12402
rect 2322 12350 2324 12402
rect 2268 12348 2324 12350
rect 1036 10780 1092 10836
rect 924 9772 980 9828
rect 1036 10332 1092 10388
rect 812 9436 868 9492
rect 364 8316 420 8372
rect 140 5404 196 5460
rect 588 6860 644 6916
rect 1036 5180 1092 5236
rect 1596 10332 1652 10388
rect 1484 9660 1540 9716
rect 1484 8092 1540 8148
rect 2044 11506 2100 11508
rect 2044 11454 2046 11506
rect 2046 11454 2098 11506
rect 2098 11454 2100 11506
rect 2044 11452 2100 11454
rect 2268 11788 2324 11844
rect 1820 9436 1876 9492
rect 2380 10668 2436 10724
rect 2380 8988 2436 9044
rect 2492 10556 2548 10612
rect 1820 7532 1876 7588
rect 2044 8876 2100 8932
rect 1708 5068 1764 5124
rect 1820 5180 1876 5236
rect 1484 4844 1540 4900
rect 1596 4956 1652 5012
rect 588 3612 644 3668
rect 1148 3724 1204 3780
rect 1036 3388 1092 3444
rect 1036 924 1092 980
rect 1260 924 1316 980
rect 1596 2940 1652 2996
rect 1708 4284 1764 4340
rect 2604 8540 2660 8596
rect 2940 12124 2996 12180
rect 3164 13916 3220 13972
rect 2268 8258 2324 8260
rect 2268 8206 2270 8258
rect 2270 8206 2322 8258
rect 2322 8206 2324 8258
rect 2268 8204 2324 8206
rect 2940 10444 2996 10500
rect 3052 9826 3108 9828
rect 3052 9774 3054 9826
rect 3054 9774 3106 9826
rect 3106 9774 3108 9826
rect 3052 9772 3108 9774
rect 3388 12348 3444 12404
rect 3612 13468 3668 13524
rect 3724 13186 3780 13188
rect 3724 13134 3726 13186
rect 3726 13134 3778 13186
rect 3778 13134 3780 13186
rect 3724 13132 3780 13134
rect 4732 13468 4788 13524
rect 4284 13356 4340 13412
rect 4464 13354 4520 13356
rect 4464 13302 4466 13354
rect 4466 13302 4518 13354
rect 4518 13302 4520 13354
rect 4464 13300 4520 13302
rect 4568 13354 4624 13356
rect 4568 13302 4570 13354
rect 4570 13302 4622 13354
rect 4622 13302 4624 13354
rect 4568 13300 4624 13302
rect 4672 13354 4728 13356
rect 4672 13302 4674 13354
rect 4674 13302 4726 13354
rect 4726 13302 4728 13354
rect 4672 13300 4728 13302
rect 4284 12962 4340 12964
rect 4284 12910 4286 12962
rect 4286 12910 4338 12962
rect 4338 12910 4340 12962
rect 4284 12908 4340 12910
rect 4956 12908 5012 12964
rect 3804 12570 3860 12572
rect 3804 12518 3806 12570
rect 3806 12518 3858 12570
rect 3858 12518 3860 12570
rect 3804 12516 3860 12518
rect 3908 12570 3964 12572
rect 3908 12518 3910 12570
rect 3910 12518 3962 12570
rect 3962 12518 3964 12570
rect 3908 12516 3964 12518
rect 4012 12570 4068 12572
rect 4012 12518 4014 12570
rect 4014 12518 4066 12570
rect 4066 12518 4068 12570
rect 4012 12516 4068 12518
rect 3388 12124 3444 12180
rect 3612 11116 3668 11172
rect 3804 11002 3860 11004
rect 3804 10950 3806 11002
rect 3806 10950 3858 11002
rect 3858 10950 3860 11002
rect 3804 10948 3860 10950
rect 3908 11002 3964 11004
rect 3908 10950 3910 11002
rect 3910 10950 3962 11002
rect 3962 10950 3964 11002
rect 3908 10948 3964 10950
rect 4012 11002 4068 11004
rect 4012 10950 4014 11002
rect 4014 10950 4066 11002
rect 4066 10950 4068 11002
rect 4012 10948 4068 10950
rect 4464 11786 4520 11788
rect 4464 11734 4466 11786
rect 4466 11734 4518 11786
rect 4518 11734 4520 11786
rect 4464 11732 4520 11734
rect 4568 11786 4624 11788
rect 4568 11734 4570 11786
rect 4570 11734 4622 11786
rect 4622 11734 4624 11786
rect 4568 11732 4624 11734
rect 4672 11786 4728 11788
rect 4672 11734 4674 11786
rect 4674 11734 4726 11786
rect 4726 11734 4728 11786
rect 4672 11732 4728 11734
rect 4620 11618 4676 11620
rect 4620 11566 4622 11618
rect 4622 11566 4674 11618
rect 4674 11566 4676 11618
rect 4620 11564 4676 11566
rect 4464 10218 4520 10220
rect 4464 10166 4466 10218
rect 4466 10166 4518 10218
rect 4518 10166 4520 10218
rect 4464 10164 4520 10166
rect 4568 10218 4624 10220
rect 4568 10166 4570 10218
rect 4570 10166 4622 10218
rect 4622 10166 4624 10218
rect 4568 10164 4624 10166
rect 4672 10218 4728 10220
rect 4672 10166 4674 10218
rect 4674 10166 4726 10218
rect 4726 10166 4728 10218
rect 4672 10164 4728 10166
rect 3804 9434 3860 9436
rect 3804 9382 3806 9434
rect 3806 9382 3858 9434
rect 3858 9382 3860 9434
rect 3804 9380 3860 9382
rect 3908 9434 3964 9436
rect 3908 9382 3910 9434
rect 3910 9382 3962 9434
rect 3962 9382 3964 9434
rect 3908 9380 3964 9382
rect 4012 9434 4068 9436
rect 4012 9382 4014 9434
rect 4014 9382 4066 9434
rect 4066 9382 4068 9434
rect 4172 9436 4228 9492
rect 4012 9380 4068 9382
rect 3388 8652 3444 8708
rect 2828 6076 2884 6132
rect 2940 7644 2996 7700
rect 2716 5628 2772 5684
rect 2604 5346 2660 5348
rect 2604 5294 2606 5346
rect 2606 5294 2658 5346
rect 2658 5294 2660 5346
rect 2604 5292 2660 5294
rect 2492 2492 2548 2548
rect 2940 5346 2996 5348
rect 2940 5294 2942 5346
rect 2942 5294 2994 5346
rect 2994 5294 2996 5346
rect 2940 5292 2996 5294
rect 4464 8650 4520 8652
rect 4464 8598 4466 8650
rect 4466 8598 4518 8650
rect 4518 8598 4520 8650
rect 4464 8596 4520 8598
rect 4568 8650 4624 8652
rect 4568 8598 4570 8650
rect 4570 8598 4622 8650
rect 4622 8598 4624 8650
rect 4568 8596 4624 8598
rect 4672 8650 4728 8652
rect 4672 8598 4674 8650
rect 4674 8598 4726 8650
rect 4726 8598 4728 8650
rect 4672 8596 4728 8598
rect 3724 8316 3780 8372
rect 3804 7866 3860 7868
rect 3804 7814 3806 7866
rect 3806 7814 3858 7866
rect 3858 7814 3860 7866
rect 3804 7812 3860 7814
rect 3908 7866 3964 7868
rect 3908 7814 3910 7866
rect 3910 7814 3962 7866
rect 3962 7814 3964 7866
rect 3908 7812 3964 7814
rect 4012 7866 4068 7868
rect 4012 7814 4014 7866
rect 4014 7814 4066 7866
rect 4066 7814 4068 7866
rect 4012 7812 4068 7814
rect 3500 7308 3556 7364
rect 4464 7082 4520 7084
rect 4464 7030 4466 7082
rect 4466 7030 4518 7082
rect 4518 7030 4520 7082
rect 4464 7028 4520 7030
rect 4568 7082 4624 7084
rect 4568 7030 4570 7082
rect 4570 7030 4622 7082
rect 4622 7030 4624 7082
rect 4568 7028 4624 7030
rect 4672 7082 4728 7084
rect 4672 7030 4674 7082
rect 4674 7030 4726 7082
rect 4726 7030 4728 7082
rect 4672 7028 4728 7030
rect 3612 6578 3668 6580
rect 3612 6526 3614 6578
rect 3614 6526 3666 6578
rect 3666 6526 3668 6578
rect 3612 6524 3668 6526
rect 3804 6298 3860 6300
rect 3804 6246 3806 6298
rect 3806 6246 3858 6298
rect 3858 6246 3860 6298
rect 3804 6244 3860 6246
rect 3908 6298 3964 6300
rect 3908 6246 3910 6298
rect 3910 6246 3962 6298
rect 3962 6246 3964 6298
rect 3908 6244 3964 6246
rect 4012 6298 4068 6300
rect 4012 6246 4014 6298
rect 4014 6246 4066 6298
rect 4066 6246 4068 6298
rect 4012 6244 4068 6246
rect 3804 4730 3860 4732
rect 3804 4678 3806 4730
rect 3806 4678 3858 4730
rect 3858 4678 3860 4730
rect 3804 4676 3860 4678
rect 3908 4730 3964 4732
rect 3908 4678 3910 4730
rect 3910 4678 3962 4730
rect 3962 4678 3964 4730
rect 3908 4676 3964 4678
rect 4012 4730 4068 4732
rect 4012 4678 4014 4730
rect 4014 4678 4066 4730
rect 4066 4678 4068 4730
rect 4012 4676 4068 4678
rect 4464 5514 4520 5516
rect 4464 5462 4466 5514
rect 4466 5462 4518 5514
rect 4518 5462 4520 5514
rect 4464 5460 4520 5462
rect 4568 5514 4624 5516
rect 4568 5462 4570 5514
rect 4570 5462 4622 5514
rect 4622 5462 4624 5514
rect 4568 5460 4624 5462
rect 4672 5514 4728 5516
rect 4672 5462 4674 5514
rect 4674 5462 4726 5514
rect 4726 5462 4728 5514
rect 4672 5460 4728 5462
rect 5628 13132 5684 13188
rect 5964 13244 6020 13300
rect 5964 12796 6020 12852
rect 5068 11564 5124 11620
rect 4956 9212 5012 9268
rect 4956 6860 5012 6916
rect 4956 5180 5012 5236
rect 4172 4620 4228 4676
rect 4396 4844 4452 4900
rect 3388 4396 3444 4452
rect 3276 4060 3332 4116
rect 5740 9996 5796 10052
rect 5292 8540 5348 8596
rect 5180 5516 5236 5572
rect 5068 4956 5124 5012
rect 4844 4844 4900 4900
rect 4844 4450 4900 4452
rect 4844 4398 4846 4450
rect 4846 4398 4898 4450
rect 4898 4398 4900 4450
rect 4844 4396 4900 4398
rect 5180 4396 5236 4452
rect 4396 4060 4452 4116
rect 4464 3946 4520 3948
rect 4464 3894 4466 3946
rect 4466 3894 4518 3946
rect 4518 3894 4520 3946
rect 4464 3892 4520 3894
rect 4568 3946 4624 3948
rect 4568 3894 4570 3946
rect 4570 3894 4622 3946
rect 4622 3894 4624 3946
rect 4568 3892 4624 3894
rect 4672 3946 4728 3948
rect 4672 3894 4674 3946
rect 4674 3894 4726 3946
rect 4726 3894 4728 3946
rect 4672 3892 4728 3894
rect 3804 3162 3860 3164
rect 3804 3110 3806 3162
rect 3806 3110 3858 3162
rect 3858 3110 3860 3162
rect 3804 3108 3860 3110
rect 3908 3162 3964 3164
rect 3908 3110 3910 3162
rect 3910 3110 3962 3162
rect 3962 3110 3964 3162
rect 3908 3108 3964 3110
rect 4012 3162 4068 3164
rect 4012 3110 4014 3162
rect 4014 3110 4066 3162
rect 4066 3110 4068 3162
rect 4012 3108 4068 3110
rect 3276 2828 3332 2884
rect 3836 2658 3892 2660
rect 3836 2606 3838 2658
rect 3838 2606 3890 2658
rect 3890 2606 3892 2658
rect 3836 2604 3892 2606
rect 4396 2546 4452 2548
rect 4396 2494 4398 2546
rect 4398 2494 4450 2546
rect 4450 2494 4452 2546
rect 4396 2492 4452 2494
rect 4956 2546 5012 2548
rect 4956 2494 4958 2546
rect 4958 2494 5010 2546
rect 5010 2494 5012 2546
rect 4956 2492 5012 2494
rect 4464 2378 4520 2380
rect 4464 2326 4466 2378
rect 4466 2326 4518 2378
rect 4518 2326 4520 2378
rect 4464 2324 4520 2326
rect 4568 2378 4624 2380
rect 4568 2326 4570 2378
rect 4570 2326 4622 2378
rect 4622 2326 4624 2378
rect 4568 2324 4624 2326
rect 4672 2378 4728 2380
rect 4672 2326 4674 2378
rect 4674 2326 4726 2378
rect 4726 2326 4728 2378
rect 4672 2324 4728 2326
rect 3388 1986 3444 1988
rect 3388 1934 3390 1986
rect 3390 1934 3442 1986
rect 3442 1934 3444 1986
rect 3388 1932 3444 1934
rect 3724 1986 3780 1988
rect 3724 1934 3726 1986
rect 3726 1934 3778 1986
rect 3778 1934 3780 1986
rect 3724 1932 3780 1934
rect 2716 1820 2772 1876
rect 3804 1594 3860 1596
rect 3804 1542 3806 1594
rect 3806 1542 3858 1594
rect 3858 1542 3860 1594
rect 3804 1540 3860 1542
rect 3908 1594 3964 1596
rect 3908 1542 3910 1594
rect 3910 1542 3962 1594
rect 3962 1542 3964 1594
rect 3908 1540 3964 1542
rect 4012 1594 4068 1596
rect 4012 1542 4014 1594
rect 4014 1542 4066 1594
rect 4066 1542 4068 1594
rect 5068 1596 5124 1652
rect 4012 1540 4068 1542
rect 2492 1260 2548 1316
rect 2828 1314 2884 1316
rect 2828 1262 2830 1314
rect 2830 1262 2882 1314
rect 2882 1262 2884 1314
rect 2828 1260 2884 1262
rect 1820 1036 1876 1092
rect 4464 810 4520 812
rect 4464 758 4466 810
rect 4466 758 4518 810
rect 4518 758 4520 810
rect 4464 756 4520 758
rect 4568 810 4624 812
rect 4568 758 4570 810
rect 4570 758 4622 810
rect 4622 758 4624 810
rect 4568 756 4624 758
rect 4672 810 4728 812
rect 4672 758 4674 810
rect 4674 758 4726 810
rect 4726 758 4728 810
rect 4672 756 4728 758
rect 1596 476 1652 532
rect 4508 588 4564 644
rect 1372 140 1428 196
rect 1820 140 1876 196
rect 5740 4226 5796 4228
rect 5740 4174 5742 4226
rect 5742 4174 5794 4226
rect 5794 4174 5796 4226
rect 5740 4172 5796 4174
rect 5964 11788 6020 11844
rect 6636 13692 6692 13748
rect 6524 12962 6580 12964
rect 6524 12910 6526 12962
rect 6526 12910 6578 12962
rect 6578 12910 6580 12962
rect 6524 12908 6580 12910
rect 7420 13244 7476 13300
rect 7532 13186 7588 13188
rect 7532 13134 7534 13186
rect 7534 13134 7586 13186
rect 7586 13134 7588 13186
rect 7532 13132 7588 13134
rect 6972 12402 7028 12404
rect 6972 12350 6974 12402
rect 6974 12350 7026 12402
rect 7026 12350 7028 12402
rect 6972 12348 7028 12350
rect 6524 11788 6580 11844
rect 6636 12012 6692 12068
rect 8092 13074 8148 13076
rect 8092 13022 8094 13074
rect 8094 13022 8146 13074
rect 8146 13022 8148 13074
rect 8092 13020 8148 13022
rect 8652 12460 8708 12516
rect 7868 12348 7924 12404
rect 8540 12402 8596 12404
rect 8540 12350 8542 12402
rect 8542 12350 8594 12402
rect 8594 12350 8596 12402
rect 8540 12348 8596 12350
rect 7532 12178 7588 12180
rect 7532 12126 7534 12178
rect 7534 12126 7586 12178
rect 7586 12126 7588 12178
rect 7532 12124 7588 12126
rect 6188 9548 6244 9604
rect 6076 9154 6132 9156
rect 6076 9102 6078 9154
rect 6078 9102 6130 9154
rect 6130 9102 6132 9154
rect 6076 9100 6132 9102
rect 6524 8818 6580 8820
rect 6524 8766 6526 8818
rect 6526 8766 6578 8818
rect 6578 8766 6580 8818
rect 6524 8764 6580 8766
rect 6412 8316 6468 8372
rect 6188 7420 6244 7476
rect 5964 7308 6020 7364
rect 6300 6748 6356 6804
rect 6188 6524 6244 6580
rect 6076 5740 6132 5796
rect 6300 6188 6356 6244
rect 6300 4284 6356 4340
rect 6188 4060 6244 4116
rect 6076 3724 6132 3780
rect 5852 1148 5908 1204
rect 6524 6860 6580 6916
rect 6524 4508 6580 4564
rect 6748 8818 6804 8820
rect 6748 8766 6750 8818
rect 6750 8766 6802 8818
rect 6802 8766 6804 8818
rect 6748 8764 6804 8766
rect 7532 10332 7588 10388
rect 6860 6412 6916 6468
rect 6972 10220 7028 10276
rect 7196 9660 7252 9716
rect 6860 5852 6916 5908
rect 6860 4508 6916 4564
rect 6636 3388 6692 3444
rect 6748 4396 6804 4452
rect 6748 3276 6804 3332
rect 7532 9212 7588 9268
rect 7980 9324 8036 9380
rect 7868 8764 7924 8820
rect 7644 4284 7700 4340
rect 7420 2604 7476 2660
rect 6524 1874 6580 1876
rect 6524 1822 6526 1874
rect 6526 1822 6578 1874
rect 6578 1822 6580 1874
rect 6524 1820 6580 1822
rect 6412 812 6468 868
rect 7196 1596 7252 1652
rect 5404 588 5460 644
rect 7420 1260 7476 1316
rect 8540 10668 8596 10724
rect 8092 8652 8148 8708
rect 7980 5740 8036 5796
rect 8316 9436 8372 9492
rect 8316 8204 8372 8260
rect 8428 7420 8484 7476
rect 8988 14028 9044 14084
rect 9212 13132 9268 13188
rect 9212 12908 9268 12964
rect 8988 11900 9044 11956
rect 8652 9100 8708 9156
rect 8876 8764 8932 8820
rect 9436 12908 9492 12964
rect 9212 11452 9268 11508
rect 9324 12572 9380 12628
rect 9212 10444 9268 10500
rect 9324 10108 9380 10164
rect 9548 12684 9604 12740
rect 9772 13186 9828 13188
rect 9772 13134 9774 13186
rect 9774 13134 9826 13186
rect 9826 13134 9828 13186
rect 9772 13132 9828 13134
rect 10332 13244 10388 13300
rect 9660 12348 9716 12404
rect 10780 13468 10836 13524
rect 10668 12348 10724 12404
rect 10108 11900 10164 11956
rect 10108 11340 10164 11396
rect 10332 11340 10388 11396
rect 11340 13356 11396 13412
rect 11452 13132 11508 13188
rect 12236 13804 12292 13860
rect 11564 13020 11620 13076
rect 11116 12236 11172 12292
rect 10332 10220 10388 10276
rect 9996 10108 10052 10164
rect 10332 9826 10388 9828
rect 10332 9774 10334 9826
rect 10334 9774 10386 9826
rect 10386 9774 10388 9826
rect 10332 9772 10388 9774
rect 10108 9212 10164 9268
rect 9548 8764 9604 8820
rect 10108 8876 10164 8932
rect 9212 7980 9268 8036
rect 9100 7868 9156 7924
rect 9660 7586 9716 7588
rect 9660 7534 9662 7586
rect 9662 7534 9714 7586
rect 9714 7534 9716 7586
rect 9660 7532 9716 7534
rect 9660 6860 9716 6916
rect 9324 6748 9380 6804
rect 8764 6636 8820 6692
rect 8764 6076 8820 6132
rect 9212 6300 9268 6356
rect 9212 5964 9268 6020
rect 8428 3836 8484 3892
rect 8652 4508 8708 4564
rect 8092 2044 8148 2100
rect 9212 5404 9268 5460
rect 9212 4732 9268 4788
rect 8876 3724 8932 3780
rect 8764 3276 8820 3332
rect 10332 8930 10388 8932
rect 10332 8878 10334 8930
rect 10334 8878 10386 8930
rect 10386 8878 10388 8930
rect 10332 8876 10388 8878
rect 10108 8092 10164 8148
rect 11116 10220 11172 10276
rect 10668 7756 10724 7812
rect 9996 7532 10052 7588
rect 10556 7362 10612 7364
rect 10556 7310 10558 7362
rect 10558 7310 10610 7362
rect 10610 7310 10612 7362
rect 10556 7308 10612 7310
rect 9772 6300 9828 6356
rect 9660 5740 9716 5796
rect 10220 6076 10276 6132
rect 9884 5180 9940 5236
rect 9884 4508 9940 4564
rect 10108 5180 10164 5236
rect 10220 4172 10276 4228
rect 10668 4172 10724 4228
rect 9996 3948 10052 4004
rect 9324 2828 9380 2884
rect 8652 1372 8708 1428
rect 7868 588 7924 644
rect 10668 3388 10724 3444
rect 10556 1596 10612 1652
rect 10892 8092 10948 8148
rect 11564 10498 11620 10500
rect 11564 10446 11566 10498
rect 11566 10446 11618 10498
rect 11618 10446 11620 10498
rect 11564 10444 11620 10446
rect 11900 9660 11956 9716
rect 12012 12124 12068 12180
rect 11676 8764 11732 8820
rect 11788 9100 11844 9156
rect 11452 8092 11508 8148
rect 12684 13132 12740 13188
rect 13244 13356 13300 13412
rect 13692 13074 13748 13076
rect 13692 13022 13694 13074
rect 13694 13022 13746 13074
rect 13746 13022 13748 13074
rect 13692 13020 13748 13022
rect 12908 12962 12964 12964
rect 12908 12910 12910 12962
rect 12910 12910 12962 12962
rect 12962 12910 12964 12962
rect 12908 12908 12964 12910
rect 13580 12460 13636 12516
rect 13356 12236 13412 12292
rect 13468 12124 13524 12180
rect 13804 12348 13860 12404
rect 13692 12290 13748 12292
rect 13692 12238 13694 12290
rect 13694 12238 13746 12290
rect 13746 12238 13748 12290
rect 13692 12236 13748 12238
rect 13580 11676 13636 11732
rect 13692 12012 13748 12068
rect 12572 10668 12628 10724
rect 12460 10108 12516 10164
rect 12460 9884 12516 9940
rect 12012 7756 12068 7812
rect 11900 7420 11956 7476
rect 11900 6076 11956 6132
rect 11676 5852 11732 5908
rect 11788 5964 11844 6020
rect 11228 5628 11284 5684
rect 13244 10220 13300 10276
rect 13132 9548 13188 9604
rect 13020 8876 13076 8932
rect 12796 7308 12852 7364
rect 11788 3948 11844 4004
rect 12572 4620 12628 4676
rect 11004 3442 11060 3444
rect 11004 3390 11006 3442
rect 11006 3390 11058 3442
rect 11058 3390 11060 3442
rect 11004 3388 11060 3390
rect 10892 2716 10948 2772
rect 11116 3276 11172 3332
rect 11116 1484 11172 1540
rect 10780 364 10836 420
rect 13244 8876 13300 8932
rect 13468 8316 13524 8372
rect 13468 7532 13524 7588
rect 13132 7308 13188 7364
rect 13020 7196 13076 7252
rect 12908 7084 12964 7140
rect 12908 6076 12964 6132
rect 14028 12348 14084 12404
rect 14028 12124 14084 12180
rect 14588 13020 14644 13076
rect 14924 13074 14980 13076
rect 14924 13022 14926 13074
rect 14926 13022 14978 13074
rect 14978 13022 14980 13074
rect 14924 13020 14980 13022
rect 14140 10780 14196 10836
rect 14252 12460 14308 12516
rect 13804 10332 13860 10388
rect 13692 10220 13748 10276
rect 14028 10108 14084 10164
rect 15260 13804 15316 13860
rect 15148 13692 15204 13748
rect 15148 11788 15204 11844
rect 14252 9996 14308 10052
rect 14252 8876 14308 8932
rect 13692 8652 13748 8708
rect 13692 6972 13748 7028
rect 14140 6972 14196 7028
rect 13804 6748 13860 6804
rect 13580 5292 13636 5348
rect 13468 4844 13524 4900
rect 13132 4172 13188 4228
rect 12796 3276 12852 3332
rect 13244 3836 13300 3892
rect 13356 3052 13412 3108
rect 13244 2492 13300 2548
rect 13580 2828 13636 2884
rect 13132 2380 13188 2436
rect 13356 2268 13412 2324
rect 13356 1820 13412 1876
rect 13132 588 13188 644
rect 13916 5628 13972 5684
rect 14924 11116 14980 11172
rect 14588 10834 14644 10836
rect 14588 10782 14590 10834
rect 14590 10782 14642 10834
rect 14642 10782 14644 10834
rect 14588 10780 14644 10782
rect 14924 8764 14980 8820
rect 14812 8428 14868 8484
rect 15148 11116 15204 11172
rect 15372 12066 15428 12068
rect 15372 12014 15374 12066
rect 15374 12014 15426 12066
rect 15426 12014 15428 12066
rect 15372 12012 15428 12014
rect 15820 13468 15876 13524
rect 16380 13020 16436 13076
rect 17500 13074 17556 13076
rect 17500 13022 17502 13074
rect 17502 13022 17554 13074
rect 17554 13022 17556 13074
rect 17500 13020 17556 13022
rect 16940 12460 16996 12516
rect 17164 12236 17220 12292
rect 15932 10780 15988 10836
rect 16268 12124 16324 12180
rect 16156 10668 16212 10724
rect 15820 9884 15876 9940
rect 15148 8316 15204 8372
rect 15260 8876 15316 8932
rect 15036 7980 15092 8036
rect 14924 6412 14980 6468
rect 15260 6300 15316 6356
rect 14476 5852 14532 5908
rect 14924 5964 14980 6020
rect 14252 5404 14308 5460
rect 14812 5628 14868 5684
rect 14028 2828 14084 2884
rect 14028 1372 14084 1428
rect 14140 2380 14196 2436
rect 13916 924 13972 980
rect 14252 2210 14308 2212
rect 14252 2158 14254 2210
rect 14254 2158 14306 2210
rect 14306 2158 14308 2210
rect 14252 2156 14308 2158
rect 14252 1708 14308 1764
rect 14252 1372 14308 1428
rect 14140 812 14196 868
rect 13580 476 13636 532
rect 14812 4620 14868 4676
rect 15484 8204 15540 8260
rect 15484 6524 15540 6580
rect 15596 8092 15652 8148
rect 15484 5740 15540 5796
rect 15148 5682 15204 5684
rect 15148 5630 15150 5682
rect 15150 5630 15202 5682
rect 15202 5630 15204 5682
rect 15148 5628 15204 5630
rect 14924 4508 14980 4564
rect 15260 4508 15316 4564
rect 15484 4172 15540 4228
rect 15036 4060 15092 4116
rect 15148 3836 15204 3892
rect 15932 8428 15988 8484
rect 16044 8204 16100 8260
rect 16156 9212 16212 9268
rect 16940 12012 16996 12068
rect 16828 11676 16884 11732
rect 16716 10834 16772 10836
rect 16716 10782 16718 10834
rect 16718 10782 16770 10834
rect 16770 10782 16772 10834
rect 16716 10780 16772 10782
rect 16268 7644 16324 7700
rect 16604 10332 16660 10388
rect 16156 6748 16212 6804
rect 16492 6972 16548 7028
rect 16380 6636 16436 6692
rect 15820 3836 15876 3892
rect 14700 3724 14756 3780
rect 14588 2210 14644 2212
rect 14588 2158 14590 2210
rect 14590 2158 14642 2210
rect 14642 2158 14644 2210
rect 14588 2156 14644 2158
rect 14476 1484 14532 1540
rect 14476 812 14532 868
rect 14364 140 14420 196
rect 16156 5852 16212 5908
rect 16044 5068 16100 5124
rect 16828 10332 16884 10388
rect 16716 10108 16772 10164
rect 17276 12178 17332 12180
rect 17276 12126 17278 12178
rect 17278 12126 17330 12178
rect 17330 12126 17332 12178
rect 17276 12124 17332 12126
rect 17724 12236 17780 12292
rect 17948 12684 18004 12740
rect 17724 11788 17780 11844
rect 17164 10108 17220 10164
rect 18284 13916 18340 13972
rect 18396 13468 18452 13524
rect 18396 13244 18452 13300
rect 18620 13020 18676 13076
rect 18956 13020 19012 13076
rect 18844 12908 18900 12964
rect 18732 12460 18788 12516
rect 18620 12236 18676 12292
rect 17948 11676 18004 11732
rect 18508 11452 18564 11508
rect 17948 10892 18004 10948
rect 17836 10780 17892 10836
rect 16828 9548 16884 9604
rect 16716 7532 16772 7588
rect 16604 5852 16660 5908
rect 16492 5292 16548 5348
rect 16716 5516 16772 5572
rect 16716 4844 16772 4900
rect 16156 4396 16212 4452
rect 16492 3836 16548 3892
rect 16044 2604 16100 2660
rect 16156 3500 16212 3556
rect 16380 3500 16436 3556
rect 18172 10892 18228 10948
rect 18060 10668 18116 10724
rect 18060 8988 18116 9044
rect 18396 9996 18452 10052
rect 18284 9436 18340 9492
rect 18732 9884 18788 9940
rect 18396 8652 18452 8708
rect 18508 9660 18564 9716
rect 18172 7084 18228 7140
rect 18284 7644 18340 7700
rect 18172 6748 18228 6804
rect 17836 3388 17892 3444
rect 18060 4732 18116 4788
rect 16940 2604 16996 2660
rect 16492 1932 16548 1988
rect 16828 2492 16884 2548
rect 17388 1874 17444 1876
rect 17388 1822 17390 1874
rect 17390 1822 17442 1874
rect 17442 1822 17444 1874
rect 17388 1820 17444 1822
rect 16940 1596 16996 1652
rect 18508 8092 18564 8148
rect 19292 12850 19348 12852
rect 19292 12798 19294 12850
rect 19294 12798 19346 12850
rect 19346 12798 19348 12850
rect 19292 12796 19348 12798
rect 19964 12796 20020 12852
rect 19740 12684 19796 12740
rect 19292 12012 19348 12068
rect 18396 7084 18452 7140
rect 19180 7756 19236 7812
rect 18284 4620 18340 4676
rect 18396 5404 18452 5460
rect 18732 4396 18788 4452
rect 18956 7586 19012 7588
rect 18956 7534 18958 7586
rect 18958 7534 19010 7586
rect 19010 7534 19012 7586
rect 18956 7532 19012 7534
rect 19180 6188 19236 6244
rect 19180 3442 19236 3444
rect 19180 3390 19182 3442
rect 19182 3390 19234 3442
rect 19234 3390 19236 3442
rect 19180 3388 19236 3390
rect 18844 3052 18900 3108
rect 18732 2492 18788 2548
rect 19628 11228 19684 11284
rect 20300 12572 20356 12628
rect 20188 12236 20244 12292
rect 19740 10332 19796 10388
rect 19404 9436 19460 9492
rect 20636 12572 20692 12628
rect 20188 11340 20244 11396
rect 20412 11340 20468 11396
rect 20412 11116 20468 11172
rect 20636 11116 20692 11172
rect 20636 10780 20692 10836
rect 20860 10780 20916 10836
rect 20972 13580 21028 13636
rect 20300 10444 20356 10500
rect 20076 10386 20132 10388
rect 20076 10334 20078 10386
rect 20078 10334 20130 10386
rect 20130 10334 20132 10386
rect 20076 10332 20132 10334
rect 19852 9212 19908 9268
rect 19964 10220 20020 10276
rect 20076 10108 20132 10164
rect 20636 10386 20692 10388
rect 20636 10334 20638 10386
rect 20638 10334 20690 10386
rect 20690 10334 20692 10386
rect 20636 10332 20692 10334
rect 20860 9660 20916 9716
rect 20076 9212 20132 9268
rect 19964 8988 20020 9044
rect 19628 8428 19684 8484
rect 19516 7474 19572 7476
rect 19516 7422 19518 7474
rect 19518 7422 19570 7474
rect 19570 7422 19572 7474
rect 19516 7420 19572 7422
rect 19740 8316 19796 8372
rect 19964 7868 20020 7924
rect 20524 7868 20580 7924
rect 19740 7420 19796 7476
rect 20412 7644 20468 7700
rect 20412 6860 20468 6916
rect 20860 7420 20916 7476
rect 20860 7196 20916 7252
rect 20860 6860 20916 6916
rect 21196 13186 21252 13188
rect 21196 13134 21198 13186
rect 21198 13134 21250 13186
rect 21250 13134 21252 13186
rect 21196 13132 21252 13134
rect 21084 11676 21140 11732
rect 21756 13132 21812 13188
rect 21756 12962 21812 12964
rect 21756 12910 21758 12962
rect 21758 12910 21810 12962
rect 21810 12910 21812 12962
rect 21756 12908 21812 12910
rect 22092 12460 22148 12516
rect 22428 12684 22484 12740
rect 21756 11788 21812 11844
rect 21980 11564 22036 11620
rect 21644 10834 21700 10836
rect 21644 10782 21646 10834
rect 21646 10782 21698 10834
rect 21698 10782 21700 10834
rect 21644 10780 21700 10782
rect 21868 10668 21924 10724
rect 22092 11116 22148 11172
rect 21756 10332 21812 10388
rect 20636 6690 20692 6692
rect 20636 6638 20638 6690
rect 20638 6638 20690 6690
rect 20690 6638 20692 6690
rect 20636 6636 20692 6638
rect 21644 9884 21700 9940
rect 19964 5516 20020 5572
rect 20412 4172 20468 4228
rect 20076 3948 20132 4004
rect 19404 2828 19460 2884
rect 19292 2268 19348 2324
rect 20188 2268 20244 2324
rect 18172 1484 18228 1540
rect 21196 9714 21252 9716
rect 21196 9662 21198 9714
rect 21198 9662 21250 9714
rect 21250 9662 21252 9714
rect 21196 9660 21252 9662
rect 21532 8258 21588 8260
rect 21532 8206 21534 8258
rect 21534 8206 21586 8258
rect 21586 8206 21588 8258
rect 21532 8204 21588 8206
rect 21532 7084 21588 7140
rect 21084 6524 21140 6580
rect 20860 6300 20916 6356
rect 21532 6300 21588 6356
rect 21420 5852 21476 5908
rect 20860 4396 20916 4452
rect 20972 5180 21028 5236
rect 21196 4620 21252 4676
rect 20972 4060 21028 4116
rect 21084 4172 21140 4228
rect 20412 2828 20468 2884
rect 20748 2098 20804 2100
rect 20748 2046 20750 2098
rect 20750 2046 20802 2098
rect 20802 2046 20804 2098
rect 20748 2044 20804 2046
rect 20860 1708 20916 1764
rect 20972 2156 21028 2212
rect 20300 1484 20356 1540
rect 16828 1372 16884 1428
rect 16380 1260 16436 1316
rect 20748 1260 20804 1316
rect 20636 924 20692 980
rect 20972 1260 21028 1316
rect 21196 2268 21252 2324
rect 21868 9100 21924 9156
rect 21868 8316 21924 8372
rect 21868 7756 21924 7812
rect 22092 9996 22148 10052
rect 23100 12348 23156 12404
rect 23436 13356 23492 13412
rect 23324 12066 23380 12068
rect 23324 12014 23326 12066
rect 23326 12014 23378 12066
rect 23378 12014 23380 12066
rect 23324 12012 23380 12014
rect 23548 13020 23604 13076
rect 23660 13132 23716 13188
rect 23996 13132 24052 13188
rect 24108 13020 24164 13076
rect 23804 12570 23860 12572
rect 23804 12518 23806 12570
rect 23806 12518 23858 12570
rect 23858 12518 23860 12570
rect 23804 12516 23860 12518
rect 23908 12570 23964 12572
rect 23908 12518 23910 12570
rect 23910 12518 23962 12570
rect 23962 12518 23964 12570
rect 23908 12516 23964 12518
rect 24012 12570 24068 12572
rect 24012 12518 24014 12570
rect 24014 12518 24066 12570
rect 24066 12518 24068 12570
rect 24012 12516 24068 12518
rect 23884 12402 23940 12404
rect 23884 12350 23886 12402
rect 23886 12350 23938 12402
rect 23938 12350 23940 12402
rect 23884 12348 23940 12350
rect 24464 13354 24520 13356
rect 24332 13244 24388 13300
rect 24464 13302 24466 13354
rect 24466 13302 24518 13354
rect 24518 13302 24520 13354
rect 24464 13300 24520 13302
rect 24568 13354 24624 13356
rect 24568 13302 24570 13354
rect 24570 13302 24622 13354
rect 24622 13302 24624 13354
rect 24568 13300 24624 13302
rect 24672 13354 24728 13356
rect 24672 13302 24674 13354
rect 24674 13302 24726 13354
rect 24726 13302 24728 13354
rect 24672 13300 24728 13302
rect 24556 13020 24612 13076
rect 24220 12348 24276 12404
rect 24892 12908 24948 12964
rect 23772 12124 23828 12180
rect 24332 11788 24388 11844
rect 22764 9996 22820 10052
rect 22428 9436 22484 9492
rect 22428 8764 22484 8820
rect 23436 9324 23492 9380
rect 23100 8540 23156 8596
rect 24464 11786 24520 11788
rect 24464 11734 24466 11786
rect 24466 11734 24518 11786
rect 24518 11734 24520 11786
rect 24464 11732 24520 11734
rect 24568 11786 24624 11788
rect 24568 11734 24570 11786
rect 24570 11734 24622 11786
rect 24622 11734 24624 11786
rect 24568 11732 24624 11734
rect 24672 11786 24728 11788
rect 24672 11734 24674 11786
rect 24674 11734 24726 11786
rect 24726 11734 24728 11786
rect 24672 11732 24728 11734
rect 25788 13804 25844 13860
rect 25676 13580 25732 13636
rect 25900 13580 25956 13636
rect 25452 13074 25508 13076
rect 25452 13022 25454 13074
rect 25454 13022 25506 13074
rect 25506 13022 25508 13074
rect 25452 13020 25508 13022
rect 25004 12460 25060 12516
rect 24892 11676 24948 11732
rect 23996 11116 24052 11172
rect 23804 11002 23860 11004
rect 23804 10950 23806 11002
rect 23806 10950 23858 11002
rect 23858 10950 23860 11002
rect 23804 10948 23860 10950
rect 23908 11002 23964 11004
rect 23908 10950 23910 11002
rect 23910 10950 23962 11002
rect 23962 10950 23964 11002
rect 23908 10948 23964 10950
rect 24012 11002 24068 11004
rect 24012 10950 24014 11002
rect 24014 10950 24066 11002
rect 24066 10950 24068 11002
rect 24012 10948 24068 10950
rect 24556 11116 24612 11172
rect 24444 10892 24500 10948
rect 25004 10780 25060 10836
rect 24464 10218 24520 10220
rect 24464 10166 24466 10218
rect 24466 10166 24518 10218
rect 24518 10166 24520 10218
rect 24464 10164 24520 10166
rect 24568 10218 24624 10220
rect 24568 10166 24570 10218
rect 24570 10166 24622 10218
rect 24622 10166 24624 10218
rect 24568 10164 24624 10166
rect 24672 10218 24728 10220
rect 24672 10166 24674 10218
rect 24674 10166 24726 10218
rect 24726 10166 24728 10218
rect 24672 10164 24728 10166
rect 25004 9884 25060 9940
rect 25228 9772 25284 9828
rect 23548 9100 23604 9156
rect 23660 9548 23716 9604
rect 23436 8540 23492 8596
rect 22092 8092 22148 8148
rect 22316 8204 22372 8260
rect 21980 7196 22036 7252
rect 21868 7084 21924 7140
rect 21868 6076 21924 6132
rect 21868 5628 21924 5684
rect 22092 5740 22148 5796
rect 22092 5516 22148 5572
rect 23212 8204 23268 8260
rect 22428 8146 22484 8148
rect 22428 8094 22430 8146
rect 22430 8094 22482 8146
rect 22482 8094 22484 8146
rect 22428 8092 22484 8094
rect 23212 7980 23268 8036
rect 23996 9548 24052 9604
rect 23804 9434 23860 9436
rect 23804 9382 23806 9434
rect 23806 9382 23858 9434
rect 23858 9382 23860 9434
rect 23804 9380 23860 9382
rect 23908 9434 23964 9436
rect 23908 9382 23910 9434
rect 23910 9382 23962 9434
rect 23962 9382 23964 9434
rect 23908 9380 23964 9382
rect 24012 9434 24068 9436
rect 24012 9382 24014 9434
rect 24014 9382 24066 9434
rect 24066 9382 24068 9434
rect 24012 9380 24068 9382
rect 25228 8876 25284 8932
rect 24464 8650 24520 8652
rect 24332 8540 24388 8596
rect 24464 8598 24466 8650
rect 24466 8598 24518 8650
rect 24518 8598 24520 8650
rect 24464 8596 24520 8598
rect 24568 8650 24624 8652
rect 24568 8598 24570 8650
rect 24570 8598 24622 8650
rect 24622 8598 24624 8650
rect 24568 8596 24624 8598
rect 24672 8650 24728 8652
rect 24672 8598 24674 8650
rect 24674 8598 24726 8650
rect 24726 8598 24728 8650
rect 24672 8596 24728 8598
rect 23804 7866 23860 7868
rect 23804 7814 23806 7866
rect 23806 7814 23858 7866
rect 23858 7814 23860 7866
rect 23804 7812 23860 7814
rect 23908 7866 23964 7868
rect 23908 7814 23910 7866
rect 23910 7814 23962 7866
rect 23962 7814 23964 7866
rect 23908 7812 23964 7814
rect 24012 7866 24068 7868
rect 24012 7814 24014 7866
rect 24014 7814 24066 7866
rect 24066 7814 24068 7866
rect 24012 7812 24068 7814
rect 24556 7980 24612 8036
rect 24444 7644 24500 7700
rect 23436 7420 23492 7476
rect 23660 7420 23716 7476
rect 22764 6524 22820 6580
rect 21756 3276 21812 3332
rect 22092 3276 22148 3332
rect 21756 2940 21812 2996
rect 21868 3052 21924 3108
rect 21868 2380 21924 2436
rect 21532 1932 21588 1988
rect 21644 1708 21700 1764
rect 21084 1036 21140 1092
rect 21308 1148 21364 1204
rect 20860 924 20916 980
rect 19964 476 20020 532
rect 16156 252 16212 308
rect 17948 364 18004 420
rect 1148 28 1204 84
rect 19964 28 20020 84
rect 21532 1148 21588 1204
rect 21644 812 21700 868
rect 21532 252 21588 308
rect 23324 6412 23380 6468
rect 23324 4732 23380 4788
rect 23436 5180 23492 5236
rect 23660 6972 23716 7028
rect 25340 8764 25396 8820
rect 25340 7308 25396 7364
rect 24464 7082 24520 7084
rect 24464 7030 24466 7082
rect 24466 7030 24518 7082
rect 24518 7030 24520 7082
rect 24464 7028 24520 7030
rect 24568 7082 24624 7084
rect 24568 7030 24570 7082
rect 24570 7030 24622 7082
rect 24622 7030 24624 7082
rect 24568 7028 24624 7030
rect 24672 7082 24728 7084
rect 24672 7030 24674 7082
rect 24674 7030 24726 7082
rect 24726 7030 24728 7082
rect 25228 7084 25284 7140
rect 24672 7028 24728 7030
rect 25452 6972 25508 7028
rect 25116 6748 25172 6804
rect 23772 6524 23828 6580
rect 23996 6578 24052 6580
rect 23996 6526 23998 6578
rect 23998 6526 24050 6578
rect 24050 6526 24052 6578
rect 23996 6524 24052 6526
rect 23804 6298 23860 6300
rect 23804 6246 23806 6298
rect 23806 6246 23858 6298
rect 23858 6246 23860 6298
rect 23804 6244 23860 6246
rect 23908 6298 23964 6300
rect 23908 6246 23910 6298
rect 23910 6246 23962 6298
rect 23962 6246 23964 6298
rect 23908 6244 23964 6246
rect 24012 6298 24068 6300
rect 24012 6246 24014 6298
rect 24014 6246 24066 6298
rect 24066 6246 24068 6298
rect 24012 6244 24068 6246
rect 24220 6300 24276 6356
rect 24108 5964 24164 6020
rect 24556 5852 24612 5908
rect 24220 5516 24276 5572
rect 24332 5404 24388 5460
rect 24464 5514 24520 5516
rect 24464 5462 24466 5514
rect 24466 5462 24518 5514
rect 24518 5462 24520 5514
rect 24464 5460 24520 5462
rect 24568 5514 24624 5516
rect 24568 5462 24570 5514
rect 24570 5462 24622 5514
rect 24622 5462 24624 5514
rect 24568 5460 24624 5462
rect 24672 5514 24728 5516
rect 24672 5462 24674 5514
rect 24674 5462 24726 5514
rect 24726 5462 24728 5514
rect 24672 5460 24728 5462
rect 24892 5516 24948 5572
rect 23660 5180 23716 5236
rect 23548 4956 23604 5012
rect 25004 5404 25060 5460
rect 24892 4844 24948 4900
rect 25228 4844 25284 4900
rect 23804 4730 23860 4732
rect 22764 3276 22820 3332
rect 23660 4620 23716 4676
rect 23804 4678 23806 4730
rect 23806 4678 23858 4730
rect 23858 4678 23860 4730
rect 23804 4676 23860 4678
rect 23908 4730 23964 4732
rect 23908 4678 23910 4730
rect 23910 4678 23962 4730
rect 23962 4678 23964 4730
rect 23908 4676 23964 4678
rect 24012 4730 24068 4732
rect 24012 4678 24014 4730
rect 24014 4678 24066 4730
rect 24066 4678 24068 4730
rect 24012 4676 24068 4678
rect 24220 4620 24276 4676
rect 25228 4172 25284 4228
rect 24220 3948 24276 4004
rect 25452 4620 25508 4676
rect 24464 3946 24520 3948
rect 24464 3894 24466 3946
rect 24466 3894 24518 3946
rect 24518 3894 24520 3946
rect 24464 3892 24520 3894
rect 24568 3946 24624 3948
rect 24568 3894 24570 3946
rect 24570 3894 24622 3946
rect 24622 3894 24624 3946
rect 24568 3892 24624 3894
rect 24672 3946 24728 3948
rect 24672 3894 24674 3946
rect 24674 3894 24726 3946
rect 24726 3894 24728 3946
rect 25340 3948 25396 4004
rect 25564 4396 25620 4452
rect 24672 3892 24728 3894
rect 25564 3612 25620 3668
rect 25788 13132 25844 13188
rect 26236 13244 26292 13300
rect 26348 13468 26404 13524
rect 25900 11564 25956 11620
rect 26012 12908 26068 12964
rect 27244 13244 27300 13300
rect 27132 12572 27188 12628
rect 27356 11900 27412 11956
rect 27804 13916 27860 13972
rect 27580 11900 27636 11956
rect 27692 13692 27748 13748
rect 27356 11116 27412 11172
rect 26796 10556 26852 10612
rect 26348 10220 26404 10276
rect 27020 10332 27076 10388
rect 26012 10108 26068 10164
rect 26012 9212 26068 9268
rect 25788 8204 25844 8260
rect 26236 8428 26292 8484
rect 26796 8540 26852 8596
rect 26348 8316 26404 8372
rect 26236 8204 26292 8260
rect 26908 8204 26964 8260
rect 27020 7980 27076 8036
rect 26012 7644 26068 7700
rect 25788 5180 25844 5236
rect 25788 4620 25844 4676
rect 25900 4396 25956 4452
rect 23548 3052 23604 3108
rect 23660 3164 23716 3220
rect 23804 3162 23860 3164
rect 23804 3110 23806 3162
rect 23806 3110 23858 3162
rect 23858 3110 23860 3162
rect 23804 3108 23860 3110
rect 23908 3162 23964 3164
rect 23908 3110 23910 3162
rect 23910 3110 23962 3162
rect 23962 3110 23964 3162
rect 23908 3108 23964 3110
rect 24012 3162 24068 3164
rect 24012 3110 24014 3162
rect 24014 3110 24066 3162
rect 24066 3110 24068 3162
rect 24012 3108 24068 3110
rect 25788 3836 25844 3892
rect 24220 3052 24276 3108
rect 25228 3164 25284 3220
rect 24892 2770 24948 2772
rect 24892 2718 24894 2770
rect 24894 2718 24946 2770
rect 24946 2718 24948 2770
rect 24892 2716 24948 2718
rect 25788 3276 25844 3332
rect 24220 2380 24276 2436
rect 24464 2378 24520 2380
rect 24332 2268 24388 2324
rect 24464 2326 24466 2378
rect 24466 2326 24518 2378
rect 24518 2326 24520 2378
rect 24464 2324 24520 2326
rect 24568 2378 24624 2380
rect 24568 2326 24570 2378
rect 24570 2326 24622 2378
rect 24622 2326 24624 2378
rect 24568 2324 24624 2326
rect 24672 2378 24728 2380
rect 24672 2326 24674 2378
rect 24674 2326 24726 2378
rect 24726 2326 24728 2378
rect 24672 2324 24728 2326
rect 23772 1932 23828 1988
rect 23884 1708 23940 1764
rect 23324 1596 23380 1652
rect 23804 1594 23860 1596
rect 23804 1542 23806 1594
rect 23806 1542 23858 1594
rect 23858 1542 23860 1594
rect 23804 1540 23860 1542
rect 23908 1594 23964 1596
rect 23908 1542 23910 1594
rect 23910 1542 23962 1594
rect 23962 1542 23964 1594
rect 23908 1540 23964 1542
rect 24012 1594 24068 1596
rect 24012 1542 24014 1594
rect 24014 1542 24066 1594
rect 24066 1542 24068 1594
rect 24012 1540 24068 1542
rect 24668 1708 24724 1764
rect 23548 1372 23604 1428
rect 24444 1372 24500 1428
rect 23996 1148 24052 1204
rect 23324 924 23380 980
rect 22428 252 22484 308
rect 23324 700 23380 756
rect 24332 812 24388 868
rect 24464 810 24520 812
rect 23436 476 23492 532
rect 24220 700 24276 756
rect 24464 758 24466 810
rect 24466 758 24518 810
rect 24518 758 24520 810
rect 24464 756 24520 758
rect 24568 810 24624 812
rect 24568 758 24570 810
rect 24570 758 24622 810
rect 24622 758 24624 810
rect 24568 756 24624 758
rect 24672 810 24728 812
rect 24672 758 24674 810
rect 24674 758 24726 810
rect 24726 758 24728 810
rect 24892 812 24948 868
rect 24672 756 24728 758
rect 25228 2492 25284 2548
rect 25116 2098 25172 2100
rect 25116 2046 25118 2098
rect 25118 2046 25170 2098
rect 25170 2046 25172 2098
rect 25116 2044 25172 2046
rect 25004 700 25060 756
rect 25228 1708 25284 1764
rect 25676 1372 25732 1428
rect 25676 1036 25732 1092
rect 25228 588 25284 644
rect 27468 7196 27524 7252
rect 27468 6636 27524 6692
rect 26908 6524 26964 6580
rect 26796 6188 26852 6244
rect 26908 5740 26964 5796
rect 26572 5404 26628 5460
rect 26796 5404 26852 5460
rect 26796 4956 26852 5012
rect 26124 3276 26180 3332
rect 26124 2940 26180 2996
rect 27020 4956 27076 5012
rect 27132 5404 27188 5460
rect 26908 2940 26964 2996
rect 27020 3500 27076 3556
rect 27244 4172 27300 4228
rect 27244 2828 27300 2884
rect 27916 12572 27972 12628
rect 28028 11788 28084 11844
rect 28140 12460 28196 12516
rect 27804 11228 27860 11284
rect 27916 10220 27972 10276
rect 27916 7196 27972 7252
rect 28028 9772 28084 9828
rect 27916 6076 27972 6132
rect 28252 12348 28308 12404
rect 28252 11004 28308 11060
rect 28364 12236 28420 12292
rect 28140 9100 28196 9156
rect 28252 10668 28308 10724
rect 28924 13916 28980 13972
rect 28700 12796 28756 12852
rect 28588 11676 28644 11732
rect 28364 9772 28420 9828
rect 28924 12572 28980 12628
rect 29260 12572 29316 12628
rect 28924 10108 28980 10164
rect 29148 11116 29204 11172
rect 29372 11116 29428 11172
rect 29484 13356 29540 13412
rect 29148 9660 29204 9716
rect 28700 9324 28756 9380
rect 29260 9212 29316 9268
rect 28252 8092 28308 8148
rect 28476 8428 28532 8484
rect 28364 6748 28420 6804
rect 28364 6188 28420 6244
rect 28028 5964 28084 6020
rect 28812 8204 28868 8260
rect 28924 8316 28980 8372
rect 28476 5628 28532 5684
rect 28700 5852 28756 5908
rect 28476 5234 28532 5236
rect 28476 5182 28478 5234
rect 28478 5182 28530 5234
rect 28530 5182 28532 5234
rect 28476 5180 28532 5182
rect 28476 4620 28532 4676
rect 27804 4508 27860 4564
rect 27804 4172 27860 4228
rect 27692 2604 27748 2660
rect 28140 2828 28196 2884
rect 28028 2044 28084 2100
rect 27244 1596 27300 1652
rect 27132 1148 27188 1204
rect 28028 1148 28084 1204
rect 28588 4172 28644 4228
rect 28588 3276 28644 3332
rect 28812 5346 28868 5348
rect 28812 5294 28814 5346
rect 28814 5294 28866 5346
rect 28866 5294 28868 5346
rect 28812 5292 28868 5294
rect 28924 4620 28980 4676
rect 29148 6636 29204 6692
rect 29036 2828 29092 2884
rect 28476 2604 28532 2660
rect 28252 2492 28308 2548
rect 28700 2492 28756 2548
rect 28252 2044 28308 2100
rect 28588 2156 28644 2212
rect 28588 1036 28644 1092
rect 28140 588 28196 644
rect 26796 476 26852 532
rect 27020 364 27076 420
rect 28140 364 28196 420
rect 26796 252 26852 308
rect 29820 13356 29876 13412
rect 30716 14028 30772 14084
rect 30268 12460 30324 12516
rect 30380 13692 30436 13748
rect 30156 12012 30212 12068
rect 30156 11676 30212 11732
rect 30268 10444 30324 10500
rect 29484 7532 29540 7588
rect 29596 9548 29652 9604
rect 29260 4508 29316 4564
rect 29372 7420 29428 7476
rect 29260 2882 29316 2884
rect 29260 2830 29262 2882
rect 29262 2830 29314 2882
rect 29314 2830 29316 2882
rect 29260 2828 29316 2830
rect 29372 2492 29428 2548
rect 29484 5180 29540 5236
rect 29708 7420 29764 7476
rect 30044 9100 30100 9156
rect 30156 8988 30212 9044
rect 30156 8316 30212 8372
rect 30044 8092 30100 8148
rect 30044 7084 30100 7140
rect 30044 6524 30100 6580
rect 30156 6748 30212 6804
rect 29820 6412 29876 6468
rect 30044 5740 30100 5796
rect 29708 2716 29764 2772
rect 29820 4508 29876 4564
rect 30156 5068 30212 5124
rect 31052 12012 31108 12068
rect 30716 11788 30772 11844
rect 31052 10668 31108 10724
rect 31388 13468 31444 13524
rect 31500 11564 31556 11620
rect 31388 10668 31444 10724
rect 31836 13020 31892 13076
rect 31836 12124 31892 12180
rect 31612 9996 31668 10052
rect 31724 11900 31780 11956
rect 31500 9212 31556 9268
rect 30380 6636 30436 6692
rect 30716 7196 30772 7252
rect 30380 5794 30436 5796
rect 30380 5742 30382 5794
rect 30382 5742 30434 5794
rect 30434 5742 30436 5794
rect 30380 5740 30436 5742
rect 30268 4844 30324 4900
rect 30716 4844 30772 4900
rect 30828 7084 30884 7140
rect 30044 3276 30100 3332
rect 30492 3388 30548 3444
rect 30940 5794 30996 5796
rect 30940 5742 30942 5794
rect 30942 5742 30994 5794
rect 30994 5742 30996 5794
rect 30940 5740 30996 5742
rect 31164 7196 31220 7252
rect 31052 5292 31108 5348
rect 31164 6412 31220 6468
rect 31052 5068 31108 5124
rect 31052 4284 31108 4340
rect 29820 1932 29876 1988
rect 30380 1986 30436 1988
rect 30380 1934 30382 1986
rect 30382 1934 30434 1986
rect 30434 1934 30436 1986
rect 30380 1932 30436 1934
rect 29596 1484 29652 1540
rect 30940 4060 30996 4116
rect 30716 2828 30772 2884
rect 30604 2716 30660 2772
rect 32060 10780 32116 10836
rect 32284 12124 32340 12180
rect 31836 10668 31892 10724
rect 33292 13132 33348 13188
rect 32956 12796 33012 12852
rect 33180 12796 33236 12852
rect 32508 11900 32564 11956
rect 32844 11788 32900 11844
rect 32284 9548 32340 9604
rect 32508 9548 32564 9604
rect 31836 8764 31892 8820
rect 31612 7644 31668 7700
rect 31612 7084 31668 7140
rect 31724 7532 31780 7588
rect 31500 6300 31556 6356
rect 32508 8988 32564 9044
rect 33068 11788 33124 11844
rect 32956 10556 33012 10612
rect 32956 8652 33012 8708
rect 31948 7084 32004 7140
rect 32844 7644 32900 7700
rect 31836 6300 31892 6356
rect 32060 6412 32116 6468
rect 31836 6018 31892 6020
rect 31836 5966 31838 6018
rect 31838 5966 31890 6018
rect 31890 5966 31892 6018
rect 31836 5964 31892 5966
rect 31724 4284 31780 4340
rect 32172 5852 32228 5908
rect 32396 5068 32452 5124
rect 31164 3388 31220 3444
rect 31052 3276 31108 3332
rect 31052 2828 31108 2884
rect 31276 2716 31332 2772
rect 31948 2770 32004 2772
rect 31948 2718 31950 2770
rect 31950 2718 32002 2770
rect 32002 2718 32004 2770
rect 31948 2716 32004 2718
rect 30940 2156 30996 2212
rect 30604 1708 30660 1764
rect 31164 1596 31220 1652
rect 30492 1372 30548 1428
rect 31836 1484 31892 1540
rect 31836 1036 31892 1092
rect 32060 1036 32116 1092
rect 32172 700 32228 756
rect 31388 140 31444 196
rect 32396 2770 32452 2772
rect 32396 2718 32398 2770
rect 32398 2718 32450 2770
rect 32450 2718 32452 2770
rect 32396 2716 32452 2718
rect 32396 2380 32452 2436
rect 32396 2156 32452 2212
rect 32956 5852 33012 5908
rect 32844 4396 32900 4452
rect 32956 5516 33012 5572
rect 33180 9548 33236 9604
rect 33404 12012 33460 12068
rect 33628 13020 33684 13076
rect 33404 11564 33460 11620
rect 33628 11228 33684 11284
rect 33740 12012 33796 12068
rect 33628 10444 33684 10500
rect 33852 11788 33908 11844
rect 33964 13804 34020 13860
rect 33740 10220 33796 10276
rect 34076 13356 34132 13412
rect 33964 10892 34020 10948
rect 33964 10220 34020 10276
rect 33628 9884 33684 9940
rect 33628 9660 33684 9716
rect 33404 7980 33460 8036
rect 33516 8092 33572 8148
rect 33292 7868 33348 7924
rect 33180 7308 33236 7364
rect 33068 5068 33124 5124
rect 33404 7308 33460 7364
rect 33852 9548 33908 9604
rect 33628 7868 33684 7924
rect 33740 9324 33796 9380
rect 33516 5852 33572 5908
rect 33628 7532 33684 7588
rect 33404 5180 33460 5236
rect 33292 5068 33348 5124
rect 33740 6860 33796 6916
rect 33740 6636 33796 6692
rect 34748 13580 34804 13636
rect 35084 13580 35140 13636
rect 34300 12684 34356 12740
rect 34860 12236 34916 12292
rect 34524 11900 34580 11956
rect 34188 11506 34244 11508
rect 34188 11454 34190 11506
rect 34190 11454 34242 11506
rect 34242 11454 34244 11506
rect 34188 11452 34244 11454
rect 34076 9884 34132 9940
rect 34300 11116 34356 11172
rect 33852 5404 33908 5460
rect 34076 5180 34132 5236
rect 33628 4956 33684 5012
rect 33292 4284 33348 4340
rect 33516 3500 33572 3556
rect 33516 3164 33572 3220
rect 34748 11900 34804 11956
rect 34748 9212 34804 9268
rect 34972 11394 35028 11396
rect 34972 11342 34974 11394
rect 34974 11342 35026 11394
rect 35026 11342 35028 11394
rect 34972 11340 35028 11342
rect 36092 12348 36148 12404
rect 36204 12684 36260 12740
rect 35644 12124 35700 12180
rect 35980 12124 36036 12180
rect 35196 10108 35252 10164
rect 35644 11788 35700 11844
rect 34972 8764 35028 8820
rect 35084 9212 35140 9268
rect 34860 8092 34916 8148
rect 35532 8876 35588 8932
rect 35308 8764 35364 8820
rect 35196 8370 35252 8372
rect 35196 8318 35198 8370
rect 35198 8318 35250 8370
rect 35250 8318 35252 8370
rect 35196 8316 35252 8318
rect 35084 5964 35140 6020
rect 35196 7084 35252 7140
rect 34636 4844 34692 4900
rect 34188 2380 34244 2436
rect 32732 1148 32788 1204
rect 32396 476 32452 532
rect 32844 364 32900 420
rect 34076 1596 34132 1652
rect 32284 140 32340 196
rect 34972 4732 35028 4788
rect 34972 4396 35028 4452
rect 35420 7420 35476 7476
rect 35420 7084 35476 7140
rect 35532 6748 35588 6804
rect 35308 6076 35364 6132
rect 35196 4396 35252 4452
rect 35308 5292 35364 5348
rect 35196 3948 35252 4004
rect 34636 1484 34692 1540
rect 34524 700 34580 756
rect 35308 3836 35364 3892
rect 35868 10050 35924 10052
rect 35868 9998 35870 10050
rect 35870 9998 35922 10050
rect 35922 9998 35924 10050
rect 35868 9996 35924 9998
rect 35756 9660 35812 9716
rect 35868 9548 35924 9604
rect 35868 6412 35924 6468
rect 35756 5516 35812 5572
rect 35868 5964 35924 6020
rect 35756 4844 35812 4900
rect 35196 2828 35252 2884
rect 35308 2940 35364 2996
rect 35308 2268 35364 2324
rect 36092 10050 36148 10052
rect 36092 9998 36094 10050
rect 36094 9998 36146 10050
rect 36146 9998 36148 10050
rect 36092 9996 36148 9998
rect 36316 12066 36372 12068
rect 36316 12014 36318 12066
rect 36318 12014 36370 12066
rect 36370 12014 36372 12066
rect 36316 12012 36372 12014
rect 37324 13244 37380 13300
rect 36652 11564 36708 11620
rect 36764 12460 36820 12516
rect 37100 12290 37156 12292
rect 37100 12238 37102 12290
rect 37102 12238 37154 12290
rect 37154 12238 37156 12290
rect 37100 12236 37156 12238
rect 38780 13244 38836 13300
rect 38556 12684 38612 12740
rect 39676 13468 39732 13524
rect 39340 13244 39396 13300
rect 39340 12124 39396 12180
rect 38332 12012 38388 12068
rect 38220 11900 38276 11956
rect 38780 11900 38836 11956
rect 37884 11788 37940 11844
rect 36764 11116 36820 11172
rect 37100 10722 37156 10724
rect 37100 10670 37102 10722
rect 37102 10670 37154 10722
rect 37154 10670 37156 10722
rect 37100 10668 37156 10670
rect 37212 9884 37268 9940
rect 36652 9826 36708 9828
rect 36652 9774 36654 9826
rect 36654 9774 36706 9826
rect 36706 9774 36708 9826
rect 36652 9772 36708 9774
rect 36540 8876 36596 8932
rect 37100 8428 37156 8484
rect 36204 6860 36260 6916
rect 36876 6972 36932 7028
rect 36540 5404 36596 5460
rect 36316 4732 36372 4788
rect 36204 4450 36260 4452
rect 36204 4398 36206 4450
rect 36206 4398 36258 4450
rect 36258 4398 36260 4450
rect 36204 4396 36260 4398
rect 35980 4284 36036 4340
rect 36204 3948 36260 4004
rect 36540 4732 36596 4788
rect 36540 4396 36596 4452
rect 36988 6860 37044 6916
rect 36988 6524 37044 6580
rect 37772 9436 37828 9492
rect 37772 8540 37828 8596
rect 38332 11228 38388 11284
rect 38108 10108 38164 10164
rect 38108 9548 38164 9604
rect 37996 9436 38052 9492
rect 39676 11228 39732 11284
rect 39340 11004 39396 11060
rect 39340 10780 39396 10836
rect 39676 10556 39732 10612
rect 40236 12908 40292 12964
rect 40236 10892 40292 10948
rect 40348 11564 40404 11620
rect 40236 10332 40292 10388
rect 40236 9772 40292 9828
rect 39788 8370 39844 8372
rect 39788 8318 39790 8370
rect 39790 8318 39842 8370
rect 39842 8318 39844 8370
rect 39788 8316 39844 8318
rect 38780 8092 38836 8148
rect 38612 7980 38668 8036
rect 38780 7868 38836 7924
rect 38444 7420 38500 7476
rect 38612 7420 38668 7476
rect 37884 6972 37940 7028
rect 37212 6524 37268 6580
rect 37100 6412 37156 6468
rect 36988 6076 37044 6132
rect 37996 6300 38052 6356
rect 37324 5852 37380 5908
rect 36988 4620 37044 4676
rect 37548 5180 37604 5236
rect 36652 4284 36708 4340
rect 35868 2604 35924 2660
rect 35756 2268 35812 2324
rect 37100 3724 37156 3780
rect 36652 2940 36708 2996
rect 36876 3388 36932 3444
rect 36876 2044 36932 2100
rect 36092 1708 36148 1764
rect 38220 5180 38276 5236
rect 38556 6188 38612 6244
rect 39004 6524 39060 6580
rect 39228 6578 39284 6580
rect 39228 6526 39230 6578
rect 39230 6526 39282 6578
rect 39282 6526 39284 6578
rect 39228 6524 39284 6526
rect 39004 6300 39060 6356
rect 38780 5068 38836 5124
rect 39900 4508 39956 4564
rect 38668 4172 38724 4228
rect 40236 8370 40292 8372
rect 40236 8318 40238 8370
rect 40238 8318 40290 8370
rect 40290 8318 40292 8370
rect 40236 8316 40292 8318
rect 41468 13132 41524 13188
rect 41020 13020 41076 13076
rect 40572 10780 40628 10836
rect 42140 12684 42196 12740
rect 40684 7084 40740 7140
rect 40460 6972 40516 7028
rect 40124 6860 40180 6916
rect 40348 6860 40404 6916
rect 40236 6748 40292 6804
rect 40460 5292 40516 5348
rect 40572 5852 40628 5908
rect 40348 4508 40404 4564
rect 40236 4396 40292 4452
rect 40012 3948 40068 4004
rect 38220 3276 38276 3332
rect 37660 2882 37716 2884
rect 37660 2830 37662 2882
rect 37662 2830 37714 2882
rect 37714 2830 37716 2882
rect 37660 2828 37716 2830
rect 38332 2604 38388 2660
rect 38444 2492 38500 2548
rect 41692 11676 41748 11732
rect 41132 10498 41188 10500
rect 41132 10446 41134 10498
rect 41134 10446 41186 10498
rect 41186 10446 41188 10498
rect 41132 10444 41188 10446
rect 41356 10498 41412 10500
rect 41356 10446 41358 10498
rect 41358 10446 41410 10498
rect 41410 10446 41412 10498
rect 41356 10444 41412 10446
rect 41132 10108 41188 10164
rect 41468 10108 41524 10164
rect 41244 9660 41300 9716
rect 41244 7980 41300 8036
rect 41580 7644 41636 7700
rect 41580 6972 41636 7028
rect 41020 4060 41076 4116
rect 41244 6524 41300 6580
rect 40572 2716 40628 2772
rect 40348 2604 40404 2660
rect 38556 1708 38612 1764
rect 38668 2044 38724 2100
rect 37548 1596 37604 1652
rect 38668 1484 38724 1540
rect 40236 1708 40292 1764
rect 39452 1260 39508 1316
rect 34748 252 34804 308
rect 36764 364 36820 420
rect 40348 1372 40404 1428
rect 41804 11116 41860 11172
rect 42028 10556 42084 10612
rect 41916 10498 41972 10500
rect 41916 10446 41918 10498
rect 41918 10446 41970 10498
rect 41970 10446 41972 10498
rect 41916 10444 41972 10446
rect 42364 12572 42420 12628
rect 42812 12236 42868 12292
rect 43036 12124 43092 12180
rect 42252 10610 42308 10612
rect 42252 10558 42254 10610
rect 42254 10558 42306 10610
rect 42306 10558 42308 10610
rect 42252 10556 42308 10558
rect 42700 10556 42756 10612
rect 42140 10220 42196 10276
rect 41804 9884 41860 9940
rect 42700 9548 42756 9604
rect 42252 9100 42308 9156
rect 42364 9436 42420 9492
rect 41916 8988 41972 9044
rect 41692 6524 41748 6580
rect 41916 7644 41972 7700
rect 41356 6300 41412 6356
rect 42028 6412 42084 6468
rect 41916 6076 41972 6132
rect 42140 5292 42196 5348
rect 41804 4956 41860 5012
rect 41356 4450 41412 4452
rect 41356 4398 41358 4450
rect 41358 4398 41410 4450
rect 41410 4398 41412 4450
rect 41356 4396 41412 4398
rect 41692 4396 41748 4452
rect 41692 4060 41748 4116
rect 41692 3500 41748 3556
rect 41916 3612 41972 3668
rect 42028 2828 42084 2884
rect 41804 2380 41860 2436
rect 41916 2156 41972 2212
rect 41244 1372 41300 1428
rect 42028 1036 42084 1092
rect 40236 476 40292 532
rect 40460 476 40516 532
rect 40460 140 40516 196
rect 42924 9548 42980 9604
rect 42924 8540 42980 8596
rect 42812 4956 42868 5012
rect 42364 3836 42420 3892
rect 42252 3612 42308 3668
rect 42364 3388 42420 3444
rect 42252 2940 42308 2996
rect 42364 2268 42420 2324
rect 43596 13916 43652 13972
rect 43260 11564 43316 11620
rect 43484 12236 43540 12292
rect 43148 9100 43204 9156
rect 43708 13580 43764 13636
rect 44604 13804 44660 13860
rect 44156 13132 44212 13188
rect 43804 12570 43860 12572
rect 43804 12518 43806 12570
rect 43806 12518 43858 12570
rect 43858 12518 43860 12570
rect 43804 12516 43860 12518
rect 43908 12570 43964 12572
rect 43908 12518 43910 12570
rect 43910 12518 43962 12570
rect 43962 12518 43964 12570
rect 43908 12516 43964 12518
rect 44012 12570 44068 12572
rect 44012 12518 44014 12570
rect 44014 12518 44066 12570
rect 44066 12518 44068 12570
rect 44012 12516 44068 12518
rect 44044 11452 44100 11508
rect 44156 11228 44212 11284
rect 44044 11116 44100 11172
rect 44464 13354 44520 13356
rect 44464 13302 44466 13354
rect 44466 13302 44518 13354
rect 44518 13302 44520 13354
rect 44464 13300 44520 13302
rect 44568 13354 44624 13356
rect 44568 13302 44570 13354
rect 44570 13302 44622 13354
rect 44622 13302 44624 13354
rect 44568 13300 44624 13302
rect 44672 13354 44728 13356
rect 44672 13302 44674 13354
rect 44674 13302 44726 13354
rect 44726 13302 44728 13354
rect 44672 13300 44728 13302
rect 44940 12962 44996 12964
rect 44940 12910 44942 12962
rect 44942 12910 44994 12962
rect 44994 12910 44996 12962
rect 44940 12908 44996 12910
rect 44492 12290 44548 12292
rect 44492 12238 44494 12290
rect 44494 12238 44546 12290
rect 44546 12238 44548 12290
rect 44492 12236 44548 12238
rect 44464 11786 44520 11788
rect 44464 11734 44466 11786
rect 44466 11734 44518 11786
rect 44518 11734 44520 11786
rect 44464 11732 44520 11734
rect 44568 11786 44624 11788
rect 44568 11734 44570 11786
rect 44570 11734 44622 11786
rect 44622 11734 44624 11786
rect 44568 11732 44624 11734
rect 44672 11786 44728 11788
rect 44672 11734 44674 11786
rect 44674 11734 44726 11786
rect 44726 11734 44728 11786
rect 44672 11732 44728 11734
rect 43804 11002 43860 11004
rect 43804 10950 43806 11002
rect 43806 10950 43858 11002
rect 43858 10950 43860 11002
rect 43804 10948 43860 10950
rect 43908 11002 43964 11004
rect 43908 10950 43910 11002
rect 43910 10950 43962 11002
rect 43962 10950 43964 11002
rect 43908 10948 43964 10950
rect 44012 11002 44068 11004
rect 44012 10950 44014 11002
rect 44014 10950 44066 11002
rect 44066 10950 44068 11002
rect 44012 10948 44068 10950
rect 43708 10780 43764 10836
rect 44268 10220 44324 10276
rect 44464 10218 44520 10220
rect 44464 10166 44466 10218
rect 44466 10166 44518 10218
rect 44518 10166 44520 10218
rect 44464 10164 44520 10166
rect 44568 10218 44624 10220
rect 44568 10166 44570 10218
rect 44570 10166 44622 10218
rect 44622 10166 44624 10218
rect 44568 10164 44624 10166
rect 44672 10218 44728 10220
rect 44672 10166 44674 10218
rect 44674 10166 44726 10218
rect 44726 10166 44728 10218
rect 44672 10164 44728 10166
rect 44156 9660 44212 9716
rect 43804 9434 43860 9436
rect 43804 9382 43806 9434
rect 43806 9382 43858 9434
rect 43858 9382 43860 9434
rect 43804 9380 43860 9382
rect 43908 9434 43964 9436
rect 43908 9382 43910 9434
rect 43910 9382 43962 9434
rect 43962 9382 43964 9434
rect 43908 9380 43964 9382
rect 44012 9434 44068 9436
rect 44012 9382 44014 9434
rect 44014 9382 44066 9434
rect 44066 9382 44068 9434
rect 44012 9380 44068 9382
rect 44044 8652 44100 8708
rect 43596 8428 43652 8484
rect 43596 7980 43652 8036
rect 44464 8650 44520 8652
rect 44464 8598 44466 8650
rect 44466 8598 44518 8650
rect 44518 8598 44520 8650
rect 44464 8596 44520 8598
rect 44568 8650 44624 8652
rect 44568 8598 44570 8650
rect 44570 8598 44622 8650
rect 44622 8598 44624 8650
rect 44568 8596 44624 8598
rect 44672 8650 44728 8652
rect 44672 8598 44674 8650
rect 44674 8598 44726 8650
rect 44726 8598 44728 8650
rect 44672 8596 44728 8598
rect 44268 8092 44324 8148
rect 43804 7866 43860 7868
rect 43804 7814 43806 7866
rect 43806 7814 43858 7866
rect 43858 7814 43860 7866
rect 43804 7812 43860 7814
rect 43908 7866 43964 7868
rect 43908 7814 43910 7866
rect 43910 7814 43962 7866
rect 43962 7814 43964 7866
rect 43908 7812 43964 7814
rect 44012 7866 44068 7868
rect 44012 7814 44014 7866
rect 44014 7814 44066 7866
rect 44066 7814 44068 7866
rect 44156 7868 44212 7924
rect 44012 7812 44068 7814
rect 43820 7420 43876 7476
rect 43820 7196 43876 7252
rect 44464 7082 44520 7084
rect 44268 6972 44324 7028
rect 44464 7030 44466 7082
rect 44466 7030 44518 7082
rect 44518 7030 44520 7082
rect 44464 7028 44520 7030
rect 44568 7082 44624 7084
rect 44568 7030 44570 7082
rect 44570 7030 44622 7082
rect 44622 7030 44624 7082
rect 44568 7028 44624 7030
rect 44672 7082 44728 7084
rect 44672 7030 44674 7082
rect 44674 7030 44726 7082
rect 44726 7030 44728 7082
rect 44672 7028 44728 7030
rect 43484 6188 43540 6244
rect 43804 6298 43860 6300
rect 43804 6246 43806 6298
rect 43806 6246 43858 6298
rect 43858 6246 43860 6298
rect 43804 6244 43860 6246
rect 43908 6298 43964 6300
rect 43908 6246 43910 6298
rect 43910 6246 43962 6298
rect 43962 6246 43964 6298
rect 43908 6244 43964 6246
rect 44012 6298 44068 6300
rect 44012 6246 44014 6298
rect 44014 6246 44066 6298
rect 44066 6246 44068 6298
rect 44012 6244 44068 6246
rect 43596 6076 43652 6132
rect 43596 5628 43652 5684
rect 44268 5628 44324 5684
rect 44464 5514 44520 5516
rect 44464 5462 44466 5514
rect 44466 5462 44518 5514
rect 44518 5462 44520 5514
rect 44464 5460 44520 5462
rect 44568 5514 44624 5516
rect 44568 5462 44570 5514
rect 44570 5462 44622 5514
rect 44622 5462 44624 5514
rect 44568 5460 44624 5462
rect 44672 5514 44728 5516
rect 44672 5462 44674 5514
rect 44674 5462 44726 5514
rect 44726 5462 44728 5514
rect 44672 5460 44728 5462
rect 43484 4620 43540 4676
rect 43804 4730 43860 4732
rect 43804 4678 43806 4730
rect 43806 4678 43858 4730
rect 43858 4678 43860 4730
rect 43804 4676 43860 4678
rect 43908 4730 43964 4732
rect 43908 4678 43910 4730
rect 43910 4678 43962 4730
rect 43962 4678 43964 4730
rect 43908 4676 43964 4678
rect 44012 4730 44068 4732
rect 44012 4678 44014 4730
rect 44014 4678 44066 4730
rect 44066 4678 44068 4730
rect 44156 4732 44212 4788
rect 44012 4676 44068 4678
rect 43596 4508 43652 4564
rect 43484 4396 43540 4452
rect 43484 3276 43540 3332
rect 44464 3946 44520 3948
rect 43708 3836 43764 3892
rect 44464 3894 44466 3946
rect 44466 3894 44518 3946
rect 44518 3894 44520 3946
rect 44464 3892 44520 3894
rect 44568 3946 44624 3948
rect 44568 3894 44570 3946
rect 44570 3894 44622 3946
rect 44622 3894 44624 3946
rect 44568 3892 44624 3894
rect 44672 3946 44728 3948
rect 44672 3894 44674 3946
rect 44674 3894 44726 3946
rect 44726 3894 44728 3946
rect 44672 3892 44728 3894
rect 44380 3442 44436 3444
rect 44380 3390 44382 3442
rect 44382 3390 44434 3442
rect 44434 3390 44436 3442
rect 44380 3388 44436 3390
rect 45724 14028 45780 14084
rect 45388 12796 45444 12852
rect 45500 12908 45556 12964
rect 45276 12290 45332 12292
rect 45276 12238 45278 12290
rect 45278 12238 45330 12290
rect 45330 12238 45332 12290
rect 45276 12236 45332 12238
rect 45164 9714 45220 9716
rect 45164 9662 45166 9714
rect 45166 9662 45218 9714
rect 45218 9662 45220 9714
rect 45164 9660 45220 9662
rect 45052 9548 45108 9604
rect 45276 8764 45332 8820
rect 45276 7644 45332 7700
rect 45388 6972 45444 7028
rect 45276 5180 45332 5236
rect 45388 6188 45444 6244
rect 45388 3948 45444 4004
rect 43596 3052 43652 3108
rect 43804 3162 43860 3164
rect 43804 3110 43806 3162
rect 43806 3110 43858 3162
rect 43858 3110 43860 3162
rect 43804 3108 43860 3110
rect 43908 3162 43964 3164
rect 43908 3110 43910 3162
rect 43910 3110 43962 3162
rect 43962 3110 43964 3162
rect 43908 3108 43964 3110
rect 44012 3162 44068 3164
rect 44012 3110 44014 3162
rect 44014 3110 44066 3162
rect 44066 3110 44068 3162
rect 44012 3108 44068 3110
rect 44464 2378 44520 2380
rect 44464 2326 44466 2378
rect 44466 2326 44518 2378
rect 44518 2326 44520 2378
rect 44464 2324 44520 2326
rect 44568 2378 44624 2380
rect 44568 2326 44570 2378
rect 44570 2326 44622 2378
rect 44622 2326 44624 2378
rect 44568 2324 44624 2326
rect 44672 2378 44728 2380
rect 44672 2326 44674 2378
rect 44674 2326 44726 2378
rect 44726 2326 44728 2378
rect 44672 2324 44728 2326
rect 43036 2044 43092 2100
rect 42252 1596 42308 1652
rect 44268 1820 44324 1876
rect 43804 1594 43860 1596
rect 43804 1542 43806 1594
rect 43806 1542 43858 1594
rect 43858 1542 43860 1594
rect 43804 1540 43860 1542
rect 43908 1594 43964 1596
rect 43908 1542 43910 1594
rect 43910 1542 43962 1594
rect 43962 1542 43964 1594
rect 43908 1540 43964 1542
rect 44012 1594 44068 1596
rect 44012 1542 44014 1594
rect 44014 1542 44066 1594
rect 44066 1542 44068 1594
rect 44012 1540 44068 1542
rect 44268 812 44324 868
rect 44828 1036 44884 1092
rect 44464 810 44520 812
rect 44464 758 44466 810
rect 44466 758 44518 810
rect 44518 758 44520 810
rect 44464 756 44520 758
rect 44568 810 44624 812
rect 44568 758 44570 810
rect 44570 758 44622 810
rect 44622 758 44624 810
rect 44568 756 44624 758
rect 44672 810 44728 812
rect 44672 758 44674 810
rect 44674 758 44726 810
rect 44726 758 44728 810
rect 44672 756 44728 758
rect 45612 11788 45668 11844
rect 45948 12460 46004 12516
rect 46060 12066 46116 12068
rect 46060 12014 46062 12066
rect 46062 12014 46114 12066
rect 46114 12014 46116 12066
rect 46060 12012 46116 12014
rect 45724 11676 45780 11732
rect 45948 11564 46004 11620
rect 45612 4396 45668 4452
rect 45724 8988 45780 9044
rect 45500 2940 45556 2996
rect 45836 3164 45892 3220
rect 44940 812 44996 868
rect 45276 1708 45332 1764
rect 45948 3052 46004 3108
rect 45836 1148 45892 1204
rect 46060 1148 46116 1204
rect 46844 13132 46900 13188
rect 46844 12962 46900 12964
rect 46844 12910 46846 12962
rect 46846 12910 46898 12962
rect 46898 12910 46900 12962
rect 46844 12908 46900 12910
rect 46956 12178 47012 12180
rect 46956 12126 46958 12178
rect 46958 12126 47010 12178
rect 47010 12126 47012 12178
rect 46956 12124 47012 12126
rect 46508 12012 46564 12068
rect 46732 12012 46788 12068
rect 46620 7868 46676 7924
rect 47852 13356 47908 13412
rect 48188 13132 48244 13188
rect 47964 13020 48020 13076
rect 47852 12348 47908 12404
rect 46956 10780 47012 10836
rect 47740 10556 47796 10612
rect 47180 9884 47236 9940
rect 47292 10444 47348 10500
rect 46956 9548 47012 9604
rect 46844 8818 46900 8820
rect 46844 8766 46846 8818
rect 46846 8766 46898 8818
rect 46898 8766 46900 8818
rect 46844 8764 46900 8766
rect 47068 8818 47124 8820
rect 47068 8766 47070 8818
rect 47070 8766 47122 8818
rect 47122 8766 47124 8818
rect 47068 8764 47124 8766
rect 46732 6748 46788 6804
rect 47068 7868 47124 7924
rect 47068 4732 47124 4788
rect 46620 1260 46676 1316
rect 47404 10108 47460 10164
rect 48076 12236 48132 12292
rect 47852 8988 47908 9044
rect 47964 10220 48020 10276
rect 47404 6076 47460 6132
rect 47516 6636 47572 6692
rect 47628 2940 47684 2996
rect 47740 8764 47796 8820
rect 49084 13580 49140 13636
rect 48972 13186 49028 13188
rect 48972 13134 48974 13186
rect 48974 13134 49026 13186
rect 49026 13134 49028 13186
rect 48972 13132 49028 13134
rect 48636 12348 48692 12404
rect 49420 12402 49476 12404
rect 49420 12350 49422 12402
rect 49422 12350 49474 12402
rect 49474 12350 49476 12402
rect 49420 12348 49476 12350
rect 48412 11788 48468 11844
rect 48188 11394 48244 11396
rect 48188 11342 48190 11394
rect 48190 11342 48242 11394
rect 48242 11342 48244 11394
rect 48188 11340 48244 11342
rect 48076 10108 48132 10164
rect 48076 8316 48132 8372
rect 48300 9548 48356 9604
rect 47964 6972 48020 7028
rect 48412 8370 48468 8372
rect 48412 8318 48414 8370
rect 48414 8318 48466 8370
rect 48466 8318 48468 8370
rect 48412 8316 48468 8318
rect 48300 5516 48356 5572
rect 48524 6748 48580 6804
rect 47740 2604 47796 2660
rect 48300 4172 48356 4228
rect 47292 1260 47348 1316
rect 47516 1596 47572 1652
rect 46396 588 46452 644
rect 46172 364 46228 420
rect 45276 252 45332 308
rect 49980 13468 50036 13524
rect 49532 11564 49588 11620
rect 49644 11900 49700 11956
rect 50428 12348 50484 12404
rect 49196 11340 49252 11396
rect 50316 11618 50372 11620
rect 50316 11566 50318 11618
rect 50318 11566 50370 11618
rect 50370 11566 50372 11618
rect 50316 11564 50372 11566
rect 49756 11506 49812 11508
rect 49756 11454 49758 11506
rect 49758 11454 49810 11506
rect 49810 11454 49812 11506
rect 49756 11452 49812 11454
rect 49644 11004 49700 11060
rect 49420 10332 49476 10388
rect 49532 10108 49588 10164
rect 48972 8876 49028 8932
rect 48972 8370 49028 8372
rect 48972 8318 48974 8370
rect 48974 8318 49026 8370
rect 49026 8318 49028 8370
rect 48972 8316 49028 8318
rect 48860 7196 48916 7252
rect 48972 6972 49028 7028
rect 48972 6188 49028 6244
rect 48748 5852 48804 5908
rect 48860 6076 48916 6132
rect 48636 5180 48692 5236
rect 48748 5628 48804 5684
rect 48748 4844 48804 4900
rect 48524 4172 48580 4228
rect 48972 4114 49028 4116
rect 48972 4062 48974 4114
rect 48974 4062 49026 4114
rect 49026 4062 49028 4114
rect 48972 4060 49028 4062
rect 49308 4114 49364 4116
rect 49308 4062 49310 4114
rect 49310 4062 49362 4114
rect 49362 4062 49364 4114
rect 49308 4060 49364 4062
rect 48860 924 48916 980
rect 48300 700 48356 756
rect 49532 4732 49588 4788
rect 49644 9100 49700 9156
rect 50204 10668 50260 10724
rect 50204 10220 50260 10276
rect 49868 8930 49924 8932
rect 49868 8878 49870 8930
rect 49870 8878 49922 8930
rect 49922 8878 49924 8930
rect 49868 8876 49924 8878
rect 51100 13580 51156 13636
rect 50988 12066 51044 12068
rect 50988 12014 50990 12066
rect 50990 12014 51042 12066
rect 51042 12014 51044 12066
rect 50988 12012 51044 12014
rect 50876 11564 50932 11620
rect 51212 11788 51268 11844
rect 52220 13132 52276 13188
rect 51772 13020 51828 13076
rect 51324 11676 51380 11732
rect 51884 11618 51940 11620
rect 51884 11566 51886 11618
rect 51886 11566 51938 11618
rect 51938 11566 51940 11618
rect 51884 11564 51940 11566
rect 50988 10444 51044 10500
rect 51100 9660 51156 9716
rect 50764 8428 50820 8484
rect 50316 7868 50372 7924
rect 50988 8370 51044 8372
rect 50988 8318 50990 8370
rect 50990 8318 51042 8370
rect 51042 8318 51044 8370
rect 50988 8316 51044 8318
rect 50988 6076 51044 6132
rect 51212 9324 51268 9380
rect 52892 13468 52948 13524
rect 52556 12402 52612 12404
rect 52556 12350 52558 12402
rect 52558 12350 52610 12402
rect 52610 12350 52612 12402
rect 52556 12348 52612 12350
rect 52108 10610 52164 10612
rect 52108 10558 52110 10610
rect 52110 10558 52162 10610
rect 52162 10558 52164 10610
rect 52108 10556 52164 10558
rect 51772 9938 51828 9940
rect 51772 9886 51774 9938
rect 51774 9886 51826 9938
rect 51826 9886 51828 9938
rect 51772 9884 51828 9886
rect 51324 9212 51380 9268
rect 51996 8146 52052 8148
rect 51996 8094 51998 8146
rect 51998 8094 52050 8146
rect 52050 8094 52052 8146
rect 51996 8092 52052 8094
rect 50428 4508 50484 4564
rect 50540 4620 50596 4676
rect 49756 3276 49812 3332
rect 49644 2716 49700 2772
rect 52108 6860 52164 6916
rect 52332 7532 52388 7588
rect 52220 6636 52276 6692
rect 51884 5404 51940 5460
rect 51436 4450 51492 4452
rect 51436 4398 51438 4450
rect 51438 4398 51490 4450
rect 51490 4398 51492 4450
rect 51436 4396 51492 4398
rect 51996 5234 52052 5236
rect 51996 5182 51998 5234
rect 51998 5182 52050 5234
rect 52050 5182 52052 5234
rect 51996 5180 52052 5182
rect 51436 4172 51492 4228
rect 51324 3164 51380 3220
rect 52556 11676 52612 11732
rect 53116 12348 53172 12404
rect 53900 12572 53956 12628
rect 52556 9826 52612 9828
rect 52556 9774 52558 9826
rect 52558 9774 52610 9826
rect 52610 9774 52612 9826
rect 52556 9772 52612 9774
rect 52780 8988 52836 9044
rect 52668 8876 52724 8932
rect 52556 8258 52612 8260
rect 52556 8206 52558 8258
rect 52558 8206 52610 8258
rect 52610 8206 52612 8258
rect 52556 8204 52612 8206
rect 52444 5628 52500 5684
rect 52332 5404 52388 5460
rect 52668 4956 52724 5012
rect 53004 9266 53060 9268
rect 53004 9214 53006 9266
rect 53006 9214 53058 9266
rect 53058 9214 53060 9266
rect 53004 9212 53060 9214
rect 53340 8370 53396 8372
rect 53340 8318 53342 8370
rect 53342 8318 53394 8370
rect 53394 8318 53396 8370
rect 53340 8316 53396 8318
rect 53564 10332 53620 10388
rect 53788 11900 53844 11956
rect 53564 8652 53620 8708
rect 53452 7980 53508 8036
rect 53004 7756 53060 7812
rect 52892 6972 52948 7028
rect 54236 13468 54292 13524
rect 54124 13020 54180 13076
rect 54908 13356 54964 13412
rect 55356 13244 55412 13300
rect 54908 13186 54964 13188
rect 54908 13134 54910 13186
rect 54910 13134 54962 13186
rect 54962 13134 54964 13186
rect 54908 13132 54964 13134
rect 55468 13020 55524 13076
rect 54460 11788 54516 11844
rect 54348 11116 54404 11172
rect 54236 10220 54292 10276
rect 54012 9212 54068 9268
rect 53900 8092 53956 8148
rect 53004 6130 53060 6132
rect 53004 6078 53006 6130
rect 53006 6078 53058 6130
rect 53058 6078 53060 6130
rect 53004 6076 53060 6078
rect 53564 5964 53620 6020
rect 54124 7420 54180 7476
rect 54124 5740 54180 5796
rect 52892 5234 52948 5236
rect 52892 5182 52894 5234
rect 52894 5182 52946 5234
rect 52946 5182 52948 5234
rect 52892 5180 52948 5182
rect 54124 5516 54180 5572
rect 53228 5122 53284 5124
rect 53228 5070 53230 5122
rect 53230 5070 53282 5122
rect 53282 5070 53284 5122
rect 53228 5068 53284 5070
rect 52892 4956 52948 5012
rect 52444 4844 52500 4900
rect 52220 4396 52276 4452
rect 52220 3052 52276 3108
rect 52108 2044 52164 2100
rect 52220 2380 52276 2436
rect 52108 1874 52164 1876
rect 52108 1822 52110 1874
rect 52110 1822 52162 1874
rect 52162 1822 52164 1874
rect 52108 1820 52164 1822
rect 51436 1708 51492 1764
rect 51100 1596 51156 1652
rect 51996 924 52052 980
rect 53676 5010 53732 5012
rect 53676 4958 53678 5010
rect 53678 4958 53730 5010
rect 53730 4958 53732 5010
rect 53676 4956 53732 4958
rect 53564 4620 53620 4676
rect 54348 8540 54404 8596
rect 54236 4284 54292 4340
rect 52556 3836 52612 3892
rect 53564 3612 53620 3668
rect 54572 10108 54628 10164
rect 54572 7196 54628 7252
rect 54572 5852 54628 5908
rect 55692 12402 55748 12404
rect 55692 12350 55694 12402
rect 55694 12350 55746 12402
rect 55746 12350 55748 12402
rect 55692 12348 55748 12350
rect 55804 11900 55860 11956
rect 55916 13916 55972 13972
rect 55468 11004 55524 11060
rect 55692 11228 55748 11284
rect 55580 10780 55636 10836
rect 54908 6412 54964 6468
rect 55468 10332 55524 10388
rect 55132 9436 55188 9492
rect 55132 8764 55188 8820
rect 55580 9884 55636 9940
rect 56252 12460 56308 12516
rect 55916 9324 55972 9380
rect 56028 12124 56084 12180
rect 55692 8316 55748 8372
rect 55916 8092 55972 8148
rect 56140 8988 56196 9044
rect 56028 7756 56084 7812
rect 56140 7698 56196 7700
rect 56140 7646 56142 7698
rect 56142 7646 56194 7698
rect 56194 7646 56196 7698
rect 56140 7644 56196 7646
rect 55132 7362 55188 7364
rect 55132 7310 55134 7362
rect 55134 7310 55186 7362
rect 55186 7310 55188 7362
rect 55132 7308 55188 7310
rect 56140 6748 56196 6804
rect 55132 6300 55188 6356
rect 56700 6076 56756 6132
rect 55020 5180 55076 5236
rect 54908 5122 54964 5124
rect 54908 5070 54910 5122
rect 54910 5070 54962 5122
rect 54962 5070 54964 5122
rect 54908 5068 54964 5070
rect 54796 4844 54852 4900
rect 54572 4562 54628 4564
rect 54572 4510 54574 4562
rect 54574 4510 54626 4562
rect 54626 4510 54628 4562
rect 54572 4508 54628 4510
rect 55132 3724 55188 3780
rect 54908 3666 54964 3668
rect 54908 3614 54910 3666
rect 54910 3614 54962 3666
rect 54962 3614 54964 3666
rect 54908 3612 54964 3614
rect 53564 3442 53620 3444
rect 53564 3390 53566 3442
rect 53566 3390 53618 3442
rect 53618 3390 53620 3442
rect 53564 3388 53620 3390
rect 54572 3164 54628 3220
rect 52444 2156 52500 2212
rect 52556 2940 52612 2996
rect 53564 2770 53620 2772
rect 53564 2718 53566 2770
rect 53566 2718 53618 2770
rect 53618 2718 53620 2770
rect 53564 2716 53620 2718
rect 52780 2658 52836 2660
rect 52780 2606 52782 2658
rect 52782 2606 52834 2658
rect 52834 2606 52836 2658
rect 52780 2604 52836 2606
rect 54124 2492 54180 2548
rect 54908 2268 54964 2324
rect 53564 1874 53620 1876
rect 53564 1822 53566 1874
rect 53566 1822 53618 1874
rect 53618 1822 53620 1874
rect 53564 1820 53620 1822
rect 56140 5404 56196 5460
rect 55244 2380 55300 2436
rect 55356 4732 55412 4788
rect 55132 1484 55188 1540
rect 53564 1426 53620 1428
rect 53564 1374 53566 1426
rect 53566 1374 53618 1426
rect 53618 1374 53620 1426
rect 53564 1372 53620 1374
rect 52332 1148 52388 1204
rect 52556 1260 52612 1316
rect 56140 4060 56196 4116
rect 56812 3388 56868 3444
rect 56140 2716 56196 2772
rect 56476 2604 56532 2660
rect 52220 476 52276 532
rect 52892 812 52948 868
rect 49420 140 49476 196
rect 50204 140 50260 196
rect 55580 700 55636 756
rect 21308 28 21364 84
rect 56812 476 56868 532
rect 56476 28 56532 84
<< metal3 >>
rect 10210 14140 10220 14196
rect 10276 14140 20972 14196
rect 21028 14140 21038 14196
rect 21186 14140 21196 14196
rect 21252 14140 29484 14196
rect 29540 14140 29550 14196
rect 29708 14140 31836 14196
rect 31892 14140 31902 14196
rect 32050 14140 32060 14196
rect 32116 14140 35420 14196
rect 35476 14140 35486 14196
rect 29708 14084 29764 14140
rect 8978 14028 8988 14084
rect 9044 14028 29764 14084
rect 30706 14028 30716 14084
rect 30772 14028 45724 14084
rect 45780 14028 45790 14084
rect 0 13972 112 14000
rect 57344 13972 57456 14000
rect 0 13916 1484 13972
rect 1540 13916 1550 13972
rect 3154 13916 3164 13972
rect 3220 13916 18284 13972
rect 18340 13916 18350 13972
rect 20962 13916 20972 13972
rect 21028 13916 27804 13972
rect 27860 13916 27870 13972
rect 28914 13916 28924 13972
rect 28980 13916 43596 13972
rect 43652 13916 43662 13972
rect 55906 13916 55916 13972
rect 55972 13916 57456 13972
rect 0 13888 112 13916
rect 57344 13888 57456 13916
rect 12226 13804 12236 13860
rect 12292 13804 13748 13860
rect 15250 13804 15260 13860
rect 15316 13804 24892 13860
rect 24948 13804 24958 13860
rect 25778 13804 25788 13860
rect 25844 13804 33964 13860
rect 34020 13804 34030 13860
rect 35410 13804 35420 13860
rect 35476 13804 44604 13860
rect 44660 13804 44670 13860
rect 6626 13692 6636 13748
rect 6692 13692 13636 13748
rect 0 13524 112 13552
rect 13580 13524 13636 13692
rect 13692 13636 13748 13804
rect 15138 13692 15148 13748
rect 15204 13692 25116 13748
rect 25172 13692 25182 13748
rect 27682 13692 27692 13748
rect 27748 13692 30156 13748
rect 30212 13692 30222 13748
rect 30370 13692 30380 13748
rect 30436 13692 36316 13748
rect 36372 13692 36382 13748
rect 13692 13580 20972 13636
rect 21028 13580 21038 13636
rect 24210 13580 24220 13636
rect 24276 13580 25676 13636
rect 25732 13580 25742 13636
rect 25890 13580 25900 13636
rect 25956 13580 34748 13636
rect 34804 13580 34814 13636
rect 35074 13580 35084 13636
rect 35140 13580 43708 13636
rect 43764 13580 43774 13636
rect 49074 13580 49084 13636
rect 49140 13580 51100 13636
rect 51156 13580 51166 13636
rect 57344 13524 57456 13552
rect 0 13468 1596 13524
rect 1652 13468 1662 13524
rect 3602 13468 3612 13524
rect 3668 13468 4732 13524
rect 4788 13468 4798 13524
rect 10770 13468 10780 13524
rect 10836 13468 13524 13524
rect 13580 13468 15820 13524
rect 15876 13468 15886 13524
rect 18386 13468 18396 13524
rect 18452 13468 26348 13524
rect 26404 13468 26414 13524
rect 26852 13468 31164 13524
rect 31220 13468 31230 13524
rect 31378 13468 31388 13524
rect 31444 13468 39676 13524
rect 39732 13468 39742 13524
rect 49970 13468 49980 13524
rect 50036 13468 52892 13524
rect 52948 13468 52958 13524
rect 54226 13468 54236 13524
rect 54292 13468 57456 13524
rect 0 13440 112 13468
rect 13468 13412 13524 13468
rect 26852 13412 26908 13468
rect 57344 13440 57456 13468
rect 2146 13356 2156 13412
rect 2212 13356 4284 13412
rect 4340 13356 4350 13412
rect 11330 13356 11340 13412
rect 11396 13356 13244 13412
rect 13300 13356 13310 13412
rect 13468 13356 23436 13412
rect 23492 13356 23502 13412
rect 24994 13356 25004 13412
rect 25060 13356 26908 13412
rect 27020 13356 29484 13412
rect 29540 13356 29550 13412
rect 29810 13356 29820 13412
rect 29876 13356 34076 13412
rect 34132 13356 34142 13412
rect 47842 13356 47852 13412
rect 47908 13356 54908 13412
rect 54964 13356 54974 13412
rect 4454 13300 4464 13356
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4728 13300 4738 13356
rect 24454 13300 24464 13356
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24728 13300 24738 13356
rect 27020 13300 27076 13356
rect 44454 13300 44464 13356
rect 44520 13300 44568 13356
rect 44624 13300 44672 13356
rect 44728 13300 44738 13356
rect 5954 13244 5964 13300
rect 6020 13244 7420 13300
rect 7476 13244 7486 13300
rect 10322 13244 10332 13300
rect 10388 13244 18396 13300
rect 18452 13244 18462 13300
rect 18610 13244 18620 13300
rect 18676 13244 24332 13300
rect 24388 13244 24398 13300
rect 26226 13244 26236 13300
rect 26292 13244 27076 13300
rect 27234 13244 27244 13300
rect 27300 13244 37324 13300
rect 37380 13244 37390 13300
rect 38770 13244 38780 13300
rect 38836 13244 39340 13300
rect 39396 13244 39406 13300
rect 50372 13244 55356 13300
rect 55412 13244 55422 13300
rect 3714 13132 3724 13188
rect 3780 13132 5628 13188
rect 5684 13132 5694 13188
rect 7522 13132 7532 13188
rect 7588 13132 9212 13188
rect 9268 13132 9278 13188
rect 9762 13132 9772 13188
rect 9828 13132 11452 13188
rect 11508 13132 11518 13188
rect 12674 13132 12684 13188
rect 12740 13132 19852 13188
rect 19908 13132 19918 13188
rect 21186 13132 21196 13188
rect 21252 13132 21756 13188
rect 21812 13132 21822 13188
rect 21980 13132 23660 13188
rect 23716 13132 23726 13188
rect 23986 13132 23996 13188
rect 24052 13132 25508 13188
rect 25778 13132 25788 13188
rect 25844 13132 32788 13188
rect 33282 13132 33292 13188
rect 33348 13132 41468 13188
rect 41524 13132 41534 13188
rect 44146 13132 44156 13188
rect 44212 13132 46844 13188
rect 46900 13132 46910 13188
rect 48178 13132 48188 13188
rect 48244 13132 48972 13188
rect 49028 13132 49038 13188
rect 0 13076 112 13104
rect 21980 13076 22036 13132
rect 25452 13076 25508 13132
rect 0 13020 364 13076
rect 420 13020 430 13076
rect 8082 13020 8092 13076
rect 8148 13020 11564 13076
rect 11620 13020 11630 13076
rect 13682 13020 13692 13076
rect 13748 13020 14588 13076
rect 14644 13020 14654 13076
rect 14914 13020 14924 13076
rect 14980 13020 16380 13076
rect 16436 13020 16446 13076
rect 17490 13020 17500 13076
rect 17556 13020 18620 13076
rect 18676 13020 18686 13076
rect 18946 13020 18956 13076
rect 19012 13020 22036 13076
rect 23538 13020 23548 13076
rect 23604 13020 24108 13076
rect 24164 13020 24174 13076
rect 24546 13020 24556 13076
rect 24612 13020 25172 13076
rect 25442 13020 25452 13076
rect 25508 13020 25518 13076
rect 25676 13020 31052 13076
rect 31108 13020 31118 13076
rect 31826 13020 31836 13076
rect 31892 13020 32508 13076
rect 32564 13020 32574 13076
rect 0 12992 112 13020
rect 25116 12964 25172 13020
rect 25676 12964 25732 13020
rect 32732 12964 32788 13132
rect 50372 13076 50428 13244
rect 52210 13132 52220 13188
rect 52276 13132 54908 13188
rect 54964 13132 54974 13188
rect 57344 13076 57456 13104
rect 33618 13020 33628 13076
rect 33684 13020 41020 13076
rect 41076 13020 41086 13076
rect 47954 13020 47964 13076
rect 48020 13020 50428 13076
rect 51762 13020 51772 13076
rect 51828 13020 54124 13076
rect 54180 13020 54190 13076
rect 55458 13020 55468 13076
rect 55524 13020 57456 13076
rect 57344 12992 57456 13020
rect 4274 12908 4284 12964
rect 4340 12908 4956 12964
rect 5012 12908 5022 12964
rect 6514 12908 6524 12964
rect 6580 12908 9212 12964
rect 9268 12908 9278 12964
rect 9426 12908 9436 12964
rect 9492 12908 12908 12964
rect 12964 12908 12974 12964
rect 15092 12908 18844 12964
rect 18900 12908 18910 12964
rect 21746 12908 21756 12964
rect 21812 12908 24892 12964
rect 24948 12908 24958 12964
rect 25116 12908 25732 12964
rect 26002 12908 26012 12964
rect 26068 12908 32676 12964
rect 32732 12908 40068 12964
rect 40226 12908 40236 12964
rect 40292 12908 44940 12964
rect 44996 12908 45006 12964
rect 45490 12908 45500 12964
rect 45556 12908 46844 12964
rect 46900 12908 46910 12964
rect 15092 12852 15148 12908
rect 32620 12852 32676 12908
rect 40012 12852 40068 12908
rect 5954 12796 5964 12852
rect 6020 12796 15148 12852
rect 16930 12796 16940 12852
rect 16996 12796 18620 12852
rect 18676 12796 18686 12852
rect 19282 12796 19292 12852
rect 19348 12796 19964 12852
rect 20020 12796 20030 12852
rect 20860 12796 28700 12852
rect 28756 12796 28766 12852
rect 29474 12796 29484 12852
rect 29540 12796 30940 12852
rect 30996 12796 31006 12852
rect 31154 12796 31164 12852
rect 31220 12796 31836 12852
rect 31892 12796 31902 12852
rect 32620 12796 32956 12852
rect 33012 12796 33022 12852
rect 33170 12796 33180 12852
rect 33236 12796 39788 12852
rect 39844 12796 39854 12852
rect 40012 12796 45388 12852
rect 45444 12796 45454 12852
rect 20860 12740 20916 12796
rect 9538 12684 9548 12740
rect 9604 12684 17948 12740
rect 18004 12684 18014 12740
rect 19730 12684 19740 12740
rect 19796 12684 20916 12740
rect 22418 12684 22428 12740
rect 22484 12684 24276 12740
rect 24882 12684 24892 12740
rect 24948 12684 34300 12740
rect 34356 12684 34366 12740
rect 36194 12684 36204 12740
rect 36260 12684 38556 12740
rect 38612 12684 38622 12740
rect 38882 12684 38892 12740
rect 38948 12684 42140 12740
rect 42196 12684 42206 12740
rect 0 12628 112 12656
rect 24220 12628 24276 12684
rect 57344 12628 57456 12656
rect 0 12572 924 12628
rect 980 12572 990 12628
rect 9314 12572 9324 12628
rect 9380 12572 20300 12628
rect 20356 12572 20636 12628
rect 20692 12572 20702 12628
rect 24220 12572 27132 12628
rect 27188 12572 27198 12628
rect 27906 12572 27916 12628
rect 27972 12572 28924 12628
rect 28980 12572 28990 12628
rect 29250 12572 29260 12628
rect 29316 12572 42364 12628
rect 42420 12572 42430 12628
rect 53890 12572 53900 12628
rect 53956 12572 57456 12628
rect 0 12544 112 12572
rect 3794 12516 3804 12572
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 4068 12516 4078 12572
rect 23794 12516 23804 12572
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 24068 12516 24078 12572
rect 43794 12516 43804 12572
rect 43860 12516 43908 12572
rect 43964 12516 44012 12572
rect 44068 12516 44078 12572
rect 57344 12544 57456 12572
rect 8642 12460 8652 12516
rect 8708 12460 13580 12516
rect 13636 12460 13646 12516
rect 14242 12460 14252 12516
rect 14308 12460 16940 12516
rect 16996 12460 17006 12516
rect 18722 12460 18732 12516
rect 18788 12460 22092 12516
rect 22148 12460 22158 12516
rect 24994 12460 25004 12516
rect 25060 12460 28140 12516
rect 28196 12460 28206 12516
rect 30258 12460 30268 12516
rect 30324 12460 36764 12516
rect 36820 12460 36830 12516
rect 38770 12460 38780 12516
rect 38836 12460 38846 12516
rect 39778 12460 39788 12516
rect 39844 12460 43484 12516
rect 43540 12460 43550 12516
rect 45938 12460 45948 12516
rect 46004 12460 56252 12516
rect 56308 12460 56318 12516
rect 38780 12404 38836 12460
rect 2258 12348 2268 12404
rect 2324 12348 3388 12404
rect 3444 12348 3454 12404
rect 6962 12348 6972 12404
rect 7028 12348 7868 12404
rect 7924 12348 7934 12404
rect 8530 12348 8540 12404
rect 8596 12348 9660 12404
rect 9716 12348 9726 12404
rect 10658 12348 10668 12404
rect 10724 12348 13804 12404
rect 13860 12348 13870 12404
rect 14018 12348 14028 12404
rect 14084 12348 21196 12404
rect 21252 12348 21262 12404
rect 23090 12348 23100 12404
rect 23156 12348 23884 12404
rect 23940 12348 23950 12404
rect 24210 12348 24220 12404
rect 24276 12348 28028 12404
rect 28084 12348 28094 12404
rect 28242 12348 28252 12404
rect 28308 12348 36092 12404
rect 36148 12348 36158 12404
rect 36306 12348 36316 12404
rect 36372 12348 38836 12404
rect 38994 12348 39004 12404
rect 39060 12348 47852 12404
rect 47908 12348 47918 12404
rect 48626 12348 48636 12404
rect 48692 12348 49420 12404
rect 49476 12348 49486 12404
rect 50418 12348 50428 12404
rect 50484 12348 52556 12404
rect 52612 12348 52622 12404
rect 53106 12348 53116 12404
rect 53172 12348 55692 12404
rect 55748 12348 55758 12404
rect 6412 12236 11116 12292
rect 11172 12236 11182 12292
rect 13346 12236 13356 12292
rect 13412 12236 13692 12292
rect 13748 12236 15708 12292
rect 15764 12236 15774 12292
rect 16146 12236 16156 12292
rect 16212 12236 17164 12292
rect 17220 12236 17230 12292
rect 17714 12236 17724 12292
rect 17780 12236 18620 12292
rect 18676 12236 18686 12292
rect 20178 12236 20188 12292
rect 20244 12236 28364 12292
rect 28420 12236 28430 12292
rect 28578 12236 28588 12292
rect 28644 12236 34860 12292
rect 34916 12236 34926 12292
rect 37090 12236 37100 12292
rect 37156 12236 42812 12292
rect 42868 12236 42878 12292
rect 43474 12236 43484 12292
rect 43540 12236 44492 12292
rect 44548 12236 44558 12292
rect 45266 12236 45276 12292
rect 45332 12236 48076 12292
rect 48132 12236 48142 12292
rect 0 12180 112 12208
rect 0 12124 1036 12180
rect 1092 12124 1102 12180
rect 2930 12124 2940 12180
rect 2996 12124 3388 12180
rect 3444 12124 3454 12180
rect 0 12096 112 12124
rect 6412 12068 6468 12236
rect 57344 12180 57456 12208
rect 7522 12124 7532 12180
rect 7588 12124 12012 12180
rect 12068 12124 12078 12180
rect 13458 12124 13468 12180
rect 13524 12124 14028 12180
rect 14084 12124 14094 12180
rect 16258 12124 16268 12180
rect 16324 12124 17276 12180
rect 17332 12124 17342 12180
rect 17490 12124 17500 12180
rect 17556 12124 23604 12180
rect 23762 12124 23772 12180
rect 23828 12124 31836 12180
rect 31892 12124 31902 12180
rect 32274 12124 32284 12180
rect 32340 12124 35644 12180
rect 35700 12124 35710 12180
rect 35970 12124 35980 12180
rect 36036 12124 39340 12180
rect 39396 12124 39406 12180
rect 43026 12124 43036 12180
rect 43092 12124 46956 12180
rect 47012 12124 47022 12180
rect 56018 12124 56028 12180
rect 56084 12124 57456 12180
rect 23548 12068 23604 12124
rect 57344 12096 57456 12124
rect 242 12012 252 12068
rect 308 12012 6468 12068
rect 6626 12012 6636 12068
rect 6692 12012 13692 12068
rect 13748 12012 13758 12068
rect 15362 12012 15372 12068
rect 15428 12012 16940 12068
rect 16996 12012 17006 12068
rect 19282 12012 19292 12068
rect 19348 12012 23324 12068
rect 23380 12012 23390 12068
rect 23548 12012 30156 12068
rect 30212 12012 30222 12068
rect 31042 12012 31052 12068
rect 31108 12012 33404 12068
rect 33460 12012 33470 12068
rect 33730 12012 33740 12068
rect 33796 12012 36316 12068
rect 36372 12012 36382 12068
rect 38322 12012 38332 12068
rect 38388 12012 46060 12068
rect 46116 12012 46508 12068
rect 46564 12012 46574 12068
rect 46722 12012 46732 12068
rect 46788 12012 50988 12068
rect 51044 12012 51054 12068
rect 1586 11900 1596 11956
rect 1652 11900 8988 11956
rect 9044 11900 9054 11956
rect 10098 11900 10108 11956
rect 10164 11900 15148 11956
rect 15204 11900 15214 11956
rect 15474 11900 15484 11956
rect 15540 11900 27356 11956
rect 27412 11900 27422 11956
rect 27570 11900 27580 11956
rect 27636 11900 31724 11956
rect 31780 11900 31790 11956
rect 32498 11900 32508 11956
rect 32564 11900 34524 11956
rect 34580 11900 34590 11956
rect 34738 11900 34748 11956
rect 34804 11900 38220 11956
rect 38276 11900 38286 11956
rect 38770 11900 38780 11956
rect 38836 11900 49644 11956
rect 49700 11900 49710 11956
rect 53778 11900 53788 11956
rect 53844 11900 55804 11956
rect 55860 11900 55870 11956
rect 1138 11788 1148 11844
rect 1204 11788 2268 11844
rect 2324 11788 2334 11844
rect 5954 11788 5964 11844
rect 6020 11788 6524 11844
rect 6580 11788 6590 11844
rect 8372 11788 15148 11844
rect 15204 11788 15214 11844
rect 15362 11788 15372 11844
rect 15428 11788 17108 11844
rect 17714 11788 17724 11844
rect 17780 11788 21756 11844
rect 21812 11788 21822 11844
rect 22082 11788 22092 11844
rect 22148 11788 24332 11844
rect 24388 11788 24398 11844
rect 28018 11788 28028 11844
rect 28084 11788 30716 11844
rect 30772 11788 30782 11844
rect 30930 11788 30940 11844
rect 30996 11788 32844 11844
rect 32900 11788 32910 11844
rect 33058 11788 33068 11844
rect 33124 11788 33852 11844
rect 33908 11788 33918 11844
rect 35634 11788 35644 11844
rect 35700 11788 37884 11844
rect 37940 11788 37950 11844
rect 38612 11788 41972 11844
rect 45602 11788 45612 11844
rect 45668 11788 48412 11844
rect 48468 11788 48478 11844
rect 51202 11788 51212 11844
rect 51268 11788 54460 11844
rect 54516 11788 54526 11844
rect 0 11732 112 11760
rect 4454 11732 4464 11788
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4728 11732 4738 11788
rect 0 11676 4284 11732
rect 4340 11676 4350 11732
rect 0 11648 112 11676
rect 3332 11564 4452 11620
rect 4610 11564 4620 11620
rect 4676 11564 5068 11620
rect 5124 11564 5134 11620
rect 3332 11508 3388 11564
rect 2034 11452 2044 11508
rect 2100 11452 3388 11508
rect 4396 11508 4452 11564
rect 8372 11508 8428 11788
rect 13570 11676 13580 11732
rect 13636 11676 16828 11732
rect 16884 11676 16894 11732
rect 17052 11620 17108 11788
rect 24454 11732 24464 11788
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24728 11732 24738 11788
rect 38612 11732 38668 11788
rect 41916 11732 41972 11788
rect 44454 11732 44464 11788
rect 44520 11732 44568 11788
rect 44624 11732 44672 11788
rect 44728 11732 44738 11788
rect 57344 11732 57456 11760
rect 17938 11676 17948 11732
rect 18004 11676 21084 11732
rect 21140 11676 21150 11732
rect 21522 11676 21532 11732
rect 21588 11676 24220 11732
rect 24276 11676 24286 11732
rect 24882 11676 24892 11732
rect 24948 11676 28588 11732
rect 28644 11676 28654 11732
rect 30146 11676 30156 11732
rect 30212 11676 38668 11732
rect 38882 11676 38892 11732
rect 38948 11676 41692 11732
rect 41748 11676 41758 11732
rect 41916 11676 44268 11732
rect 44324 11676 44334 11732
rect 45714 11676 45724 11732
rect 45780 11676 51100 11732
rect 51156 11676 51166 11732
rect 51314 11676 51324 11732
rect 51380 11676 52556 11732
rect 52612 11676 52622 11732
rect 53900 11676 57456 11732
rect 14578 11564 14588 11620
rect 14644 11564 15484 11620
rect 15540 11564 15550 11620
rect 17052 11564 18788 11620
rect 19058 11564 19068 11620
rect 19124 11564 21644 11620
rect 21700 11564 21710 11620
rect 21970 11564 21980 11620
rect 22036 11564 25900 11620
rect 25956 11564 25966 11620
rect 26114 11564 26124 11620
rect 26180 11564 31500 11620
rect 31556 11564 31566 11620
rect 31826 11564 31836 11620
rect 31892 11564 33180 11620
rect 33236 11564 33246 11620
rect 33394 11564 33404 11620
rect 33460 11564 36652 11620
rect 36708 11564 36718 11620
rect 40338 11564 40348 11620
rect 40404 11564 43260 11620
rect 43316 11564 43326 11620
rect 43474 11564 43484 11620
rect 43540 11564 45948 11620
rect 46004 11564 46014 11620
rect 49522 11564 49532 11620
rect 49588 11564 50316 11620
rect 50372 11564 50382 11620
rect 50866 11564 50876 11620
rect 50932 11564 51884 11620
rect 51940 11564 51950 11620
rect 18732 11508 18788 11564
rect 53900 11508 53956 11676
rect 57344 11648 57456 11676
rect 4396 11452 8428 11508
rect 9202 11452 9212 11508
rect 9268 11452 14700 11508
rect 14756 11452 14766 11508
rect 14924 11452 18508 11508
rect 18564 11452 18574 11508
rect 18732 11452 34188 11508
rect 34244 11452 34254 11508
rect 34748 11452 44044 11508
rect 44100 11452 44110 11508
rect 44258 11452 44268 11508
rect 44324 11452 49756 11508
rect 49812 11452 49822 11508
rect 50372 11452 53956 11508
rect 14924 11396 14980 11452
rect 34748 11396 34804 11452
rect 50372 11396 50428 11452
rect 4274 11340 4284 11396
rect 4340 11340 10108 11396
rect 10164 11340 10174 11396
rect 10322 11340 10332 11396
rect 10388 11340 14980 11396
rect 15138 11340 15148 11396
rect 15204 11340 20188 11396
rect 20244 11340 20254 11396
rect 20402 11340 20412 11396
rect 20468 11340 26124 11396
rect 26180 11340 26190 11396
rect 26852 11340 34804 11396
rect 34962 11340 34972 11396
rect 35028 11340 48188 11396
rect 48244 11340 48254 11396
rect 49186 11340 49196 11396
rect 49252 11340 50428 11396
rect 0 11284 112 11312
rect 26852 11284 26908 11340
rect 57344 11284 57456 11312
rect 0 11228 9268 11284
rect 10098 11228 10108 11284
rect 10164 11228 17052 11284
rect 17108 11228 17118 11284
rect 19618 11228 19628 11284
rect 19684 11228 26908 11284
rect 27794 11228 27804 11284
rect 27860 11228 33628 11284
rect 33684 11228 33694 11284
rect 33842 11228 33852 11284
rect 33908 11228 38332 11284
rect 38388 11228 38398 11284
rect 39666 11228 39676 11284
rect 39732 11228 44156 11284
rect 44212 11228 44222 11284
rect 55682 11228 55692 11284
rect 55748 11228 57456 11284
rect 0 11200 112 11228
rect 9212 11172 9268 11228
rect 57344 11200 57456 11228
rect 3602 11116 3612 11172
rect 3668 11116 6636 11172
rect 6692 11116 6702 11172
rect 9212 11116 14924 11172
rect 14980 11116 14990 11172
rect 15138 11116 15148 11172
rect 15204 11116 20412 11172
rect 20468 11116 20478 11172
rect 20626 11116 20636 11172
rect 20692 11116 21532 11172
rect 21588 11116 21598 11172
rect 22082 11116 22092 11172
rect 22148 11116 23996 11172
rect 24052 11116 24556 11172
rect 24612 11116 24622 11172
rect 27346 11116 27356 11172
rect 27412 11116 29148 11172
rect 29204 11116 29214 11172
rect 29362 11116 29372 11172
rect 29428 11116 34300 11172
rect 34356 11116 34366 11172
rect 36754 11116 36764 11172
rect 36820 11116 38892 11172
rect 38948 11116 38958 11172
rect 39116 11116 41804 11172
rect 41860 11116 41870 11172
rect 44034 11116 44044 11172
rect 44100 11116 54348 11172
rect 54404 11116 54414 11172
rect 39116 11060 39172 11116
rect 10220 11004 19068 11060
rect 19124 11004 19134 11060
rect 20402 11004 20412 11060
rect 20468 11004 22092 11060
rect 22148 11004 22158 11060
rect 24220 11004 28252 11060
rect 28308 11004 28318 11060
rect 28690 11004 28700 11060
rect 28756 11004 30828 11060
rect 30884 11004 30894 11060
rect 31042 11004 31052 11060
rect 31108 11004 39172 11060
rect 39330 11004 39340 11060
rect 39396 11004 41916 11060
rect 41972 11004 41982 11060
rect 49634 11004 49644 11060
rect 49700 11004 55468 11060
rect 55524 11004 55534 11060
rect 3794 10948 3804 11004
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 4068 10948 4078 11004
rect 0 10836 112 10864
rect 10220 10836 10276 11004
rect 23794 10948 23804 11004
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 24068 10948 24078 11004
rect 0 10780 812 10836
rect 868 10780 878 10836
rect 1026 10780 1036 10836
rect 1092 10780 10276 10836
rect 10332 10892 17948 10948
rect 18004 10892 18014 10948
rect 18162 10892 18172 10948
rect 18228 10892 21924 10948
rect 0 10752 112 10780
rect 2370 10668 2380 10724
rect 2436 10668 8540 10724
rect 8596 10668 8606 10724
rect 10332 10612 10388 10892
rect 21868 10836 21924 10892
rect 24220 10836 24276 11004
rect 43794 10948 43804 11004
rect 43860 10948 43908 11004
rect 43964 10948 44012 11004
rect 44068 10948 44078 11004
rect 24434 10892 24444 10948
rect 24500 10892 26572 10948
rect 26628 10892 26638 10948
rect 26898 10892 26908 10948
rect 26964 10892 30156 10948
rect 30212 10892 30222 10948
rect 30370 10892 30380 10948
rect 30436 10892 33964 10948
rect 34020 10892 34030 10948
rect 34188 10892 40236 10948
rect 40292 10892 40302 10948
rect 34188 10836 34244 10892
rect 57344 10836 57456 10864
rect 14130 10780 14140 10836
rect 14196 10780 14588 10836
rect 14644 10780 14654 10836
rect 15922 10780 15932 10836
rect 15988 10780 16716 10836
rect 16772 10780 16782 10836
rect 17826 10780 17836 10836
rect 17892 10780 20636 10836
rect 20692 10780 20702 10836
rect 20850 10780 20860 10836
rect 20916 10780 21644 10836
rect 21700 10780 21710 10836
rect 21868 10780 24276 10836
rect 24994 10780 25004 10836
rect 25060 10780 32060 10836
rect 32116 10780 32126 10836
rect 32722 10780 32732 10836
rect 32788 10780 34244 10836
rect 34300 10780 39340 10836
rect 39396 10780 39406 10836
rect 39554 10780 39564 10836
rect 39620 10780 40572 10836
rect 40628 10780 40638 10836
rect 43698 10780 43708 10836
rect 43764 10780 46956 10836
rect 47012 10780 47022 10836
rect 55570 10780 55580 10836
rect 55636 10780 57456 10836
rect 34300 10724 34356 10780
rect 57344 10752 57456 10780
rect 12562 10668 12572 10724
rect 12628 10668 16156 10724
rect 16212 10668 16222 10724
rect 18050 10668 18060 10724
rect 18116 10668 21868 10724
rect 21924 10668 21934 10724
rect 22082 10668 22092 10724
rect 22148 10668 27132 10724
rect 27188 10668 27198 10724
rect 28242 10668 28252 10724
rect 28308 10668 31052 10724
rect 31108 10668 31118 10724
rect 31266 10668 31276 10724
rect 31332 10668 31388 10724
rect 31444 10668 31454 10724
rect 31826 10668 31836 10724
rect 31892 10668 33236 10724
rect 34066 10668 34076 10724
rect 34132 10668 34356 10724
rect 37090 10668 37100 10724
rect 37156 10668 50204 10724
rect 50260 10668 50270 10724
rect 33180 10612 33236 10668
rect 2482 10556 2492 10612
rect 2548 10556 10388 10612
rect 10444 10556 26460 10612
rect 26516 10556 26526 10612
rect 26786 10556 26796 10612
rect 26852 10556 32956 10612
rect 33012 10556 33022 10612
rect 33180 10556 39676 10612
rect 39732 10556 39742 10612
rect 39900 10556 42028 10612
rect 42084 10556 42252 10612
rect 42308 10556 42318 10612
rect 42690 10556 42700 10612
rect 42756 10556 47572 10612
rect 47730 10556 47740 10612
rect 47796 10556 52108 10612
rect 52164 10556 52174 10612
rect 2930 10444 2940 10500
rect 2996 10444 9212 10500
rect 9268 10444 9278 10500
rect 0 10388 112 10416
rect 10444 10388 10500 10556
rect 39900 10500 39956 10556
rect 47516 10500 47572 10556
rect 11554 10444 11564 10500
rect 11620 10444 20300 10500
rect 20356 10444 20366 10500
rect 22306 10444 22316 10500
rect 22372 10444 27356 10500
rect 27412 10444 27422 10500
rect 30258 10444 30268 10500
rect 30324 10444 32732 10500
rect 32788 10444 32798 10500
rect 33618 10444 33628 10500
rect 33684 10444 39956 10500
rect 40226 10444 40236 10500
rect 40292 10444 41132 10500
rect 41188 10444 41356 10500
rect 41412 10444 41422 10500
rect 41906 10444 41916 10500
rect 41972 10444 47292 10500
rect 47348 10444 47358 10500
rect 47516 10444 50988 10500
rect 51044 10444 51054 10500
rect 57344 10388 57456 10416
rect 0 10332 1036 10388
rect 1092 10332 1102 10388
rect 1586 10332 1596 10388
rect 1652 10332 7308 10388
rect 7364 10332 7374 10388
rect 7522 10332 7532 10388
rect 7588 10332 10500 10388
rect 13794 10332 13804 10388
rect 13860 10332 16604 10388
rect 16660 10332 16670 10388
rect 16818 10332 16828 10388
rect 16884 10332 19740 10388
rect 19796 10332 19806 10388
rect 20066 10332 20076 10388
rect 20132 10332 20636 10388
rect 20692 10332 21756 10388
rect 21812 10332 21822 10388
rect 22194 10332 22204 10388
rect 22260 10332 26852 10388
rect 26908 10332 26918 10388
rect 27010 10332 27020 10388
rect 27076 10332 39564 10388
rect 39620 10332 39630 10388
rect 40226 10332 40236 10388
rect 40292 10332 49420 10388
rect 49476 10332 49486 10388
rect 49644 10332 53564 10388
rect 53620 10332 53630 10388
rect 55458 10332 55468 10388
rect 55524 10332 57456 10388
rect 0 10304 112 10332
rect 49644 10276 49700 10332
rect 57344 10304 57456 10332
rect 6962 10220 6972 10276
rect 7028 10220 10332 10276
rect 10388 10220 10398 10276
rect 11106 10220 11116 10276
rect 11172 10220 13244 10276
rect 13300 10220 13310 10276
rect 13682 10220 13692 10276
rect 13748 10220 19964 10276
rect 20020 10220 20030 10276
rect 20178 10220 20188 10276
rect 20244 10220 21980 10276
rect 22036 10220 22046 10276
rect 26338 10220 26348 10276
rect 26404 10220 27916 10276
rect 27972 10220 27982 10276
rect 28140 10220 33740 10276
rect 33796 10220 33806 10276
rect 33954 10220 33964 10276
rect 34020 10220 41972 10276
rect 42130 10220 42140 10276
rect 42196 10220 44268 10276
rect 44324 10220 44334 10276
rect 47954 10220 47964 10276
rect 48020 10220 49700 10276
rect 50194 10220 50204 10276
rect 50260 10220 54236 10276
rect 54292 10220 54302 10276
rect 4454 10164 4464 10220
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4728 10164 4738 10220
rect 24454 10164 24464 10220
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24728 10164 24738 10220
rect 4844 10108 9324 10164
rect 9380 10108 9390 10164
rect 9986 10108 9996 10164
rect 10052 10108 12460 10164
rect 12516 10108 12526 10164
rect 14018 10108 14028 10164
rect 14084 10108 16716 10164
rect 16772 10108 16782 10164
rect 17154 10108 17164 10164
rect 17220 10108 20076 10164
rect 20132 10108 20142 10164
rect 20290 10108 20300 10164
rect 20356 10108 24220 10164
rect 24276 10108 24286 10164
rect 26002 10108 26012 10164
rect 26068 10108 27916 10164
rect 27972 10108 27982 10164
rect 4844 10052 4900 10108
rect 28140 10052 28196 10220
rect 28914 10108 28924 10164
rect 28980 10108 31836 10164
rect 31892 10108 31902 10164
rect 32050 10108 32060 10164
rect 32116 10108 35196 10164
rect 35252 10108 35262 10164
rect 35634 10108 35644 10164
rect 35700 10108 38108 10164
rect 38164 10108 38174 10164
rect 38612 10108 41132 10164
rect 41188 10108 41468 10164
rect 41524 10108 41534 10164
rect 38612 10052 38668 10108
rect 1596 9996 4900 10052
rect 5730 9996 5740 10052
rect 5796 9996 14252 10052
rect 14308 9996 14318 10052
rect 14466 9996 14476 10052
rect 14532 9996 18172 10052
rect 18228 9996 18238 10052
rect 18386 9996 18396 10052
rect 18452 9996 22092 10052
rect 22148 9996 22158 10052
rect 22754 9996 22764 10052
rect 22820 9996 28196 10052
rect 28578 9996 28588 10052
rect 28644 9996 31388 10052
rect 31444 9996 31454 10052
rect 31602 9996 31612 10052
rect 31668 9996 35868 10052
rect 35924 9996 36092 10052
rect 36148 9996 36158 10052
rect 37314 9996 37324 10052
rect 37380 9996 38668 10052
rect 41916 10052 41972 10220
rect 44454 10164 44464 10220
rect 44520 10164 44568 10220
rect 44624 10164 44672 10220
rect 44728 10164 44738 10220
rect 47068 10108 47404 10164
rect 47460 10108 47470 10164
rect 48066 10108 48076 10164
rect 48132 10108 49532 10164
rect 49588 10108 49598 10164
rect 54562 10108 54572 10164
rect 54628 10108 55860 10164
rect 47068 10052 47124 10108
rect 41916 9996 47124 10052
rect 0 9940 112 9968
rect 1596 9940 1652 9996
rect 55804 9940 55860 10108
rect 57344 9940 57456 9968
rect 0 9884 1652 9940
rect 1708 9884 10108 9940
rect 10164 9884 10174 9940
rect 12450 9884 12460 9940
rect 12516 9884 15260 9940
rect 15316 9884 15326 9940
rect 15810 9884 15820 9940
rect 15876 9884 18732 9940
rect 18788 9884 18798 9940
rect 21634 9884 21644 9940
rect 21700 9884 25004 9940
rect 25060 9884 25070 9940
rect 25218 9884 25228 9940
rect 25284 9884 33628 9940
rect 33684 9884 33694 9940
rect 34066 9884 34076 9940
rect 34132 9884 37212 9940
rect 37268 9884 37278 9940
rect 37436 9884 40236 9940
rect 40292 9884 40302 9940
rect 41794 9884 41804 9940
rect 41860 9884 47180 9940
rect 47236 9884 47246 9940
rect 51762 9884 51772 9940
rect 51828 9884 55580 9940
rect 55636 9884 55646 9940
rect 55804 9884 57456 9940
rect 0 9856 112 9884
rect 1708 9828 1764 9884
rect 37436 9828 37492 9884
rect 57344 9856 57456 9884
rect 914 9772 924 9828
rect 980 9772 1764 9828
rect 3042 9772 3052 9828
rect 3108 9772 7028 9828
rect 10322 9772 10332 9828
rect 10388 9772 14588 9828
rect 14644 9772 14654 9828
rect 15138 9772 15148 9828
rect 15204 9772 21756 9828
rect 21812 9772 21822 9828
rect 21970 9772 21980 9828
rect 22036 9772 25004 9828
rect 25060 9772 25070 9828
rect 25218 9772 25228 9828
rect 25284 9772 28028 9828
rect 28084 9772 28094 9828
rect 28354 9772 28364 9828
rect 28420 9772 36652 9828
rect 36708 9772 36718 9828
rect 36866 9772 36876 9828
rect 36932 9772 37492 9828
rect 38612 9772 40236 9828
rect 40292 9772 40302 9828
rect 40562 9772 40572 9828
rect 40628 9772 52556 9828
rect 52612 9772 52622 9828
rect 690 9660 700 9716
rect 756 9660 1484 9716
rect 1540 9660 1550 9716
rect 6972 9604 7028 9772
rect 38612 9716 38668 9772
rect 7186 9660 7196 9716
rect 7252 9660 10220 9716
rect 10276 9660 10286 9716
rect 11890 9660 11900 9716
rect 11956 9660 18508 9716
rect 18564 9660 18574 9716
rect 20850 9660 20860 9716
rect 20916 9660 21196 9716
rect 21252 9660 28700 9716
rect 28756 9660 28766 9716
rect 29138 9660 29148 9716
rect 29204 9660 33628 9716
rect 33684 9660 33694 9716
rect 35746 9660 35756 9716
rect 35812 9660 38668 9716
rect 41234 9660 41244 9716
rect 41300 9660 44156 9716
rect 44212 9660 44222 9716
rect 45154 9660 45164 9716
rect 45220 9660 51100 9716
rect 51156 9660 51166 9716
rect 252 9548 6188 9604
rect 6244 9548 6254 9604
rect 6972 9548 13132 9604
rect 13188 9548 13198 9604
rect 15698 9548 15708 9604
rect 15764 9548 16828 9604
rect 16884 9548 16894 9604
rect 18162 9548 18172 9604
rect 18228 9548 23660 9604
rect 23716 9548 23726 9604
rect 23986 9548 23996 9604
rect 24052 9548 29596 9604
rect 29652 9548 29662 9604
rect 29810 9548 29820 9604
rect 29876 9548 30828 9604
rect 30884 9548 30894 9604
rect 31042 9548 31052 9604
rect 31108 9548 32284 9604
rect 32340 9548 32350 9604
rect 32498 9548 32508 9604
rect 32564 9548 33180 9604
rect 33236 9548 33246 9604
rect 33842 9548 33852 9604
rect 33908 9548 35644 9604
rect 35700 9548 35710 9604
rect 35858 9548 35868 9604
rect 35924 9548 37884 9604
rect 37940 9548 37950 9604
rect 38098 9548 38108 9604
rect 38164 9548 42700 9604
rect 42756 9548 42766 9604
rect 42914 9548 42924 9604
rect 42980 9548 45052 9604
rect 45108 9548 45118 9604
rect 46946 9548 46956 9604
rect 47012 9548 48300 9604
rect 48356 9548 48366 9604
rect 0 9492 112 9520
rect 252 9492 308 9548
rect 57344 9492 57456 9520
rect 0 9436 308 9492
rect 802 9436 812 9492
rect 868 9436 1820 9492
rect 1876 9436 1886 9492
rect 4162 9436 4172 9492
rect 4228 9436 8316 9492
rect 8372 9436 8382 9492
rect 8540 9436 14476 9492
rect 14532 9436 14542 9492
rect 15922 9436 15932 9492
rect 15988 9436 18284 9492
rect 18340 9436 18350 9492
rect 19394 9436 19404 9492
rect 19460 9436 22428 9492
rect 22484 9436 22494 9492
rect 27122 9436 27132 9492
rect 27188 9436 31724 9492
rect 31780 9436 31790 9492
rect 31938 9436 31948 9492
rect 32004 9436 37772 9492
rect 37828 9436 37838 9492
rect 37986 9436 37996 9492
rect 38052 9436 42364 9492
rect 42420 9436 42430 9492
rect 55122 9436 55132 9492
rect 55188 9436 57456 9492
rect 0 9408 112 9436
rect 3794 9380 3804 9436
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 4068 9380 4078 9436
rect 8540 9380 8596 9436
rect 23794 9380 23804 9436
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 24068 9380 24078 9436
rect 43794 9380 43804 9436
rect 43860 9380 43908 9436
rect 43964 9380 44012 9436
rect 44068 9380 44078 9436
rect 57344 9408 57456 9436
rect 7970 9324 7980 9380
rect 8036 9324 8596 9380
rect 8866 9324 8876 9380
rect 8932 9324 20860 9380
rect 20916 9324 20926 9380
rect 21084 9324 23436 9380
rect 23492 9324 23502 9380
rect 24210 9324 24220 9380
rect 24276 9324 26292 9380
rect 28690 9324 28700 9380
rect 28756 9324 32396 9380
rect 32452 9324 32462 9380
rect 33730 9324 33740 9380
rect 33796 9324 40852 9380
rect 51202 9324 51212 9380
rect 51268 9324 55916 9380
rect 55972 9324 55982 9380
rect 21084 9268 21140 9324
rect 26236 9268 26292 9324
rect 40796 9268 40852 9324
rect 4946 9212 4956 9268
rect 5012 9212 7532 9268
rect 7588 9212 7598 9268
rect 10098 9212 10108 9268
rect 10164 9212 15932 9268
rect 15988 9212 15998 9268
rect 16146 9212 16156 9268
rect 16212 9212 19852 9268
rect 19908 9212 19918 9268
rect 20066 9212 20076 9268
rect 20132 9212 21140 9268
rect 21298 9212 21308 9268
rect 21364 9212 26012 9268
rect 26068 9212 26078 9268
rect 26236 9212 27244 9268
rect 27300 9212 27310 9268
rect 29250 9212 29260 9268
rect 29316 9212 30660 9268
rect 31490 9212 31500 9268
rect 31556 9212 34748 9268
rect 34804 9212 34814 9268
rect 35074 9212 35084 9268
rect 35140 9212 40572 9268
rect 40628 9212 40638 9268
rect 40796 9212 51324 9268
rect 51380 9212 51390 9268
rect 52994 9212 53004 9268
rect 53060 9212 54012 9268
rect 54068 9212 54078 9268
rect 6066 9100 6076 9156
rect 6132 9100 8652 9156
rect 8708 9100 8718 9156
rect 11778 9100 11788 9156
rect 11844 9100 21868 9156
rect 21924 9100 21934 9156
rect 23538 9100 23548 9156
rect 23604 9100 27132 9156
rect 27188 9100 27198 9156
rect 28130 9100 28140 9156
rect 28196 9100 30044 9156
rect 30100 9100 30110 9156
rect 0 9044 112 9072
rect 0 8988 2380 9044
rect 2436 8988 2446 9044
rect 3332 8988 18060 9044
rect 18116 8988 18126 9044
rect 19954 8988 19964 9044
rect 20020 8988 30156 9044
rect 30212 8988 30222 9044
rect 0 8960 112 8988
rect 3332 8932 3388 8988
rect 30604 8932 30660 9212
rect 31154 9100 31164 9156
rect 31220 9100 42252 9156
rect 42308 9100 42318 9156
rect 43138 9100 43148 9156
rect 43204 9100 49644 9156
rect 49700 9100 49710 9156
rect 57344 9044 57456 9072
rect 30818 8988 30828 9044
rect 30884 8988 32508 9044
rect 32564 8988 32574 9044
rect 32722 8988 32732 9044
rect 32788 8988 40236 9044
rect 40292 8988 40302 9044
rect 41906 8988 41916 9044
rect 41972 8988 45724 9044
rect 45780 8988 45790 9044
rect 47842 8988 47852 9044
rect 47908 8988 52780 9044
rect 52836 8988 52846 9044
rect 56130 8988 56140 9044
rect 56196 8988 57456 9044
rect 57344 8960 57456 8988
rect 2034 8876 2044 8932
rect 2100 8876 3388 8932
rect 5068 8876 10108 8932
rect 10164 8876 10174 8932
rect 10322 8876 10332 8932
rect 10388 8876 13020 8932
rect 13076 8876 13086 8932
rect 13234 8876 13244 8932
rect 13300 8876 14252 8932
rect 14308 8876 14318 8932
rect 15250 8876 15260 8932
rect 15316 8876 25228 8932
rect 25284 8876 25294 8932
rect 26898 8876 26908 8932
rect 26964 8876 30380 8932
rect 30436 8876 30446 8932
rect 30604 8876 35532 8932
rect 35588 8876 35598 8932
rect 36530 8876 36540 8932
rect 36596 8876 37716 8932
rect 37874 8876 37884 8932
rect 37940 8876 48972 8932
rect 49028 8876 49038 8932
rect 49858 8876 49868 8932
rect 49924 8876 52668 8932
rect 52724 8876 52734 8932
rect 2156 8652 3388 8708
rect 3444 8652 3454 8708
rect 0 8596 112 8624
rect 2156 8596 2212 8652
rect 4454 8596 4464 8652
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4728 8596 4738 8652
rect 0 8540 2212 8596
rect 2594 8540 2604 8596
rect 2660 8540 2670 8596
rect 0 8512 112 8540
rect 2604 8484 2660 8540
rect 5068 8484 5124 8876
rect 37660 8820 37716 8876
rect 6514 8764 6524 8820
rect 6580 8764 6748 8820
rect 6804 8764 7868 8820
rect 7924 8764 7934 8820
rect 8866 8764 8876 8820
rect 8932 8764 9548 8820
rect 9604 8764 9614 8820
rect 11666 8764 11676 8820
rect 11732 8764 14700 8820
rect 14756 8764 14766 8820
rect 14914 8764 14924 8820
rect 14980 8764 22428 8820
rect 22484 8764 22494 8820
rect 23660 8764 24948 8820
rect 25330 8764 25340 8820
rect 25396 8764 31836 8820
rect 31892 8764 31902 8820
rect 32050 8764 32060 8820
rect 32116 8764 34972 8820
rect 35028 8764 35038 8820
rect 35298 8764 35308 8820
rect 35364 8764 37604 8820
rect 37660 8764 44324 8820
rect 45266 8764 45276 8820
rect 45332 8764 46844 8820
rect 46900 8764 47068 8820
rect 47124 8764 47134 8820
rect 47730 8764 47740 8820
rect 47796 8764 55132 8820
rect 55188 8764 55198 8820
rect 23660 8708 23716 8764
rect 8082 8652 8092 8708
rect 8148 8652 13132 8708
rect 13188 8652 13198 8708
rect 13682 8652 13692 8708
rect 13748 8652 18396 8708
rect 18452 8652 18462 8708
rect 18610 8652 18620 8708
rect 18676 8652 21532 8708
rect 21588 8652 21598 8708
rect 21746 8652 21756 8708
rect 21812 8652 23716 8708
rect 24892 8708 24948 8764
rect 24892 8652 32732 8708
rect 32788 8652 32798 8708
rect 32946 8652 32956 8708
rect 33012 8652 37492 8708
rect 24454 8596 24464 8652
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24728 8596 24738 8652
rect 5282 8540 5292 8596
rect 5348 8540 14140 8596
rect 14196 8540 14206 8596
rect 15708 8540 23100 8596
rect 23156 8540 23166 8596
rect 23426 8540 23436 8596
rect 23492 8540 24332 8596
rect 24388 8540 24398 8596
rect 26786 8540 26796 8596
rect 15708 8484 15764 8540
rect 26852 8484 26908 8596
rect 27010 8540 27020 8596
rect 27076 8540 37380 8596
rect 2604 8428 5124 8484
rect 6636 8428 13524 8484
rect 14802 8428 14812 8484
rect 14868 8428 15764 8484
rect 15922 8428 15932 8484
rect 15988 8428 19628 8484
rect 19684 8428 19694 8484
rect 21644 8428 26236 8484
rect 26292 8428 26302 8484
rect 26852 8428 27300 8484
rect 28466 8428 28476 8484
rect 28532 8428 37100 8484
rect 37156 8428 37166 8484
rect 354 8316 364 8372
rect 420 8316 3388 8372
rect 3714 8316 3724 8372
rect 3780 8316 6412 8372
rect 6468 8316 6478 8372
rect 3332 8260 3388 8316
rect 6636 8260 6692 8428
rect 13468 8372 13524 8428
rect 21644 8372 21700 8428
rect 27244 8372 27300 8428
rect 8306 8316 8316 8372
rect 8372 8316 13244 8372
rect 13300 8316 13310 8372
rect 13458 8316 13468 8372
rect 13524 8316 13534 8372
rect 14130 8316 14140 8372
rect 14196 8316 15148 8372
rect 15204 8316 15214 8372
rect 17042 8316 17052 8372
rect 17108 8316 19516 8372
rect 19572 8316 19582 8372
rect 19730 8316 19740 8372
rect 19796 8316 21700 8372
rect 21858 8316 21868 8372
rect 21924 8316 26348 8372
rect 26404 8316 26414 8372
rect 27244 8316 28924 8372
rect 28980 8316 28990 8372
rect 30146 8316 30156 8372
rect 30212 8316 35196 8372
rect 35252 8316 35262 8372
rect 37324 8260 37380 8540
rect 37436 8372 37492 8652
rect 37548 8484 37604 8764
rect 40226 8652 40236 8708
rect 40292 8652 44044 8708
rect 44100 8652 44110 8708
rect 37762 8540 37772 8596
rect 37828 8540 42924 8596
rect 42980 8540 42990 8596
rect 44268 8484 44324 8764
rect 47618 8652 47628 8708
rect 47684 8652 53564 8708
rect 53620 8652 53630 8708
rect 44454 8596 44464 8652
rect 44520 8596 44568 8652
rect 44624 8596 44672 8652
rect 44728 8596 44738 8652
rect 57344 8596 57456 8624
rect 54338 8540 54348 8596
rect 54404 8540 57456 8596
rect 57344 8512 57456 8540
rect 37548 8428 43596 8484
rect 43652 8428 43662 8484
rect 44268 8428 50764 8484
rect 50820 8428 50830 8484
rect 37436 8316 39788 8372
rect 39844 8316 40236 8372
rect 40292 8316 40302 8372
rect 41906 8316 41916 8372
rect 41972 8316 48076 8372
rect 48132 8316 48412 8372
rect 48468 8316 48478 8372
rect 48962 8316 48972 8372
rect 49028 8316 50988 8372
rect 51044 8316 51054 8372
rect 53330 8316 53340 8372
rect 53396 8316 55692 8372
rect 55748 8316 55758 8372
rect 2230 8204 2268 8260
rect 2324 8204 2334 8260
rect 3332 8204 6692 8260
rect 8306 8204 8316 8260
rect 8372 8204 13692 8260
rect 13748 8204 13758 8260
rect 13906 8204 13916 8260
rect 13972 8204 15484 8260
rect 15540 8204 15550 8260
rect 16034 8204 16044 8260
rect 16100 8204 21532 8260
rect 21588 8204 21598 8260
rect 21756 8204 22316 8260
rect 22372 8204 22382 8260
rect 23202 8204 23212 8260
rect 23268 8204 25788 8260
rect 25844 8204 25854 8260
rect 26226 8204 26236 8260
rect 26292 8204 26908 8260
rect 26964 8204 26974 8260
rect 28802 8204 28812 8260
rect 28868 8204 30380 8260
rect 30436 8204 30446 8260
rect 30706 8204 30716 8260
rect 30772 8204 35644 8260
rect 35700 8204 35710 8260
rect 37324 8204 38780 8260
rect 38836 8204 38846 8260
rect 43362 8204 43372 8260
rect 43428 8204 52556 8260
rect 52612 8204 52622 8260
rect 0 8148 112 8176
rect 21756 8148 21812 8204
rect 57344 8148 57456 8176
rect 0 8092 1484 8148
rect 1540 8092 1550 8148
rect 10098 8092 10108 8148
rect 10164 8092 10892 8148
rect 10948 8092 10958 8148
rect 11442 8092 11452 8148
rect 11508 8092 15372 8148
rect 15428 8092 15438 8148
rect 15586 8092 15596 8148
rect 15652 8092 17500 8148
rect 17556 8092 17566 8148
rect 18498 8092 18508 8148
rect 18564 8092 21812 8148
rect 22082 8092 22092 8148
rect 22148 8092 22428 8148
rect 22484 8092 28252 8148
rect 28308 8092 28318 8148
rect 30034 8092 30044 8148
rect 30100 8092 33516 8148
rect 33572 8092 33582 8148
rect 34850 8092 34860 8148
rect 34916 8092 38780 8148
rect 38836 8092 38846 8148
rect 39218 8092 39228 8148
rect 39284 8092 44268 8148
rect 44324 8092 44334 8148
rect 51986 8092 51996 8148
rect 52052 8092 53900 8148
rect 53956 8092 53966 8148
rect 55906 8092 55916 8148
rect 55972 8092 57456 8148
rect 0 8064 112 8092
rect 57344 8064 57456 8092
rect 1596 7980 6804 8036
rect 9202 7980 9212 8036
rect 9268 7980 14812 8036
rect 14868 7980 14878 8036
rect 15026 7980 15036 8036
rect 15092 7980 23212 8036
rect 23268 7980 23278 8036
rect 23436 7980 24388 8036
rect 24546 7980 24556 8036
rect 24612 7980 26796 8036
rect 26852 7980 26862 8036
rect 27010 7980 27020 8036
rect 27076 7980 33404 8036
rect 33460 7980 33470 8036
rect 34962 7980 34972 8036
rect 35028 7980 38444 8036
rect 38500 7980 38510 8036
rect 38602 7980 38612 8036
rect 38668 7980 41244 8036
rect 41300 7980 41310 8036
rect 43586 7980 43596 8036
rect 43652 7980 53452 8036
rect 53508 7980 53518 8036
rect 0 7700 112 7728
rect 1596 7700 1652 7980
rect 3794 7812 3804 7868
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 4068 7812 4078 7868
rect 6748 7812 6804 7980
rect 23436 7924 23492 7980
rect 9090 7868 9100 7924
rect 9156 7868 19964 7924
rect 20020 7868 20030 7924
rect 20514 7868 20524 7924
rect 20580 7868 23492 7924
rect 24332 7924 24388 7980
rect 24332 7868 31052 7924
rect 31108 7868 31118 7924
rect 31490 7868 31500 7924
rect 31556 7868 33292 7924
rect 33348 7868 33358 7924
rect 33618 7868 33628 7924
rect 33684 7868 38780 7924
rect 38836 7868 38846 7924
rect 44146 7868 44156 7924
rect 44212 7868 46620 7924
rect 46676 7868 46686 7924
rect 47058 7868 47068 7924
rect 47124 7868 50316 7924
rect 50372 7868 50382 7924
rect 23794 7812 23804 7868
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 24068 7812 24078 7868
rect 43794 7812 43804 7868
rect 43860 7812 43908 7868
rect 43964 7812 44012 7868
rect 44068 7812 44078 7868
rect 6748 7756 10668 7812
rect 10724 7756 10734 7812
rect 12002 7756 12012 7812
rect 12068 7756 19180 7812
rect 19236 7756 19246 7812
rect 19506 7756 19516 7812
rect 19572 7756 21868 7812
rect 21924 7756 21934 7812
rect 24220 7756 26684 7812
rect 26740 7756 26750 7812
rect 30258 7756 30268 7812
rect 30324 7756 43148 7812
rect 43204 7756 43214 7812
rect 52994 7756 53004 7812
rect 53060 7756 56028 7812
rect 56084 7756 56094 7812
rect 24220 7700 24276 7756
rect 57344 7700 57456 7728
rect 0 7644 1652 7700
rect 2930 7644 2940 7700
rect 2996 7644 16268 7700
rect 16324 7644 16334 7700
rect 16492 7644 18284 7700
rect 18340 7644 18350 7700
rect 20402 7644 20412 7700
rect 20468 7644 24276 7700
rect 24434 7644 24444 7700
rect 24500 7644 26012 7700
rect 26068 7644 26078 7700
rect 26786 7644 26796 7700
rect 26852 7644 31276 7700
rect 31332 7644 31342 7700
rect 31602 7644 31612 7700
rect 31668 7644 32004 7700
rect 32834 7644 32844 7700
rect 32900 7644 41580 7700
rect 41636 7644 41646 7700
rect 41906 7644 41916 7700
rect 41972 7644 45276 7700
rect 45332 7644 45342 7700
rect 56130 7644 56140 7700
rect 56196 7644 57456 7700
rect 0 7616 112 7644
rect 16492 7588 16548 7644
rect 31948 7588 32004 7644
rect 57344 7616 57456 7644
rect 1810 7532 1820 7588
rect 1876 7532 9660 7588
rect 9716 7532 9996 7588
rect 10052 7532 10062 7588
rect 13458 7532 13468 7588
rect 13524 7532 16548 7588
rect 16706 7532 16716 7588
rect 16772 7532 18956 7588
rect 19012 7532 19022 7588
rect 19292 7532 26908 7588
rect 26964 7532 26974 7588
rect 29474 7532 29484 7588
rect 29540 7532 31724 7588
rect 31780 7532 31790 7588
rect 31948 7532 33404 7588
rect 33460 7532 33470 7588
rect 33618 7532 33628 7588
rect 33684 7532 43372 7588
rect 43428 7532 43438 7588
rect 43596 7532 52332 7588
rect 52388 7532 52398 7588
rect 19292 7476 19348 7532
rect 43596 7476 43652 7532
rect 6178 7420 6188 7476
rect 6244 7420 8428 7476
rect 8484 7420 8494 7476
rect 11890 7420 11900 7476
rect 11956 7420 14924 7476
rect 14980 7420 14990 7476
rect 15082 7420 15092 7476
rect 15148 7420 16716 7476
rect 16772 7420 16782 7476
rect 18386 7420 18396 7476
rect 18452 7420 19348 7476
rect 19506 7420 19516 7476
rect 19572 7420 19740 7476
rect 19796 7420 19806 7476
rect 20850 7420 20860 7476
rect 20916 7420 23436 7476
rect 23492 7420 23502 7476
rect 23650 7420 23660 7476
rect 23716 7420 25620 7476
rect 26674 7420 26684 7476
rect 26740 7420 29372 7476
rect 29428 7420 29438 7476
rect 29698 7420 29708 7476
rect 29764 7420 35420 7476
rect 35476 7420 35486 7476
rect 35634 7420 35644 7476
rect 35700 7420 38444 7476
rect 38500 7420 38510 7476
rect 38602 7420 38612 7476
rect 38668 7420 43652 7476
rect 43810 7420 43820 7476
rect 43876 7420 54124 7476
rect 54180 7420 54190 7476
rect 25564 7364 25620 7420
rect 3490 7308 3500 7364
rect 3556 7308 5964 7364
rect 6020 7308 6030 7364
rect 7298 7308 7308 7364
rect 7364 7308 10276 7364
rect 10546 7308 10556 7364
rect 10612 7308 12796 7364
rect 12852 7308 12862 7364
rect 13122 7308 13132 7364
rect 13188 7308 25340 7364
rect 25396 7308 25406 7364
rect 25564 7308 30044 7364
rect 30100 7308 30110 7364
rect 30370 7308 30380 7364
rect 30436 7308 33180 7364
rect 33236 7308 33246 7364
rect 33394 7308 33404 7364
rect 33460 7308 55132 7364
rect 55188 7308 55198 7364
rect 0 7252 112 7280
rect 10220 7252 10276 7308
rect 57344 7252 57456 7280
rect 0 7196 9268 7252
rect 10220 7196 12124 7252
rect 12180 7196 12190 7252
rect 13010 7196 13020 7252
rect 13076 7196 20860 7252
rect 20916 7196 20926 7252
rect 21970 7196 21980 7252
rect 22036 7196 27468 7252
rect 27524 7196 27534 7252
rect 27906 7196 27916 7252
rect 27972 7196 30716 7252
rect 30772 7196 30782 7252
rect 31154 7196 31164 7252
rect 31220 7196 43820 7252
rect 43876 7196 43886 7252
rect 44044 7196 48860 7252
rect 48916 7196 48926 7252
rect 54562 7196 54572 7252
rect 54628 7196 57456 7252
rect 0 7168 112 7196
rect 9212 7140 9268 7196
rect 44044 7140 44100 7196
rect 57344 7168 57456 7196
rect 9212 7084 12908 7140
rect 12964 7084 12974 7140
rect 13682 7084 13692 7140
rect 13748 7084 16044 7140
rect 16100 7084 16110 7140
rect 16268 7084 18172 7140
rect 18228 7084 18238 7140
rect 18386 7084 18396 7140
rect 18452 7084 21532 7140
rect 21588 7084 21598 7140
rect 21858 7084 21868 7140
rect 21924 7084 24220 7140
rect 24276 7084 24286 7140
rect 25218 7084 25228 7140
rect 25284 7084 30044 7140
rect 30100 7084 30110 7140
rect 30818 7084 30828 7140
rect 30884 7084 31612 7140
rect 31668 7084 31678 7140
rect 31938 7084 31948 7140
rect 32004 7084 35196 7140
rect 35252 7084 35262 7140
rect 35410 7084 35420 7140
rect 35476 7084 40684 7140
rect 40740 7084 40750 7140
rect 43586 7084 43596 7140
rect 43652 7084 44100 7140
rect 4454 7028 4464 7084
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4728 7028 4738 7084
rect 16268 7028 16324 7084
rect 24454 7028 24464 7084
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 24728 7028 24738 7084
rect 44454 7028 44464 7084
rect 44520 7028 44568 7084
rect 44624 7028 44672 7084
rect 44728 7028 44738 7084
rect 5964 6972 13692 7028
rect 13748 6972 13758 7028
rect 14130 6972 14140 7028
rect 14196 6972 16324 7028
rect 16482 6972 16492 7028
rect 16548 6972 23660 7028
rect 23716 6972 23726 7028
rect 25442 6972 25452 7028
rect 25508 6972 36876 7028
rect 36932 6972 36942 7028
rect 37874 6972 37884 7028
rect 37940 6972 40460 7028
rect 40516 6972 40526 7028
rect 41570 6972 41580 7028
rect 41636 6972 44268 7028
rect 44324 6972 44334 7028
rect 45378 6972 45388 7028
rect 45444 6972 47964 7028
rect 48020 6972 48030 7028
rect 48962 6972 48972 7028
rect 49028 6972 52892 7028
rect 52948 6972 52958 7028
rect 578 6860 588 6916
rect 644 6860 4956 6916
rect 5012 6860 5022 6916
rect 0 6804 112 6832
rect 5964 6804 6020 6972
rect 6514 6860 6524 6916
rect 6580 6860 9660 6916
rect 9716 6860 9726 6916
rect 9996 6860 20412 6916
rect 20468 6860 20478 6916
rect 20850 6860 20860 6916
rect 20916 6860 33740 6916
rect 33796 6860 33806 6916
rect 33954 6860 33964 6916
rect 34020 6860 36204 6916
rect 36260 6860 36270 6916
rect 36978 6860 36988 6916
rect 37044 6860 40124 6916
rect 40180 6860 40190 6916
rect 40338 6860 40348 6916
rect 40404 6860 52108 6916
rect 52164 6860 52174 6916
rect 9996 6804 10052 6860
rect 57344 6804 57456 6832
rect 0 6748 6020 6804
rect 6290 6748 6300 6804
rect 6356 6748 8428 6804
rect 9314 6748 9324 6804
rect 9380 6748 10052 6804
rect 10108 6748 13412 6804
rect 13794 6748 13804 6804
rect 13860 6748 16156 6804
rect 16212 6748 16222 6804
rect 16604 6748 17948 6804
rect 18004 6748 18014 6804
rect 18162 6748 18172 6804
rect 18228 6748 25116 6804
rect 25172 6748 25182 6804
rect 25330 6748 25340 6804
rect 25396 6748 28364 6804
rect 28420 6748 28430 6804
rect 30146 6748 30156 6804
rect 30212 6748 33516 6804
rect 33572 6748 33582 6804
rect 35522 6748 35532 6804
rect 35588 6748 40236 6804
rect 40292 6748 40302 6804
rect 42028 6748 46732 6804
rect 46788 6748 46798 6804
rect 46956 6748 48524 6804
rect 48580 6748 48590 6804
rect 56130 6748 56140 6804
rect 56196 6748 57456 6804
rect 0 6720 112 6748
rect 8372 6580 8428 6748
rect 10108 6692 10164 6748
rect 8754 6636 8764 6692
rect 8820 6636 10164 6692
rect 13356 6692 13412 6748
rect 16604 6692 16660 6748
rect 42028 6692 42084 6748
rect 13356 6636 16156 6692
rect 16212 6636 16222 6692
rect 16370 6636 16380 6692
rect 16436 6636 16660 6692
rect 20626 6636 20636 6692
rect 20692 6636 27300 6692
rect 27458 6636 27468 6692
rect 27524 6636 29148 6692
rect 29204 6636 29214 6692
rect 29372 6636 30380 6692
rect 30436 6636 30446 6692
rect 31378 6636 31388 6692
rect 31444 6636 33740 6692
rect 33796 6636 33806 6692
rect 33954 6636 33964 6692
rect 34020 6636 42084 6692
rect 3602 6524 3612 6580
rect 3668 6524 6188 6580
rect 6244 6524 6254 6580
rect 8372 6524 15148 6580
rect 15474 6524 15484 6580
rect 15540 6524 19740 6580
rect 19796 6524 19806 6580
rect 21074 6524 21084 6580
rect 21140 6524 22764 6580
rect 22820 6524 22830 6580
rect 23650 6524 23660 6580
rect 23716 6524 23772 6580
rect 23828 6524 23838 6580
rect 23986 6524 23996 6580
rect 24052 6524 26908 6580
rect 26964 6524 26974 6580
rect 15092 6468 15148 6524
rect 27244 6468 27300 6636
rect 29372 6580 29428 6636
rect 46956 6580 47012 6748
rect 57344 6720 57456 6748
rect 47506 6636 47516 6692
rect 47572 6636 52220 6692
rect 52276 6636 52286 6692
rect 28466 6524 28476 6580
rect 28532 6524 29428 6580
rect 30034 6524 30044 6580
rect 30100 6524 36988 6580
rect 37044 6524 37054 6580
rect 37202 6524 37212 6580
rect 37268 6524 39004 6580
rect 39060 6524 39070 6580
rect 39218 6524 39228 6580
rect 39284 6524 41244 6580
rect 41300 6524 41310 6580
rect 41682 6524 41692 6580
rect 41748 6524 47012 6580
rect 3276 6412 4900 6468
rect 6850 6412 6860 6468
rect 6916 6412 14924 6468
rect 14980 6412 14990 6468
rect 15092 6412 16548 6468
rect 16706 6412 16716 6468
rect 16772 6412 21756 6468
rect 21812 6412 21822 6468
rect 23314 6412 23324 6468
rect 23380 6412 25340 6468
rect 25396 6412 25406 6468
rect 27244 6412 29820 6468
rect 29876 6412 29886 6468
rect 30034 6412 30044 6468
rect 30100 6412 31164 6468
rect 31220 6412 31230 6468
rect 32050 6412 32060 6468
rect 32116 6412 35868 6468
rect 35924 6412 35934 6468
rect 37090 6412 37100 6468
rect 37156 6412 42028 6468
rect 42084 6412 42094 6468
rect 43138 6412 43148 6468
rect 43204 6412 54908 6468
rect 54964 6412 54974 6468
rect 0 6356 112 6384
rect 3276 6356 3332 6412
rect 0 6300 3332 6356
rect 4844 6356 4900 6412
rect 16492 6356 16548 6412
rect 57344 6356 57456 6384
rect 4844 6300 9212 6356
rect 9268 6300 9278 6356
rect 9762 6300 9772 6356
rect 9828 6300 15260 6356
rect 15316 6300 15326 6356
rect 16492 6300 20860 6356
rect 20916 6300 20926 6356
rect 21522 6300 21532 6356
rect 21588 6300 22260 6356
rect 24210 6300 24220 6356
rect 24276 6300 31500 6356
rect 31556 6300 31566 6356
rect 31826 6300 31836 6356
rect 31892 6300 37996 6356
rect 38052 6300 38062 6356
rect 38994 6300 39004 6356
rect 39060 6300 41356 6356
rect 41412 6300 41422 6356
rect 55122 6300 55132 6356
rect 55188 6300 57456 6356
rect 0 6272 112 6300
rect 3794 6244 3804 6300
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 4068 6244 4078 6300
rect 22204 6244 22260 6300
rect 23794 6244 23804 6300
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 24068 6244 24078 6300
rect 43794 6244 43804 6300
rect 43860 6244 43908 6300
rect 43964 6244 44012 6300
rect 44068 6244 44078 6300
rect 57344 6272 57456 6300
rect 6290 6188 6300 6244
rect 6356 6188 18284 6244
rect 18340 6188 18350 6244
rect 19170 6188 19180 6244
rect 19236 6188 22148 6244
rect 22204 6188 23660 6244
rect 23716 6188 23726 6244
rect 26786 6188 26796 6244
rect 26852 6188 28196 6244
rect 28354 6188 28364 6244
rect 28420 6188 38556 6244
rect 38612 6188 38622 6244
rect 40338 6188 40348 6244
rect 40404 6188 43484 6244
rect 43540 6188 43550 6244
rect 45378 6188 45388 6244
rect 45444 6188 48972 6244
rect 49028 6188 49038 6244
rect 22092 6132 22148 6188
rect 28140 6132 28196 6188
rect 2818 6076 2828 6132
rect 2884 6076 8764 6132
rect 8820 6076 8830 6132
rect 10210 6076 10220 6132
rect 10276 6076 11900 6132
rect 11956 6076 11966 6132
rect 12898 6076 12908 6132
rect 12964 6076 14812 6132
rect 14868 6076 14878 6132
rect 15026 6076 15036 6132
rect 15092 6076 21868 6132
rect 21924 6076 21934 6132
rect 22092 6076 27916 6132
rect 27972 6076 27982 6132
rect 28140 6076 35308 6132
rect 35364 6076 35374 6132
rect 36978 6076 36988 6132
rect 37044 6076 41916 6132
rect 41972 6076 41982 6132
rect 43586 6076 43596 6132
rect 43652 6076 47404 6132
rect 47460 6076 47470 6132
rect 48850 6076 48860 6132
rect 48916 6076 50988 6132
rect 51044 6076 51054 6132
rect 52994 6076 53004 6132
rect 53060 6076 56700 6132
rect 56756 6076 56766 6132
rect 9202 5964 9212 6020
rect 9268 5964 11788 6020
rect 11844 5964 11854 6020
rect 12002 5964 12012 6020
rect 12068 5964 14756 6020
rect 14914 5964 14924 6020
rect 14980 5964 24108 6020
rect 24164 5964 24174 6020
rect 24332 5964 27804 6020
rect 27860 5964 27870 6020
rect 28018 5964 28028 6020
rect 28084 5964 28980 6020
rect 29138 5964 29148 6020
rect 29204 5964 31500 6020
rect 31556 5964 31566 6020
rect 31826 5964 31836 6020
rect 31892 5964 35084 6020
rect 35140 5964 35150 6020
rect 35858 5964 35868 6020
rect 35924 5964 37324 6020
rect 37380 5964 37390 6020
rect 37538 5964 37548 6020
rect 37604 5964 53564 6020
rect 53620 5964 53630 6020
rect 0 5908 112 5936
rect 14700 5908 14756 5964
rect 24332 5908 24388 5964
rect 28924 5908 28980 5964
rect 57344 5908 57456 5936
rect 0 5852 6860 5908
rect 6916 5852 6926 5908
rect 9100 5852 11676 5908
rect 11732 5852 11742 5908
rect 11890 5852 11900 5908
rect 11956 5852 14476 5908
rect 14532 5852 14542 5908
rect 14700 5852 16156 5908
rect 16212 5852 16222 5908
rect 16594 5852 16604 5908
rect 16660 5852 18060 5908
rect 18116 5852 18126 5908
rect 18274 5852 18284 5908
rect 18340 5852 20972 5908
rect 21028 5852 21038 5908
rect 21410 5852 21420 5908
rect 21476 5852 24388 5908
rect 24546 5852 24556 5908
rect 24612 5852 28700 5908
rect 28756 5852 28766 5908
rect 28924 5852 32172 5908
rect 32228 5852 32238 5908
rect 32946 5852 32956 5908
rect 33012 5852 33292 5908
rect 33348 5852 33358 5908
rect 33506 5852 33516 5908
rect 33572 5852 37324 5908
rect 37380 5852 37390 5908
rect 40562 5852 40572 5908
rect 40628 5852 48748 5908
rect 48804 5852 48814 5908
rect 54562 5852 54572 5908
rect 54628 5852 57456 5908
rect 0 5824 112 5852
rect 6066 5740 6076 5796
rect 6132 5740 7980 5796
rect 8036 5740 8046 5796
rect 9100 5684 9156 5852
rect 57344 5824 57456 5852
rect 9650 5740 9660 5796
rect 9716 5740 15484 5796
rect 15540 5740 15550 5796
rect 16146 5740 16156 5796
rect 16212 5740 21532 5796
rect 21588 5740 21598 5796
rect 22082 5740 22092 5796
rect 22148 5740 25228 5796
rect 25284 5740 25294 5796
rect 26898 5740 26908 5796
rect 26964 5740 29092 5796
rect 30034 5740 30044 5796
rect 30100 5740 30380 5796
rect 30436 5740 30446 5796
rect 30930 5740 30940 5796
rect 30996 5740 54124 5796
rect 54180 5740 54190 5796
rect 29036 5684 29092 5740
rect 2706 5628 2716 5684
rect 2772 5628 9156 5684
rect 11218 5628 11228 5684
rect 11284 5628 13916 5684
rect 13972 5628 13982 5684
rect 14802 5628 14812 5684
rect 14868 5628 15148 5684
rect 15204 5628 15214 5684
rect 15362 5628 15372 5684
rect 15428 5628 16268 5684
rect 16324 5628 16334 5684
rect 16492 5628 18396 5684
rect 18452 5628 18462 5684
rect 18722 5628 18732 5684
rect 18788 5628 19964 5684
rect 20020 5628 20030 5684
rect 20178 5628 20188 5684
rect 20244 5628 21644 5684
rect 21700 5628 21710 5684
rect 21858 5628 21868 5684
rect 21924 5628 28476 5684
rect 28532 5628 28542 5684
rect 29036 5628 31556 5684
rect 31826 5628 31836 5684
rect 31892 5628 37548 5684
rect 37604 5628 37614 5684
rect 38658 5628 38668 5684
rect 38724 5628 43596 5684
rect 43652 5628 43662 5684
rect 44258 5628 44268 5684
rect 44324 5628 44884 5684
rect 48738 5628 48748 5684
rect 48804 5628 52444 5684
rect 52500 5628 52510 5684
rect 16492 5572 16548 5628
rect 5170 5516 5180 5572
rect 5236 5516 11452 5572
rect 11508 5516 11518 5572
rect 11666 5516 11676 5572
rect 11732 5516 16548 5572
rect 16706 5516 16716 5572
rect 16772 5516 19964 5572
rect 20020 5516 20030 5572
rect 20962 5516 20972 5572
rect 21028 5516 22092 5572
rect 22148 5516 22158 5572
rect 22306 5516 22316 5572
rect 22372 5516 24220 5572
rect 24276 5516 24286 5572
rect 24882 5516 24892 5572
rect 24948 5516 31164 5572
rect 31220 5516 31230 5572
rect 0 5460 112 5488
rect 4454 5460 4464 5516
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4728 5460 4738 5516
rect 24454 5460 24464 5516
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24728 5460 24738 5516
rect 31500 5460 31556 5628
rect 32946 5516 32956 5572
rect 33012 5516 35756 5572
rect 35812 5516 35822 5572
rect 37090 5516 37100 5572
rect 37156 5516 44324 5572
rect 0 5404 140 5460
rect 196 5404 206 5460
rect 9202 5404 9212 5460
rect 9268 5404 13580 5460
rect 13636 5404 13646 5460
rect 14242 5404 14252 5460
rect 14308 5404 18396 5460
rect 18452 5404 18462 5460
rect 18610 5404 18620 5460
rect 18676 5404 24332 5460
rect 24388 5404 24398 5460
rect 24994 5404 25004 5460
rect 25060 5404 26572 5460
rect 26628 5404 26638 5460
rect 26786 5404 26796 5460
rect 26852 5404 27132 5460
rect 27188 5404 27198 5460
rect 28354 5404 28364 5460
rect 28420 5404 28430 5460
rect 31500 5404 33852 5460
rect 33908 5404 33918 5460
rect 34076 5404 36540 5460
rect 36596 5404 36606 5460
rect 0 5376 112 5404
rect 28364 5348 28420 5404
rect 34076 5348 34132 5404
rect 44268 5348 44324 5516
rect 44454 5460 44464 5516
rect 44520 5460 44568 5516
rect 44624 5460 44672 5516
rect 44728 5460 44738 5516
rect 44828 5460 44884 5628
rect 48290 5516 48300 5572
rect 48356 5516 54124 5572
rect 54180 5516 54190 5572
rect 57344 5460 57456 5488
rect 44828 5404 51884 5460
rect 51940 5404 52332 5460
rect 52388 5404 52398 5460
rect 56130 5404 56140 5460
rect 56196 5404 57456 5460
rect 57344 5376 57456 5404
rect 2594 5292 2604 5348
rect 2660 5292 2940 5348
rect 2996 5292 13356 5348
rect 13412 5292 13422 5348
rect 13570 5292 13580 5348
rect 13636 5292 16492 5348
rect 16548 5292 16558 5348
rect 16706 5292 16716 5348
rect 16772 5292 28420 5348
rect 28476 5292 28812 5348
rect 28868 5292 31052 5348
rect 31108 5292 31118 5348
rect 31714 5292 31724 5348
rect 31780 5292 33404 5348
rect 33460 5292 33470 5348
rect 33852 5292 34132 5348
rect 35298 5292 35308 5348
rect 35364 5292 40292 5348
rect 40450 5292 40460 5348
rect 40516 5292 42140 5348
rect 42196 5292 42206 5348
rect 44268 5292 45388 5348
rect 45444 5292 45454 5348
rect 28476 5236 28532 5292
rect 33852 5236 33908 5292
rect 40236 5236 40292 5292
rect 1026 5180 1036 5236
rect 1092 5180 1820 5236
rect 1876 5180 1886 5236
rect 4946 5180 4956 5236
rect 5012 5180 9884 5236
rect 9940 5180 9950 5236
rect 10098 5180 10108 5236
rect 10164 5180 11564 5236
rect 11620 5180 11630 5236
rect 11778 5180 11788 5236
rect 11844 5180 14924 5236
rect 14980 5180 14990 5236
rect 15092 5180 20972 5236
rect 21028 5180 21038 5236
rect 21196 5180 23436 5236
rect 23492 5180 23502 5236
rect 23650 5180 23660 5236
rect 23716 5180 25788 5236
rect 25844 5180 25854 5236
rect 28466 5180 28476 5236
rect 28532 5180 28542 5236
rect 29474 5180 29484 5236
rect 29540 5180 33404 5236
rect 33460 5180 33470 5236
rect 33740 5180 33908 5236
rect 34066 5180 34076 5236
rect 34132 5180 37548 5236
rect 37604 5180 37614 5236
rect 38210 5180 38220 5236
rect 38276 5180 38668 5236
rect 38724 5180 38734 5236
rect 40236 5180 45276 5236
rect 45332 5180 45342 5236
rect 48626 5180 48636 5236
rect 48692 5180 51996 5236
rect 52052 5180 52062 5236
rect 52882 5180 52892 5236
rect 52948 5180 55020 5236
rect 55076 5180 55086 5236
rect 15092 5124 15148 5180
rect 21196 5124 21252 5180
rect 33740 5124 33796 5180
rect 1698 5068 1708 5124
rect 1764 5068 13412 5124
rect 13570 5068 13580 5124
rect 13636 5068 15148 5124
rect 16034 5068 16044 5124
rect 16100 5068 21252 5124
rect 21756 5068 30156 5124
rect 30212 5068 30222 5124
rect 31042 5068 31052 5124
rect 31108 5068 31948 5124
rect 32004 5068 32014 5124
rect 32358 5068 32396 5124
rect 32452 5068 32462 5124
rect 32946 5068 32956 5124
rect 33012 5068 33068 5124
rect 33124 5068 33134 5124
rect 33282 5068 33292 5124
rect 33348 5068 33796 5124
rect 33954 5068 33964 5124
rect 34020 5068 35252 5124
rect 38770 5068 38780 5124
rect 38836 5068 40516 5124
rect 0 5012 112 5040
rect 13356 5012 13412 5068
rect 21756 5012 21812 5068
rect 35196 5012 35252 5068
rect 0 4956 1596 5012
rect 1652 4956 1662 5012
rect 2258 4956 2268 5012
rect 2324 4956 4676 5012
rect 5058 4956 5068 5012
rect 5124 4956 13188 5012
rect 13356 4956 21812 5012
rect 23538 4956 23548 5012
rect 23604 4956 26796 5012
rect 26852 4956 26862 5012
rect 27010 4956 27020 5012
rect 27076 4956 33628 5012
rect 33684 4956 33694 5012
rect 33842 4956 33852 5012
rect 33908 4956 34916 5012
rect 35196 4956 40404 5012
rect 0 4928 112 4956
rect 1474 4844 1484 4900
rect 1540 4844 4396 4900
rect 4452 4844 4462 4900
rect 4620 4788 4676 4956
rect 13132 4900 13188 4956
rect 34860 4900 34916 4956
rect 4834 4844 4844 4900
rect 4900 4844 11788 4900
rect 11844 4844 11854 4900
rect 13132 4844 13244 4900
rect 13300 4844 13310 4900
rect 13458 4844 13468 4900
rect 13524 4844 16716 4900
rect 16772 4844 16782 4900
rect 16940 4844 24892 4900
rect 24948 4844 24958 4900
rect 25218 4844 25228 4900
rect 25284 4844 30268 4900
rect 30324 4844 30334 4900
rect 30706 4844 30716 4900
rect 30772 4844 34636 4900
rect 34692 4844 34702 4900
rect 34860 4844 35756 4900
rect 35812 4844 35822 4900
rect 4620 4732 9212 4788
rect 9268 4732 9278 4788
rect 11900 4732 16716 4788
rect 16772 4732 16782 4788
rect 3794 4676 3804 4732
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 4068 4676 4078 4732
rect 11900 4676 11956 4732
rect 16940 4676 16996 4844
rect 40348 4788 40404 4956
rect 40460 4900 40516 5068
rect 42028 5068 53228 5124
rect 53284 5068 53294 5124
rect 54898 5068 54908 5124
rect 54964 5068 56084 5124
rect 42028 5012 42084 5068
rect 56028 5012 56084 5068
rect 57344 5012 57456 5040
rect 41794 4956 41804 5012
rect 41860 4956 42084 5012
rect 42802 4956 42812 5012
rect 42868 4956 45164 5012
rect 45220 4956 45230 5012
rect 45378 4956 45388 5012
rect 45444 4956 52668 5012
rect 52724 4956 52734 5012
rect 52882 4956 52892 5012
rect 52948 4956 53676 5012
rect 53732 4956 53742 5012
rect 56028 4956 57456 5012
rect 57344 4928 57456 4956
rect 40460 4844 48748 4900
rect 48804 4844 48814 4900
rect 52434 4844 52444 4900
rect 52500 4844 54796 4900
rect 54852 4844 54862 4900
rect 18050 4732 18060 4788
rect 18116 4732 23324 4788
rect 23380 4732 23390 4788
rect 25106 4732 25116 4788
rect 25172 4732 33628 4788
rect 33684 4732 33694 4788
rect 34962 4732 34972 4788
rect 35028 4732 36316 4788
rect 36372 4732 36382 4788
rect 36530 4732 36540 4788
rect 36596 4732 38668 4788
rect 40348 4732 43596 4788
rect 43652 4732 43662 4788
rect 44146 4732 44156 4788
rect 44212 4732 47068 4788
rect 47124 4732 47134 4788
rect 49522 4732 49532 4788
rect 49588 4732 55356 4788
rect 55412 4732 55422 4788
rect 23794 4676 23804 4732
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 24068 4676 24078 4732
rect 38612 4676 38668 4732
rect 43794 4676 43804 4732
rect 43860 4676 43908 4732
rect 43964 4676 44012 4732
rect 44068 4676 44078 4732
rect 4162 4620 4172 4676
rect 4228 4620 11956 4676
rect 12562 4620 12572 4676
rect 12628 4620 14812 4676
rect 14868 4620 14878 4676
rect 15092 4620 16996 4676
rect 18274 4620 18284 4676
rect 18340 4620 21196 4676
rect 21252 4620 21262 4676
rect 21858 4620 21868 4676
rect 21924 4620 23660 4676
rect 23716 4620 23726 4676
rect 24210 4620 24220 4676
rect 24276 4620 25452 4676
rect 25508 4620 25518 4676
rect 25778 4620 25788 4676
rect 25844 4620 28476 4676
rect 28532 4620 28542 4676
rect 28914 4620 28924 4676
rect 28980 4620 36988 4676
rect 37044 4620 37054 4676
rect 38612 4620 43484 4676
rect 43540 4620 43550 4676
rect 50530 4620 50540 4676
rect 50596 4620 53564 4676
rect 53620 4620 53630 4676
rect 0 4564 112 4592
rect 0 4508 6524 4564
rect 6580 4508 6590 4564
rect 6850 4508 6860 4564
rect 6916 4508 8652 4564
rect 8708 4508 8718 4564
rect 9874 4508 9884 4564
rect 9940 4508 14924 4564
rect 14980 4508 14990 4564
rect 0 4480 112 4508
rect 15092 4452 15148 4620
rect 57344 4564 57456 4592
rect 15250 4508 15260 4564
rect 15316 4508 27580 4564
rect 27636 4508 27646 4564
rect 27794 4508 27804 4564
rect 27860 4508 29260 4564
rect 29316 4508 29326 4564
rect 29810 4508 29820 4564
rect 29876 4508 36876 4564
rect 36932 4508 36942 4564
rect 39890 4508 39900 4564
rect 39956 4508 40348 4564
rect 40404 4508 40414 4564
rect 43586 4508 43596 4564
rect 43652 4508 50428 4564
rect 50484 4508 50494 4564
rect 54562 4508 54572 4564
rect 54628 4508 57456 4564
rect 57344 4480 57456 4508
rect 3378 4396 3388 4452
rect 3444 4396 4844 4452
rect 4900 4396 5180 4452
rect 5236 4396 5246 4452
rect 6738 4396 6748 4452
rect 6804 4396 15148 4452
rect 16146 4396 16156 4452
rect 16212 4396 18732 4452
rect 18788 4396 18798 4452
rect 18946 4396 18956 4452
rect 19012 4396 20412 4452
rect 20468 4396 20478 4452
rect 20850 4396 20860 4452
rect 20916 4396 25564 4452
rect 25620 4396 25630 4452
rect 25890 4396 25900 4452
rect 25956 4396 32844 4452
rect 32900 4396 32910 4452
rect 33068 4396 34972 4452
rect 35028 4396 35038 4452
rect 35186 4396 35196 4452
rect 35252 4396 36204 4452
rect 36260 4396 36540 4452
rect 36596 4396 36606 4452
rect 40226 4396 40236 4452
rect 40292 4396 41356 4452
rect 41412 4396 41692 4452
rect 41748 4396 41758 4452
rect 43474 4396 43484 4452
rect 43540 4396 45612 4452
rect 45668 4396 45678 4452
rect 51090 4396 51100 4452
rect 51156 4396 51436 4452
rect 51492 4396 52220 4452
rect 52276 4396 52286 4452
rect 33068 4340 33124 4396
rect 1698 4284 1708 4340
rect 1764 4284 6300 4340
rect 6356 4284 6366 4340
rect 7634 4284 7644 4340
rect 7700 4284 31052 4340
rect 31108 4284 31118 4340
rect 31714 4284 31724 4340
rect 31780 4284 33124 4340
rect 33282 4284 33292 4340
rect 33348 4284 35980 4340
rect 36036 4284 36046 4340
rect 36642 4284 36652 4340
rect 36708 4284 54236 4340
rect 54292 4284 54302 4340
rect 5730 4172 5740 4228
rect 5796 4172 10220 4228
rect 10276 4172 10286 4228
rect 10658 4172 10668 4228
rect 10724 4172 12572 4228
rect 12628 4172 12638 4228
rect 13122 4172 13132 4228
rect 13188 4172 15316 4228
rect 15474 4172 15484 4228
rect 15540 4172 20412 4228
rect 20468 4172 20478 4228
rect 21074 4172 21084 4228
rect 21140 4172 25228 4228
rect 25284 4172 25294 4228
rect 27234 4172 27244 4228
rect 27300 4172 27804 4228
rect 27860 4172 27870 4228
rect 28578 4172 28588 4228
rect 28644 4172 37324 4228
rect 37380 4172 37390 4228
rect 38658 4172 38668 4228
rect 38724 4172 48300 4228
rect 48356 4172 48366 4228
rect 48514 4172 48524 4228
rect 48580 4172 51436 4228
rect 51492 4172 51502 4228
rect 0 4116 112 4144
rect 15260 4116 15316 4172
rect 57344 4116 57456 4144
rect 0 4060 3276 4116
rect 3332 4060 3342 4116
rect 4386 4060 4396 4116
rect 4452 4060 4900 4116
rect 6178 4060 6188 4116
rect 6244 4060 15036 4116
rect 15092 4060 15102 4116
rect 15260 4060 20356 4116
rect 20962 4060 20972 4116
rect 21028 4060 28588 4116
rect 28644 4060 28654 4116
rect 28802 4060 28812 4116
rect 28868 4060 30716 4116
rect 30772 4060 30782 4116
rect 30930 4060 30940 4116
rect 30996 4060 35476 4116
rect 0 4032 112 4060
rect 4844 4004 4900 4060
rect 20300 4004 20356 4060
rect 35420 4004 35476 4060
rect 35980 4060 41020 4116
rect 41076 4060 41086 4116
rect 41682 4060 41692 4116
rect 41748 4060 44884 4116
rect 45378 4060 45388 4116
rect 45444 4060 48972 4116
rect 49028 4060 49308 4116
rect 49364 4060 49374 4116
rect 56130 4060 56140 4116
rect 56196 4060 57456 4116
rect 35980 4004 36036 4060
rect 44828 4004 44884 4060
rect 57344 4032 57456 4060
rect 4844 3948 9996 4004
rect 10052 3948 10062 4004
rect 11778 3948 11788 4004
rect 11844 3948 20076 4004
rect 20132 3948 20142 4004
rect 20300 3948 24220 4004
rect 24276 3948 24286 4004
rect 25330 3948 25340 4004
rect 25396 3948 35196 4004
rect 35252 3948 35262 4004
rect 35420 3948 36036 4004
rect 36194 3948 36204 4004
rect 36260 3948 40012 4004
rect 40068 3948 40078 4004
rect 44828 3948 45388 4004
rect 45444 3948 45454 4004
rect 4454 3892 4464 3948
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4728 3892 4738 3948
rect 24454 3892 24464 3948
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24728 3892 24738 3948
rect 44454 3892 44464 3948
rect 44520 3892 44568 3948
rect 44624 3892 44672 3948
rect 44728 3892 44738 3948
rect 8418 3836 8428 3892
rect 8484 3836 13244 3892
rect 13300 3836 13310 3892
rect 13458 3836 13468 3892
rect 13524 3836 14980 3892
rect 15138 3836 15148 3892
rect 15204 3836 15820 3892
rect 15876 3836 15886 3892
rect 16482 3836 16492 3892
rect 16548 3836 23660 3892
rect 23716 3836 23726 3892
rect 25778 3836 25788 3892
rect 25844 3836 35308 3892
rect 35364 3836 35374 3892
rect 42354 3836 42364 3892
rect 42420 3836 43708 3892
rect 43764 3836 43774 3892
rect 45154 3836 45164 3892
rect 45220 3836 52556 3892
rect 52612 3836 52622 3892
rect 14924 3780 14980 3836
rect 1138 3724 1148 3780
rect 1204 3724 6076 3780
rect 6132 3724 6142 3780
rect 8838 3724 8876 3780
rect 8932 3724 8942 3780
rect 12114 3724 12124 3780
rect 12180 3724 14700 3780
rect 14756 3724 14766 3780
rect 14924 3724 37100 3780
rect 37156 3724 37166 3780
rect 37314 3724 37324 3780
rect 37380 3724 55132 3780
rect 55188 3724 55198 3780
rect 0 3668 112 3696
rect 57344 3668 57456 3696
rect 0 3612 588 3668
rect 644 3612 654 3668
rect 3332 3612 12348 3668
rect 12404 3612 12414 3668
rect 12562 3612 12572 3668
rect 12628 3612 13244 3668
rect 13300 3612 13310 3668
rect 14018 3612 14028 3668
rect 14084 3612 19460 3668
rect 19618 3612 19628 3668
rect 19684 3612 25340 3668
rect 25396 3612 25406 3668
rect 25554 3612 25564 3668
rect 25620 3612 27300 3668
rect 27570 3612 27580 3668
rect 27636 3612 41916 3668
rect 41972 3612 41982 3668
rect 42242 3612 42252 3668
rect 42308 3612 53564 3668
rect 53620 3612 53630 3668
rect 54898 3612 54908 3668
rect 54964 3612 57456 3668
rect 0 3584 112 3612
rect 3332 3444 3388 3612
rect 19404 3556 19460 3612
rect 27244 3556 27300 3612
rect 57344 3584 57456 3612
rect 6626 3500 6636 3556
rect 6692 3500 9380 3556
rect 9538 3500 9548 3556
rect 9604 3500 13916 3556
rect 13972 3500 13982 3556
rect 14130 3500 14140 3556
rect 14196 3500 16156 3556
rect 16212 3500 16222 3556
rect 16370 3500 16380 3556
rect 16436 3500 18396 3556
rect 18452 3500 18462 3556
rect 19404 3500 20300 3556
rect 20356 3500 20366 3556
rect 23650 3500 23660 3556
rect 23716 3500 27020 3556
rect 27076 3500 27086 3556
rect 27244 3500 33516 3556
rect 33572 3500 33582 3556
rect 33740 3500 41692 3556
rect 41748 3500 41758 3556
rect 41916 3500 45332 3556
rect 9324 3444 9380 3500
rect 33740 3444 33796 3500
rect 41916 3444 41972 3500
rect 1026 3388 1036 3444
rect 1092 3388 3388 3444
rect 6626 3388 6636 3444
rect 6692 3388 8428 3444
rect 9324 3388 10668 3444
rect 10724 3388 10734 3444
rect 10994 3388 11004 3444
rect 11060 3388 13356 3444
rect 13412 3388 13422 3444
rect 13580 3388 16604 3444
rect 16660 3388 16670 3444
rect 16940 3388 17836 3444
rect 17892 3388 17902 3444
rect 19170 3388 19180 3444
rect 19236 3388 21812 3444
rect 3612 3276 6748 3332
rect 6804 3276 6814 3332
rect 0 3220 112 3248
rect 3612 3220 3668 3276
rect 0 3164 3668 3220
rect 8372 3220 8428 3388
rect 13580 3332 13636 3388
rect 8754 3276 8764 3332
rect 8820 3276 11116 3332
rect 11172 3276 11182 3332
rect 12786 3276 12796 3332
rect 12852 3276 13636 3332
rect 15474 3276 15484 3332
rect 15540 3276 16716 3332
rect 16772 3276 16782 3332
rect 16940 3220 16996 3388
rect 21756 3332 21812 3388
rect 22092 3388 30268 3444
rect 30324 3388 30334 3444
rect 30482 3388 30492 3444
rect 30548 3388 30940 3444
rect 30996 3388 31006 3444
rect 31154 3388 31164 3444
rect 31220 3388 33796 3444
rect 36866 3388 36876 3444
rect 36932 3388 41972 3444
rect 42354 3388 42364 3444
rect 42420 3388 44380 3444
rect 44436 3388 44446 3444
rect 22092 3332 22148 3388
rect 45276 3332 45332 3500
rect 53554 3388 53564 3444
rect 53620 3388 56812 3444
rect 56868 3388 56878 3444
rect 21746 3276 21756 3332
rect 21812 3276 21822 3332
rect 22082 3276 22092 3332
rect 22148 3276 22158 3332
rect 22754 3276 22764 3332
rect 22820 3276 25788 3332
rect 25844 3276 25854 3332
rect 26114 3276 26124 3332
rect 26180 3276 28588 3332
rect 28644 3276 28654 3332
rect 29362 3276 29372 3332
rect 29428 3276 30044 3332
rect 30100 3276 30110 3332
rect 30258 3276 30268 3332
rect 30324 3276 31052 3332
rect 31108 3276 31118 3332
rect 33618 3276 33628 3332
rect 33684 3276 38220 3332
rect 38276 3276 38286 3332
rect 38612 3276 43484 3332
rect 43540 3276 43550 3332
rect 45276 3276 49756 3332
rect 49812 3276 49822 3332
rect 38612 3220 38668 3276
rect 57344 3220 57456 3248
rect 8372 3164 16996 3220
rect 17154 3164 17164 3220
rect 17220 3164 19124 3220
rect 23622 3164 23660 3220
rect 23716 3164 23726 3220
rect 25218 3164 25228 3220
rect 25284 3164 28252 3220
rect 28308 3164 28318 3220
rect 33506 3164 33516 3220
rect 33572 3164 38668 3220
rect 45826 3164 45836 3220
rect 45892 3164 51324 3220
rect 51380 3164 51390 3220
rect 54562 3164 54572 3220
rect 54628 3164 57456 3220
rect 0 3136 112 3164
rect 3794 3108 3804 3164
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 4068 3108 4078 3164
rect 19068 3108 19124 3164
rect 23794 3108 23804 3164
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 24068 3108 24078 3164
rect 43794 3108 43804 3164
rect 43860 3108 43908 3164
rect 43964 3108 44012 3164
rect 44068 3108 44078 3164
rect 57344 3136 57456 3164
rect 4162 3052 4172 3108
rect 4228 3052 13356 3108
rect 13412 3052 13422 3108
rect 13682 3052 13692 3108
rect 13748 3052 18844 3108
rect 18900 3052 18910 3108
rect 19068 3052 21868 3108
rect 21924 3052 21934 3108
rect 23510 3052 23548 3108
rect 23604 3052 23614 3108
rect 24210 3052 24220 3108
rect 24276 3052 43596 3108
rect 43652 3052 43662 3108
rect 45938 3052 45948 3108
rect 46004 3052 52220 3108
rect 52276 3052 52286 3108
rect 1586 2940 1596 2996
rect 1652 2940 11676 2996
rect 11732 2940 11742 2996
rect 12338 2940 12348 2996
rect 12404 2940 18284 2996
rect 18340 2940 18350 2996
rect 20178 2940 20188 2996
rect 20244 2940 21420 2996
rect 21476 2940 21486 2996
rect 21746 2940 21756 2996
rect 21812 2940 26124 2996
rect 26180 2940 26190 2996
rect 26338 2940 26348 2996
rect 26404 2940 26908 2996
rect 26964 2940 26974 2996
rect 27122 2940 27132 2996
rect 27188 2940 28364 2996
rect 28420 2940 28430 2996
rect 28578 2940 28588 2996
rect 28644 2940 34972 2996
rect 35028 2940 35038 2996
rect 35298 2940 35308 2996
rect 35364 2940 36652 2996
rect 36708 2940 36718 2996
rect 42242 2940 42252 2996
rect 42308 2940 45500 2996
rect 45556 2940 45566 2996
rect 47618 2940 47628 2996
rect 47684 2940 52556 2996
rect 52612 2940 52622 2996
rect 3266 2828 3276 2884
rect 3332 2828 9324 2884
rect 9380 2828 9390 2884
rect 13122 2828 13132 2884
rect 13188 2828 13580 2884
rect 13636 2828 13646 2884
rect 14018 2828 14028 2884
rect 14084 2828 19404 2884
rect 19460 2828 19470 2884
rect 20402 2828 20412 2884
rect 20468 2828 27244 2884
rect 27300 2828 27310 2884
rect 28130 2828 28140 2884
rect 28196 2828 28812 2884
rect 28868 2828 28878 2884
rect 29026 2828 29036 2884
rect 29092 2828 29260 2884
rect 29316 2828 30716 2884
rect 30772 2828 30782 2884
rect 31042 2828 31052 2884
rect 31108 2828 32900 2884
rect 33058 2828 33068 2884
rect 33124 2828 34076 2884
rect 34132 2828 34142 2884
rect 35186 2828 35196 2884
rect 35252 2828 37660 2884
rect 37716 2828 37726 2884
rect 42018 2828 42028 2884
rect 42084 2828 45276 2884
rect 45332 2828 45342 2884
rect 0 2772 112 2800
rect 32844 2772 32900 2828
rect 57344 2772 57456 2800
rect 0 2716 8316 2772
rect 8372 2716 8382 2772
rect 10882 2716 10892 2772
rect 10948 2716 24892 2772
rect 24948 2716 24958 2772
rect 25116 2716 29708 2772
rect 29764 2716 29774 2772
rect 30594 2716 30604 2772
rect 30660 2716 31276 2772
rect 31332 2716 31342 2772
rect 31938 2716 31948 2772
rect 32004 2716 32396 2772
rect 32452 2716 32620 2772
rect 32676 2716 32686 2772
rect 32844 2716 40572 2772
rect 40628 2716 40638 2772
rect 49634 2716 49644 2772
rect 49700 2716 53564 2772
rect 53620 2716 53630 2772
rect 56130 2716 56140 2772
rect 56196 2716 57456 2772
rect 0 2688 112 2716
rect 25116 2660 25172 2716
rect 57344 2688 57456 2716
rect 3826 2604 3836 2660
rect 3892 2604 6748 2660
rect 6804 2604 6814 2660
rect 7410 2604 7420 2660
rect 7476 2604 16044 2660
rect 16100 2604 16110 2660
rect 16930 2604 16940 2660
rect 16996 2604 19628 2660
rect 19684 2604 19694 2660
rect 19852 2604 25172 2660
rect 26002 2604 26012 2660
rect 26068 2604 27692 2660
rect 27748 2604 27758 2660
rect 28466 2604 28476 2660
rect 28532 2604 35868 2660
rect 35924 2604 35934 2660
rect 36092 2604 38332 2660
rect 38388 2604 38398 2660
rect 40338 2604 40348 2660
rect 40404 2604 47740 2660
rect 47796 2604 47806 2660
rect 52770 2604 52780 2660
rect 52836 2604 56476 2660
rect 56532 2604 56542 2660
rect 19852 2548 19908 2604
rect 36092 2548 36148 2604
rect 2482 2492 2492 2548
rect 2548 2492 4172 2548
rect 4228 2492 4238 2548
rect 4386 2492 4396 2548
rect 4452 2492 4956 2548
rect 5012 2492 5022 2548
rect 13234 2492 13244 2548
rect 13300 2492 16828 2548
rect 16884 2492 16894 2548
rect 18722 2492 18732 2548
rect 18788 2492 19908 2548
rect 20636 2492 25228 2548
rect 25284 2492 25294 2548
rect 25442 2492 25452 2548
rect 25508 2492 28252 2548
rect 28308 2492 28318 2548
rect 28690 2492 28700 2548
rect 28756 2492 28794 2548
rect 29362 2492 29372 2548
rect 29428 2492 36148 2548
rect 38434 2492 38444 2548
rect 38500 2492 54124 2548
rect 54180 2492 54190 2548
rect 20636 2436 20692 2492
rect 13122 2380 13132 2436
rect 13188 2380 13692 2436
rect 13748 2380 13758 2436
rect 14130 2380 14140 2436
rect 14196 2380 20692 2436
rect 21858 2380 21868 2436
rect 21924 2380 24220 2436
rect 24276 2380 24286 2436
rect 25330 2380 25340 2436
rect 25396 2380 32396 2436
rect 32452 2380 32462 2436
rect 32834 2380 32844 2436
rect 32900 2380 33348 2436
rect 34178 2380 34188 2436
rect 34244 2380 41804 2436
rect 41860 2380 41870 2436
rect 52210 2380 52220 2436
rect 52276 2380 55244 2436
rect 55300 2380 55310 2436
rect 0 2324 112 2352
rect 4454 2324 4464 2380
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4728 2324 4738 2380
rect 24454 2324 24464 2380
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24728 2324 24738 2380
rect 33292 2324 33348 2380
rect 44454 2324 44464 2380
rect 44520 2324 44568 2380
rect 44624 2324 44672 2380
rect 44728 2324 44738 2380
rect 57344 2324 57456 2352
rect 0 2268 3220 2324
rect 13346 2268 13356 2324
rect 13412 2268 19292 2324
rect 19348 2268 19358 2324
rect 20178 2268 20188 2324
rect 20244 2268 21196 2324
rect 21252 2268 21262 2324
rect 21410 2268 21420 2324
rect 21476 2268 24332 2324
rect 24388 2268 24398 2324
rect 24882 2268 24892 2324
rect 24948 2268 32956 2324
rect 33012 2268 33022 2324
rect 33292 2268 35308 2324
rect 35364 2268 35374 2324
rect 35746 2268 35756 2324
rect 35812 2268 42364 2324
rect 42420 2268 42430 2324
rect 54898 2268 54908 2324
rect 54964 2268 57456 2324
rect 0 2240 112 2268
rect 0 1876 112 1904
rect 0 1820 2716 1876
rect 2772 1820 2782 1876
rect 0 1792 112 1820
rect 3164 1764 3220 2268
rect 57344 2240 57456 2268
rect 14242 2156 14252 2212
rect 14308 2156 14588 2212
rect 14644 2156 20972 2212
rect 21028 2156 21038 2212
rect 21196 2156 26348 2212
rect 26404 2156 26414 2212
rect 26562 2156 26572 2212
rect 26628 2156 28364 2212
rect 28420 2156 28430 2212
rect 28578 2156 28588 2212
rect 28644 2156 30940 2212
rect 30996 2156 31006 2212
rect 32386 2156 32396 2212
rect 32452 2156 41916 2212
rect 41972 2156 41982 2212
rect 43652 2156 52444 2212
rect 52500 2156 52510 2212
rect 8082 2044 8092 2100
rect 8148 2044 20748 2100
rect 20804 2044 20814 2100
rect 21196 1988 21252 2156
rect 22092 2044 24892 2100
rect 24948 2044 24958 2100
rect 25106 2044 25116 2100
rect 25172 2044 28028 2100
rect 28084 2044 28094 2100
rect 28242 2044 28252 2100
rect 28308 2044 36876 2100
rect 36932 2044 36942 2100
rect 38658 2044 38668 2100
rect 38724 2044 43036 2100
rect 43092 2044 43102 2100
rect 22092 1988 22148 2044
rect 43652 1988 43708 2156
rect 3378 1932 3388 1988
rect 3444 1932 3724 1988
rect 3780 1932 16492 1988
rect 16548 1932 16558 1988
rect 16930 1932 16940 1988
rect 16996 1932 21252 1988
rect 21522 1932 21532 1988
rect 21588 1932 22148 1988
rect 23762 1932 23772 1988
rect 23828 1932 29820 1988
rect 29876 1932 29886 1988
rect 30370 1932 30380 1988
rect 30436 1932 43708 1988
rect 43820 2044 52108 2100
rect 52164 2044 52174 2100
rect 43820 1876 43876 2044
rect 57344 1876 57456 1904
rect 6514 1820 6524 1876
rect 6580 1820 13356 1876
rect 13412 1820 13422 1876
rect 13906 1820 13916 1876
rect 13972 1820 17220 1876
rect 17378 1820 17388 1876
rect 17444 1820 23548 1876
rect 3164 1708 14252 1764
rect 14308 1708 14318 1764
rect 14802 1708 14812 1764
rect 14868 1708 16940 1764
rect 16996 1708 17006 1764
rect 17164 1652 17220 1820
rect 23492 1764 23548 1820
rect 23660 1820 43876 1876
rect 44258 1820 44268 1876
rect 44324 1820 52108 1876
rect 52164 1820 52174 1876
rect 53554 1820 53564 1876
rect 53620 1820 57456 1876
rect 23660 1764 23716 1820
rect 57344 1792 57456 1820
rect 20850 1708 20860 1764
rect 20916 1708 21644 1764
rect 21700 1708 21710 1764
rect 23492 1708 23716 1764
rect 23874 1708 23884 1764
rect 23940 1708 24500 1764
rect 24658 1708 24668 1764
rect 24724 1708 25060 1764
rect 25218 1708 25228 1764
rect 25284 1708 30604 1764
rect 30660 1708 30670 1764
rect 30940 1708 36092 1764
rect 36148 1708 36158 1764
rect 36316 1708 38556 1764
rect 38612 1708 38622 1764
rect 40226 1708 40236 1764
rect 40292 1708 45108 1764
rect 45266 1708 45276 1764
rect 45332 1708 51436 1764
rect 51492 1708 51502 1764
rect 5058 1596 5068 1652
rect 5124 1596 7196 1652
rect 7252 1596 7262 1652
rect 10546 1596 10556 1652
rect 10612 1596 16940 1652
rect 16996 1596 17006 1652
rect 17164 1596 23324 1652
rect 23380 1596 23390 1652
rect 23492 1596 23660 1652
rect 23716 1596 23726 1652
rect 3794 1540 3804 1596
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 4068 1540 4078 1596
rect 23492 1540 23548 1596
rect 23794 1540 23804 1596
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 24068 1540 24078 1596
rect 24444 1540 24500 1708
rect 25004 1652 25060 1708
rect 30940 1652 30996 1708
rect 36316 1652 36372 1708
rect 45052 1652 45108 1708
rect 25004 1596 27020 1652
rect 27076 1596 27086 1652
rect 27234 1596 27244 1652
rect 27300 1596 30996 1652
rect 31154 1596 31164 1652
rect 31220 1596 34076 1652
rect 34132 1596 34142 1652
rect 34412 1596 36372 1652
rect 37538 1596 37548 1652
rect 37604 1596 42252 1652
rect 42308 1596 42318 1652
rect 45052 1596 45556 1652
rect 47506 1596 47516 1652
rect 47572 1596 51100 1652
rect 51156 1596 51166 1652
rect 34412 1540 34468 1596
rect 43794 1540 43804 1596
rect 43860 1540 43908 1596
rect 43964 1540 44012 1596
rect 44068 1540 44078 1596
rect 45500 1540 45556 1596
rect 4172 1484 9548 1540
rect 9604 1484 9614 1540
rect 11106 1484 11116 1540
rect 11172 1484 14476 1540
rect 14532 1484 14542 1540
rect 15092 1484 18172 1540
rect 18228 1484 18238 1540
rect 20290 1484 20300 1540
rect 20356 1484 23548 1540
rect 24444 1484 29372 1540
rect 29428 1484 29438 1540
rect 29586 1484 29596 1540
rect 29652 1484 30772 1540
rect 31826 1484 31836 1540
rect 31892 1484 34468 1540
rect 34626 1484 34636 1540
rect 34692 1484 38668 1540
rect 38724 1484 38734 1540
rect 38882 1484 38892 1540
rect 38948 1484 40236 1540
rect 40292 1484 40302 1540
rect 45500 1484 47628 1540
rect 47684 1484 47694 1540
rect 49420 1484 55132 1540
rect 55188 1484 55198 1540
rect 0 1428 112 1456
rect 4172 1428 4228 1484
rect 15092 1428 15148 1484
rect 30716 1428 30772 1484
rect 49420 1428 49476 1484
rect 57344 1428 57456 1456
rect 0 1372 4228 1428
rect 6738 1372 6748 1428
rect 6804 1372 8428 1428
rect 8642 1372 8652 1428
rect 8708 1372 14028 1428
rect 14084 1372 14094 1428
rect 14242 1372 14252 1428
rect 14308 1372 15148 1428
rect 16034 1372 16044 1428
rect 16100 1372 16660 1428
rect 16818 1372 16828 1428
rect 16884 1372 23548 1428
rect 23604 1372 23614 1428
rect 24434 1372 24444 1428
rect 24500 1372 25676 1428
rect 25732 1372 25742 1428
rect 26852 1372 30492 1428
rect 30548 1372 30558 1428
rect 30716 1372 40348 1428
rect 40404 1372 40414 1428
rect 41234 1372 41244 1428
rect 41300 1372 49476 1428
rect 53554 1372 53564 1428
rect 53620 1372 57456 1428
rect 0 1344 112 1372
rect 8372 1316 8428 1372
rect 16604 1316 16660 1372
rect 26852 1316 26908 1372
rect 57344 1344 57456 1372
rect 2482 1260 2492 1316
rect 2548 1260 2828 1316
rect 2884 1260 7420 1316
rect 7476 1260 7486 1316
rect 8372 1260 16380 1316
rect 16436 1260 16446 1316
rect 16604 1260 20748 1316
rect 20804 1260 20814 1316
rect 20962 1260 20972 1316
rect 21028 1260 26908 1316
rect 27122 1260 27132 1316
rect 27188 1260 38892 1316
rect 38948 1260 38958 1316
rect 39442 1260 39452 1316
rect 39508 1260 46620 1316
rect 46676 1260 46686 1316
rect 47282 1260 47292 1316
rect 47348 1260 52556 1316
rect 52612 1260 52622 1316
rect 5842 1148 5852 1204
rect 5908 1148 21308 1204
rect 21364 1148 21374 1204
rect 21522 1148 21532 1204
rect 21588 1148 23996 1204
rect 24052 1148 24062 1204
rect 24210 1148 24220 1204
rect 24276 1148 26908 1204
rect 26964 1148 26974 1204
rect 27122 1148 27132 1204
rect 27188 1148 27804 1204
rect 27860 1148 27870 1204
rect 28018 1148 28028 1204
rect 28084 1148 32508 1204
rect 32564 1148 32574 1204
rect 32722 1148 32732 1204
rect 32788 1148 45836 1204
rect 45892 1148 45902 1204
rect 46050 1148 46060 1204
rect 46116 1148 52332 1204
rect 52388 1148 52398 1204
rect 1810 1036 1820 1092
rect 1876 1036 21084 1092
rect 21140 1036 21150 1092
rect 21298 1036 21308 1092
rect 21364 1036 25452 1092
rect 25508 1036 25518 1092
rect 25666 1036 25676 1092
rect 25732 1036 28588 1092
rect 28644 1036 28654 1092
rect 28802 1036 28812 1092
rect 28868 1036 31836 1092
rect 31892 1036 31902 1092
rect 32050 1036 32060 1092
rect 32116 1036 33012 1092
rect 33170 1036 33180 1092
rect 33236 1036 37100 1092
rect 37156 1036 37166 1092
rect 42018 1036 42028 1092
rect 42084 1036 44828 1092
rect 44884 1036 44894 1092
rect 0 980 112 1008
rect 32956 980 33012 1036
rect 57344 980 57456 1008
rect 0 924 1036 980
rect 1092 924 1102 980
rect 1250 924 1260 980
rect 1316 924 4900 980
rect 13906 924 13916 980
rect 13972 924 20636 980
rect 20692 924 20702 980
rect 20850 924 20860 980
rect 20916 924 23324 980
rect 23380 924 23390 980
rect 23538 924 23548 980
rect 23604 924 32788 980
rect 32956 924 48860 980
rect 48916 924 48926 980
rect 51986 924 51996 980
rect 52052 924 57456 980
rect 0 896 112 924
rect 4454 756 4464 812
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4728 756 4738 812
rect 4844 756 4900 924
rect 6402 812 6412 868
rect 6468 812 14140 868
rect 14196 812 14206 868
rect 14466 812 14476 868
rect 14532 812 15148 868
rect 15204 812 15214 868
rect 16930 812 16940 868
rect 16996 812 21308 868
rect 21364 812 21374 868
rect 21634 812 21644 868
rect 21700 812 24332 868
rect 24388 812 24398 868
rect 24882 812 24892 868
rect 24948 812 26684 868
rect 26740 812 26750 868
rect 26898 812 26908 868
rect 26964 812 32508 868
rect 32564 812 32574 868
rect 24454 756 24464 812
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24728 756 24738 812
rect 4844 700 23324 756
rect 23380 700 23390 756
rect 23538 700 23548 756
rect 23604 700 24220 756
rect 24276 700 24286 756
rect 24994 700 25004 756
rect 25060 700 25340 756
rect 25396 700 25406 756
rect 25676 700 32172 756
rect 32228 700 32238 756
rect 4498 588 4508 644
rect 4564 588 5404 644
rect 5460 588 5470 644
rect 7858 588 7868 644
rect 7924 588 13132 644
rect 13188 588 13198 644
rect 13346 588 13356 644
rect 13412 588 25228 644
rect 25284 588 25294 644
rect 0 532 112 560
rect 25676 532 25732 700
rect 32732 644 32788 924
rect 57344 896 57456 924
rect 34300 812 34972 868
rect 35028 812 35038 868
rect 36978 812 36988 868
rect 37044 812 44268 868
rect 44324 812 44334 868
rect 44930 812 44940 868
rect 44996 812 52892 868
rect 52948 812 52958 868
rect 34300 756 34356 812
rect 44454 756 44464 812
rect 44520 756 44568 812
rect 44624 756 44672 812
rect 44728 756 44738 812
rect 33058 700 33068 756
rect 33124 700 34356 756
rect 34514 700 34524 756
rect 34580 700 40684 756
rect 40740 700 40750 756
rect 48290 700 48300 756
rect 48356 700 55580 756
rect 55636 700 55646 756
rect 25890 588 25900 644
rect 25956 588 28140 644
rect 28196 588 28206 644
rect 28354 588 28364 644
rect 28420 588 32676 644
rect 32732 588 46396 644
rect 46452 588 46462 644
rect 32620 532 32676 588
rect 57344 532 57456 560
rect 0 476 1596 532
rect 1652 476 1662 532
rect 13570 476 13580 532
rect 13636 476 19796 532
rect 19954 476 19964 532
rect 20020 476 23212 532
rect 23268 476 23278 532
rect 23426 476 23436 532
rect 23492 476 25732 532
rect 26786 476 26796 532
rect 26852 476 32396 532
rect 32452 476 32462 532
rect 32620 476 40236 532
rect 40292 476 40302 532
rect 40450 476 40460 532
rect 40516 476 52220 532
rect 52276 476 52286 532
rect 56802 476 56812 532
rect 56868 476 57456 532
rect 0 448 112 476
rect 19740 420 19796 476
rect 57344 448 57456 476
rect 10770 364 10780 420
rect 10836 364 17948 420
rect 18004 364 18014 420
rect 19740 364 27020 420
rect 27076 364 27086 420
rect 27234 364 27244 420
rect 27300 364 27916 420
rect 27972 364 27982 420
rect 28130 364 28140 420
rect 28196 364 32620 420
rect 32676 364 32686 420
rect 32834 364 32844 420
rect 32900 364 36764 420
rect 36820 364 36830 420
rect 40460 364 46172 420
rect 46228 364 46238 420
rect 40460 308 40516 364
rect 16146 252 16156 308
rect 16212 252 21532 308
rect 21588 252 21598 308
rect 22418 252 22428 308
rect 22484 252 26796 308
rect 26852 252 26862 308
rect 27010 252 27020 308
rect 27076 252 34748 308
rect 34804 252 34814 308
rect 34962 252 34972 308
rect 35028 252 40516 308
rect 40674 252 40684 308
rect 40740 252 45276 308
rect 45332 252 45342 308
rect 1362 140 1372 196
rect 1428 140 1820 196
rect 1876 140 1886 196
rect 14354 140 14364 196
rect 14420 140 31388 196
rect 31444 140 31454 196
rect 32274 140 32284 196
rect 32340 140 40460 196
rect 40516 140 40526 196
rect 49410 140 49420 196
rect 49476 140 50204 196
rect 50260 140 50270 196
rect 0 84 112 112
rect 57344 84 57456 112
rect 0 28 1148 84
rect 1204 28 1214 84
rect 15138 28 15148 84
rect 15204 28 19964 84
rect 20020 28 20030 84
rect 21298 28 21308 84
rect 21364 28 26012 84
rect 26068 28 26078 84
rect 27906 28 27916 84
rect 27972 28 36988 84
rect 37044 28 37054 84
rect 56466 28 56476 84
rect 56532 28 57456 84
rect 0 0 112 28
rect 57344 0 57456 28
<< via3 >>
rect 10220 14140 10276 14196
rect 20972 14140 21028 14196
rect 21196 14140 21252 14196
rect 29484 14140 29540 14196
rect 32060 14140 32116 14196
rect 35420 14140 35476 14196
rect 20972 13916 21028 13972
rect 24892 13804 24948 13860
rect 35420 13804 35476 13860
rect 25116 13692 25172 13748
rect 30156 13692 30212 13748
rect 36316 13692 36372 13748
rect 24220 13580 24276 13636
rect 1596 13468 1652 13524
rect 31164 13468 31220 13524
rect 25004 13356 25060 13412
rect 4464 13300 4520 13356
rect 4568 13300 4624 13356
rect 4672 13300 4728 13356
rect 24464 13300 24520 13356
rect 24568 13300 24624 13356
rect 24672 13300 24728 13356
rect 44464 13300 44520 13356
rect 44568 13300 44624 13356
rect 44672 13300 44728 13356
rect 18620 13244 18676 13300
rect 19852 13132 19908 13188
rect 31052 13020 31108 13076
rect 32508 13020 32564 13076
rect 16940 12796 16996 12852
rect 18620 12796 18676 12852
rect 29484 12796 29540 12852
rect 30940 12796 30996 12852
rect 31164 12796 31220 12852
rect 31836 12796 31892 12852
rect 39788 12796 39844 12852
rect 24892 12684 24948 12740
rect 38892 12684 38948 12740
rect 3804 12516 3860 12572
rect 3908 12516 3964 12572
rect 4012 12516 4068 12572
rect 23804 12516 23860 12572
rect 23908 12516 23964 12572
rect 24012 12516 24068 12572
rect 43804 12516 43860 12572
rect 43908 12516 43964 12572
rect 44012 12516 44068 12572
rect 38780 12460 38836 12516
rect 39788 12460 39844 12516
rect 43484 12460 43540 12516
rect 21196 12348 21252 12404
rect 28028 12348 28084 12404
rect 36316 12348 36372 12404
rect 39004 12348 39060 12404
rect 15708 12236 15764 12292
rect 16156 12236 16212 12292
rect 28588 12236 28644 12292
rect 17500 12124 17556 12180
rect 1596 11900 1652 11956
rect 15148 11900 15204 11956
rect 15484 11900 15540 11956
rect 15372 11788 15428 11844
rect 22092 11788 22148 11844
rect 30940 11788 30996 11844
rect 4464 11732 4520 11788
rect 4568 11732 4624 11788
rect 4672 11732 4728 11788
rect 4284 11676 4340 11732
rect 24464 11732 24520 11788
rect 24568 11732 24624 11788
rect 24672 11732 24728 11788
rect 44464 11732 44520 11788
rect 44568 11732 44624 11788
rect 44672 11732 44728 11788
rect 21532 11676 21588 11732
rect 24220 11676 24276 11732
rect 38892 11676 38948 11732
rect 44268 11676 44324 11732
rect 51100 11676 51156 11732
rect 14588 11564 14644 11620
rect 15484 11564 15540 11620
rect 19068 11564 19124 11620
rect 21644 11564 21700 11620
rect 26124 11564 26180 11620
rect 31836 11564 31892 11620
rect 33180 11564 33236 11620
rect 43484 11564 43540 11620
rect 14700 11452 14756 11508
rect 44268 11452 44324 11508
rect 4284 11340 4340 11396
rect 15148 11340 15204 11396
rect 26124 11340 26180 11396
rect 10108 11228 10164 11284
rect 17052 11228 17108 11284
rect 33852 11228 33908 11284
rect 6636 11116 6692 11172
rect 21532 11116 21588 11172
rect 38892 11116 38948 11172
rect 19068 11004 19124 11060
rect 20412 11004 20468 11060
rect 22092 11004 22148 11060
rect 28700 11004 28756 11060
rect 30828 11004 30884 11060
rect 31052 11004 31108 11060
rect 41916 11004 41972 11060
rect 3804 10948 3860 11004
rect 3908 10948 3964 11004
rect 4012 10948 4068 11004
rect 23804 10948 23860 11004
rect 23908 10948 23964 11004
rect 24012 10948 24068 11004
rect 43804 10948 43860 11004
rect 43908 10948 43964 11004
rect 44012 10948 44068 11004
rect 26572 10892 26628 10948
rect 26908 10892 26964 10948
rect 30156 10892 30212 10948
rect 30380 10892 30436 10948
rect 32732 10780 32788 10836
rect 39564 10780 39620 10836
rect 22092 10668 22148 10724
rect 27132 10668 27188 10724
rect 31276 10668 31332 10724
rect 34076 10668 34132 10724
rect 26460 10556 26516 10612
rect 22316 10444 22372 10500
rect 27356 10444 27412 10500
rect 32732 10444 32788 10500
rect 40236 10444 40292 10500
rect 7308 10332 7364 10388
rect 22204 10332 22260 10388
rect 26852 10332 26908 10388
rect 39564 10332 39620 10388
rect 20188 10220 20244 10276
rect 21980 10220 22036 10276
rect 4464 10164 4520 10220
rect 4568 10164 4624 10220
rect 4672 10164 4728 10220
rect 24464 10164 24520 10220
rect 24568 10164 24624 10220
rect 24672 10164 24728 10220
rect 20300 10108 20356 10164
rect 24220 10108 24276 10164
rect 27916 10108 27972 10164
rect 31836 10108 31892 10164
rect 32060 10108 32116 10164
rect 35644 10108 35700 10164
rect 14476 9996 14532 10052
rect 18172 9996 18228 10052
rect 28588 9996 28644 10052
rect 31388 9996 31444 10052
rect 37324 9996 37380 10052
rect 44464 10164 44520 10220
rect 44568 10164 44624 10220
rect 44672 10164 44728 10220
rect 10108 9884 10164 9940
rect 15260 9884 15316 9940
rect 25228 9884 25284 9940
rect 40236 9884 40292 9940
rect 14588 9772 14644 9828
rect 15148 9772 15204 9828
rect 21756 9772 21812 9828
rect 21980 9772 22036 9828
rect 25004 9772 25060 9828
rect 36876 9772 36932 9828
rect 40572 9772 40628 9828
rect 10220 9660 10276 9716
rect 28700 9660 28756 9716
rect 15708 9548 15764 9604
rect 18172 9548 18228 9604
rect 29820 9548 29876 9604
rect 30828 9548 30884 9604
rect 31052 9548 31108 9604
rect 35644 9548 35700 9604
rect 37884 9548 37940 9604
rect 14476 9436 14532 9492
rect 15932 9436 15988 9492
rect 27132 9436 27188 9492
rect 31724 9436 31780 9492
rect 31948 9436 32004 9492
rect 3804 9380 3860 9436
rect 3908 9380 3964 9436
rect 4012 9380 4068 9436
rect 23804 9380 23860 9436
rect 23908 9380 23964 9436
rect 24012 9380 24068 9436
rect 43804 9380 43860 9436
rect 43908 9380 43964 9436
rect 44012 9380 44068 9436
rect 8876 9324 8932 9380
rect 20860 9324 20916 9380
rect 24220 9324 24276 9380
rect 32396 9324 32452 9380
rect 15932 9212 15988 9268
rect 21308 9212 21364 9268
rect 27244 9212 27300 9268
rect 40572 9212 40628 9268
rect 27132 9100 27188 9156
rect 31164 9100 31220 9156
rect 30828 8988 30884 9044
rect 32732 8988 32788 9044
rect 40236 8988 40292 9044
rect 26908 8876 26964 8932
rect 30380 8876 30436 8932
rect 37884 8876 37940 8932
rect 4464 8596 4520 8652
rect 4568 8596 4624 8652
rect 4672 8596 4728 8652
rect 14700 8764 14756 8820
rect 32060 8764 32116 8820
rect 13132 8652 13188 8708
rect 18620 8652 18676 8708
rect 21532 8652 21588 8708
rect 21756 8652 21812 8708
rect 32732 8652 32788 8708
rect 24464 8596 24520 8652
rect 24568 8596 24624 8652
rect 24672 8596 24728 8652
rect 14140 8540 14196 8596
rect 27020 8540 27076 8596
rect 8316 8316 8372 8372
rect 13244 8316 13300 8372
rect 14140 8316 14196 8372
rect 17052 8316 17108 8372
rect 19516 8316 19572 8372
rect 40236 8652 40292 8708
rect 47628 8652 47684 8708
rect 44464 8596 44520 8652
rect 44568 8596 44624 8652
rect 44672 8596 44728 8652
rect 41916 8316 41972 8372
rect 2268 8204 2324 8260
rect 13692 8204 13748 8260
rect 13916 8204 13972 8260
rect 30380 8204 30436 8260
rect 30716 8204 30772 8260
rect 35644 8204 35700 8260
rect 38780 8204 38836 8260
rect 43372 8204 43428 8260
rect 15372 8092 15428 8148
rect 17500 8092 17556 8148
rect 39228 8092 39284 8148
rect 14812 7980 14868 8036
rect 26796 7980 26852 8036
rect 34972 7980 35028 8036
rect 38444 7980 38500 8036
rect 3804 7812 3860 7868
rect 3908 7812 3964 7868
rect 4012 7812 4068 7868
rect 31052 7868 31108 7924
rect 31500 7868 31556 7924
rect 23804 7812 23860 7868
rect 23908 7812 23964 7868
rect 24012 7812 24068 7868
rect 43804 7812 43860 7868
rect 43908 7812 43964 7868
rect 44012 7812 44068 7868
rect 19516 7756 19572 7812
rect 26684 7756 26740 7812
rect 30268 7756 30324 7812
rect 43148 7756 43204 7812
rect 26796 7644 26852 7700
rect 31276 7644 31332 7700
rect 26908 7532 26964 7588
rect 33404 7532 33460 7588
rect 43372 7532 43428 7588
rect 14924 7420 14980 7476
rect 15092 7420 15148 7476
rect 16716 7420 16772 7476
rect 18396 7420 18452 7476
rect 26684 7420 26740 7476
rect 35644 7420 35700 7476
rect 7308 7308 7364 7364
rect 30044 7308 30100 7364
rect 30380 7308 30436 7364
rect 12124 7196 12180 7252
rect 13692 7084 13748 7140
rect 16044 7084 16100 7140
rect 24220 7084 24276 7140
rect 43596 7084 43652 7140
rect 4464 7028 4520 7084
rect 4568 7028 4624 7084
rect 4672 7028 4728 7084
rect 24464 7028 24520 7084
rect 24568 7028 24624 7084
rect 24672 7028 24728 7084
rect 44464 7028 44520 7084
rect 44568 7028 44624 7084
rect 44672 7028 44728 7084
rect 33964 6860 34020 6916
rect 17948 6748 18004 6804
rect 25340 6748 25396 6804
rect 33516 6748 33572 6804
rect 16156 6636 16212 6692
rect 31388 6636 31444 6692
rect 33964 6636 34020 6692
rect 19740 6524 19796 6580
rect 23660 6524 23716 6580
rect 28476 6524 28532 6580
rect 16716 6412 16772 6468
rect 21756 6412 21812 6468
rect 25340 6412 25396 6468
rect 30044 6412 30100 6468
rect 43148 6412 43204 6468
rect 3804 6244 3860 6300
rect 3908 6244 3964 6300
rect 4012 6244 4068 6300
rect 23804 6244 23860 6300
rect 23908 6244 23964 6300
rect 24012 6244 24068 6300
rect 43804 6244 43860 6300
rect 43908 6244 43964 6300
rect 44012 6244 44068 6300
rect 18284 6188 18340 6244
rect 23660 6188 23716 6244
rect 40348 6188 40404 6244
rect 14812 6076 14868 6132
rect 15036 6076 15092 6132
rect 12012 5964 12068 6020
rect 27804 5964 27860 6020
rect 29148 5964 29204 6020
rect 31500 5964 31556 6020
rect 37324 5964 37380 6020
rect 37548 5964 37604 6020
rect 11900 5852 11956 5908
rect 18060 5852 18116 5908
rect 18284 5852 18340 5908
rect 20972 5852 21028 5908
rect 33292 5852 33348 5908
rect 16156 5740 16212 5796
rect 21532 5740 21588 5796
rect 25228 5740 25284 5796
rect 15372 5628 15428 5684
rect 16268 5628 16324 5684
rect 18396 5628 18452 5684
rect 18732 5628 18788 5684
rect 19964 5628 20020 5684
rect 20188 5628 20244 5684
rect 21644 5628 21700 5684
rect 31836 5628 31892 5684
rect 37548 5628 37604 5684
rect 38668 5628 38724 5684
rect 11452 5516 11508 5572
rect 11676 5516 11732 5572
rect 20972 5516 21028 5572
rect 22316 5516 22372 5572
rect 31164 5516 31220 5572
rect 4464 5460 4520 5516
rect 4568 5460 4624 5516
rect 4672 5460 4728 5516
rect 24464 5460 24520 5516
rect 24568 5460 24624 5516
rect 24672 5460 24728 5516
rect 37100 5516 37156 5572
rect 13580 5404 13636 5460
rect 18620 5404 18676 5460
rect 28364 5404 28420 5460
rect 44464 5460 44520 5516
rect 44568 5460 44624 5516
rect 44672 5460 44728 5516
rect 13356 5292 13412 5348
rect 16716 5292 16772 5348
rect 31724 5292 31780 5348
rect 33404 5292 33460 5348
rect 45388 5292 45444 5348
rect 11564 5180 11620 5236
rect 11788 5180 11844 5236
rect 14924 5180 14980 5236
rect 38668 5180 38724 5236
rect 13580 5068 13636 5124
rect 31948 5068 32004 5124
rect 32396 5068 32452 5124
rect 32956 5068 33012 5124
rect 33964 5068 34020 5124
rect 2268 4956 2324 5012
rect 33852 4956 33908 5012
rect 11788 4844 11844 4900
rect 13244 4844 13300 4900
rect 16716 4732 16772 4788
rect 3804 4676 3860 4732
rect 3908 4676 3964 4732
rect 4012 4676 4068 4732
rect 45164 4956 45220 5012
rect 45388 4956 45444 5012
rect 25116 4732 25172 4788
rect 33628 4732 33684 4788
rect 43596 4732 43652 4788
rect 23804 4676 23860 4732
rect 23908 4676 23964 4732
rect 24012 4676 24068 4732
rect 43804 4676 43860 4732
rect 43908 4676 43964 4732
rect 44012 4676 44068 4732
rect 21868 4620 21924 4676
rect 27580 4508 27636 4564
rect 36876 4508 36932 4564
rect 18956 4396 19012 4452
rect 20412 4396 20468 4452
rect 51100 4396 51156 4452
rect 12572 4172 12628 4228
rect 37324 4172 37380 4228
rect 28588 4060 28644 4116
rect 28812 4060 28868 4116
rect 30716 4060 30772 4116
rect 45388 4060 45444 4116
rect 4464 3892 4520 3948
rect 4568 3892 4624 3948
rect 4672 3892 4728 3948
rect 24464 3892 24520 3948
rect 24568 3892 24624 3948
rect 24672 3892 24728 3948
rect 44464 3892 44520 3948
rect 44568 3892 44624 3948
rect 44672 3892 44728 3948
rect 13468 3836 13524 3892
rect 23660 3836 23716 3892
rect 45164 3836 45220 3892
rect 8876 3724 8932 3780
rect 12124 3724 12180 3780
rect 37324 3724 37380 3780
rect 12348 3612 12404 3668
rect 12572 3612 12628 3668
rect 13244 3612 13300 3668
rect 14028 3612 14084 3668
rect 19628 3612 19684 3668
rect 25340 3612 25396 3668
rect 27580 3612 27636 3668
rect 6636 3500 6692 3556
rect 9548 3500 9604 3556
rect 13916 3500 13972 3556
rect 14140 3500 14196 3556
rect 18396 3500 18452 3556
rect 20300 3500 20356 3556
rect 23660 3500 23716 3556
rect 13356 3388 13412 3444
rect 16604 3388 16660 3444
rect 15484 3276 15540 3332
rect 16716 3276 16772 3332
rect 30268 3388 30324 3444
rect 30940 3388 30996 3444
rect 29372 3276 29428 3332
rect 30268 3276 30324 3332
rect 33628 3276 33684 3332
rect 17164 3164 17220 3220
rect 23660 3164 23716 3220
rect 28252 3164 28308 3220
rect 3804 3108 3860 3164
rect 3908 3108 3964 3164
rect 4012 3108 4068 3164
rect 23804 3108 23860 3164
rect 23908 3108 23964 3164
rect 24012 3108 24068 3164
rect 43804 3108 43860 3164
rect 43908 3108 43964 3164
rect 44012 3108 44068 3164
rect 4172 3052 4228 3108
rect 13692 3052 13748 3108
rect 23548 3052 23604 3108
rect 11676 2940 11732 2996
rect 12348 2940 12404 2996
rect 18284 2940 18340 2996
rect 20188 2940 20244 2996
rect 21420 2940 21476 2996
rect 26348 2940 26404 2996
rect 27132 2940 27188 2996
rect 28364 2940 28420 2996
rect 28588 2940 28644 2996
rect 34972 2940 35028 2996
rect 13132 2828 13188 2884
rect 28812 2828 28868 2884
rect 33068 2828 33124 2884
rect 34076 2828 34132 2884
rect 45276 2828 45332 2884
rect 8316 2716 8372 2772
rect 32620 2716 32676 2772
rect 6748 2604 6804 2660
rect 19628 2604 19684 2660
rect 26012 2604 26068 2660
rect 4172 2492 4228 2548
rect 25452 2492 25508 2548
rect 28700 2492 28756 2548
rect 13692 2380 13748 2436
rect 25340 2380 25396 2436
rect 32844 2380 32900 2436
rect 4464 2324 4520 2380
rect 4568 2324 4624 2380
rect 4672 2324 4728 2380
rect 24464 2324 24520 2380
rect 24568 2324 24624 2380
rect 24672 2324 24728 2380
rect 44464 2324 44520 2380
rect 44568 2324 44624 2380
rect 44672 2324 44728 2380
rect 21420 2268 21476 2324
rect 24892 2268 24948 2324
rect 32956 2268 33012 2324
rect 26348 2156 26404 2212
rect 26572 2156 26628 2212
rect 28364 2156 28420 2212
rect 24892 2044 24948 2100
rect 16940 1932 16996 1988
rect 13916 1820 13972 1876
rect 14812 1708 14868 1764
rect 16940 1708 16996 1764
rect 23660 1596 23716 1652
rect 3804 1540 3860 1596
rect 3908 1540 3964 1596
rect 4012 1540 4068 1596
rect 23804 1540 23860 1596
rect 23908 1540 23964 1596
rect 24012 1540 24068 1596
rect 27020 1596 27076 1652
rect 43804 1540 43860 1596
rect 43908 1540 43964 1596
rect 44012 1540 44068 1596
rect 9548 1484 9604 1540
rect 29372 1484 29428 1540
rect 38892 1484 38948 1540
rect 40236 1484 40292 1540
rect 47628 1484 47684 1540
rect 6748 1372 6804 1428
rect 16044 1372 16100 1428
rect 27132 1260 27188 1316
rect 38892 1260 38948 1316
rect 24220 1148 24276 1204
rect 26908 1148 26964 1204
rect 27804 1148 27860 1204
rect 32508 1148 32564 1204
rect 21308 1036 21364 1092
rect 25452 1036 25508 1092
rect 28812 1036 28868 1092
rect 33180 1036 33236 1092
rect 37100 1036 37156 1092
rect 23548 924 23604 980
rect 4464 756 4520 812
rect 4568 756 4624 812
rect 4672 756 4728 812
rect 15148 812 15204 868
rect 16940 812 16996 868
rect 21308 812 21364 868
rect 26684 812 26740 868
rect 26908 812 26964 868
rect 32508 812 32564 868
rect 24464 756 24520 812
rect 24568 756 24624 812
rect 24672 756 24728 812
rect 23548 700 23604 756
rect 25340 700 25396 756
rect 13356 588 13412 644
rect 34972 812 35028 868
rect 36988 812 37044 868
rect 44464 756 44520 812
rect 44568 756 44624 812
rect 44672 756 44728 812
rect 33068 700 33124 756
rect 40684 700 40740 756
rect 25900 588 25956 644
rect 28364 588 28420 644
rect 23212 476 23268 532
rect 27244 364 27300 420
rect 27916 364 27972 420
rect 32620 364 32676 420
rect 27020 252 27076 308
rect 34972 252 35028 308
rect 40684 252 40740 308
rect 15148 28 15204 84
rect 26012 28 26068 84
rect 27916 28 27972 84
rect 36988 28 37044 84
<< metal4 >>
rect 1596 13524 1652 13534
rect 1596 11956 1652 13468
rect 1596 11890 1652 11900
rect 3776 12572 4096 14224
rect 3776 12516 3804 12572
rect 3860 12516 3908 12572
rect 3964 12516 4012 12572
rect 4068 12516 4096 12572
rect 3776 11004 4096 12516
rect 4436 13356 4756 14224
rect 4436 13300 4464 13356
rect 4520 13300 4568 13356
rect 4624 13300 4672 13356
rect 4728 13300 4756 13356
rect 4436 11788 4756 13300
rect 4284 11732 4340 11742
rect 4284 11396 4340 11676
rect 4284 11330 4340 11340
rect 4436 11732 4464 11788
rect 4520 11732 4568 11788
rect 4624 11732 4672 11788
rect 4728 11732 4756 11788
rect 3776 10948 3804 11004
rect 3860 10948 3908 11004
rect 3964 10948 4012 11004
rect 4068 10948 4096 11004
rect 3776 9436 4096 10948
rect 3776 9380 3804 9436
rect 3860 9380 3908 9436
rect 3964 9380 4012 9436
rect 4068 9380 4096 9436
rect 2268 8260 2324 8270
rect 2268 5012 2324 8204
rect 2268 4946 2324 4956
rect 3776 7868 4096 9380
rect 3776 7812 3804 7868
rect 3860 7812 3908 7868
rect 3964 7812 4012 7868
rect 4068 7812 4096 7868
rect 3776 6300 4096 7812
rect 3776 6244 3804 6300
rect 3860 6244 3908 6300
rect 3964 6244 4012 6300
rect 4068 6244 4096 6300
rect 3776 4732 4096 6244
rect 3776 4676 3804 4732
rect 3860 4676 3908 4732
rect 3964 4676 4012 4732
rect 4068 4676 4096 4732
rect 3776 3164 4096 4676
rect 3776 3108 3804 3164
rect 3860 3108 3908 3164
rect 3964 3108 4012 3164
rect 4068 3108 4096 3164
rect 4436 10220 4756 11732
rect 10220 14196 10276 14206
rect 10108 11284 10164 11294
rect 4436 10164 4464 10220
rect 4520 10164 4568 10220
rect 4624 10164 4672 10220
rect 4728 10164 4756 10220
rect 4436 8652 4756 10164
rect 4436 8596 4464 8652
rect 4520 8596 4568 8652
rect 4624 8596 4672 8652
rect 4728 8596 4756 8652
rect 4436 7084 4756 8596
rect 4436 7028 4464 7084
rect 4520 7028 4568 7084
rect 4624 7028 4672 7084
rect 4728 7028 4756 7084
rect 4436 5516 4756 7028
rect 4436 5460 4464 5516
rect 4520 5460 4568 5516
rect 4624 5460 4672 5516
rect 4728 5460 4756 5516
rect 4436 3948 4756 5460
rect 4436 3892 4464 3948
rect 4520 3892 4568 3948
rect 4624 3892 4672 3948
rect 4728 3892 4756 3948
rect 3776 1596 4096 3108
rect 4172 3108 4228 3118
rect 4172 2548 4228 3052
rect 4172 2482 4228 2492
rect 3776 1540 3804 1596
rect 3860 1540 3908 1596
rect 3964 1540 4012 1596
rect 4068 1540 4096 1596
rect 3776 0 4096 1540
rect 4436 2380 4756 3892
rect 6636 11172 6692 11182
rect 6636 3556 6692 11116
rect 7308 10388 7364 10398
rect 7308 7364 7364 10332
rect 10108 9940 10164 11228
rect 10108 9874 10164 9884
rect 10220 9716 10276 14140
rect 20972 14196 21028 14206
rect 20972 13972 21028 14140
rect 20972 13906 21028 13916
rect 21196 14196 21252 14206
rect 18620 13300 18676 13310
rect 16940 12852 16996 12862
rect 15708 12302 16212 12358
rect 15708 12292 15764 12302
rect 15708 12226 15764 12236
rect 16156 12292 16212 12302
rect 16156 12226 16212 12236
rect 15148 11956 15204 11966
rect 15148 11818 15204 11900
rect 15484 11956 15540 11966
rect 15372 11844 15428 11854
rect 15148 11788 15372 11818
rect 15148 11762 15428 11788
rect 14588 11620 14644 11630
rect 10220 9650 10276 9660
rect 14476 10052 14532 10062
rect 14476 9492 14532 9996
rect 14588 9828 14644 11564
rect 15484 11620 15540 11900
rect 15484 11554 15540 11564
rect 14700 11508 14756 11518
rect 14756 11452 15092 11458
rect 14700 11402 15092 11452
rect 15036 11278 15092 11402
rect 15148 11396 15204 11406
rect 15148 11278 15204 11340
rect 15036 11222 15204 11278
rect 15260 9940 15316 9950
rect 14588 9762 14644 9772
rect 15148 9828 15204 9838
rect 14476 9426 14532 9436
rect 8876 9380 8932 9390
rect 7308 7298 7364 7308
rect 8316 8372 8372 8382
rect 6636 3490 6692 3500
rect 8316 2772 8372 8316
rect 8876 3780 8932 9324
rect 15148 9118 15204 9772
rect 14924 9062 15204 9118
rect 14700 8820 14756 8830
rect 13132 8708 13188 8718
rect 12124 7252 12180 7262
rect 11452 6020 12068 6058
rect 11452 6002 12012 6020
rect 11452 5572 11508 6002
rect 12012 5954 12068 5964
rect 11900 5908 11956 5918
rect 11452 5506 11508 5516
rect 11564 5852 11900 5878
rect 11564 5822 11956 5852
rect 11564 5236 11620 5822
rect 11564 5170 11620 5180
rect 11676 5572 11732 5582
rect 8876 3714 8932 3724
rect 8316 2706 8372 2716
rect 9548 3556 9604 3566
rect 4436 2324 4464 2380
rect 4520 2324 4568 2380
rect 4624 2324 4672 2380
rect 4728 2324 4756 2380
rect 4436 812 4756 2324
rect 6748 2660 6804 2670
rect 6748 1428 6804 2604
rect 9548 1540 9604 3500
rect 11676 2996 11732 5516
rect 11788 5236 11844 5246
rect 11788 4900 11844 5180
rect 11788 4834 11844 4844
rect 12124 3780 12180 7196
rect 12124 3714 12180 3724
rect 12572 4228 12628 4238
rect 11676 2930 11732 2940
rect 12348 3668 12404 3678
rect 12348 2996 12404 3612
rect 12572 3668 12628 4172
rect 12572 3602 12628 3612
rect 12348 2930 12404 2940
rect 13132 2884 13188 8652
rect 14140 8596 14196 8606
rect 13244 8372 13972 8398
rect 13300 8342 13972 8372
rect 13244 8306 13300 8316
rect 13692 8260 13748 8270
rect 13692 7140 13748 8204
rect 13916 8260 13972 8342
rect 14140 8372 14196 8540
rect 14140 8306 14196 8316
rect 13916 8194 13972 8204
rect 13692 7074 13748 7084
rect 14700 7138 14756 8764
rect 14812 8036 14868 8046
rect 14812 7318 14868 7980
rect 14924 7476 14980 9062
rect 15260 8938 15316 9884
rect 15148 8882 15316 8938
rect 15708 9604 15764 9614
rect 15148 7678 15204 8882
rect 15708 8218 15764 9548
rect 15932 9492 15988 9502
rect 15932 9268 15988 9436
rect 15932 9202 15988 9212
rect 15372 8162 15764 8218
rect 15372 8148 15428 8162
rect 15372 8082 15428 8092
rect 15148 7622 15540 7678
rect 14924 7410 14980 7420
rect 15036 7476 15148 7498
rect 15036 7420 15092 7476
rect 15036 7410 15148 7420
rect 15036 7318 15092 7410
rect 14812 7262 15092 7318
rect 14700 7082 15092 7138
rect 14812 6132 14868 6142
rect 13580 5460 13636 5470
rect 13356 5348 13412 5358
rect 13412 5292 13524 5338
rect 13356 5282 13524 5292
rect 13468 4978 13524 5282
rect 13580 5124 13636 5404
rect 13580 5058 13636 5068
rect 13468 4922 14196 4978
rect 13244 4900 13300 4910
rect 13244 4078 13300 4844
rect 13244 4022 13524 4078
rect 13468 3892 13524 4022
rect 13468 3826 13524 3836
rect 13244 3668 14084 3718
rect 13300 3662 14028 3668
rect 13244 3602 13300 3612
rect 14028 3602 14084 3612
rect 13916 3556 13972 3566
rect 13132 2818 13188 2828
rect 13356 3444 13412 3454
rect 9548 1474 9604 1484
rect 6748 1362 6804 1372
rect 4436 756 4464 812
rect 4520 756 4568 812
rect 4624 756 4672 812
rect 4728 756 4756 812
rect 4436 0 4756 756
rect 13356 644 13412 3388
rect 13692 3108 13748 3118
rect 13692 2436 13748 3052
rect 13692 2370 13748 2380
rect 13916 1876 13972 3500
rect 14140 3556 14196 4922
rect 14140 3490 14196 3500
rect 13916 1810 13972 1820
rect 14812 1764 14868 6076
rect 15036 6132 15092 7082
rect 15036 6066 15092 6076
rect 15372 5684 15428 5694
rect 15372 5518 15428 5628
rect 15148 5462 15428 5518
rect 15148 5338 15204 5462
rect 14924 5282 15204 5338
rect 14924 5236 14980 5282
rect 14924 5170 14980 5180
rect 15484 3332 15540 7622
rect 16716 7476 16772 7486
rect 15484 3266 15540 3276
rect 16044 7140 16100 7150
rect 14812 1698 14868 1708
rect 16044 1428 16100 7084
rect 16156 6692 16212 6702
rect 16156 5796 16212 6636
rect 16716 6468 16772 7420
rect 16716 6402 16772 6412
rect 16940 6058 16996 12796
rect 18620 12852 18676 13244
rect 18620 12786 18676 12796
rect 19852 13188 19908 13198
rect 17500 12180 17556 12190
rect 17052 11284 17108 11294
rect 17052 8372 17108 11228
rect 17052 8306 17108 8316
rect 17500 8148 17556 12124
rect 19068 11620 19124 11630
rect 19068 11060 19124 11564
rect 19068 10994 19124 11004
rect 18172 10052 18228 10062
rect 18172 9604 18228 9996
rect 18172 9538 18228 9548
rect 18620 8708 18676 8718
rect 18620 8578 18676 8652
rect 17500 8082 17556 8092
rect 18284 8522 18676 8578
rect 18284 7498 18340 8522
rect 19516 8372 19572 8382
rect 19516 7812 19572 8316
rect 19516 7746 19572 7756
rect 17948 7442 18340 7498
rect 18396 7476 18452 7486
rect 17948 6804 18004 7442
rect 17948 6738 18004 6748
rect 16156 5730 16212 5740
rect 16828 6002 16996 6058
rect 18284 6244 18340 6254
rect 16828 5698 16884 6002
rect 16268 5684 16884 5698
rect 16324 5642 16884 5684
rect 18060 5908 18116 5918
rect 16268 5618 16324 5628
rect 18060 5518 18116 5852
rect 18284 5908 18340 6188
rect 18284 5842 18340 5852
rect 18396 5684 18452 7420
rect 19740 6580 19796 6590
rect 18396 5618 18452 5628
rect 18732 5684 18788 5694
rect 18060 5462 18676 5518
rect 18620 5460 18676 5462
rect 18620 5394 18676 5404
rect 16716 5348 16772 5358
rect 18732 5338 18788 5628
rect 16716 4788 16772 5292
rect 16716 4722 16772 4732
rect 18284 5282 18788 5338
rect 16604 3444 16660 3454
rect 16604 2998 16660 3388
rect 16716 3332 16772 3342
rect 16716 3178 16772 3276
rect 17164 3220 17220 3230
rect 16716 3164 17164 3178
rect 16716 3122 17220 3164
rect 16604 2942 16996 2998
rect 16940 1988 16996 2942
rect 18284 2996 18340 5282
rect 19740 4978 19796 6524
rect 19852 5518 19908 13132
rect 21196 12404 21252 14140
rect 21196 12338 21252 12348
rect 23776 12572 24096 14224
rect 23776 12516 23804 12572
rect 23860 12516 23908 12572
rect 23964 12516 24012 12572
rect 24068 12516 24096 12572
rect 22092 11844 22148 11854
rect 21532 11732 21588 11742
rect 21532 11172 21588 11676
rect 22092 11638 22148 11788
rect 21644 11620 22148 11638
rect 21700 11582 22148 11620
rect 21644 11554 21700 11564
rect 21532 11106 21588 11116
rect 20412 11060 20468 11070
rect 20188 10276 20244 10286
rect 20188 10198 20244 10220
rect 19964 10142 20244 10198
rect 20300 10164 20356 10174
rect 19964 5684 20020 10142
rect 19964 5618 20020 5628
rect 20188 5684 20244 5694
rect 20188 5518 20244 5628
rect 19852 5462 20244 5518
rect 19740 4922 20244 4978
rect 18956 4452 19012 4462
rect 18396 4396 18956 4438
rect 18396 4382 19012 4396
rect 18396 3556 18452 4382
rect 18396 3490 18452 3500
rect 19628 3668 19684 3678
rect 18284 2930 18340 2940
rect 19628 2660 19684 3612
rect 20188 2996 20244 4922
rect 20300 3556 20356 10108
rect 20412 4452 20468 11004
rect 22092 11060 22148 11070
rect 22092 10724 22148 11004
rect 22092 10658 22148 10668
rect 23776 11004 24096 12516
rect 24220 13636 24276 13646
rect 24220 11732 24276 13580
rect 24220 11666 24276 11676
rect 24436 13356 24756 14224
rect 29484 14196 29540 14206
rect 32060 14196 32116 14206
rect 24436 13300 24464 13356
rect 24520 13300 24568 13356
rect 24624 13300 24672 13356
rect 24728 13300 24756 13356
rect 24436 11788 24756 13300
rect 24892 13860 24948 13870
rect 24892 12740 24948 13804
rect 25116 13748 25172 13758
rect 24892 12674 24948 12684
rect 25004 13412 25060 13422
rect 24436 11732 24464 11788
rect 24520 11732 24568 11788
rect 24624 11732 24672 11788
rect 24728 11732 24756 11788
rect 23776 10948 23804 11004
rect 23860 10948 23908 11004
rect 23964 10948 24012 11004
rect 24068 10948 24096 11004
rect 22316 10500 22372 10510
rect 22204 10388 22260 10398
rect 21980 10332 22204 10378
rect 21980 10322 22260 10332
rect 21980 10276 22036 10322
rect 21980 10210 22036 10220
rect 22316 10018 22372 10444
rect 21756 9962 22372 10018
rect 21756 9828 21812 9962
rect 21756 9762 21812 9772
rect 21980 9828 22036 9838
rect 21980 9658 22036 9772
rect 21532 9602 22036 9658
rect 20860 9380 20916 9390
rect 20860 9298 20916 9324
rect 20860 9268 21364 9298
rect 20860 9242 21308 9268
rect 21308 9202 21364 9212
rect 21532 8708 21588 9602
rect 23776 9436 24096 10948
rect 24436 10220 24756 11732
rect 23776 9380 23804 9436
rect 23860 9380 23908 9436
rect 23964 9380 24012 9436
rect 24068 9380 24096 9436
rect 21532 8642 21588 8652
rect 21756 8708 21812 8718
rect 21756 6468 21812 8652
rect 23776 7868 24096 9380
rect 24220 10164 24276 10174
rect 24220 9380 24276 10108
rect 24220 9314 24276 9324
rect 24436 10164 24464 10220
rect 24520 10164 24568 10220
rect 24624 10164 24672 10220
rect 24728 10164 24756 10220
rect 23776 7812 23804 7868
rect 23860 7812 23908 7868
rect 23964 7812 24012 7868
rect 24068 7812 24096 7868
rect 21756 6402 21812 6412
rect 23660 6580 23716 6590
rect 23660 6244 23716 6524
rect 23660 6178 23716 6188
rect 23776 6300 24096 7812
rect 24436 8652 24756 10164
rect 25004 9828 25060 13356
rect 25004 9762 25060 9772
rect 24436 8596 24464 8652
rect 24520 8596 24568 8652
rect 24624 8596 24672 8652
rect 24728 8596 24756 8652
rect 23776 6244 23804 6300
rect 23860 6244 23908 6300
rect 23964 6244 24012 6300
rect 24068 6244 24096 6300
rect 20972 5908 21028 5918
rect 20972 5572 21028 5852
rect 20972 5506 21028 5516
rect 21532 5796 21588 5806
rect 21532 5518 21588 5740
rect 21644 5684 22372 5698
rect 21700 5642 22372 5684
rect 21644 5618 21700 5628
rect 22316 5572 22372 5642
rect 21532 5462 21924 5518
rect 22316 5506 22372 5516
rect 21868 4676 21924 5462
rect 21868 4610 21924 4620
rect 23776 4732 24096 6244
rect 23776 4676 23804 4732
rect 23860 4676 23908 4732
rect 23964 4676 24012 4732
rect 24068 4676 24096 4732
rect 20412 4386 20468 4396
rect 20300 3490 20356 3500
rect 23660 3892 23716 3902
rect 23660 3556 23716 3836
rect 23660 3490 23716 3500
rect 23660 3220 23716 3230
rect 23548 3108 23604 3118
rect 20188 2930 20244 2940
rect 21420 2996 21476 3006
rect 19628 2594 19684 2604
rect 21420 2324 21476 2940
rect 21420 2258 21476 2268
rect 16940 1922 16996 1932
rect 16044 1362 16100 1372
rect 16940 1764 16996 1774
rect 13356 578 13412 588
rect 15148 868 15204 878
rect 15148 84 15204 812
rect 16940 868 16996 1708
rect 16940 802 16996 812
rect 21308 1092 21364 1102
rect 21308 868 21364 1036
rect 23548 980 23604 3052
rect 23660 1652 23716 3164
rect 23660 1586 23716 1596
rect 23776 3164 24096 4676
rect 23776 3108 23804 3164
rect 23860 3108 23908 3164
rect 23964 3108 24012 3164
rect 24068 3108 24096 3164
rect 23776 1596 24096 3108
rect 23548 914 23604 924
rect 23776 1540 23804 1596
rect 23860 1540 23908 1596
rect 23964 1540 24012 1596
rect 24068 1540 24096 1596
rect 21308 802 21364 812
rect 23548 756 23604 766
rect 23548 658 23604 700
rect 23212 602 23604 658
rect 23212 532 23268 602
rect 23212 466 23268 476
rect 15148 18 15204 28
rect 23776 0 24096 1540
rect 24220 7140 24276 7150
rect 24220 1204 24276 7084
rect 24220 1138 24276 1148
rect 24436 7084 24756 8596
rect 24436 7028 24464 7084
rect 24520 7028 24568 7084
rect 24624 7028 24672 7084
rect 24728 7028 24756 7084
rect 24436 5516 24756 7028
rect 24436 5460 24464 5516
rect 24520 5460 24568 5516
rect 24624 5460 24672 5516
rect 24728 5460 24756 5516
rect 24436 3948 24756 5460
rect 25116 4788 25172 13692
rect 29484 12852 29540 14140
rect 30156 14140 32060 14158
rect 30156 14102 32116 14140
rect 35420 14196 35476 14206
rect 30156 13748 30212 14102
rect 35420 13860 35476 14140
rect 35420 13794 35476 13804
rect 30156 13682 30212 13692
rect 36316 13748 36372 13758
rect 31164 13524 31220 13534
rect 31052 13076 31108 13086
rect 29484 12786 29540 12796
rect 30940 12852 30996 12862
rect 28028 12404 28084 12414
rect 28084 12348 28644 12358
rect 28028 12302 28644 12348
rect 28588 12292 28644 12302
rect 28588 12226 28644 12236
rect 30940 11844 30996 12796
rect 30940 11778 30996 11788
rect 26124 11620 26180 11630
rect 26124 11396 26180 11564
rect 26124 11330 26180 11340
rect 26460 11042 26740 11098
rect 26460 10612 26516 11042
rect 26460 10546 26516 10556
rect 26572 10948 26628 10958
rect 25228 9940 25284 9950
rect 25228 5796 25284 9884
rect 25340 6804 25396 6814
rect 25340 6468 25396 6748
rect 25340 6402 25396 6412
rect 25228 5730 25284 5740
rect 25116 4722 25172 4732
rect 24436 3892 24464 3948
rect 24520 3892 24568 3948
rect 24624 3892 24672 3948
rect 24728 3892 24756 3948
rect 24436 2380 24756 3892
rect 24436 2324 24464 2380
rect 24520 2324 24568 2380
rect 24624 2324 24672 2380
rect 24728 2324 24756 2380
rect 25340 3668 25396 3678
rect 25340 2436 25396 3612
rect 26348 2996 26404 3006
rect 26012 2660 26068 2670
rect 25340 2370 25396 2380
rect 25452 2548 25508 2558
rect 24436 812 24756 2324
rect 24892 2324 24948 2334
rect 24892 2100 24948 2268
rect 24892 2034 24948 2044
rect 25452 1092 25508 2492
rect 25452 1026 25508 1036
rect 24436 756 24464 812
rect 24520 756 24568 812
rect 24624 756 24672 812
rect 24728 756 24756 812
rect 24436 0 24756 756
rect 25340 756 25396 766
rect 25340 658 25396 700
rect 25340 644 25956 658
rect 25340 602 25900 644
rect 25900 578 25956 588
rect 26012 84 26068 2604
rect 26348 2212 26404 2940
rect 26348 2146 26404 2156
rect 26572 2212 26628 10892
rect 26684 10918 26740 11042
rect 28700 11060 28756 11070
rect 26908 10948 26964 10958
rect 26684 10892 26908 10918
rect 26684 10862 26964 10892
rect 27132 10724 27188 10734
rect 26852 10388 26908 10398
rect 26908 10332 27076 10378
rect 26852 10322 27076 10332
rect 26908 8932 26964 8942
rect 26796 8036 26852 8046
rect 26684 7812 26740 7822
rect 26684 7476 26740 7756
rect 26796 7700 26852 7980
rect 26796 7634 26852 7644
rect 26908 7588 26964 8876
rect 27020 8596 27076 10322
rect 27132 9492 27188 10668
rect 27132 9426 27188 9436
rect 27356 10500 27412 10510
rect 27244 9268 27300 9278
rect 27020 8530 27076 8540
rect 27132 9156 27188 9166
rect 26908 7522 26964 7532
rect 26684 7410 26740 7420
rect 27132 2996 27188 9100
rect 27132 2930 27188 2940
rect 26572 2146 26628 2156
rect 27020 1652 27076 1662
rect 27020 1558 27076 1596
rect 27020 1502 27188 1558
rect 27132 1316 27188 1502
rect 27132 1250 27188 1260
rect 26908 1204 26964 1214
rect 26684 868 26740 878
rect 26684 298 26740 812
rect 26908 868 26964 1148
rect 26908 802 26964 812
rect 27244 420 27300 9212
rect 27356 1018 27412 10444
rect 27916 10164 28644 10198
rect 27972 10142 28644 10164
rect 27916 10098 27972 10108
rect 28588 10052 28644 10142
rect 28588 9986 28644 9996
rect 28700 9716 28756 11004
rect 30828 11060 30884 11070
rect 30156 10948 30212 10958
rect 30156 10738 30212 10892
rect 30380 10948 30436 10958
rect 30156 10682 30324 10738
rect 28700 9650 28756 9660
rect 29820 9604 29876 9614
rect 28476 6580 28532 6590
rect 28476 6418 28532 6524
rect 27804 6362 28532 6418
rect 27804 6020 27860 6362
rect 27804 5954 27860 5964
rect 29148 6020 29204 6030
rect 29148 5878 29204 5964
rect 28364 5822 29204 5878
rect 28364 5460 28420 5822
rect 28364 5394 28420 5404
rect 27580 4564 27636 4574
rect 27580 3668 27636 4508
rect 27580 3602 27636 3612
rect 28252 4202 28868 4258
rect 28252 3220 28308 4202
rect 28252 3154 28308 3164
rect 28588 4116 28644 4126
rect 28364 2996 28420 3006
rect 28364 2818 28420 2940
rect 28588 2996 28644 4060
rect 28812 4116 28868 4202
rect 28812 4050 28868 4060
rect 29820 3898 29876 9548
rect 30268 7812 30324 10682
rect 30380 8932 30436 10892
rect 30828 10918 30884 11004
rect 31052 11060 31108 13020
rect 31164 12852 31220 13468
rect 32508 13076 32564 13086
rect 32508 12898 32564 13020
rect 31164 12786 31220 12796
rect 31836 12852 31892 12862
rect 32508 12842 32676 12898
rect 31836 11620 31892 12796
rect 31836 11554 31892 11564
rect 31052 10994 31108 11004
rect 30828 10862 31332 10918
rect 31276 10724 31332 10862
rect 31276 10658 31332 10668
rect 31276 10322 32116 10378
rect 30828 9604 30884 9614
rect 30828 9044 30884 9548
rect 30828 8978 30884 8988
rect 31052 9604 31108 9614
rect 30380 8866 30436 8876
rect 30268 7746 30324 7756
rect 30380 8260 30436 8270
rect 30044 7364 30100 7374
rect 30044 6468 30100 7308
rect 30380 7364 30436 8204
rect 30380 7298 30436 7308
rect 30716 8260 30772 8270
rect 30044 6402 30100 6412
rect 30716 4116 30772 8204
rect 31052 7924 31108 9548
rect 31052 7858 31108 7868
rect 31164 9156 31220 9166
rect 31164 5572 31220 9100
rect 31276 7700 31332 10322
rect 31836 10164 31892 10174
rect 31276 7634 31332 7644
rect 31388 10052 31444 10062
rect 31388 6692 31444 9996
rect 31724 9492 31780 9502
rect 31388 6626 31444 6636
rect 31500 7924 31556 7934
rect 31500 6020 31556 7868
rect 31500 5954 31556 5964
rect 31164 5506 31220 5516
rect 31724 5348 31780 9436
rect 31836 5684 31892 10108
rect 32060 10164 32116 10322
rect 32060 10098 32116 10108
rect 31836 5618 31892 5628
rect 31948 9492 32004 9502
rect 31724 5282 31780 5292
rect 31948 5124 32004 9436
rect 32396 9380 32452 9390
rect 31948 5058 32004 5068
rect 32060 8820 32116 8830
rect 30716 4050 30772 4060
rect 28588 2930 28644 2940
rect 28812 3842 29876 3898
rect 28812 2884 28868 3842
rect 32060 3538 32116 8764
rect 32396 5124 32452 9324
rect 32396 5058 32452 5068
rect 30940 3482 32116 3538
rect 30268 3444 30324 3454
rect 28812 2818 28868 2828
rect 29372 3332 29428 3342
rect 28364 2762 28756 2818
rect 28700 2548 28756 2762
rect 28700 2482 28756 2492
rect 28364 2212 28420 2222
rect 28364 2098 28420 2156
rect 28364 2042 28868 2098
rect 27804 1204 27860 1214
rect 27860 1148 28532 1198
rect 27804 1142 28532 1148
rect 27804 1138 27860 1142
rect 27356 962 28420 1018
rect 28364 644 28420 962
rect 28476 658 28532 1142
rect 28812 1092 28868 2042
rect 29372 1540 29428 3276
rect 30268 3332 30324 3388
rect 30940 3444 30996 3482
rect 30940 3378 30996 3388
rect 30268 3266 30324 3276
rect 32620 2772 32676 12842
rect 36316 12404 36372 13692
rect 39788 12852 39844 12862
rect 38892 12740 38948 12750
rect 38780 12684 38892 12718
rect 38780 12662 38948 12684
rect 38780 12516 38836 12662
rect 38780 12450 38836 12460
rect 39788 12516 39844 12796
rect 43776 12572 44096 14224
rect 39788 12450 39844 12460
rect 43484 12516 43540 12526
rect 39004 12404 39060 12414
rect 36316 12338 36372 12348
rect 38668 12348 39004 12358
rect 38668 12302 39060 12348
rect 38668 11998 38724 12302
rect 38444 11942 38724 11998
rect 33180 11620 33236 11630
rect 33180 11458 33236 11564
rect 33180 11402 33908 11458
rect 33852 11284 33908 11402
rect 33852 11218 33908 11228
rect 32732 10836 32788 10846
rect 32732 10500 32788 10780
rect 32732 10434 32788 10444
rect 34076 10724 34132 10734
rect 32732 9044 32788 9054
rect 32732 8708 32788 8988
rect 32732 8642 32788 8652
rect 33404 7588 33460 7598
rect 33404 6958 33460 7532
rect 33404 6916 34020 6958
rect 33404 6902 33964 6916
rect 33964 6850 34020 6860
rect 33516 6804 33572 6814
rect 33572 6748 34020 6778
rect 33516 6722 34020 6748
rect 33964 6692 34020 6722
rect 33964 6626 34020 6636
rect 33292 5908 33348 5918
rect 32620 2706 32676 2716
rect 32956 5124 33012 5134
rect 32844 2436 32900 2446
rect 32844 2278 32900 2380
rect 29372 1474 29428 1484
rect 32508 2222 32900 2278
rect 32956 2324 33012 5068
rect 33292 4978 33348 5852
rect 33404 5348 33460 5358
rect 33404 5158 33460 5292
rect 33404 5124 34020 5158
rect 33404 5102 33964 5124
rect 33964 5058 34020 5068
rect 33852 5012 33908 5022
rect 33292 4956 33852 4978
rect 33292 4922 33908 4956
rect 33628 4788 33684 4798
rect 33628 3332 33684 4732
rect 33628 3266 33684 3276
rect 32956 2258 33012 2268
rect 33068 2884 33124 2894
rect 32508 1204 32564 2222
rect 33068 1738 33124 2828
rect 34076 2884 34132 10668
rect 35644 10164 35700 10174
rect 35644 9604 35700 10108
rect 37324 10052 37380 10062
rect 35644 9538 35700 9548
rect 36876 9828 36932 9838
rect 35644 8260 35700 8270
rect 34972 8036 35028 8046
rect 34972 2996 35028 7980
rect 35644 7476 35700 8204
rect 35644 7410 35700 7420
rect 36876 4564 36932 9772
rect 37324 6020 37380 9996
rect 37884 9604 37940 9614
rect 37884 8932 37940 9548
rect 37884 8866 37940 8876
rect 38444 8036 38500 11942
rect 38892 11732 38948 11742
rect 38892 11172 38948 11676
rect 43484 11620 43540 12460
rect 43484 11554 43540 11564
rect 43776 12516 43804 12572
rect 43860 12516 43908 12572
rect 43964 12516 44012 12572
rect 44068 12516 44096 12572
rect 38892 11106 38948 11116
rect 41916 11060 41972 11070
rect 39564 10836 39620 10846
rect 39564 10388 39620 10780
rect 39564 10322 39620 10332
rect 40236 10500 40292 10510
rect 40236 9940 40292 10444
rect 40236 9874 40292 9884
rect 40572 9828 40628 9838
rect 40572 9268 40628 9772
rect 40572 9202 40628 9212
rect 40236 9044 40292 9054
rect 40236 8708 40292 8988
rect 40236 8642 40292 8652
rect 41916 8372 41972 11004
rect 41916 8306 41972 8316
rect 43776 11004 44096 12516
rect 44436 13356 44756 14224
rect 44436 13300 44464 13356
rect 44520 13300 44568 13356
rect 44624 13300 44672 13356
rect 44728 13300 44756 13356
rect 44436 11788 44756 13300
rect 44268 11732 44324 11742
rect 44268 11508 44324 11676
rect 44268 11442 44324 11452
rect 44436 11732 44464 11788
rect 44520 11732 44568 11788
rect 44624 11732 44672 11788
rect 44728 11732 44756 11788
rect 43776 10948 43804 11004
rect 43860 10948 43908 11004
rect 43964 10948 44012 11004
rect 44068 10948 44096 11004
rect 43776 9436 44096 10948
rect 43776 9380 43804 9436
rect 43860 9380 43908 9436
rect 43964 9380 44012 9436
rect 44068 9380 44096 9436
rect 38780 8260 38836 8270
rect 43372 8260 43428 8270
rect 38836 8204 39284 8218
rect 38780 8162 39284 8204
rect 39228 8148 39284 8162
rect 39228 8082 39284 8092
rect 38444 7970 38500 7980
rect 43148 7812 43204 7822
rect 43148 6468 43204 7756
rect 43372 7588 43428 8204
rect 43372 7522 43428 7532
rect 43776 7868 44096 9380
rect 43776 7812 43804 7868
rect 43860 7812 43908 7868
rect 43964 7812 44012 7868
rect 44068 7812 44096 7868
rect 43148 6402 43204 6412
rect 43596 7140 43652 7150
rect 40348 6244 40404 6254
rect 40236 6188 40348 6238
rect 40236 6182 40404 6188
rect 37324 5954 37380 5964
rect 37548 6020 37604 6030
rect 37548 5684 37604 5964
rect 37548 5618 37604 5628
rect 38668 5684 38724 5694
rect 36876 4498 36932 4508
rect 37100 5572 37156 5582
rect 34972 2930 35028 2940
rect 34076 2818 34132 2828
rect 32508 1138 32564 1148
rect 32620 1682 33124 1738
rect 28812 1026 28868 1036
rect 32620 1018 32676 1682
rect 32508 962 32676 1018
rect 33180 1092 33236 1102
rect 32508 868 32564 962
rect 32508 802 32564 812
rect 33068 756 33124 766
rect 33068 658 33124 700
rect 28476 602 33124 658
rect 28364 578 28420 588
rect 33180 478 33236 1036
rect 37100 1092 37156 5516
rect 38668 5236 38724 5628
rect 38668 5170 38724 5180
rect 37324 4228 37380 4238
rect 37324 3780 37380 4172
rect 37324 3714 37380 3724
rect 38892 1540 38948 1550
rect 38892 1316 38948 1484
rect 40236 1540 40292 6182
rect 40348 6178 40404 6182
rect 43596 4788 43652 7084
rect 43596 4722 43652 4732
rect 43776 6300 44096 7812
rect 43776 6244 43804 6300
rect 43860 6244 43908 6300
rect 43964 6244 44012 6300
rect 44068 6244 44096 6300
rect 43776 4732 44096 6244
rect 40236 1474 40292 1484
rect 43776 4676 43804 4732
rect 43860 4676 43908 4732
rect 43964 4676 44012 4732
rect 44068 4676 44096 4732
rect 43776 3164 44096 4676
rect 43776 3108 43804 3164
rect 43860 3108 43908 3164
rect 43964 3108 44012 3164
rect 44068 3108 44096 3164
rect 43776 1596 44096 3108
rect 43776 1540 43804 1596
rect 43860 1540 43908 1596
rect 43964 1540 44012 1596
rect 44068 1540 44096 1596
rect 38892 1250 38948 1260
rect 37100 1026 37156 1036
rect 27244 354 27300 364
rect 27916 420 27972 430
rect 27020 308 27076 318
rect 26684 252 27020 298
rect 26684 242 27076 252
rect 26012 18 26068 28
rect 27916 84 27972 364
rect 32620 422 33236 478
rect 34972 868 35028 878
rect 32620 420 32676 422
rect 32620 354 32676 364
rect 34972 308 35028 812
rect 34972 242 35028 252
rect 36988 868 37044 878
rect 27916 18 27972 28
rect 36988 84 37044 812
rect 40684 756 40740 766
rect 40684 308 40740 700
rect 40684 242 40740 252
rect 36988 18 37044 28
rect 43776 0 44096 1540
rect 44436 10220 44756 11732
rect 44436 10164 44464 10220
rect 44520 10164 44568 10220
rect 44624 10164 44672 10220
rect 44728 10164 44756 10220
rect 44436 8652 44756 10164
rect 51100 11732 51156 11742
rect 44436 8596 44464 8652
rect 44520 8596 44568 8652
rect 44624 8596 44672 8652
rect 44728 8596 44756 8652
rect 44436 7084 44756 8596
rect 44436 7028 44464 7084
rect 44520 7028 44568 7084
rect 44624 7028 44672 7084
rect 44728 7028 44756 7084
rect 44436 5516 44756 7028
rect 44436 5460 44464 5516
rect 44520 5460 44568 5516
rect 44624 5460 44672 5516
rect 44728 5460 44756 5516
rect 44436 3948 44756 5460
rect 47628 8708 47684 8718
rect 45388 5348 45444 5358
rect 44436 3892 44464 3948
rect 44520 3892 44568 3948
rect 44624 3892 44672 3948
rect 44728 3892 44756 3948
rect 44436 2380 44756 3892
rect 45164 5012 45220 5022
rect 45164 3892 45220 4956
rect 45388 5012 45444 5292
rect 45388 4946 45444 4956
rect 45388 4116 45444 4126
rect 45164 3826 45220 3836
rect 45276 4060 45388 4078
rect 45276 4022 45444 4060
rect 45276 2884 45332 4022
rect 45276 2818 45332 2828
rect 44436 2324 44464 2380
rect 44520 2324 44568 2380
rect 44624 2324 44672 2380
rect 44728 2324 44756 2380
rect 44436 812 44756 2324
rect 47628 1540 47684 8652
rect 51100 4452 51156 11676
rect 51100 4386 51156 4396
rect 47628 1474 47684 1484
rect 44436 756 44464 812
rect 44520 756 44568 812
rect 44624 756 44672 812
rect 44728 756 44756 812
rect 44436 0 44756 756
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _001_
timestamp 1486834041
transform 1 0 41328 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _002_
timestamp 1486834041
transform 1 0 42112 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _003_
timestamp 1486834041
transform 1 0 44464 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _004_
timestamp 1486834041
transform 1 0 41216 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _005_
timestamp 1486834041
transform 1 0 46928 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _006_
timestamp 1486834041
transform 1 0 37744 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _007_
timestamp 1486834041
transform 1 0 44576 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _008_
timestamp 1486834041
transform 1 0 42448 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _009_
timestamp 1486834041
transform -1 0 55216 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _010_
timestamp 1486834041
transform 1 0 38528 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _011_
timestamp 1486834041
transform 1 0 41552 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _012_
timestamp 1486834041
transform 1 0 47488 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _013_
timestamp 1486834041
transform 1 0 18480 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _014_
timestamp 1486834041
transform 1 0 27216 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _015_
timestamp 1486834041
transform 1 0 30240 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _016_
timestamp 1486834041
transform 1 0 24416 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _017_
timestamp 1486834041
transform 1 0 49840 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _018_
timestamp 1486834041
transform 1 0 28784 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _019_
timestamp 1486834041
transform 1 0 23296 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _020_
timestamp 1486834041
transform 1 0 5040 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _021_
timestamp 1486834041
transform 1 0 52192 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _022_
timestamp 1486834041
transform 1 0 24416 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _023_
timestamp 1486834041
transform 1 0 20496 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _024_
timestamp 1486834041
transform 1 0 30464 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _025_
timestamp 1486834041
transform 1 0 9856 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _026_
timestamp 1486834041
transform 1 0 23296 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _027_
timestamp 1486834041
transform 1 0 34272 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _028_
timestamp 1486834041
transform 1 0 39200 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _029_
timestamp 1486834041
transform 1 0 48272 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _030_
timestamp 1486834041
transform 1 0 21392 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _031_
timestamp 1486834041
transform 1 0 32144 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _032_
timestamp 1486834041
transform 1 0 49168 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _033_
timestamp 1486834041
transform 1 0 5600 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _034_
timestamp 1486834041
transform -1 0 4592 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _035_
timestamp 1486834041
transform 1 0 10304 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _036_
timestamp 1486834041
transform 1 0 15008 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _037_
timestamp 1486834041
transform 1 0 14896 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _038_
timestamp 1486834041
transform -1 0 11088 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _039_
timestamp 1486834041
transform -1 0 11088 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _040_
timestamp 1486834041
transform 1 0 1344 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _041_
timestamp 1486834041
transform -1 0 13552 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _042_
timestamp 1486834041
transform -1 0 20272 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _043_
timestamp 1486834041
transform -1 0 14336 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _044_
timestamp 1486834041
transform -1 0 31136 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _045_
timestamp 1486834041
transform -1 0 32480 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _046_
timestamp 1486834041
transform 1 0 46816 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _047_
timestamp 1486834041
transform -1 0 37744 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _048_
timestamp 1486834041
transform -1 0 9632 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _049_
timestamp 1486834041
transform 1 0 51296 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _050_
timestamp 1486834041
transform 1 0 49168 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _051_
timestamp 1486834041
transform -1 0 21392 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _052_
timestamp 1486834041
transform -1 0 18032 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _053_
timestamp 1486834041
transform 1 0 53088 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _054_
timestamp 1486834041
transform -1 0 25648 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _055_
timestamp 1486834041
transform 1 0 37408 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _056_
timestamp 1486834041
transform 1 0 49952 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _057_
timestamp 1486834041
transform 1 0 51520 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _058_
timestamp 1486834041
transform 1 0 48384 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _059_
timestamp 1486834041
transform 1 0 50288 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _060_
timestamp 1486834041
transform 1 0 30800 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _061_
timestamp 1486834041
transform 1 0 36400 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _062_
timestamp 1486834041
transform 1 0 37520 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _063_
timestamp 1486834041
transform 1 0 40096 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _064_
timestamp 1486834041
transform 1 0 36400 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _065_
timestamp 1486834041
transform -1 0 23184 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _066_
timestamp 1486834041
transform 1 0 34496 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _067_
timestamp 1486834041
transform -1 0 21504 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _068_
timestamp 1486834041
transform 1 0 35952 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _069_
timestamp 1486834041
transform -1 0 28672 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _070_
timestamp 1486834041
transform 1 0 52080 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _071_
timestamp 1486834041
transform 1 0 51520 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _072_
timestamp 1486834041
transform 1 0 41440 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _073_
timestamp 1486834041
transform -1 0 20720 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _074_
timestamp 1486834041
transform -1 0 21056 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _075_
timestamp 1486834041
transform -1 0 29232 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _076_
timestamp 1486834041
transform -1 0 33152 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _077_
timestamp 1486834041
transform 1 0 46256 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _078_
timestamp 1486834041
transform -1 0 35504 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _079_
timestamp 1486834041
transform 1 0 43792 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _080_
timestamp 1486834041
transform -1 0 19712 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _081_
timestamp 1486834041
transform 1 0 50736 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _082_
timestamp 1486834041
transform -1 0 14112 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _083_
timestamp 1486834041
transform -1 0 20272 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _084_
timestamp 1486834041
transform -1 0 10192 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _085_
timestamp 1486834041
transform -1 0 17584 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _086_
timestamp 1486834041
transform -1 0 15008 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _087_
timestamp 1486834041
transform -1 0 13328 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _088_
timestamp 1486834041
transform -1 0 22288 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _089_
timestamp 1486834041
transform -1 0 4704 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _090_
timestamp 1486834041
transform -1 0 6720 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _091_
timestamp 1486834041
transform -1 0 2688 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _092_
timestamp 1486834041
transform -1 0 3584 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _093_
timestamp 1486834041
transform -1 0 6496 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _094_
timestamp 1486834041
transform -1 0 7504 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _095_
timestamp 1486834041
transform 1 0 5264 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _096_
timestamp 1486834041
transform -1 0 3696 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _097_
timestamp 1486834041
transform -1 0 14448 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _098_
timestamp 1486834041
transform -1 0 9632 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _099_
timestamp 1486834041
transform -1 0 37072 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _100_
timestamp 1486834041
transform -1 0 29232 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _101_
timestamp 1486834041
transform -1 0 2800 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _102_
timestamp 1486834041
transform -1 0 4256 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _103_
timestamp 1486834041
transform -1 0 7168 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _104_
timestamp 1486834041
transform -1 0 26320 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _105_
timestamp 1486834041
transform 1 0 1008 0 -1 10192
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_1
timestamp 1486834041
transform 1 0 46816 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__001__I
timestamp 1486834041
transform 1 0 41104 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__002__I
timestamp 1486834041
transform -1 0 42112 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__003__I
timestamp 1486834041
transform 1 0 44240 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__004__I
timestamp 1486834041
transform -1 0 41216 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__005__I
timestamp 1486834041
transform -1 0 46928 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__006__I
timestamp 1486834041
transform -1 0 37744 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__007__I
timestamp 1486834041
transform -1 0 44576 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__008__I
timestamp 1486834041
transform 1 0 42224 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__009__I
timestamp 1486834041
transform 1 0 55216 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__010__I
timestamp 1486834041
transform 1 0 38304 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__011__I
timestamp 1486834041
transform 1 0 41328 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__012__I
timestamp 1486834041
transform -1 0 47488 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__013__I
timestamp 1486834041
transform -1 0 18480 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__014__I
timestamp 1486834041
transform -1 0 27216 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__015__I
timestamp 1486834041
transform 1 0 30016 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__016__I
timestamp 1486834041
transform 1 0 23968 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__017__I
timestamp 1486834041
transform -1 0 49840 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__018__I
timestamp 1486834041
transform -1 0 28784 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__019__I
timestamp 1486834041
transform 1 0 23072 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__020__I
timestamp 1486834041
transform 1 0 4816 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__021__I
timestamp 1486834041
transform -1 0 52080 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__022__I
timestamp 1486834041
transform -1 0 24192 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__023__I
timestamp 1486834041
transform -1 0 20384 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__024__I
timestamp 1486834041
transform 1 0 30240 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__025__I
timestamp 1486834041
transform 1 0 9632 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__026__I
timestamp 1486834041
transform -1 0 23296 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__027__I
timestamp 1486834041
transform -1 0 34272 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__028__I
timestamp 1486834041
transform 1 0 38976 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__029__I
timestamp 1486834041
transform -1 0 48272 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__030__I
timestamp 1486834041
transform 1 0 21168 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__031__I
timestamp 1486834041
transform 1 0 31920 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__032__I
timestamp 1486834041
transform 1 0 48944 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__033__I
timestamp 1486834041
transform 1 0 5376 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__034__I
timestamp 1486834041
transform -1 0 5040 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__035__I
timestamp 1486834041
transform 1 0 10080 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__036__I
timestamp 1486834041
transform 1 0 14784 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__037__I
timestamp 1486834041
transform 1 0 15792 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__038__I
timestamp 1486834041
transform 1 0 11088 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__039__I
timestamp 1486834041
transform -1 0 11312 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__040__I
timestamp 1486834041
transform -1 0 1344 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__041__I
timestamp 1486834041
transform -1 0 13776 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__042__I
timestamp 1486834041
transform -1 0 20720 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__043__I
timestamp 1486834041
transform 1 0 14336 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__044__I
timestamp 1486834041
transform 1 0 31136 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__045__I
timestamp 1486834041
transform -1 0 32704 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__046__I
timestamp 1486834041
transform 1 0 46592 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__047__I
timestamp 1486834041
transform -1 0 37968 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__048__I
timestamp 1486834041
transform 1 0 9632 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__049__I
timestamp 1486834041
transform 1 0 51072 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__050__I
timestamp 1486834041
transform -1 0 49168 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__051__I
timestamp 1486834041
transform 1 0 21392 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__052__I
timestamp 1486834041
transform 1 0 18032 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__053__I
timestamp 1486834041
transform -1 0 53200 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__054__I
timestamp 1486834041
transform 1 0 25648 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__055__I
timestamp 1486834041
transform -1 0 37408 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__056__I
timestamp 1486834041
transform -1 0 49952 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__057__I
timestamp 1486834041
transform -1 0 51520 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__058__I
timestamp 1486834041
transform -1 0 48384 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__059__I
timestamp 1486834041
transform 1 0 49952 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__060__I
timestamp 1486834041
transform -1 0 30800 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__061__I
timestamp 1486834041
transform 1 0 36176 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__062__I
timestamp 1486834041
transform 1 0 37296 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__063__I
timestamp 1486834041
transform -1 0 39872 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__064__I
timestamp 1486834041
transform -1 0 36400 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__065__I
timestamp 1486834041
transform 1 0 23184 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__066__I
timestamp 1486834041
transform -1 0 34496 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__067__I
timestamp 1486834041
transform -1 0 21728 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__068__I
timestamp 1486834041
transform -1 0 35952 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__069__I
timestamp 1486834041
transform -1 0 28896 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__070__I
timestamp 1486834041
transform 1 0 51408 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__071__I
timestamp 1486834041
transform -1 0 51520 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__072__I
timestamp 1486834041
transform -1 0 41440 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__073__I
timestamp 1486834041
transform -1 0 20944 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__074__I
timestamp 1486834041
transform -1 0 21280 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__075__I
timestamp 1486834041
transform 1 0 29232 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__076__I
timestamp 1486834041
transform -1 0 33376 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__077__I
timestamp 1486834041
transform 1 0 46032 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__078__I
timestamp 1486834041
transform -1 0 35728 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__079__I
timestamp 1486834041
transform -1 0 43792 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__080__I
timestamp 1486834041
transform 1 0 19712 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__081__I
timestamp 1486834041
transform 1 0 50512 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__082__I
timestamp 1486834041
transform 1 0 14112 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__083__I
timestamp 1486834041
transform 1 0 20496 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__084__I
timestamp 1486834041
transform -1 0 10192 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__085__I
timestamp 1486834041
transform -1 0 17808 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__086__I
timestamp 1486834041
transform -1 0 15232 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__087__I
timestamp 1486834041
transform -1 0 13552 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__088__I
timestamp 1486834041
transform -1 0 22512 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__089__I
timestamp 1486834041
transform -1 0 4928 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__090__I
timestamp 1486834041
transform 1 0 6720 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__091__I
timestamp 1486834041
transform -1 0 2912 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__092__I
timestamp 1486834041
transform -1 0 3808 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__093__I
timestamp 1486834041
transform -1 0 6720 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__094__I
timestamp 1486834041
transform -1 0 7728 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__095__I
timestamp 1486834041
transform -1 0 5264 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__096__I
timestamp 1486834041
transform 1 0 3696 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__097__I
timestamp 1486834041
transform -1 0 14672 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__098__I
timestamp 1486834041
transform -1 0 9856 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__099__I
timestamp 1486834041
transform 1 0 37072 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__100__I
timestamp 1486834041
transform 1 0 29232 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__101__I
timestamp 1486834041
transform -1 0 3024 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__102__I
timestamp 1486834041
transform -1 0 4480 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__103__I
timestamp 1486834041
transform -1 0 7392 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__104__I
timestamp 1486834041
transform -1 0 26544 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__105__I
timestamp 1486834041
transform -1 0 1456 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2
timestamp 1486834041
transform 1 0 896 0 1 784
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20
timestamp 1486834041
transform 1 0 2912 0 1 784
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28
timestamp 1486834041
transform 1 0 3808 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32
timestamp 1486834041
transform 1 0 4256 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36
timestamp 1486834041
transform 1 0 4704 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_70
timestamp 1486834041
transform 1 0 8512 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_104
timestamp 1486834041
transform 1 0 12320 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_138
timestamp 1486834041
transform 1 0 16128 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_172
timestamp 1486834041
transform 1 0 19936 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_206
timestamp 1486834041
transform 1 0 23744 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_240
timestamp 1486834041
transform 1 0 27552 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_274
timestamp 1486834041
transform 1 0 31360 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_308
timestamp 1486834041
transform 1 0 35168 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_342
timestamp 1486834041
transform 1 0 38976 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_376
timestamp 1486834041
transform 1 0 42784 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_410
timestamp 1486834041
transform 1 0 46592 0 1 784
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_444
timestamp 1486834041
transform 1 0 50400 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_478
timestamp 1486834041
transform 1 0 54208 0 1 784
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_482
timestamp 1486834041
transform 1 0 54656 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_484
timestamp 1486834041
transform 1 0 54880 0 1 784
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_2
timestamp 1486834041
transform 1 0 896 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_28
timestamp 1486834041
transform 1 0 3808 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_44
timestamp 1486834041
transform 1 0 5600 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_48
timestamp 1486834041
transform 1 0 6048 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_60
timestamp 1486834041
transform 1 0 7392 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_68
timestamp 1486834041
transform 1 0 8288 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_72
timestamp 1486834041
transform 1 0 8736 0 -1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_104
timestamp 1486834041
transform 1 0 12320 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_112
timestamp 1486834041
transform 1 0 13216 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_114
timestamp 1486834041
transform 1 0 13440 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_125
timestamp 1486834041
transform 1 0 14672 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_133
timestamp 1486834041
transform 1 0 15568 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_137
timestamp 1486834041
transform 1 0 16016 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_139
timestamp 1486834041
transform 1 0 16240 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_142
timestamp 1486834041
transform 1 0 16576 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_146
timestamp 1486834041
transform 1 0 17024 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_157
timestamp 1486834041
transform 1 0 18256 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_173
timestamp 1486834041
transform 1 0 20048 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_177
timestamp 1486834041
transform 1 0 20496 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_188
timestamp 1486834041
transform 1 0 21728 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_204
timestamp 1486834041
transform 1 0 23520 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_220
timestamp 1486834041
transform 1 0 25312 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_236
timestamp 1486834041
transform 1 0 27104 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_244
timestamp 1486834041
transform 1 0 28000 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_248
timestamp 1486834041
transform 1 0 28448 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_259
timestamp 1486834041
transform 1 0 29680 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_263
timestamp 1486834041
transform 1 0 30128 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_274
timestamp 1486834041
transform 1 0 31360 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_278
timestamp 1486834041
transform 1 0 31808 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_282
timestamp 1486834041
transform 1 0 32256 0 -1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_346
timestamp 1486834041
transform 1 0 39424 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_352
timestamp 1486834041
transform 1 0 40096 0 -1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_416
timestamp 1486834041
transform 1 0 47264 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_422
timestamp 1486834041
transform 1 0 47936 0 -1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_438
timestamp 1486834041
transform 1 0 49728 0 -1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_446
timestamp 1486834041
transform 1 0 50624 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_450
timestamp 1486834041
transform 1 0 51072 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_492
timestamp 1486834041
transform 1 0 55776 0 -1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_496
timestamp 1486834041
transform 1 0 56224 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_498
timestamp 1486834041
transform 1 0 56448 0 -1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_2
timestamp 1486834041
transform 1 0 896 0 1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_18
timestamp 1486834041
transform 1 0 2688 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_26
timestamp 1486834041
transform 1 0 3584 0 1 2352
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_39
timestamp 1486834041
transform 1 0 5040 0 1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_103
timestamp 1486834041
transform 1 0 12208 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_107
timestamp 1486834041
transform 1 0 12656 0 1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_171
timestamp 1486834041
transform 1 0 19824 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_177
timestamp 1486834041
transform 1 0 20496 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_181
timestamp 1486834041
transform 1 0 20944 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_193
timestamp 1486834041
transform 1 0 22288 0 1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_209
timestamp 1486834041
transform 1 0 24080 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_213
timestamp 1486834041
transform 1 0 24528 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_225
timestamp 1486834041
transform 1 0 25872 0 1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_241
timestamp 1486834041
transform 1 0 27664 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_257
timestamp 1486834041
transform 1 0 29456 0 1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_273
timestamp 1486834041
transform 1 0 31248 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_277
timestamp 1486834041
transform 1 0 31696 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_289
timestamp 1486834041
transform 1 0 33040 0 1 2352
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_305
timestamp 1486834041
transform 1 0 34832 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_313
timestamp 1486834041
transform 1 0 35728 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_317
timestamp 1486834041
transform 1 0 36176 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_325
timestamp 1486834041
transform 1 0 37072 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_339
timestamp 1486834041
transform 1 0 38640 0 1 2352
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_371
timestamp 1486834041
transform 1 0 42224 0 1 2352
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_379
timestamp 1486834041
transform 1 0 43120 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_383
timestamp 1486834041
transform 1 0 43568 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_387
timestamp 1486834041
transform 1 0 44016 0 1 2352
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_451
timestamp 1486834041
transform 1 0 51184 0 1 2352
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_2
timestamp 1486834041
transform 1 0 896 0 -1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_66
timestamp 1486834041
transform 1 0 8064 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_82
timestamp 1486834041
transform 1 0 9856 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_94
timestamp 1486834041
transform 1 0 11200 0 -1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_126
timestamp 1486834041
transform 1 0 14784 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_137
timestamp 1486834041
transform 1 0 16016 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_139
timestamp 1486834041
transform 1 0 16240 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_142
timestamp 1486834041
transform 1 0 16576 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_150
timestamp 1486834041
transform 1 0 17472 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_154
timestamp 1486834041
transform 1 0 17920 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_156
timestamp 1486834041
transform 1 0 18144 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_167
timestamp 1486834041
transform 1 0 19376 0 -1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_199
timestamp 1486834041
transform 1 0 22960 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_207
timestamp 1486834041
transform 1 0 23856 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_209
timestamp 1486834041
transform 1 0 24080 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_212
timestamp 1486834041
transform 1 0 24416 0 -1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_276
timestamp 1486834041
transform 1 0 31584 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_292
timestamp 1486834041
transform 1 0 33376 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_300
timestamp 1486834041
transform 1 0 34272 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_302
timestamp 1486834041
transform 1 0 34496 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_313
timestamp 1486834041
transform 1 0 35728 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_327
timestamp 1486834041
transform 1 0 37296 0 -1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_343
timestamp 1486834041
transform 1 0 39088 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_347
timestamp 1486834041
transform 1 0 39536 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_349
timestamp 1486834041
transform 1 0 39760 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_352
timestamp 1486834041
transform 1 0 40096 0 -1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_368
timestamp 1486834041
transform 1 0 41888 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_376
timestamp 1486834041
transform 1 0 42784 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_380
timestamp 1486834041
transform 1 0 43232 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_382
timestamp 1486834041
transform 1 0 43456 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_393
timestamp 1486834041
transform 1 0 44688 0 -1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_409
timestamp 1486834041
transform 1 0 46480 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_417
timestamp 1486834041
transform 1 0 47376 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_419
timestamp 1486834041
transform 1 0 47600 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_422
timestamp 1486834041
transform 1 0 47936 0 -1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_430
timestamp 1486834041
transform 1 0 48832 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_434
timestamp 1486834041
transform 1 0 49280 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_436
timestamp 1486834041
transform 1 0 49504 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_447
timestamp 1486834041
transform 1 0 50736 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_451
timestamp 1486834041
transform 1 0 51184 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_492
timestamp 1486834041
transform 1 0 55776 0 -1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_496
timestamp 1486834041
transform 1 0 56224 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_498
timestamp 1486834041
transform 1 0 56448 0 -1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_2
timestamp 1486834041
transform 1 0 896 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1486834041
transform 1 0 4480 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_47
timestamp 1486834041
transform 1 0 5936 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_79
timestamp 1486834041
transform 1 0 9520 0 1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_95
timestamp 1486834041
transform 1 0 11312 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_103
timestamp 1486834041
transform 1 0 12208 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_107
timestamp 1486834041
transform 1 0 12656 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_111
timestamp 1486834041
transform 1 0 13104 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_115
timestamp 1486834041
transform 1 0 13552 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_147
timestamp 1486834041
transform 1 0 17136 0 1 3920
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_163
timestamp 1486834041
transform 1 0 18928 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_171
timestamp 1486834041
transform 1 0 19824 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_177
timestamp 1486834041
transform 1 0 20496 0 1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_241
timestamp 1486834041
transform 1 0 27664 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_247
timestamp 1486834041
transform 1 0 28336 0 1 3920
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_311
timestamp 1486834041
transform 1 0 35504 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_327
timestamp 1486834041
transform 1 0 37296 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_335
timestamp 1486834041
transform 1 0 38192 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_339
timestamp 1486834041
transform 1 0 38640 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_341
timestamp 1486834041
transform 1 0 38864 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_352
timestamp 1486834041
transform 1 0 40096 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_360
timestamp 1486834041
transform 1 0 40992 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_362
timestamp 1486834041
transform 1 0 41216 0 1 3920
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_373
timestamp 1486834041
transform 1 0 42448 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_381
timestamp 1486834041
transform 1 0 43344 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_387
timestamp 1486834041
transform 1 0 44016 0 1 3920
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_419
timestamp 1486834041
transform 1 0 47600 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_427
timestamp 1486834041
transform 1 0 48496 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_441
timestamp 1486834041
transform 1 0 50064 0 1 3920
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_449
timestamp 1486834041
transform 1 0 50960 0 1 3920
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_469
timestamp 1486834041
transform 1 0 53200 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_2
timestamp 1486834041
transform 1 0 896 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_10
timestamp 1486834041
transform 1 0 1792 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_21
timestamp 1486834041
transform 1 0 3024 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_25
timestamp 1486834041
transform 1 0 3472 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_27
timestamp 1486834041
transform 1 0 3696 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_38
timestamp 1486834041
transform 1 0 4928 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_46
timestamp 1486834041
transform 1 0 5824 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_50
timestamp 1486834041
transform 1 0 6272 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_52
timestamp 1486834041
transform 1 0 6496 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_63
timestamp 1486834041
transform 1 0 7728 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_67
timestamp 1486834041
transform 1 0 8176 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_69
timestamp 1486834041
transform 1 0 8400 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_72
timestamp 1486834041
transform 1 0 8736 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_104
timestamp 1486834041
transform 1 0 12320 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_113
timestamp 1486834041
transform 1 0 13328 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_124
timestamp 1486834041
transform 1 0 14560 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_130
timestamp 1486834041
transform 1 0 15232 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_138
timestamp 1486834041
transform 1 0 16128 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_142
timestamp 1486834041
transform 1 0 16576 0 -1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_206
timestamp 1486834041
transform 1 0 23744 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_212
timestamp 1486834041
transform 1 0 24416 0 -1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_228
timestamp 1486834041
transform 1 0 26208 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_236
timestamp 1486834041
transform 1 0 27104 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_240
timestamp 1486834041
transform 1 0 27552 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_252
timestamp 1486834041
transform 1 0 28896 0 -1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_268
timestamp 1486834041
transform 1 0 30688 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_276
timestamp 1486834041
transform 1 0 31584 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_282
timestamp 1486834041
transform 1 0 32256 0 -1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_346
timestamp 1486834041
transform 1 0 39424 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_352
timestamp 1486834041
transform 1 0 40096 0 -1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_384
timestamp 1486834041
transform 1 0 43680 0 -1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_400
timestamp 1486834041
transform 1 0 45472 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_408
timestamp 1486834041
transform 1 0 46368 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_422
timestamp 1486834041
transform 1 0 47936 0 -1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_438
timestamp 1486834041
transform 1 0 49728 0 -1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_446
timestamp 1486834041
transform 1 0 50624 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_492
timestamp 1486834041
transform 1 0 55776 0 -1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_496
timestamp 1486834041
transform 1 0 56224 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_498
timestamp 1486834041
transform 1 0 56448 0 -1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1486834041
transform 1 0 896 0 1 5488
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1486834041
transform 1 0 4480 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_37
timestamp 1486834041
transform 1 0 4816 0 1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_101
timestamp 1486834041
transform 1 0 11984 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_107
timestamp 1486834041
transform 1 0 12656 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_111
timestamp 1486834041
transform 1 0 13104 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_136
timestamp 1486834041
transform 1 0 15904 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_152
timestamp 1486834041
transform 1 0 17696 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_160
timestamp 1486834041
transform 1 0 18592 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_164
timestamp 1486834041
transform 1 0 19040 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_166
timestamp 1486834041
transform 1 0 19264 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_179
timestamp 1486834041
transform 1 0 20720 0 1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_243
timestamp 1486834041
transform 1 0 27888 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_247
timestamp 1486834041
transform 1 0 28336 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_255
timestamp 1486834041
transform 1 0 29232 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_259
timestamp 1486834041
transform 1 0 29680 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_261
timestamp 1486834041
transform 1 0 29904 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_272
timestamp 1486834041
transform 1 0 31136 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_286
timestamp 1486834041
transform 1 0 32704 0 1 5488
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_302
timestamp 1486834041
transform 1 0 34496 0 1 5488
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_310
timestamp 1486834041
transform 1 0 35392 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_314
timestamp 1486834041
transform 1 0 35840 0 1 5488
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_317
timestamp 1486834041
transform 1 0 36176 0 1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_381
timestamp 1486834041
transform 1 0 43344 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_387
timestamp 1486834041
transform 1 0 44016 0 1 5488
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_451
timestamp 1486834041
transform 1 0 51184 0 1 5488
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_2
timestamp 1486834041
transform 1 0 896 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_18
timestamp 1486834041
transform 1 0 2688 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_22
timestamp 1486834041
transform 1 0 3136 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_34
timestamp 1486834041
transform 1 0 4480 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_66
timestamp 1486834041
transform 1 0 8064 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_72
timestamp 1486834041
transform 1 0 8736 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_104
timestamp 1486834041
transform 1 0 12320 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_122
timestamp 1486834041
transform 1 0 14336 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_138
timestamp 1486834041
transform 1 0 16128 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_142
timestamp 1486834041
transform 1 0 16576 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_174
timestamp 1486834041
transform 1 0 20160 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_176
timestamp 1486834041
transform 1 0 20384 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_187
timestamp 1486834041
transform 1 0 21616 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_195
timestamp 1486834041
transform 1 0 22512 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_199
timestamp 1486834041
transform 1 0 22960 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_212
timestamp 1486834041
transform 1 0 24416 0 -1 7056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_276
timestamp 1486834041
transform 1 0 31584 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_282
timestamp 1486834041
transform 1 0 32256 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_314
timestamp 1486834041
transform 1 0 35840 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_322
timestamp 1486834041
transform 1 0 36736 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_346
timestamp 1486834041
transform 1 0 39424 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_352
timestamp 1486834041
transform 1 0 40096 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_360
timestamp 1486834041
transform 1 0 40992 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_372
timestamp 1486834041
transform 1 0 42336 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_404
timestamp 1486834041
transform 1 0 45920 0 -1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_422
timestamp 1486834041
transform 1 0 47936 0 -1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_454
timestamp 1486834041
transform 1 0 51520 0 -1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_492
timestamp 1486834041
transform 1 0 55776 0 -1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_496
timestamp 1486834041
transform 1 0 56224 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_498
timestamp 1486834041
transform 1 0 56448 0 -1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1486834041
transform 1 0 896 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1486834041
transform 1 0 4480 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_37
timestamp 1486834041
transform 1 0 4816 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_69
timestamp 1486834041
transform 1 0 8400 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_77
timestamp 1486834041
transform 1 0 9296 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_79
timestamp 1486834041
transform 1 0 9520 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_90
timestamp 1486834041
transform 1 0 10752 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_98
timestamp 1486834041
transform 1 0 11648 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_102
timestamp 1486834041
transform 1 0 12096 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_104
timestamp 1486834041
transform 1 0 12320 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_107
timestamp 1486834041
transform 1 0 12656 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_139
timestamp 1486834041
transform 1 0 16240 0 1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_155
timestamp 1486834041
transform 1 0 18032 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_159
timestamp 1486834041
transform 1 0 18480 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_161
timestamp 1486834041
transform 1 0 18704 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_172
timestamp 1486834041
transform 1 0 19936 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_174
timestamp 1486834041
transform 1 0 20160 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_177
timestamp 1486834041
transform 1 0 20496 0 1 7056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_241
timestamp 1486834041
transform 1 0 27664 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_247
timestamp 1486834041
transform 1 0 28336 0 1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_263
timestamp 1486834041
transform 1 0 30128 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_274
timestamp 1486834041
transform 1 0 31360 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_306
timestamp 1486834041
transform 1 0 34944 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_314
timestamp 1486834041
transform 1 0 35840 0 1 7056
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_317
timestamp 1486834041
transform 1 0 36176 0 1 7056
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_381
timestamp 1486834041
transform 1 0 43344 0 1 7056
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_387
timestamp 1486834041
transform 1 0 44016 0 1 7056
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_419
timestamp 1486834041
transform 1 0 47600 0 1 7056
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_435
timestamp 1486834041
transform 1 0 49392 0 1 7056
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_443
timestamp 1486834041
transform 1 0 50288 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_16
timestamp 1486834041
transform 1 0 2464 0 -1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_32
timestamp 1486834041
transform 1 0 4256 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_40
timestamp 1486834041
transform 1 0 5152 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_52
timestamp 1486834041
transform 1 0 6496 0 -1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_68
timestamp 1486834041
transform 1 0 8288 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_82
timestamp 1486834041
transform 1 0 9856 0 -1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_114
timestamp 1486834041
transform 1 0 13440 0 -1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_130
timestamp 1486834041
transform 1 0 15232 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_138
timestamp 1486834041
transform 1 0 16128 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_142
timestamp 1486834041
transform 1 0 16576 0 -1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_158
timestamp 1486834041
transform 1 0 18368 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_166
timestamp 1486834041
transform 1 0 19264 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_170
timestamp 1486834041
transform 1 0 19712 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_181
timestamp 1486834041
transform 1 0 20944 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_195
timestamp 1486834041
transform 1 0 22512 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_203
timestamp 1486834041
transform 1 0 23408 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_207
timestamp 1486834041
transform 1 0 23856 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_209
timestamp 1486834041
transform 1 0 24080 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_212
timestamp 1486834041
transform 1 0 24416 0 -1 8624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_276
timestamp 1486834041
transform 1 0 31584 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_282
timestamp 1486834041
transform 1 0 32256 0 -1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_298
timestamp 1486834041
transform 1 0 34048 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_310
timestamp 1486834041
transform 1 0 35392 0 -1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_342
timestamp 1486834041
transform 1 0 38976 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_346
timestamp 1486834041
transform 1 0 39424 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_360
timestamp 1486834041
transform 1 0 40992 0 -1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_392
timestamp 1486834041
transform 1 0 44576 0 -1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_408
timestamp 1486834041
transform 1 0 46368 0 -1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_416
timestamp 1486834041
transform 1 0 47264 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_422
timestamp 1486834041
transform 1 0 47936 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_433
timestamp 1486834041
transform 1 0 49168 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_437
timestamp 1486834041
transform 1 0 49616 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_492
timestamp 1486834041
transform 1 0 55776 0 -1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_496
timestamp 1486834041
transform 1 0 56224 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_498
timestamp 1486834041
transform 1 0 56448 0 -1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_2
timestamp 1486834041
transform 1 0 896 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_4
timestamp 1486834041
transform 1 0 1120 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_29
timestamp 1486834041
transform 1 0 3920 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_33
timestamp 1486834041
transform 1 0 4368 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_37
timestamp 1486834041
transform 1 0 4816 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_45
timestamp 1486834041
transform 1 0 5712 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_56
timestamp 1486834041
transform 1 0 6944 0 1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_72
timestamp 1486834041
transform 1 0 8736 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_80
timestamp 1486834041
transform 1 0 9632 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_82
timestamp 1486834041
transform 1 0 9856 0 1 8624
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_95
timestamp 1486834041
transform 1 0 11312 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_103
timestamp 1486834041
transform 1 0 12208 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_107
timestamp 1486834041
transform 1 0 12656 0 1 8624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_171
timestamp 1486834041
transform 1 0 19824 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_177
timestamp 1486834041
transform 1 0 20496 0 1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_203
timestamp 1486834041
transform 1 0 23408 0 1 8624
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_235
timestamp 1486834041
transform 1 0 26992 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_243
timestamp 1486834041
transform 1 0 27888 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_247
timestamp 1486834041
transform 1 0 28336 0 1 8624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_311
timestamp 1486834041
transform 1 0 35504 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_317
timestamp 1486834041
transform 1 0 36176 0 1 8624
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_381
timestamp 1486834041
transform 1 0 43344 0 1 8624
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_387
timestamp 1486834041
transform 1 0 44016 0 1 8624
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_403
timestamp 1486834041
transform 1 0 45808 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_421
timestamp 1486834041
transform 1 0 47824 0 1 8624
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_429
timestamp 1486834041
transform 1 0 48720 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_2
timestamp 1486834041
transform 1 0 896 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_23
timestamp 1486834041
transform 1 0 3248 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_27
timestamp 1486834041
transform 1 0 3696 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_43
timestamp 1486834041
transform 1 0 5488 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_54
timestamp 1486834041
transform 1 0 6720 0 -1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_72
timestamp 1486834041
transform 1 0 8736 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_76
timestamp 1486834041
transform 1 0 9184 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_95
timestamp 1486834041
transform 1 0 11312 0 -1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_127
timestamp 1486834041
transform 1 0 14896 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_135
timestamp 1486834041
transform 1 0 15792 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_139
timestamp 1486834041
transform 1 0 16240 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_142
timestamp 1486834041
transform 1 0 16576 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_153
timestamp 1486834041
transform 1 0 17808 0 -1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_169
timestamp 1486834041
transform 1 0 19600 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_173
timestamp 1486834041
transform 1 0 20048 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_184
timestamp 1486834041
transform 1 0 21280 0 -1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_212
timestamp 1486834041
transform 1 0 24416 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_220
timestamp 1486834041
transform 1 0 25312 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_231
timestamp 1486834041
transform 1 0 26544 0 -1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_263
timestamp 1486834041
transform 1 0 30128 0 -1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_279
timestamp 1486834041
transform 1 0 31920 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_282
timestamp 1486834041
transform 1 0 32256 0 -1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_298
timestamp 1486834041
transform 1 0 34048 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_306
timestamp 1486834041
transform 1 0 34944 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_310
timestamp 1486834041
transform 1 0 35392 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_312
timestamp 1486834041
transform 1 0 35616 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_323
timestamp 1486834041
transform 1 0 36848 0 -1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_339
timestamp 1486834041
transform 1 0 38640 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_347
timestamp 1486834041
transform 1 0 39536 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_349
timestamp 1486834041
transform 1 0 39760 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_352
timestamp 1486834041
transform 1 0 40096 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_360
timestamp 1486834041
transform 1 0 40992 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_381
timestamp 1486834041
transform 1 0 43344 0 -1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_399
timestamp 1486834041
transform 1 0 45360 0 -1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_415
timestamp 1486834041
transform 1 0 47152 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_419
timestamp 1486834041
transform 1 0 47600 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_422
timestamp 1486834041
transform 1 0 47936 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_492
timestamp 1486834041
transform 1 0 55776 0 -1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_496
timestamp 1486834041
transform 1 0 56224 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_498
timestamp 1486834041
transform 1 0 56448 0 -1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_2
timestamp 1486834041
transform 1 0 896 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_4
timestamp 1486834041
transform 1 0 1120 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_37
timestamp 1486834041
transform 1 0 4816 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_41
timestamp 1486834041
transform 1 0 5264 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_99
timestamp 1486834041
transform 1 0 11760 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_103
timestamp 1486834041
transform 1 0 12208 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_135
timestamp 1486834041
transform 1 0 15792 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_151
timestamp 1486834041
transform 1 0 17584 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_179
timestamp 1486834041
transform 1 0 20720 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_195
timestamp 1486834041
transform 1 0 22512 0 1 10192
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_227
timestamp 1486834041
transform 1 0 26096 0 1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_243
timestamp 1486834041
transform 1 0 27888 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_247
timestamp 1486834041
transform 1 0 28336 0 1 10192
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_311
timestamp 1486834041
transform 1 0 35504 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_317
timestamp 1486834041
transform 1 0 36176 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_321
timestamp 1486834041
transform 1 0 36624 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_333
timestamp 1486834041
transform 1 0 37968 0 1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_349
timestamp 1486834041
transform 1 0 39760 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_357
timestamp 1486834041
transform 1 0 40656 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_359
timestamp 1486834041
transform 1 0 40880 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_378
timestamp 1486834041
transform 1 0 43008 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_382
timestamp 1486834041
transform 1 0 43456 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_384
timestamp 1486834041
transform 1 0 43680 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_387
timestamp 1486834041
transform 1 0 44016 0 1 10192
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_403
timestamp 1486834041
transform 1 0 45808 0 1 10192
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_411
timestamp 1486834041
transform 1 0 46704 0 1 10192
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_415
timestamp 1486834041
transform 1 0 47152 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_426
timestamp 1486834041
transform 1 0 48384 0 1 10192
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_2
timestamp 1486834041
transform 1 0 896 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_72
timestamp 1486834041
transform 1 0 8736 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_80
timestamp 1486834041
transform 1 0 9632 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_142
timestamp 1486834041
transform 1 0 16576 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_199
timestamp 1486834041
transform 1 0 22960 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_207
timestamp 1486834041
transform 1 0 23856 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_220
timestamp 1486834041
transform 1 0 25312 0 -1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_252
timestamp 1486834041
transform 1 0 28896 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_260
timestamp 1486834041
transform 1 0 29792 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_264
timestamp 1486834041
transform 1 0 30240 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_266
timestamp 1486834041
transform 1 0 30464 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_277
timestamp 1486834041
transform 1 0 31696 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_279
timestamp 1486834041
transform 1 0 31920 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_282
timestamp 1486834041
transform 1 0 32256 0 -1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_308
timestamp 1486834041
transform 1 0 35168 0 -1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_340
timestamp 1486834041
transform 1 0 38752 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_348
timestamp 1486834041
transform 1 0 39648 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_352
timestamp 1486834041
transform 1 0 40096 0 -1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_370
timestamp 1486834041
transform 1 0 42112 0 -1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_402
timestamp 1486834041
transform 1 0 45696 0 -1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_410
timestamp 1486834041
transform 1 0 46592 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_422
timestamp 1486834041
transform 1 0 47936 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_489
timestamp 1486834041
transform 1 0 55440 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_492
timestamp 1486834041
transform 1 0 55776 0 -1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_496
timestamp 1486834041
transform 1 0 56224 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_498
timestamp 1486834041
transform 1 0 56448 0 -1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_2
timestamp 1486834041
transform 1 0 896 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_6
timestamp 1486834041
transform 1 0 1344 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_37
timestamp 1486834041
transform 1 0 4816 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_117
timestamp 1486834041
transform 1 0 13776 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_185
timestamp 1486834041
transform 1 0 21392 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_215
timestamp 1486834041
transform 1 0 24752 0 1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_231
timestamp 1486834041
transform 1 0 26544 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_257
timestamp 1486834041
transform 1 0 29456 0 1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_289
timestamp 1486834041
transform 1 0 33040 0 1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_305
timestamp 1486834041
transform 1 0 34832 0 1 11760
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_313
timestamp 1486834041
transform 1 0 35728 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_337
timestamp 1486834041
transform 1 0 38416 0 1 11760
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_369
timestamp 1486834041
transform 1 0 42000 0 1 11760
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_387
timestamp 1486834041
transform 1 0 44016 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_389
timestamp 1486834041
transform 1 0 44240 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_400
timestamp 1486834041
transform 1 0 45472 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_404
timestamp 1486834041
transform 1 0 45920 0 1 11760
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_451
timestamp 1486834041
transform 1 0 51184 0 1 11760
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_2
timestamp 1486834041
transform 1 0 896 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_36
timestamp 1486834041
transform 1 0 4704 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_70
timestamp 1486834041
transform 1 0 8512 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_104
timestamp 1486834041
transform 1 0 12320 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_138
timestamp 1486834041
transform 1 0 16128 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_172
timestamp 1486834041
transform 1 0 19936 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_224
timestamp 1486834041
transform 1 0 25760 0 -1 13328
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_232
timestamp 1486834041
transform 1 0 26656 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_236
timestamp 1486834041
transform 1 0 27104 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_240
timestamp 1486834041
transform 1 0 27552 0 -1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_274
timestamp 1486834041
transform 1 0 31360 0 -1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_308
timestamp 1486834041
transform 1 0 35168 0 -1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_342
timestamp 1486834041
transform 1 0 38976 0 -1 13328
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_376
timestamp 1486834041
transform 1 0 42784 0 -1 13328
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_392
timestamp 1486834041
transform 1 0 44576 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_410
timestamp 1486834041
transform 1 0 46592 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_439
timestamp 1486834041
transform 1 0 49840 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_472
timestamp 1486834041
transform 1 0 53536 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_492
timestamp 1486834041
transform 1 0 55776 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_496
timestamp 1486834041
transform 1 0 56224 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_498
timestamp 1486834041
transform 1 0 56448 0 -1 13328
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output1
timestamp 1486834041
transform 1 0 51856 0 1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output2
timestamp 1486834041
transform 1 0 53424 0 1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output3
timestamp 1486834041
transform 1 0 53984 0 -1 5488
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output4
timestamp 1486834041
transform 1 0 54992 0 1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output5
timestamp 1486834041
transform 1 0 53424 0 1 5488
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output6
timestamp 1486834041
transform 1 0 53984 0 -1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output7
timestamp 1486834041
transform 1 0 54992 0 1 5488
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output8
timestamp 1486834041
transform 1 0 53424 0 1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output9
timestamp 1486834041
transform 1 0 54992 0 1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output10
timestamp 1486834041
transform 1 0 54992 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output11
timestamp 1486834041
transform 1 0 53424 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output12
timestamp 1486834041
transform 1 0 52416 0 -1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output13
timestamp 1486834041
transform 1 0 54992 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output14
timestamp 1486834041
transform 1 0 53984 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output15
timestamp 1486834041
transform 1 0 53424 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output16
timestamp 1486834041
transform 1 0 53984 0 -1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output17
timestamp 1486834041
transform 1 0 50848 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output18
timestamp 1486834041
transform 1 0 52416 0 -1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output19
timestamp 1486834041
transform 1 0 48048 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output20
timestamp 1486834041
transform 1 0 51856 0 1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output21
timestamp 1486834041
transform 1 0 50848 0 -1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output22
timestamp 1486834041
transform 1 0 48496 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output23
timestamp 1486834041
transform 1 0 50848 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output24
timestamp 1486834041
transform 1 0 49280 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output25
timestamp 1486834041
transform 1 0 50064 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output26
timestamp 1486834041
transform 1 0 52416 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output27
timestamp 1486834041
transform 1 0 52416 0 -1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output28
timestamp 1486834041
transform 1 0 53984 0 -1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output29
timestamp 1486834041
transform 1 0 54992 0 1 784
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output30
timestamp 1486834041
transform 1 0 53424 0 1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output31
timestamp 1486834041
transform 1 0 53984 0 -1 3920
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output32
timestamp 1486834041
transform 1 0 54992 0 1 2352
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output33
timestamp 1486834041
transform 1 0 48272 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output34
timestamp 1486834041
transform 1 0 52752 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output35
timestamp 1486834041
transform 1 0 54992 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output36
timestamp 1486834041
transform 1 0 52416 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output37
timestamp 1486834041
transform 1 0 51856 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output38
timestamp 1486834041
transform 1 0 50064 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output39
timestamp 1486834041
transform 1 0 46704 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output40
timestamp 1486834041
transform -1 0 48720 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output41
timestamp 1486834041
transform 1 0 52416 0 -1 7056
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output42
timestamp 1486834041
transform 1 0 44800 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output43
timestamp 1486834041
transform 1 0 51856 0 1 5488
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output44
timestamp 1486834041
transform 1 0 48720 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output45
timestamp 1486834041
transform 1 0 50400 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output46
timestamp 1486834041
transform 1 0 49616 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output47
timestamp 1486834041
transform 1 0 51968 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output48
timestamp 1486834041
transform 1 0 51856 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output49
timestamp 1486834041
transform 1 0 51184 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output50
timestamp 1486834041
transform 1 0 51856 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output51
timestamp 1486834041
transform 1 0 53424 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output52
timestamp 1486834041
transform 1 0 54208 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output53
timestamp 1486834041
transform -1 0 2464 0 -1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output54
timestamp 1486834041
transform -1 0 2800 0 1 8624
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output55
timestamp 1486834041
transform -1 0 3248 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output56
timestamp 1486834041
transform -1 0 3024 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output57
timestamp 1486834041
transform -1 0 3808 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output58
timestamp 1486834041
transform -1 0 4592 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output59
timestamp 1486834041
transform -1 0 3024 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output60
timestamp 1486834041
transform -1 0 5488 0 -1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output61
timestamp 1486834041
transform -1 0 2912 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output62
timestamp 1486834041
transform -1 0 4592 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output63
timestamp 1486834041
transform -1 0 5376 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output64
timestamp 1486834041
transform -1 0 4480 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output65
timestamp 1486834041
transform -1 0 7056 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output66
timestamp 1486834041
transform -1 0 6944 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output67
timestamp 1486834041
transform -1 0 8624 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output68
timestamp 1486834041
transform -1 0 6720 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output69
timestamp 1486834041
transform -1 0 7728 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output70
timestamp 1486834041
transform -1 0 8512 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output71
timestamp 1486834041
transform -1 0 10192 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output72
timestamp 1486834041
transform -1 0 8288 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output73
timestamp 1486834041
transform -1 0 9296 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output74
timestamp 1486834041
transform -1 0 15792 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output75
timestamp 1486834041
transform 1 0 12768 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output76
timestamp 1486834041
transform -1 0 15568 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output77
timestamp 1486834041
transform 1 0 14784 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output78
timestamp 1486834041
transform 1 0 16016 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output79
timestamp 1486834041
transform -1 0 15904 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output80
timestamp 1486834041
transform -1 0 11760 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output81
timestamp 1486834041
transform -1 0 10864 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output82
timestamp 1486834041
transform -1 0 11648 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output83
timestamp 1486834041
transform -1 0 10528 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output84
timestamp 1486834041
transform -1 0 12432 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output85
timestamp 1486834041
transform -1 0 13216 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output86
timestamp 1486834041
transform -1 0 14224 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output87
timestamp 1486834041
transform -1 0 12096 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output88
timestamp 1486834041
transform 1 0 13216 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output89
timestamp 1486834041
transform 1 0 15568 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output90
timestamp 1486834041
transform -1 0 22960 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output91
timestamp 1486834041
transform -1 0 21952 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output92
timestamp 1486834041
transform 1 0 21616 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output93
timestamp 1486834041
transform 1 0 21952 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output94
timestamp 1486834041
transform 1 0 23184 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output95
timestamp 1486834041
transform -1 0 25312 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output96
timestamp 1486834041
transform 1 0 16688 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output97
timestamp 1486834041
transform 1 0 17808 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output98
timestamp 1486834041
transform 1 0 17136 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output99
timestamp 1486834041
transform 1 0 16576 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output100
timestamp 1486834041
transform 1 0 18256 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output101
timestamp 1486834041
transform 1 0 18704 0 1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output102
timestamp 1486834041
transform 1 0 18144 0 -1 13328
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output103
timestamp 1486834041
transform 1 0 19824 0 -1 11760
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  output104
timestamp 1486834041
transform 1 0 20944 0 1 10192
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  output105
timestamp 1486834041
transform 1 0 47040 0 -1 11760
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_16
timestamp 1486834041
transform 1 0 672 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1486834041
transform -1 0 56784 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_17
timestamp 1486834041
transform 1 0 672 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1486834041
transform -1 0 56784 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_18
timestamp 1486834041
transform 1 0 672 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1486834041
transform -1 0 56784 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_19
timestamp 1486834041
transform 1 0 672 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1486834041
transform -1 0 56784 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_20
timestamp 1486834041
transform 1 0 672 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1486834041
transform -1 0 56784 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_21
timestamp 1486834041
transform 1 0 672 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1486834041
transform -1 0 56784 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_22
timestamp 1486834041
transform 1 0 672 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1486834041
transform -1 0 56784 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_23
timestamp 1486834041
transform 1 0 672 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1486834041
transform -1 0 56784 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_24
timestamp 1486834041
transform 1 0 672 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1486834041
transform -1 0 56784 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_25
timestamp 1486834041
transform 1 0 672 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1486834041
transform -1 0 56784 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_26
timestamp 1486834041
transform 1 0 672 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1486834041
transform -1 0 56784 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_27
timestamp 1486834041
transform 1 0 672 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1486834041
transform -1 0 56784 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_28
timestamp 1486834041
transform 1 0 672 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1486834041
transform -1 0 56784 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_29
timestamp 1486834041
transform 1 0 672 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1486834041
transform -1 0 56784 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_30
timestamp 1486834041
transform 1 0 672 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1486834041
transform -1 0 56784 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_31
timestamp 1486834041
transform 1 0 672 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1486834041
transform -1 0 56784 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  S_term_single_106
timestamp 1486834041
transform -1 0 25760 0 -1 13328
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_32
timestamp 1486834041
transform 1 0 4480 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_33
timestamp 1486834041
transform 1 0 8288 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_34
timestamp 1486834041
transform 1 0 12096 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_35
timestamp 1486834041
transform 1 0 15904 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_36
timestamp 1486834041
transform 1 0 19712 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_37
timestamp 1486834041
transform 1 0 23520 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_38
timestamp 1486834041
transform 1 0 27328 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_39
timestamp 1486834041
transform 1 0 31136 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_40
timestamp 1486834041
transform 1 0 34944 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_41
timestamp 1486834041
transform 1 0 38752 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_42
timestamp 1486834041
transform 1 0 42560 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_43
timestamp 1486834041
transform 1 0 46368 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_44
timestamp 1486834041
transform 1 0 50176 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_45
timestamp 1486834041
transform 1 0 53984 0 1 784
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_46
timestamp 1486834041
transform 1 0 8512 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_47
timestamp 1486834041
transform 1 0 16352 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_48
timestamp 1486834041
transform 1 0 24192 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_49
timestamp 1486834041
transform 1 0 32032 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_50
timestamp 1486834041
transform 1 0 39872 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_51
timestamp 1486834041
transform 1 0 47712 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_52
timestamp 1486834041
transform 1 0 55552 0 -1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_53
timestamp 1486834041
transform 1 0 4592 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_54
timestamp 1486834041
transform 1 0 12432 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_55
timestamp 1486834041
transform 1 0 20272 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_56
timestamp 1486834041
transform 1 0 28112 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_57
timestamp 1486834041
transform 1 0 35952 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_58
timestamp 1486834041
transform 1 0 43792 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_59
timestamp 1486834041
transform 1 0 51632 0 1 2352
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_60
timestamp 1486834041
transform 1 0 8512 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_61
timestamp 1486834041
transform 1 0 16352 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_62
timestamp 1486834041
transform 1 0 24192 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_63
timestamp 1486834041
transform 1 0 32032 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_64
timestamp 1486834041
transform 1 0 39872 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_65
timestamp 1486834041
transform 1 0 47712 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_66
timestamp 1486834041
transform 1 0 55552 0 -1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_67
timestamp 1486834041
transform 1 0 4592 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_68
timestamp 1486834041
transform 1 0 12432 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_69
timestamp 1486834041
transform 1 0 20272 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_70
timestamp 1486834041
transform 1 0 28112 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_71
timestamp 1486834041
transform 1 0 35952 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_72
timestamp 1486834041
transform 1 0 43792 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_73
timestamp 1486834041
transform 1 0 51632 0 1 3920
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_74
timestamp 1486834041
transform 1 0 8512 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_75
timestamp 1486834041
transform 1 0 16352 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_76
timestamp 1486834041
transform 1 0 24192 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_77
timestamp 1486834041
transform 1 0 32032 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_78
timestamp 1486834041
transform 1 0 39872 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_79
timestamp 1486834041
transform 1 0 47712 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_80
timestamp 1486834041
transform 1 0 55552 0 -1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_81
timestamp 1486834041
transform 1 0 4592 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_82
timestamp 1486834041
transform 1 0 12432 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_83
timestamp 1486834041
transform 1 0 20272 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_84
timestamp 1486834041
transform 1 0 28112 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_85
timestamp 1486834041
transform 1 0 35952 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_86
timestamp 1486834041
transform 1 0 43792 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_87
timestamp 1486834041
transform 1 0 51632 0 1 5488
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_88
timestamp 1486834041
transform 1 0 8512 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_89
timestamp 1486834041
transform 1 0 16352 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_90
timestamp 1486834041
transform 1 0 24192 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_91
timestamp 1486834041
transform 1 0 32032 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_92
timestamp 1486834041
transform 1 0 39872 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_93
timestamp 1486834041
transform 1 0 47712 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_94
timestamp 1486834041
transform 1 0 55552 0 -1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_95
timestamp 1486834041
transform 1 0 4592 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_96
timestamp 1486834041
transform 1 0 12432 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_97
timestamp 1486834041
transform 1 0 20272 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_98
timestamp 1486834041
transform 1 0 28112 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_99
timestamp 1486834041
transform 1 0 35952 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_100
timestamp 1486834041
transform 1 0 43792 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_101
timestamp 1486834041
transform 1 0 51632 0 1 7056
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_102
timestamp 1486834041
transform 1 0 8512 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_103
timestamp 1486834041
transform 1 0 16352 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_104
timestamp 1486834041
transform 1 0 24192 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_105
timestamp 1486834041
transform 1 0 32032 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_106
timestamp 1486834041
transform 1 0 39872 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_107
timestamp 1486834041
transform 1 0 47712 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_108
timestamp 1486834041
transform 1 0 55552 0 -1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_109
timestamp 1486834041
transform 1 0 4592 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_110
timestamp 1486834041
transform 1 0 12432 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_111
timestamp 1486834041
transform 1 0 20272 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_112
timestamp 1486834041
transform 1 0 28112 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_113
timestamp 1486834041
transform 1 0 35952 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_114
timestamp 1486834041
transform 1 0 43792 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_115
timestamp 1486834041
transform 1 0 51632 0 1 8624
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_116
timestamp 1486834041
transform 1 0 8512 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_117
timestamp 1486834041
transform 1 0 16352 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_118
timestamp 1486834041
transform 1 0 24192 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_119
timestamp 1486834041
transform 1 0 32032 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_120
timestamp 1486834041
transform 1 0 39872 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_121
timestamp 1486834041
transform 1 0 47712 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_122
timestamp 1486834041
transform 1 0 55552 0 -1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_123
timestamp 1486834041
transform 1 0 4592 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_124
timestamp 1486834041
transform 1 0 12432 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_125
timestamp 1486834041
transform 1 0 20272 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_126
timestamp 1486834041
transform 1 0 28112 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_127
timestamp 1486834041
transform 1 0 35952 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_128
timestamp 1486834041
transform 1 0 43792 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_129
timestamp 1486834041
transform 1 0 51632 0 1 10192
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_130
timestamp 1486834041
transform 1 0 8512 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_131
timestamp 1486834041
transform 1 0 16352 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_132
timestamp 1486834041
transform 1 0 24192 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_133
timestamp 1486834041
transform 1 0 32032 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_134
timestamp 1486834041
transform 1 0 39872 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_135
timestamp 1486834041
transform 1 0 47712 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_136
timestamp 1486834041
transform 1 0 55552 0 -1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_137
timestamp 1486834041
transform 1 0 4592 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_138
timestamp 1486834041
transform 1 0 12432 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_139
timestamp 1486834041
transform 1 0 20272 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_140
timestamp 1486834041
transform 1 0 28112 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_141
timestamp 1486834041
transform 1 0 35952 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_142
timestamp 1486834041
transform 1 0 43792 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_143
timestamp 1486834041
transform 1 0 51632 0 1 11760
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_144
timestamp 1486834041
transform 1 0 4480 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_145
timestamp 1486834041
transform 1 0 8288 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_146
timestamp 1486834041
transform 1 0 12096 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_147
timestamp 1486834041
transform 1 0 15904 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_148
timestamp 1486834041
transform 1 0 19712 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_149
timestamp 1486834041
transform 1 0 23520 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_150
timestamp 1486834041
transform 1 0 27328 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_151
timestamp 1486834041
transform 1 0 31136 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_152
timestamp 1486834041
transform 1 0 34944 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_153
timestamp 1486834041
transform 1 0 38752 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_154
timestamp 1486834041
transform 1 0 42560 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_155
timestamp 1486834041
transform 1 0 46368 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_156
timestamp 1486834041
transform 1 0 50176 0 -1 13328
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_157
timestamp 1486834041
transform 1 0 53984 0 -1 13328
box -86 -86 310 870
<< labels >>
flabel metal2 s 23968 14112 24080 14224 0 FreeSans 448 0 0 0 Co
port 0 nsew signal output
flabel metal3 s 0 0 112 112 0 FreeSans 448 0 0 0 FrameData[0]
port 1 nsew signal input
flabel metal3 s 0 4480 112 4592 0 FreeSans 448 0 0 0 FrameData[10]
port 2 nsew signal input
flabel metal3 s 0 4928 112 5040 0 FreeSans 448 0 0 0 FrameData[11]
port 3 nsew signal input
flabel metal3 s 0 5376 112 5488 0 FreeSans 448 0 0 0 FrameData[12]
port 4 nsew signal input
flabel metal3 s 0 5824 112 5936 0 FreeSans 448 0 0 0 FrameData[13]
port 5 nsew signal input
flabel metal3 s 0 6272 112 6384 0 FreeSans 448 0 0 0 FrameData[14]
port 6 nsew signal input
flabel metal3 s 0 6720 112 6832 0 FreeSans 448 0 0 0 FrameData[15]
port 7 nsew signal input
flabel metal3 s 0 7168 112 7280 0 FreeSans 448 0 0 0 FrameData[16]
port 8 nsew signal input
flabel metal3 s 0 7616 112 7728 0 FreeSans 448 0 0 0 FrameData[17]
port 9 nsew signal input
flabel metal3 s 0 8064 112 8176 0 FreeSans 448 0 0 0 FrameData[18]
port 10 nsew signal input
flabel metal3 s 0 8512 112 8624 0 FreeSans 448 0 0 0 FrameData[19]
port 11 nsew signal input
flabel metal3 s 0 448 112 560 0 FreeSans 448 0 0 0 FrameData[1]
port 12 nsew signal input
flabel metal3 s 0 8960 112 9072 0 FreeSans 448 0 0 0 FrameData[20]
port 13 nsew signal input
flabel metal3 s 0 9408 112 9520 0 FreeSans 448 0 0 0 FrameData[21]
port 14 nsew signal input
flabel metal3 s 0 9856 112 9968 0 FreeSans 448 0 0 0 FrameData[22]
port 15 nsew signal input
flabel metal3 s 0 10304 112 10416 0 FreeSans 448 0 0 0 FrameData[23]
port 16 nsew signal input
flabel metal3 s 0 10752 112 10864 0 FreeSans 448 0 0 0 FrameData[24]
port 17 nsew signal input
flabel metal3 s 0 11200 112 11312 0 FreeSans 448 0 0 0 FrameData[25]
port 18 nsew signal input
flabel metal3 s 0 11648 112 11760 0 FreeSans 448 0 0 0 FrameData[26]
port 19 nsew signal input
flabel metal3 s 0 12096 112 12208 0 FreeSans 448 0 0 0 FrameData[27]
port 20 nsew signal input
flabel metal3 s 0 12544 112 12656 0 FreeSans 448 0 0 0 FrameData[28]
port 21 nsew signal input
flabel metal3 s 0 12992 112 13104 0 FreeSans 448 0 0 0 FrameData[29]
port 22 nsew signal input
flabel metal3 s 0 896 112 1008 0 FreeSans 448 0 0 0 FrameData[2]
port 23 nsew signal input
flabel metal3 s 0 13440 112 13552 0 FreeSans 448 0 0 0 FrameData[30]
port 24 nsew signal input
flabel metal3 s 0 13888 112 14000 0 FreeSans 448 0 0 0 FrameData[31]
port 25 nsew signal input
flabel metal3 s 0 1344 112 1456 0 FreeSans 448 0 0 0 FrameData[3]
port 26 nsew signal input
flabel metal3 s 0 1792 112 1904 0 FreeSans 448 0 0 0 FrameData[4]
port 27 nsew signal input
flabel metal3 s 0 2240 112 2352 0 FreeSans 448 0 0 0 FrameData[5]
port 28 nsew signal input
flabel metal3 s 0 2688 112 2800 0 FreeSans 448 0 0 0 FrameData[6]
port 29 nsew signal input
flabel metal3 s 0 3136 112 3248 0 FreeSans 448 0 0 0 FrameData[7]
port 30 nsew signal input
flabel metal3 s 0 3584 112 3696 0 FreeSans 448 0 0 0 FrameData[8]
port 31 nsew signal input
flabel metal3 s 0 4032 112 4144 0 FreeSans 448 0 0 0 FrameData[9]
port 32 nsew signal input
flabel metal3 s 57344 0 57456 112 0 FreeSans 448 0 0 0 FrameData_O[0]
port 33 nsew signal output
flabel metal3 s 57344 4480 57456 4592 0 FreeSans 448 0 0 0 FrameData_O[10]
port 34 nsew signal output
flabel metal3 s 57344 4928 57456 5040 0 FreeSans 448 0 0 0 FrameData_O[11]
port 35 nsew signal output
flabel metal3 s 57344 5376 57456 5488 0 FreeSans 448 0 0 0 FrameData_O[12]
port 36 nsew signal output
flabel metal3 s 57344 5824 57456 5936 0 FreeSans 448 0 0 0 FrameData_O[13]
port 37 nsew signal output
flabel metal3 s 57344 6272 57456 6384 0 FreeSans 448 0 0 0 FrameData_O[14]
port 38 nsew signal output
flabel metal3 s 57344 6720 57456 6832 0 FreeSans 448 0 0 0 FrameData_O[15]
port 39 nsew signal output
flabel metal3 s 57344 7168 57456 7280 0 FreeSans 448 0 0 0 FrameData_O[16]
port 40 nsew signal output
flabel metal3 s 57344 7616 57456 7728 0 FreeSans 448 0 0 0 FrameData_O[17]
port 41 nsew signal output
flabel metal3 s 57344 8064 57456 8176 0 FreeSans 448 0 0 0 FrameData_O[18]
port 42 nsew signal output
flabel metal3 s 57344 8512 57456 8624 0 FreeSans 448 0 0 0 FrameData_O[19]
port 43 nsew signal output
flabel metal3 s 57344 448 57456 560 0 FreeSans 448 0 0 0 FrameData_O[1]
port 44 nsew signal output
flabel metal3 s 57344 8960 57456 9072 0 FreeSans 448 0 0 0 FrameData_O[20]
port 45 nsew signal output
flabel metal3 s 57344 9408 57456 9520 0 FreeSans 448 0 0 0 FrameData_O[21]
port 46 nsew signal output
flabel metal3 s 57344 9856 57456 9968 0 FreeSans 448 0 0 0 FrameData_O[22]
port 47 nsew signal output
flabel metal3 s 57344 10304 57456 10416 0 FreeSans 448 0 0 0 FrameData_O[23]
port 48 nsew signal output
flabel metal3 s 57344 10752 57456 10864 0 FreeSans 448 0 0 0 FrameData_O[24]
port 49 nsew signal output
flabel metal3 s 57344 11200 57456 11312 0 FreeSans 448 0 0 0 FrameData_O[25]
port 50 nsew signal output
flabel metal3 s 57344 11648 57456 11760 0 FreeSans 448 0 0 0 FrameData_O[26]
port 51 nsew signal output
flabel metal3 s 57344 12096 57456 12208 0 FreeSans 448 0 0 0 FrameData_O[27]
port 52 nsew signal output
flabel metal3 s 57344 12544 57456 12656 0 FreeSans 448 0 0 0 FrameData_O[28]
port 53 nsew signal output
flabel metal3 s 57344 12992 57456 13104 0 FreeSans 448 0 0 0 FrameData_O[29]
port 54 nsew signal output
flabel metal3 s 57344 896 57456 1008 0 FreeSans 448 0 0 0 FrameData_O[2]
port 55 nsew signal output
flabel metal3 s 57344 13440 57456 13552 0 FreeSans 448 0 0 0 FrameData_O[30]
port 56 nsew signal output
flabel metal3 s 57344 13888 57456 14000 0 FreeSans 448 0 0 0 FrameData_O[31]
port 57 nsew signal output
flabel metal3 s 57344 1344 57456 1456 0 FreeSans 448 0 0 0 FrameData_O[3]
port 58 nsew signal output
flabel metal3 s 57344 1792 57456 1904 0 FreeSans 448 0 0 0 FrameData_O[4]
port 59 nsew signal output
flabel metal3 s 57344 2240 57456 2352 0 FreeSans 448 0 0 0 FrameData_O[5]
port 60 nsew signal output
flabel metal3 s 57344 2688 57456 2800 0 FreeSans 448 0 0 0 FrameData_O[6]
port 61 nsew signal output
flabel metal3 s 57344 3136 57456 3248 0 FreeSans 448 0 0 0 FrameData_O[7]
port 62 nsew signal output
flabel metal3 s 57344 3584 57456 3696 0 FreeSans 448 0 0 0 FrameData_O[8]
port 63 nsew signal output
flabel metal3 s 57344 4032 57456 4144 0 FreeSans 448 0 0 0 FrameData_O[9]
port 64 nsew signal output
flabel metal2 s 4480 0 4592 112 0 FreeSans 448 0 0 0 FrameStrobe[0]
port 65 nsew signal input
flabel metal2 s 31360 0 31472 112 0 FreeSans 448 0 0 0 FrameStrobe[10]
port 66 nsew signal input
flabel metal2 s 34048 0 34160 112 0 FreeSans 448 0 0 0 FrameStrobe[11]
port 67 nsew signal input
flabel metal2 s 36736 0 36848 112 0 FreeSans 448 0 0 0 FrameStrobe[12]
port 68 nsew signal input
flabel metal2 s 39424 0 39536 112 0 FreeSans 448 0 0 0 FrameStrobe[13]
port 69 nsew signal input
flabel metal2 s 42112 0 42224 112 0 FreeSans 448 0 0 0 FrameStrobe[14]
port 70 nsew signal input
flabel metal2 s 44800 0 44912 112 0 FreeSans 448 0 0 0 FrameStrobe[15]
port 71 nsew signal input
flabel metal2 s 47488 0 47600 112 0 FreeSans 448 0 0 0 FrameStrobe[16]
port 72 nsew signal input
flabel metal2 s 50176 0 50288 112 0 FreeSans 448 0 0 0 FrameStrobe[17]
port 73 nsew signal input
flabel metal2 s 52864 0 52976 112 0 FreeSans 448 0 0 0 FrameStrobe[18]
port 74 nsew signal input
flabel metal2 s 55552 0 55664 112 0 FreeSans 448 0 0 0 FrameStrobe[19]
port 75 nsew signal input
flabel metal2 s 7168 0 7280 112 0 FreeSans 448 0 0 0 FrameStrobe[1]
port 76 nsew signal input
flabel metal2 s 9856 0 9968 112 0 FreeSans 448 0 0 0 FrameStrobe[2]
port 77 nsew signal input
flabel metal2 s 12544 0 12656 112 0 FreeSans 448 0 0 0 FrameStrobe[3]
port 78 nsew signal input
flabel metal2 s 15232 0 15344 112 0 FreeSans 448 0 0 0 FrameStrobe[4]
port 79 nsew signal input
flabel metal2 s 17920 0 18032 112 0 FreeSans 448 0 0 0 FrameStrobe[5]
port 80 nsew signal input
flabel metal2 s 20608 0 20720 112 0 FreeSans 448 0 0 0 FrameStrobe[6]
port 81 nsew signal input
flabel metal2 s 23296 0 23408 112 0 FreeSans 448 0 0 0 FrameStrobe[7]
port 82 nsew signal input
flabel metal2 s 25984 0 26096 112 0 FreeSans 448 0 0 0 FrameStrobe[8]
port 83 nsew signal input
flabel metal2 s 28672 0 28784 112 0 FreeSans 448 0 0 0 FrameStrobe[9]
port 84 nsew signal input
flabel metal2 s 48160 14112 48272 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[0]
port 85 nsew signal output
flabel metal2 s 52640 14112 52752 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[10]
port 86 nsew signal output
flabel metal2 s 53088 14112 53200 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[11]
port 87 nsew signal output
flabel metal2 s 53536 14112 53648 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[12]
port 88 nsew signal output
flabel metal2 s 53984 14112 54096 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[13]
port 89 nsew signal output
flabel metal2 s 54432 14112 54544 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[14]
port 90 nsew signal output
flabel metal2 s 54880 14112 54992 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[15]
port 91 nsew signal output
flabel metal2 s 55328 14112 55440 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[16]
port 92 nsew signal output
flabel metal2 s 55776 14112 55888 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[17]
port 93 nsew signal output
flabel metal2 s 56224 14112 56336 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[18]
port 94 nsew signal output
flabel metal2 s 56672 14112 56784 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[19]
port 95 nsew signal output
flabel metal2 s 48608 14112 48720 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[1]
port 96 nsew signal output
flabel metal2 s 49056 14112 49168 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[2]
port 97 nsew signal output
flabel metal2 s 49504 14112 49616 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[3]
port 98 nsew signal output
flabel metal2 s 49952 14112 50064 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[4]
port 99 nsew signal output
flabel metal2 s 50400 14112 50512 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[5]
port 100 nsew signal output
flabel metal2 s 50848 14112 50960 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[6]
port 101 nsew signal output
flabel metal2 s 51296 14112 51408 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[7]
port 102 nsew signal output
flabel metal2 s 51744 14112 51856 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[8]
port 103 nsew signal output
flabel metal2 s 52192 14112 52304 14224 0 FreeSans 448 0 0 0 FrameStrobe_O[9]
port 104 nsew signal output
flabel metal2 s 672 14112 784 14224 0 FreeSans 448 0 0 0 N1BEG[0]
port 105 nsew signal output
flabel metal2 s 1120 14112 1232 14224 0 FreeSans 448 0 0 0 N1BEG[1]
port 106 nsew signal output
flabel metal2 s 1568 14112 1680 14224 0 FreeSans 448 0 0 0 N1BEG[2]
port 107 nsew signal output
flabel metal2 s 2016 14112 2128 14224 0 FreeSans 448 0 0 0 N1BEG[3]
port 108 nsew signal output
flabel metal2 s 2464 14112 2576 14224 0 FreeSans 448 0 0 0 N2BEG[0]
port 109 nsew signal output
flabel metal2 s 2912 14112 3024 14224 0 FreeSans 448 0 0 0 N2BEG[1]
port 110 nsew signal output
flabel metal2 s 3360 14112 3472 14224 0 FreeSans 448 0 0 0 N2BEG[2]
port 111 nsew signal output
flabel metal2 s 3808 14112 3920 14224 0 FreeSans 448 0 0 0 N2BEG[3]
port 112 nsew signal output
flabel metal2 s 4256 14112 4368 14224 0 FreeSans 448 0 0 0 N2BEG[4]
port 113 nsew signal output
flabel metal2 s 4704 14112 4816 14224 0 FreeSans 448 0 0 0 N2BEG[5]
port 114 nsew signal output
flabel metal2 s 5152 14112 5264 14224 0 FreeSans 448 0 0 0 N2BEG[6]
port 115 nsew signal output
flabel metal2 s 5600 14112 5712 14224 0 FreeSans 448 0 0 0 N2BEG[7]
port 116 nsew signal output
flabel metal2 s 6048 14112 6160 14224 0 FreeSans 448 0 0 0 N2BEGb[0]
port 117 nsew signal output
flabel metal2 s 6496 14112 6608 14224 0 FreeSans 448 0 0 0 N2BEGb[1]
port 118 nsew signal output
flabel metal2 s 6944 14112 7056 14224 0 FreeSans 448 0 0 0 N2BEGb[2]
port 119 nsew signal output
flabel metal2 s 7392 14112 7504 14224 0 FreeSans 448 0 0 0 N2BEGb[3]
port 120 nsew signal output
flabel metal2 s 7840 14112 7952 14224 0 FreeSans 448 0 0 0 N2BEGb[4]
port 121 nsew signal output
flabel metal2 s 8288 14112 8400 14224 0 FreeSans 448 0 0 0 N2BEGb[5]
port 122 nsew signal output
flabel metal2 s 8736 14112 8848 14224 0 FreeSans 448 0 0 0 N2BEGb[6]
port 123 nsew signal output
flabel metal2 s 9184 14112 9296 14224 0 FreeSans 448 0 0 0 N2BEGb[7]
port 124 nsew signal output
flabel metal2 s 9632 14112 9744 14224 0 FreeSans 448 0 0 0 N4BEG[0]
port 125 nsew signal output
flabel metal2 s 14112 14112 14224 14224 0 FreeSans 448 0 0 0 N4BEG[10]
port 126 nsew signal output
flabel metal2 s 14560 14112 14672 14224 0 FreeSans 448 0 0 0 N4BEG[11]
port 127 nsew signal output
flabel metal2 s 15008 14112 15120 14224 0 FreeSans 448 0 0 0 N4BEG[12]
port 128 nsew signal output
flabel metal2 s 15456 14112 15568 14224 0 FreeSans 448 0 0 0 N4BEG[13]
port 129 nsew signal output
flabel metal2 s 15904 14112 16016 14224 0 FreeSans 448 0 0 0 N4BEG[14]
port 130 nsew signal output
flabel metal2 s 16352 14112 16464 14224 0 FreeSans 448 0 0 0 N4BEG[15]
port 131 nsew signal output
flabel metal2 s 10080 14112 10192 14224 0 FreeSans 448 0 0 0 N4BEG[1]
port 132 nsew signal output
flabel metal2 s 10528 14112 10640 14224 0 FreeSans 448 0 0 0 N4BEG[2]
port 133 nsew signal output
flabel metal2 s 10976 14112 11088 14224 0 FreeSans 448 0 0 0 N4BEG[3]
port 134 nsew signal output
flabel metal2 s 11424 14112 11536 14224 0 FreeSans 448 0 0 0 N4BEG[4]
port 135 nsew signal output
flabel metal2 s 11872 14112 11984 14224 0 FreeSans 448 0 0 0 N4BEG[5]
port 136 nsew signal output
flabel metal2 s 12320 14112 12432 14224 0 FreeSans 448 0 0 0 N4BEG[6]
port 137 nsew signal output
flabel metal2 s 12768 14112 12880 14224 0 FreeSans 448 0 0 0 N4BEG[7]
port 138 nsew signal output
flabel metal2 s 13216 14112 13328 14224 0 FreeSans 448 0 0 0 N4BEG[8]
port 139 nsew signal output
flabel metal2 s 13664 14112 13776 14224 0 FreeSans 448 0 0 0 N4BEG[9]
port 140 nsew signal output
flabel metal2 s 16800 14112 16912 14224 0 FreeSans 448 0 0 0 NN4BEG[0]
port 141 nsew signal output
flabel metal2 s 21280 14112 21392 14224 0 FreeSans 448 0 0 0 NN4BEG[10]
port 142 nsew signal output
flabel metal2 s 21728 14112 21840 14224 0 FreeSans 448 0 0 0 NN4BEG[11]
port 143 nsew signal output
flabel metal2 s 22176 14112 22288 14224 0 FreeSans 448 0 0 0 NN4BEG[12]
port 144 nsew signal output
flabel metal2 s 22624 14112 22736 14224 0 FreeSans 448 0 0 0 NN4BEG[13]
port 145 nsew signal output
flabel metal2 s 23072 14112 23184 14224 0 FreeSans 448 0 0 0 NN4BEG[14]
port 146 nsew signal output
flabel metal2 s 23520 14112 23632 14224 0 FreeSans 448 0 0 0 NN4BEG[15]
port 147 nsew signal output
flabel metal2 s 17248 14112 17360 14224 0 FreeSans 448 0 0 0 NN4BEG[1]
port 148 nsew signal output
flabel metal2 s 17696 14112 17808 14224 0 FreeSans 448 0 0 0 NN4BEG[2]
port 149 nsew signal output
flabel metal2 s 18144 14112 18256 14224 0 FreeSans 448 0 0 0 NN4BEG[3]
port 150 nsew signal output
flabel metal2 s 18592 14112 18704 14224 0 FreeSans 448 0 0 0 NN4BEG[4]
port 151 nsew signal output
flabel metal2 s 19040 14112 19152 14224 0 FreeSans 448 0 0 0 NN4BEG[5]
port 152 nsew signal output
flabel metal2 s 19488 14112 19600 14224 0 FreeSans 448 0 0 0 NN4BEG[6]
port 153 nsew signal output
flabel metal2 s 19936 14112 20048 14224 0 FreeSans 448 0 0 0 NN4BEG[7]
port 154 nsew signal output
flabel metal2 s 20384 14112 20496 14224 0 FreeSans 448 0 0 0 NN4BEG[8]
port 155 nsew signal output
flabel metal2 s 20832 14112 20944 14224 0 FreeSans 448 0 0 0 NN4BEG[9]
port 156 nsew signal output
flabel metal2 s 24416 14112 24528 14224 0 FreeSans 448 0 0 0 S1END[0]
port 157 nsew signal input
flabel metal2 s 24864 14112 24976 14224 0 FreeSans 448 0 0 0 S1END[1]
port 158 nsew signal input
flabel metal2 s 25312 14112 25424 14224 0 FreeSans 448 0 0 0 S1END[2]
port 159 nsew signal input
flabel metal2 s 25760 14112 25872 14224 0 FreeSans 448 0 0 0 S1END[3]
port 160 nsew signal input
flabel metal2 s 29792 14112 29904 14224 0 FreeSans 448 0 0 0 S2END[0]
port 161 nsew signal input
flabel metal2 s 30240 14112 30352 14224 0 FreeSans 448 0 0 0 S2END[1]
port 162 nsew signal input
flabel metal2 s 30688 14112 30800 14224 0 FreeSans 448 0 0 0 S2END[2]
port 163 nsew signal input
flabel metal2 s 31136 14112 31248 14224 0 FreeSans 448 0 0 0 S2END[3]
port 164 nsew signal input
flabel metal2 s 31584 14112 31696 14224 0 FreeSans 448 0 0 0 S2END[4]
port 165 nsew signal input
flabel metal2 s 32032 14112 32144 14224 0 FreeSans 448 0 0 0 S2END[5]
port 166 nsew signal input
flabel metal2 s 32480 14112 32592 14224 0 FreeSans 448 0 0 0 S2END[6]
port 167 nsew signal input
flabel metal2 s 32928 14112 33040 14224 0 FreeSans 448 0 0 0 S2END[7]
port 168 nsew signal input
flabel metal2 s 26208 14112 26320 14224 0 FreeSans 448 0 0 0 S2MID[0]
port 169 nsew signal input
flabel metal2 s 26656 14112 26768 14224 0 FreeSans 448 0 0 0 S2MID[1]
port 170 nsew signal input
flabel metal2 s 27104 14112 27216 14224 0 FreeSans 448 0 0 0 S2MID[2]
port 171 nsew signal input
flabel metal2 s 27552 14112 27664 14224 0 FreeSans 448 0 0 0 S2MID[3]
port 172 nsew signal input
flabel metal2 s 28000 14112 28112 14224 0 FreeSans 448 0 0 0 S2MID[4]
port 173 nsew signal input
flabel metal2 s 28448 14112 28560 14224 0 FreeSans 448 0 0 0 S2MID[5]
port 174 nsew signal input
flabel metal2 s 28896 14112 29008 14224 0 FreeSans 448 0 0 0 S2MID[6]
port 175 nsew signal input
flabel metal2 s 29344 14112 29456 14224 0 FreeSans 448 0 0 0 S2MID[7]
port 176 nsew signal input
flabel metal2 s 33376 14112 33488 14224 0 FreeSans 448 0 0 0 S4END[0]
port 177 nsew signal input
flabel metal2 s 37856 14112 37968 14224 0 FreeSans 448 0 0 0 S4END[10]
port 178 nsew signal input
flabel metal2 s 38304 14112 38416 14224 0 FreeSans 448 0 0 0 S4END[11]
port 179 nsew signal input
flabel metal2 s 38752 14112 38864 14224 0 FreeSans 448 0 0 0 S4END[12]
port 180 nsew signal input
flabel metal2 s 39200 14112 39312 14224 0 FreeSans 448 0 0 0 S4END[13]
port 181 nsew signal input
flabel metal2 s 39648 14112 39760 14224 0 FreeSans 448 0 0 0 S4END[14]
port 182 nsew signal input
flabel metal2 s 40096 14112 40208 14224 0 FreeSans 448 0 0 0 S4END[15]
port 183 nsew signal input
flabel metal2 s 33824 14112 33936 14224 0 FreeSans 448 0 0 0 S4END[1]
port 184 nsew signal input
flabel metal2 s 34272 14112 34384 14224 0 FreeSans 448 0 0 0 S4END[2]
port 185 nsew signal input
flabel metal2 s 34720 14112 34832 14224 0 FreeSans 448 0 0 0 S4END[3]
port 186 nsew signal input
flabel metal2 s 35168 14112 35280 14224 0 FreeSans 448 0 0 0 S4END[4]
port 187 nsew signal input
flabel metal2 s 35616 14112 35728 14224 0 FreeSans 448 0 0 0 S4END[5]
port 188 nsew signal input
flabel metal2 s 36064 14112 36176 14224 0 FreeSans 448 0 0 0 S4END[6]
port 189 nsew signal input
flabel metal2 s 36512 14112 36624 14224 0 FreeSans 448 0 0 0 S4END[7]
port 190 nsew signal input
flabel metal2 s 36960 14112 37072 14224 0 FreeSans 448 0 0 0 S4END[8]
port 191 nsew signal input
flabel metal2 s 37408 14112 37520 14224 0 FreeSans 448 0 0 0 S4END[9]
port 192 nsew signal input
flabel metal2 s 40544 14112 40656 14224 0 FreeSans 448 0 0 0 SS4END[0]
port 193 nsew signal input
flabel metal2 s 45024 14112 45136 14224 0 FreeSans 448 0 0 0 SS4END[10]
port 194 nsew signal input
flabel metal2 s 45472 14112 45584 14224 0 FreeSans 448 0 0 0 SS4END[11]
port 195 nsew signal input
flabel metal2 s 45920 14112 46032 14224 0 FreeSans 448 0 0 0 SS4END[12]
port 196 nsew signal input
flabel metal2 s 46368 14112 46480 14224 0 FreeSans 448 0 0 0 SS4END[13]
port 197 nsew signal input
flabel metal2 s 46816 14112 46928 14224 0 FreeSans 448 0 0 0 SS4END[14]
port 198 nsew signal input
flabel metal2 s 47264 14112 47376 14224 0 FreeSans 448 0 0 0 SS4END[15]
port 199 nsew signal input
flabel metal2 s 40992 14112 41104 14224 0 FreeSans 448 0 0 0 SS4END[1]
port 200 nsew signal input
flabel metal2 s 41440 14112 41552 14224 0 FreeSans 448 0 0 0 SS4END[2]
port 201 nsew signal input
flabel metal2 s 41888 14112 42000 14224 0 FreeSans 448 0 0 0 SS4END[3]
port 202 nsew signal input
flabel metal2 s 42336 14112 42448 14224 0 FreeSans 448 0 0 0 SS4END[4]
port 203 nsew signal input
flabel metal2 s 42784 14112 42896 14224 0 FreeSans 448 0 0 0 SS4END[5]
port 204 nsew signal input
flabel metal2 s 43232 14112 43344 14224 0 FreeSans 448 0 0 0 SS4END[6]
port 205 nsew signal input
flabel metal2 s 43680 14112 43792 14224 0 FreeSans 448 0 0 0 SS4END[7]
port 206 nsew signal input
flabel metal2 s 44128 14112 44240 14224 0 FreeSans 448 0 0 0 SS4END[8]
port 207 nsew signal input
flabel metal2 s 44576 14112 44688 14224 0 FreeSans 448 0 0 0 SS4END[9]
port 208 nsew signal input
flabel metal2 s 1792 0 1904 112 0 FreeSans 448 0 0 0 UserCLK
port 209 nsew signal input
flabel metal2 s 47712 14112 47824 14224 0 FreeSans 448 0 0 0 UserCLKo
port 210 nsew signal output
flabel metal4 s 3776 0 4096 14224 0 FreeSans 1472 90 0 0 VDD
port 211 nsew power bidirectional
flabel metal4 s 3776 0 4096 56 0 FreeSans 368 0 0 0 VDD
port 211 nsew power bidirectional
flabel metal4 s 3776 14168 4096 14224 0 FreeSans 368 0 0 0 VDD
port 211 nsew power bidirectional
flabel metal4 s 23776 0 24096 14224 0 FreeSans 1472 90 0 0 VDD
port 211 nsew power bidirectional
flabel metal4 s 23776 0 24096 56 0 FreeSans 368 0 0 0 VDD
port 211 nsew power bidirectional
flabel metal4 s 23776 14168 24096 14224 0 FreeSans 368 0 0 0 VDD
port 211 nsew power bidirectional
flabel metal4 s 43776 0 44096 14224 0 FreeSans 1472 90 0 0 VDD
port 211 nsew power bidirectional
flabel metal4 s 43776 0 44096 56 0 FreeSans 368 0 0 0 VDD
port 211 nsew power bidirectional
flabel metal4 s 43776 14168 44096 14224 0 FreeSans 368 0 0 0 VDD
port 211 nsew power bidirectional
flabel metal4 s 4436 0 4756 14224 0 FreeSans 1472 90 0 0 VSS
port 212 nsew ground bidirectional
flabel metal4 s 4436 0 4756 56 0 FreeSans 368 0 0 0 VSS
port 212 nsew ground bidirectional
flabel metal4 s 4436 14168 4756 14224 0 FreeSans 368 0 0 0 VSS
port 212 nsew ground bidirectional
flabel metal4 s 24436 0 24756 14224 0 FreeSans 1472 90 0 0 VSS
port 212 nsew ground bidirectional
flabel metal4 s 24436 0 24756 56 0 FreeSans 368 0 0 0 VSS
port 212 nsew ground bidirectional
flabel metal4 s 24436 14168 24756 14224 0 FreeSans 368 0 0 0 VSS
port 212 nsew ground bidirectional
flabel metal4 s 44436 0 44756 14224 0 FreeSans 1472 90 0 0 VSS
port 212 nsew ground bidirectional
flabel metal4 s 44436 0 44756 56 0 FreeSans 368 0 0 0 VSS
port 212 nsew ground bidirectional
flabel metal4 s 44436 14168 44756 14224 0 FreeSans 368 0 0 0 VSS
port 212 nsew ground bidirectional
rlabel metal1 28728 12544 28728 12544 0 VDD
rlabel metal1 28728 13328 28728 13328 0 VSS
rlabel metal3 630 56 630 56 0 FrameData[0]
rlabel metal2 15512 4984 15512 4984 0 FrameData[10]
rlabel metal3 854 4984 854 4984 0 FrameData[11]
rlabel metal3 126 5432 126 5432 0 FrameData[12]
rlabel metal3 11368 1400 11368 1400 0 FrameData[13]
rlabel metal3 1694 6328 1694 6328 0 FrameData[14]
rlabel metal2 24024 11200 24024 11200 0 FrameData[15]
rlabel metal3 47544 3304 47544 3304 0 FrameData[16]
rlabel metal3 854 7672 854 7672 0 FrameData[17]
rlabel metal3 798 8120 798 8120 0 FrameData[18]
rlabel metal3 1134 8568 1134 8568 0 FrameData[19]
rlabel metal3 854 504 854 504 0 FrameData[1]
rlabel metal3 1246 9016 1246 9016 0 FrameData[20]
rlabel metal3 182 9464 182 9464 0 FrameData[21]
rlabel metal3 854 9912 854 9912 0 FrameData[22]
rlabel metal3 1456 5208 1456 5208 0 FrameData[23]
rlabel metal3 462 10808 462 10808 0 FrameData[24]
rlabel metal2 23240 7336 23240 7336 0 FrameData[25]
rlabel metal4 15176 11859 15176 11859 0 FrameData[26]
rlabel metal3 574 12152 574 12152 0 FrameData[27]
rlabel metal3 518 12600 518 12600 0 FrameData[28]
rlabel metal3 238 13048 238 13048 0 FrameData[29]
rlabel metal3 574 952 574 952 0 FrameData[2]
rlabel metal3 854 13496 854 13496 0 FrameData[30]
rlabel metal3 798 13944 798 13944 0 FrameData[31]
rlabel metal3 2142 1400 2142 1400 0 FrameData[3]
rlabel metal3 1414 1848 1414 1848 0 FrameData[4]
rlabel metal3 1638 2296 1638 2296 0 FrameData[5]
rlabel metal3 4214 2744 4214 2744 0 FrameData[6]
rlabel metal3 1862 3192 1862 3192 0 FrameData[7]
rlabel metal3 350 3640 350 3640 0 FrameData[8]
rlabel metal3 1694 4088 1694 4088 0 FrameData[9]
rlabel metal3 56938 56 56938 56 0 FrameData_O[0]
rlabel metal3 55986 4536 55986 4536 0 FrameData_O[10]
rlabel metal3 56714 4984 56714 4984 0 FrameData_O[11]
rlabel metal2 56168 4984 56168 4984 0 FrameData_O[12]
rlabel metal3 55986 5880 55986 5880 0 FrameData_O[13]
rlabel metal3 56266 6328 56266 6328 0 FrameData_O[14]
rlabel metal2 56168 6440 56168 6440 0 FrameData_O[15]
rlabel metal3 55986 7224 55986 7224 0 FrameData_O[16]
rlabel metal3 56770 7672 56770 7672 0 FrameData_O[17]
rlabel metal3 56658 8120 56658 8120 0 FrameData_O[18]
rlabel metal3 55874 8568 55874 8568 0 FrameData_O[19]
rlabel metal3 57106 504 57106 504 0 FrameData_O[1]
rlabel metal3 56770 9016 56770 9016 0 FrameData_O[20]
rlabel metal3 56266 9464 56266 9464 0 FrameData_O[21]
rlabel metal3 56602 9912 56602 9912 0 FrameData_O[22]
rlabel metal2 55160 8232 55160 8232 0 FrameData_O[23]
rlabel metal3 53704 9912 53704 9912 0 FrameData_O[24]
rlabel metal3 54544 8344 54544 8344 0 FrameData_O[25]
rlabel metal2 49224 11312 49224 11312 0 FrameData_O[26]
rlabel metal2 53032 7728 53032 7728 0 FrameData_O[27]
rlabel metal3 52976 8120 52976 8120 0 FrameData_O[28]
rlabel metal2 49672 10920 49672 10920 0 FrameData_O[29]
rlabel metal2 52024 1120 52024 1120 0 FrameData_O[2]
rlabel metal2 50232 10080 50232 10080 0 FrameData_O[30]
rlabel metal2 51240 9296 51240 9296 0 FrameData_O[31]
rlabel metal3 55482 1400 55482 1400 0 FrameData_O[3]
rlabel metal3 55482 1848 55482 1848 0 FrameData_O[4]
rlabel metal2 54936 2184 54936 2184 0 FrameData_O[5]
rlabel metal2 56168 2072 56168 2072 0 FrameData_O[6]
rlabel metal2 54600 3080 54600 3080 0 FrameData_O[7]
rlabel metal3 56154 3640 56154 3640 0 FrameData_O[8]
rlabel metal3 56770 4088 56770 4088 0 FrameData_O[9]
rlabel metal3 4984 616 4984 616 0 FrameStrobe[0]
rlabel metal2 31416 126 31416 126 0 FrameStrobe[10]
rlabel metal2 31192 1736 31192 1736 0 FrameStrobe[11]
rlabel metal2 36792 238 36792 238 0 FrameStrobe[12]
rlabel metal2 39480 686 39480 686 0 FrameStrobe[13]
rlabel metal2 40488 6160 40488 6160 0 FrameStrobe[14]
rlabel metal2 44856 574 44856 574 0 FrameStrobe[15]
rlabel metal3 49336 1624 49336 1624 0 FrameStrobe[16]
rlabel metal2 50232 126 50232 126 0 FrameStrobe[17]
rlabel metal2 52920 462 52920 462 0 FrameStrobe[18]
rlabel metal2 55608 406 55608 406 0 FrameStrobe[19]
rlabel metal2 5040 2520 5040 2520 0 FrameStrobe[1]
rlabel metal2 9968 3304 9968 3304 0 FrameStrobe[2]
rlabel metal2 14840 4872 14840 4872 0 FrameStrobe[3]
rlabel metal2 15176 3584 15176 3584 0 FrameStrobe[4]
rlabel metal2 17976 238 17976 238 0 FrameStrobe[5]
rlabel metal2 20664 518 20664 518 0 FrameStrobe[6]
rlabel metal2 1232 4536 1232 4536 0 FrameStrobe[7]
rlabel metal3 18648 10136 18648 10136 0 FrameStrobe[8]
rlabel metal3 21224 10360 21224 10360 0 FrameStrobe[9]
rlabel metal2 48216 13650 48216 13650 0 FrameStrobe_O[0]
rlabel metal2 52696 13538 52696 13538 0 FrameStrobe_O[10]
rlabel metal2 53144 13258 53144 13258 0 FrameStrobe_O[11]
rlabel metal2 53648 9688 53648 9688 0 FrameStrobe_O[12]
rlabel metal3 53536 9240 53536 9240 0 FrameStrobe_O[13]
rlabel metal2 51240 11312 51240 11312 0 FrameStrobe_O[14]
rlabel metal2 47880 13104 47880 13104 0 FrameStrobe_O[15]
rlabel metal2 47992 12712 47992 12712 0 FrameStrobe_O[16]
rlabel metal2 53592 7504 53592 7504 0 FrameStrobe_O[17]
rlabel metal2 45976 12600 45976 12600 0 FrameStrobe_O[18]
rlabel metal3 54880 6104 54880 6104 0 FrameStrobe_O[19]
rlabel metal2 48664 13258 48664 13258 0 FrameStrobe_O[1]
rlabel metal2 49112 13874 49112 13874 0 FrameStrobe_O[2]
rlabel metal3 49952 11592 49952 11592 0 FrameStrobe_O[3]
rlabel metal2 50008 13818 50008 13818 0 FrameStrobe_O[4]
rlabel metal2 50456 13258 50456 13258 0 FrameStrobe_O[5]
rlabel metal2 50904 12866 50904 12866 0 FrameStrobe_O[6]
rlabel metal2 51352 12922 51352 12922 0 FrameStrobe_O[7]
rlabel metal2 51800 13594 51800 13594 0 FrameStrobe_O[8]
rlabel metal2 52248 13650 52248 13650 0 FrameStrobe_O[9]
rlabel metal2 728 11914 728 11914 0 N1BEG[0]
rlabel metal2 2072 9352 2072 9352 0 N1BEG[1]
rlabel metal2 1624 12978 1624 12978 0 N1BEG[2]
rlabel metal2 2184 11368 2184 11368 0 N1BEG[3]
rlabel metal2 2520 12698 2520 12698 0 N2BEG[0]
rlabel metal2 2968 13146 2968 13146 0 N2BEG[1]
rlabel metal2 3416 13258 3416 13258 0 N2BEG[2]
rlabel metal2 3864 13426 3864 13426 0 N2BEG[3]
rlabel metal2 2184 13272 2184 13272 0 N2BEG[4]
rlabel metal2 4760 13818 4760 13818 0 N2BEG[5]
rlabel metal3 4872 11592 4872 11592 0 N2BEG[6]
rlabel metal2 5656 13650 5656 13650 0 N2BEG[7]
rlabel metal2 6104 12418 6104 12418 0 N2BEGb[0]
rlabel metal2 6216 12376 6216 12376 0 N2BEGb[1]
rlabel metal2 7448 11704 7448 11704 0 N2BEGb[2]
rlabel metal2 5992 13216 5992 13216 0 N2BEGb[3]
rlabel metal2 7896 13258 7896 13258 0 N2BEGb[4]
rlabel metal2 7896 11592 7896 11592 0 N2BEGb[5]
rlabel metal2 9016 11299 9016 11299 0 N2BEGb[6]
rlabel metal3 8400 13160 8400 13160 0 N2BEGb[7]
rlabel metal2 9688 13258 9688 13258 0 N4BEG[0]
rlabel metal3 14392 10808 14392 10808 0 N4BEG[10]
rlabel metal3 14168 13048 14168 13048 0 N4BEG[11]
rlabel metal2 15064 13258 15064 13258 0 N4BEG[12]
rlabel metal2 15512 12866 15512 12866 0 N4BEG[13]
rlabel metal2 15960 12474 15960 12474 0 N4BEG[14]
rlabel metal2 16408 13594 16408 13594 0 N4BEG[15]
rlabel metal2 10584 11480 10584 11480 0 N4BEG[1]
rlabel metal2 10584 13258 10584 13258 0 N4BEG[2]
rlabel metal2 10976 11592 10976 11592 0 N4BEG[3]
rlabel metal3 10640 13160 10640 13160 0 N4BEG[4]
rlabel metal2 11928 13650 11928 13650 0 N4BEG[5]
rlabel metal2 12376 12698 12376 12698 0 N4BEG[6]
rlabel metal2 12992 10808 12992 10808 0 N4BEG[7]
rlabel metal2 11368 13272 11368 13272 0 N4BEG[8]
rlabel metal2 13720 13706 13720 13706 0 N4BEG[9]
rlabel metal2 16800 12376 16800 12376 0 NN4BEG[0]
rlabel metal2 21336 12698 21336 12698 0 NN4BEG[10]
rlabel metal3 21504 13160 21504 13160 0 NN4BEG[11]
rlabel metal2 22232 13258 22232 13258 0 NN4BEG[12]
rlabel metal2 22680 13650 22680 13650 0 NN4BEG[13]
rlabel metal2 23128 13258 23128 13258 0 NN4BEG[14]
rlabel metal2 23576 13594 23576 13594 0 NN4BEG[15]
rlabel metal2 17304 13538 17304 13538 0 NN4BEG[1]
rlabel metal2 17752 13202 17752 13202 0 NN4BEG[2]
rlabel metal2 18200 13202 18200 13202 0 NN4BEG[3]
rlabel metal3 18088 13048 18088 13048 0 NN4BEG[4]
rlabel metal2 19096 12698 19096 12698 0 NN4BEG[5]
rlabel metal2 19544 13202 19544 13202 0 NN4BEG[6]
rlabel metal3 19656 12824 19656 12824 0 NN4BEG[7]
rlabel metal2 20440 12866 20440 12866 0 NN4BEG[8]
rlabel metal2 20888 12474 20888 12474 0 NN4BEG[9]
rlabel metal2 24472 13818 24472 13818 0 S1END[0]
rlabel metal2 24920 13762 24920 13762 0 S1END[1]
rlabel metal2 25592 2744 25592 2744 0 S1END[2]
rlabel metal2 25816 13986 25816 13986 0 S1END[3]
rlabel metal2 41384 6440 41384 6440 0 S2END[0]
rlabel metal4 38920 11424 38920 11424 0 S2END[1]
rlabel metal2 45752 12880 45752 12880 0 S2END[2]
rlabel metal3 29960 5320 29960 5320 0 S2END[3]
rlabel metal3 33768 10024 33768 10024 0 S2END[4]
rlabel metal2 21504 2184 21504 2184 0 S2END[5]
rlabel metal2 34496 8344 34496 8344 0 S2END[6]
rlabel metal2 23240 8512 23240 8512 0 S2END[7]
rlabel metal2 26264 13706 26264 13706 0 S2MID[0]
rlabel metal2 26712 12362 26712 12362 0 S2MID[1]
rlabel metal2 37352 12768 37352 12768 0 S2MID[2]
rlabel metal3 35728 4424 35728 4424 0 S2MID[3]
rlabel metal2 30744 11704 30744 11704 0 S2MID[4]
rlabel metal2 50008 12376 50008 12376 0 S2MID[5]
rlabel metal2 48328 9632 48328 9632 0 S2MID[6]
rlabel metal2 51464 1792 51464 1792 0 S2MID[7]
rlabel metal2 22120 8176 22120 8176 0 S4END[0]
rlabel metal2 35672 7784 35672 7784 0 S4END[10]
rlabel metal2 46536 12096 46536 12096 0 S4END[11]
rlabel metal2 38808 13706 38808 13706 0 S4END[12]
rlabel metal2 39256 13314 39256 13314 0 S4END[13]
rlabel metal2 20888 9744 20888 9744 0 S4END[14]
rlabel metal2 20888 7784 20888 7784 0 S4END[15]
rlabel metal3 20720 2296 20720 2296 0 S4END[1]
rlabel metal2 15176 5936 15176 5936 0 S4END[2]
rlabel metal2 17752 10920 17752 10920 0 S4END[3]
rlabel metal4 15960 9352 15960 9352 0 S4END[4]
rlabel metal2 20552 6944 20552 6944 0 S4END[5]
rlabel metal3 16296 7056 16296 7056 0 S4END[6]
rlabel metal3 44296 8624 44296 8624 0 S4END[7]
rlabel metal2 19768 7952 19768 7952 0 S4END[8]
rlabel metal2 43736 3808 43736 3808 0 S4END[9]
rlabel metal2 26320 10024 26320 10024 0 SS4END[0]
rlabel metal2 45080 11858 45080 11858 0 SS4END[10]
rlabel metal3 12684 3192 12684 3192 0 SS4END[11]
rlabel metal3 3584 1960 3584 1960 0 SS4END[12]
rlabel metal3 5152 1288 5152 1288 0 SS4END[13]
rlabel metal2 13160 1512 13160 1512 0 SS4END[14]
rlabel metal4 15176 5400 15176 5400 0 SS4END[15]
rlabel metal2 7280 2184 7280 2184 0 SS4END[1]
rlabel metal4 16744 5040 16744 5040 0 SS4END[2]
rlabel metal3 2800 5320 2800 5320 0 SS4END[3]
rlabel metal2 42392 13370 42392 13370 0 SS4END[4]
rlabel metal2 42840 13202 42840 13202 0 SS4END[5]
rlabel metal2 15288 7616 15288 7616 0 SS4END[6]
rlabel metal3 14448 2184 14448 2184 0 SS4END[7]
rlabel metal2 14168 1624 14168 1624 0 SS4END[8]
rlabel metal2 21336 616 21336 616 0 SS4END[9]
rlabel metal2 1848 126 1848 126 0 UserCLK
rlabel metal2 47656 11592 47656 11592 0 UserCLKo
rlabel metal3 49112 3080 49112 3080 0 net1
rlabel metal2 40376 2016 40376 2016 0 net10
rlabel metal2 18536 11424 18536 11424 0 net100
rlabel metal2 18872 12544 18872 12544 0 net101
rlabel metal2 3136 9128 3136 9128 0 net102
rlabel metal2 16184 8008 16184 8008 0 net103
rlabel metal2 17976 12208 17976 12208 0 net104
rlabel metal2 1624 9912 1624 9912 0 net105
rlabel metal3 25480 13104 25480 13104 0 net106
rlabel metal3 45080 1680 45080 1680 0 net11
rlabel metal4 45192 4424 45192 4424 0 net12
rlabel metal3 53984 5208 53984 5208 0 net13
rlabel metal2 28056 1624 28056 1624 0 net14
rlabel metal3 24304 3304 24304 3304 0 net15
rlabel metal2 43848 7336 43848 7336 0 net16
rlabel metal4 26376 2576 26376 2576 0 net17
rlabel metal4 43400 7896 43400 7896 0 net18
rlabel metal3 41608 11368 41608 11368 0 net19
rlabel metal2 42280 3920 42280 3920 0 net2
rlabel metal2 39928 4480 39928 4480 0 net20
rlabel metal3 50008 8344 50008 8344 0 net21
rlabel metal2 22120 3080 22120 3080 0 net22
rlabel metal2 51128 7784 51128 7784 0 net23
rlabel metal2 40264 10080 40264 10080 0 net24
rlabel metal2 49896 5488 49896 5488 0 net25
rlabel metal3 49952 1288 49952 1288 0 net26
rlabel metal3 50120 2968 50120 2968 0 net27
rlabel metal2 54152 2296 54152 2296 0 net28
rlabel metal2 49560 7448 49560 7448 0 net29
rlabel metal2 48328 6944 48328 6944 0 net3
rlabel metal3 51632 2744 51632 2744 0 net30
rlabel metal2 54432 3528 54432 3528 0 net31
rlabel metal3 49448 1456 49448 1456 0 net32
rlabel metal3 16520 6384 16520 6384 0 net33
rlabel metal2 16520 6160 16520 6160 0 net34
rlabel metal3 48076 2184 48076 2184 0 net35
rlabel metal4 40600 9520 40600 9520 0 net36
rlabel metal2 47544 5936 47544 5936 0 net37
rlabel metal2 50232 10640 50232 10640 0 net38
rlabel metal2 42280 2296 42280 2296 0 net39
rlabel metal2 21784 3136 21784 3136 0 net4
rlabel metal2 48664 7616 48664 7616 0 net40
rlabel metal2 52696 7784 52696 7784 0 net41
rlabel metal2 40264 11928 40264 11928 0 net42
rlabel metal3 43848 1960 43848 1960 0 net43
rlabel metal4 6776 2016 6776 2016 0 net44
rlabel metal2 25256 1176 25256 1176 0 net45
rlabel metal2 15624 7056 15624 7056 0 net46
rlabel metal4 25032 11592 25032 11592 0 net47
rlabel metal4 15512 11760 15512 11760 0 net48
rlabel metal2 20888 7056 20888 7056 0 net49
rlabel metal4 37576 5824 37576 5824 0 net5
rlabel metal2 15176 12768 15176 12768 0 net50
rlabel metal4 19880 9325 19880 9325 0 net51
rlabel metal2 19656 10976 19656 10976 0 net52
rlabel metal4 2296 6608 2296 6608 0 net53
rlabel metal3 2632 8512 2632 8512 0 net54
rlabel metal2 25368 8064 25368 8064 0 net55
rlabel metal2 2856 8288 2856 8288 0 net56
rlabel metal2 44296 1344 44296 1344 0 net57
rlabel metal2 49000 9296 49000 9296 0 net58
rlabel metal2 2968 10864 2968 10864 0 net59
rlabel metal2 54152 6216 54152 6216 0 net6
rlabel metal2 15176 9744 15176 9744 0 net60
rlabel metal3 3360 2520 3360 2520 0 net61
rlabel metal2 24192 5992 24192 5992 0 net62
rlabel metal3 19320 2520 19320 2520 0 net63
rlabel metal3 14952 3808 14952 3808 0 net64
rlabel metal2 22456 8848 22456 8848 0 net65
rlabel metal2 19992 9632 19992 9632 0 net66
rlabel metal3 14448 2072 14448 2072 0 net67
rlabel metal4 15176 11309 15176 11309 0 net68
rlabel metal2 19208 7000 19208 7000 0 net69
rlabel metal2 52248 1456 52248 1456 0 net7
rlabel metal3 13384 2856 13384 2856 0 net70
rlabel metal3 49224 1176 49224 1176 0 net71
rlabel metal2 21896 5880 21896 5880 0 net72
rlabel metal2 19992 8008 19992 8008 0 net73
rlabel metal2 19656 7224 19656 7224 0 net74
rlabel metal2 9464 11424 9464 11424 0 net75
rlabel metal2 16968 10864 16968 10864 0 net76
rlabel metal2 14392 8680 14392 8680 0 net77
rlabel metal2 16184 10640 16184 10640 0 net78
rlabel metal3 18816 8232 18816 8232 0 net79
rlabel metal2 50568 4144 50568 4144 0 net8
rlabel metal2 20328 10192 20328 10192 0 net80
rlabel metal2 16632 8120 16632 8120 0 net81
rlabel metal4 15400 8155 15400 8155 0 net82
rlabel metal2 38696 1792 38696 1792 0 net83
rlabel metal3 21280 1736 21280 1736 0 net84
rlabel metal3 43400 3416 43400 3416 0 net85
rlabel metal3 17864 7560 17864 7560 0 net86
rlabel metal2 45864 2184 45864 2184 0 net87
rlabel metal2 13552 5992 13552 5992 0 net88
rlabel metal2 15848 12824 15848 12824 0 net89
rlabel metal3 31472 5208 31472 5208 0 net9
rlabel metal2 22792 10696 22792 10696 0 net90
rlabel metal2 24920 12320 24920 12320 0 net91
rlabel metal2 2072 7056 2072 7056 0 net92
rlabel metal2 15176 3976 15176 3976 0 net93
rlabel metal2 13384 2072 13384 2072 0 net94
rlabel metal2 25480 9912 25480 9912 0 net95
rlabel metal2 16856 11592 16856 11592 0 net96
rlabel metal2 2128 1848 2128 1848 0 net97
rlabel metal2 2856 3808 2856 3808 0 net98
rlabel metal2 16968 12712 16968 12712 0 net99
<< properties >>
string FIXED_BBOX 0 0 57456 14224
<< end >>
