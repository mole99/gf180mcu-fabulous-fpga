module LUT4AB (Ci,
    Co,
    UserCLK,
    UserCLKo,
    VDD,
    VSS,
    E1BEG,
    E1END,
    E2BEG,
    E2BEGb,
    E2END,
    E2MID,
    E6BEG,
    E6END,
    EE4BEG,
    EE4END,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N1END,
    N2BEG,
    N2BEGb,
    N2END,
    N2MID,
    N4BEG,
    N4END,
    NN4BEG,
    NN4END,
    S1BEG,
    S1END,
    S2BEG,
    S2BEGb,
    S2END,
    S2MID,
    S4BEG,
    S4END,
    SS4BEG,
    SS4END,
    W1BEG,
    W1END,
    W2BEG,
    W2BEGb,
    W2END,
    W2MID,
    W6BEG,
    W6END,
    WW4BEG,
    WW4END);
 input Ci;
 output Co;
 input UserCLK;
 output UserCLKo;
 inout VDD;
 inout VSS;
 output [3:0] E1BEG;
 input [3:0] E1END;
 output [7:0] E2BEG;
 output [7:0] E2BEGb;
 input [7:0] E2END;
 input [7:0] E2MID;
 output [11:0] E6BEG;
 input [11:0] E6END;
 output [15:0] EE4BEG;
 input [15:0] EE4END;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 input [3:0] N1END;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 input [7:0] N2END;
 input [7:0] N2MID;
 output [15:0] N4BEG;
 input [15:0] N4END;
 output [15:0] NN4BEG;
 input [15:0] NN4END;
 output [3:0] S1BEG;
 input [3:0] S1END;
 output [7:0] S2BEG;
 output [7:0] S2BEGb;
 input [7:0] S2END;
 input [7:0] S2MID;
 output [15:0] S4BEG;
 input [15:0] S4END;
 output [15:0] SS4BEG;
 input [15:0] SS4END;
 output [3:0] W1BEG;
 input [3:0] W1END;
 output [7:0] W2BEG;
 output [7:0] W2BEGb;
 input [7:0] W2END;
 input [7:0] W2MID;
 output [11:0] W6BEG;
 input [11:0] W6END;
 output [15:0] WW4BEG;
 input [15:0] WW4END;

 wire A;
 wire B;
 wire C;
 wire net1;
 wire D;
 wire E;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire F;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire G;
 wire H;
 wire \Inst_LA_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.c_I0mux ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.c_out_mux ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.c_reset_value ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame11_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame12_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame14_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame3_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame5_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame6_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame7_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit10.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit12.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit13.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit14.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit18.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit19.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit2.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit20.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit22.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit23.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit24.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit28.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit29.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit3.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit31.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit4.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit5.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit6.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit7.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit8.Q ;
 wire \Inst_LUT4AB_ConfigMem.Inst_frame9_bit9.Q ;
 wire \Inst_LUT4AB_switch_matrix.E1BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.E1BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.E1BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.E1BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG4 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG5 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG6 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG7 ;
 wire \Inst_LUT4AB_switch_matrix.E6BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.E6BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.EE4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.EE4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.EE4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.EE4BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG4 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG5 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG6 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG7 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG4 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG5 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG6 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG7 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG4 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG5 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG6 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG7 ;
 wire \Inst_LUT4AB_switch_matrix.M_AB ;
 wire \Inst_LUT4AB_switch_matrix.M_AD ;
 wire \Inst_LUT4AB_switch_matrix.M_AH ;
 wire \Inst_LUT4AB_switch_matrix.M_EF ;
 wire \Inst_LUT4AB_switch_matrix.N1BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.N1BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.N1BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.N1BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.N4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.N4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.N4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.N4BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.NN4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.NN4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.NN4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.NN4BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.S1BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.S1BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.S1BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.S1BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.S4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.S4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.S4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.S4BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.SS4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.SS4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.SS4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.SS4BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.W1BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.W1BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.W1BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.W1BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.W6BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.W6BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.WW4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.WW4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.WW4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.WW4BEG3 ;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire UserCLK_regs;
 wire clknet_0_UserCLK;
 wire clknet_1_0__leaf_UserCLK;
 wire clknet_0_UserCLK_regs;
 wire clknet_1_0__leaf_UserCLK_regs;
 wire clknet_1_1__leaf_UserCLK_regs;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0859_ (.I(S2MID[6]),
    .ZN(_0707_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0860_ (.I(W2MID[6]),
    .ZN(_0708_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0861_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q ),
    .ZN(_0709_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0862_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q ),
    .ZN(_0710_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0863_ (.I(N2MID[7]),
    .ZN(_0711_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0864_ (.I(S2MID[7]),
    .ZN(_0712_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0865_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q ),
    .ZN(_0713_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0866_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q ),
    .ZN(_0714_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0867_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q ),
    .ZN(_0715_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0868_ (.I(S2MID[3]),
    .ZN(_0716_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0869_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q ),
    .ZN(_0717_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0870_ (.I(E2MID[4]),
    .ZN(_0718_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0871_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q ),
    .ZN(_0719_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0872_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q ),
    .ZN(_0720_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0873_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q ),
    .ZN(_0721_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0874_ (.I(E6END[1]),
    .ZN(_0722_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0875_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q ),
    .ZN(_0723_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0876_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q ),
    .ZN(_0724_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0877_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit7.Q ),
    .ZN(_0725_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0878_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q ),
    .ZN(_0726_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0879_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q ),
    .ZN(_0727_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0880_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q ),
    .ZN(_0728_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0881_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q ),
    .ZN(_0729_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0882_ (.I(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .ZN(_0730_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0883_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q ),
    .ZN(_0731_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0884_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q ),
    .ZN(_0732_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0885_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ),
    .ZN(_0733_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0886_ (.I(\Inst_LA_LUT4c_frame_config_dffesr.LUT_flop ),
    .ZN(_0734_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0887_ (.I(\Inst_LB_LUT4c_frame_config_dffesr.c_I0mux ),
    .ZN(_0735_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0888_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit18.Q ),
    .ZN(_0736_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0889_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q ),
    .ZN(_0737_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0890_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q ),
    .ZN(_0738_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0891_ (.I(S2END[6]),
    .ZN(_0739_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0892_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q ),
    .ZN(_0740_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0893_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q ),
    .ZN(_0741_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0894_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q ),
    .ZN(_0742_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0895_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q ),
    .ZN(_0743_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0896_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q ),
    .ZN(_0744_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0897_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q ),
    .ZN(_0745_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0898_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q ),
    .ZN(_0746_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0899_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit13.Q ),
    .ZN(_0747_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0900_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q ),
    .ZN(_0748_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0901_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit5.Q ),
    .ZN(_0749_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0902_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q ),
    .ZN(_0750_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0903_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q ),
    .ZN(_0751_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0904_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q ),
    .ZN(_0752_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0905_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q ),
    .ZN(_0753_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0906_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q ),
    .ZN(_0754_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0907_ (.I(\Inst_LE_LUT4c_frame_config_dffesr.c_I0mux ),
    .ZN(_0755_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0908_ (.I(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .ZN(_0756_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0909_ (.I(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .ZN(_0757_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0910_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q ),
    .ZN(_0758_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0911_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q ),
    .ZN(_0759_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0912_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q ),
    .ZN(_0760_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0913_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q ),
    .ZN(_0761_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0914_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q ),
    .ZN(_0762_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0915_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q ),
    .ZN(_0763_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0916_ (.I(S2END[1]),
    .ZN(_0764_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0917_ (.I(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .ZN(_0765_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0918_ (.I(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .ZN(_0766_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0919_ (.I(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .ZN(_0767_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0920_ (.I(\Inst_LG_LUT4c_frame_config_dffesr.c_I0mux ),
    .ZN(_0768_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0921_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q ),
    .ZN(_0769_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0922_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q ),
    .ZN(_0770_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0923_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q ),
    .ZN(_0771_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0924_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q ),
    .ZN(_0772_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0925_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q ),
    .ZN(_0773_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0926_ (.I(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .ZN(_0774_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0927_ (.I(\Inst_LH_LUT4c_frame_config_dffesr.c_I0mux ),
    .ZN(_0775_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0928_ (.I(\Inst_LH_LUT4c_frame_config_dffesr.LUT_flop ),
    .ZN(_0776_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0929_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q ),
    .ZN(_0777_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0930_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q ),
    .ZN(_0778_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0931_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q ),
    .ZN(_0779_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0932_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q ),
    .ZN(_0780_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0933_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q ),
    .ZN(_0781_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0934_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q ),
    .ZN(_0782_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0935_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ),
    .ZN(_0783_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0936_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q ),
    .ZN(_0784_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0937_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q ),
    .ZN(_0785_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0938_ (.I(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q ),
    .ZN(_0786_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0939_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(E),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ),
    .Z(_0787_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0940_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q ),
    .A2(_0787_),
    .ZN(_0788_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0941_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ),
    .Z(_0789_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0942_ (.A1(_0715_),
    .A2(_0789_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit9.Q ),
    .ZN(_0790_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0943_ (.I0(N1END[2]),
    .I1(N2END[4]),
    .I2(N4END[0]),
    .I3(E2END[4]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ),
    .Z(_0791_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0944_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q ),
    .A2(_0791_),
    .ZN(_0792_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0945_ (.I0(E6END[0]),
    .I1(S2END[4]),
    .I2(W2END[4]),
    .I3(W6END[0]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ),
    .Z(_0793_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0946_ (.A1(_0715_),
    .A2(_0793_),
    .ZN(_0794_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _0947_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit9.Q ),
    .A2(_0792_),
    .A3(_0794_),
    .B1(_0788_),
    .B2(_0790_),
    .ZN(\Inst_LUT4AB_switch_matrix.E2BEG3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0948_ (.I0(E2MID[2]),
    .I1(S2MID[2]),
    .I2(W2MID[2]),
    .I3(\Inst_LUT4AB_switch_matrix.E2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit28.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit29.Q ),
    .Z(_0795_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0949_ (.I0(N2MID[3]),
    .I1(E2MID[3]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit28.Q ),
    .Z(_0796_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0950_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit28.Q ),
    .A2(W2MID[3]),
    .ZN(_0797_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _0951_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit28.Q ),
    .A2(_0716_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit29.Q ),
    .C(_0797_),
    .ZN(_0798_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0952_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit29.Q ),
    .A2(_0796_),
    .B(_0798_),
    .ZN(_0799_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0953_ (.I(_0799_),
    .ZN(_0800_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0954_ (.I0(A),
    .I1(D),
    .I2(C),
    .I3(E),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ),
    .Z(_0801_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0955_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q ),
    .A2(_0801_),
    .ZN(_0802_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0956_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_AB ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ),
    .Z(_0803_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0957_ (.A1(_0717_),
    .A2(_0803_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q ),
    .ZN(_0804_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0958_ (.I0(N1END[0]),
    .I1(N2END[2]),
    .I2(N4END[2]),
    .I3(E2END[2]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ),
    .Z(_0805_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0959_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q ),
    .A2(_0805_),
    .ZN(_0806_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0960_ (.I0(E6END[0]),
    .I1(S2END[2]),
    .I2(W2END[2]),
    .I3(WW4END[3]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ),
    .Z(_0807_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0961_ (.A1(_0717_),
    .A2(_0807_),
    .ZN(_0808_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _0962_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q ),
    .A2(_0806_),
    .A3(_0808_),
    .B1(_0802_),
    .B2(_0804_),
    .ZN(\Inst_LUT4AB_switch_matrix.E2BEG1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0963_ (.I0(EE4END[2]),
    .I1(S4END[2]),
    .I2(W2END[7]),
    .I3(\Inst_LUT4AB_switch_matrix.E2BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit28.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit29.Q ),
    .Z(_0809_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0964_ (.I0(NN4END[0]),
    .I1(S2END[2]),
    .I2(E2END[2]),
    .I3(W2END[2]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit29.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit28.Q ),
    .Z(_0810_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0965_ (.I0(_0795_),
    .I1(_0800_),
    .I2(_0810_),
    .I3(_0809_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit4.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit5.Q ),
    .Z(_0811_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0966_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(E),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q ),
    .Z(_0812_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0967_ (.A1(_0709_),
    .A2(_0812_),
    .ZN(_0813_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0968_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q ),
    .Z(_0814_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0969_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q ),
    .A2(_0814_),
    .B(_0710_),
    .ZN(_0815_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0970_ (.I0(E6END[0]),
    .I1(S2END[4]),
    .I2(W2END[4]),
    .I3(W6END[0]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q ),
    .Z(_0816_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0971_ (.I0(N2END[4]),
    .I1(E1END[2]),
    .I2(N4END[0]),
    .I3(E2END[4]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ),
    .Z(_0817_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0972_ (.A1(_0709_),
    .A2(_0817_),
    .ZN(_0818_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0973_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q ),
    .A2(_0816_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q ),
    .ZN(_0819_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0974_ (.A1(_0813_),
    .A2(_0815_),
    .B1(_0818_),
    .B2(_0819_),
    .ZN(\Inst_LUT4AB_switch_matrix.JN2BEG3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0975_ (.I0(N2MID[6]),
    .I1(S2MID[6]),
    .I2(W2MID[6]),
    .I3(\Inst_LUT4AB_switch_matrix.JN2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit27.Q ),
    .Z(_0820_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0976_ (.I0(N2MID[7]),
    .I1(E2MID[7]),
    .I2(S2MID[7]),
    .I3(W2MID[7]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit27.Q ),
    .Z(_0821_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0977_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_AD ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ),
    .Z(_0822_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0978_ (.I0(A),
    .I1(D),
    .I2(C),
    .I3(E),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ),
    .Z(_0823_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0979_ (.A1(_0713_),
    .A2(_0823_),
    .ZN(_0824_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0980_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q ),
    .A2(_0822_),
    .B(_0714_),
    .ZN(_0825_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0981_ (.I0(E6END[0]),
    .I1(S2END[2]),
    .I2(W2END[2]),
    .I3(W6END[0]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ),
    .Z(_0826_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0982_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q ),
    .A2(_0826_),
    .ZN(_0827_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0983_ (.I0(N2END[2]),
    .I1(E1END[0]),
    .I2(N4END[2]),
    .I3(E2END[2]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ),
    .Z(_0828_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0984_ (.A1(_0713_),
    .A2(_0828_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q ),
    .ZN(_0829_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0985_ (.A1(_0824_),
    .A2(_0825_),
    .B1(_0827_),
    .B2(_0829_),
    .ZN(\Inst_LUT4AB_switch_matrix.JN2BEG1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0986_ (.I0(NN4END[3]),
    .I1(WW4END[0]),
    .I2(S4END[3]),
    .I3(\Inst_LUT4AB_switch_matrix.JN2BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit26.Q ),
    .Z(_0830_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0987_ (.I0(N2END[6]),
    .I1(SS4END[3]),
    .I2(E2END[6]),
    .I3(W2END[6]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit26.Q ),
    .Z(_0831_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0988_ (.I(_0831_),
    .ZN(_0832_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0989_ (.I0(_0820_),
    .I1(_0821_),
    .I2(_0831_),
    .I3(_0830_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit3.Q ),
    .Z(_0833_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0990_ (.I0(_0833_),
    .I1(Ci),
    .S(\Inst_LA_LUT4c_frame_config_dffesr.c_I0mux ),
    .Z(_0834_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _0991_ (.I0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .I1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .S(_0834_),
    .Z(_0835_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0992_ (.A1(N4END[1]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q ),
    .ZN(_0836_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _0993_ (.A1(_0722_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q ),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit31.Q ),
    .C(_0836_),
    .ZN(_0837_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0994_ (.I0(A),
    .I1(D),
    .I2(C),
    .I3(E),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ),
    .Z(_0838_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0995_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ),
    .Z(_0839_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0996_ (.A1(_0723_),
    .A2(_0839_),
    .ZN(_0840_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0997_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q ),
    .A2(_0838_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q ),
    .ZN(_0841_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _0998_ (.I0(NN4END[2]),
    .I1(EE4END[2]),
    .I2(E1END[0]),
    .I3(E6END[0]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ),
    .Z(_0842_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0999_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q ),
    .A2(_0842_),
    .ZN(_0843_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1000_ (.I0(S4END[2]),
    .I1(SS4END[2]),
    .I2(W2END[2]),
    .I3(W6END[0]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ),
    .Z(_0844_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1001_ (.A1(_0723_),
    .A2(_0844_),
    .B(_0724_),
    .ZN(_0845_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1002_ (.A1(_0840_),
    .A2(_0841_),
    .B1(_0843_),
    .B2(_0845_),
    .ZN(\Inst_LUT4AB_switch_matrix.JS2BEG1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1003_ (.A1(_0840_),
    .A2(_0841_),
    .B1(_0843_),
    .B2(_0845_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q ),
    .ZN(_0846_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1004_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q ),
    .A2(W6END[1]),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit31.Q ),
    .ZN(_0847_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1005_ (.I(_0847_),
    .ZN(_0848_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1006_ (.I0(N4END[1]),
    .I1(E6END[1]),
    .I2(W6END[1]),
    .I3(\Inst_LUT4AB_switch_matrix.JS2BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit31.Q ),
    .Z(_0849_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1007_ (.A1(_0846_),
    .A2(_0848_),
    .B(_0721_),
    .C(_0837_),
    .ZN(_0850_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1008_ (.I0(N2END[4]),
    .I1(S2END[4]),
    .I2(EE4END[0]),
    .I3(W2END[4]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit30.Q ),
    .Z(_0851_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1009_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q ),
    .A2(_0851_),
    .ZN(_0852_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1010_ (.A1(_0725_),
    .A2(_0852_),
    .ZN(_0853_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1011_ (.I(_0853_),
    .ZN(_0854_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1012_ (.A1(_0850_),
    .A2(_0854_),
    .ZN(_0855_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1013_ (.A1(N2MID[4]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q ),
    .ZN(_0856_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1014_ (.A1(_0718_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q ),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q ),
    .C(_0856_),
    .ZN(_0857_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1015_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_AD ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ),
    .Z(_0858_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1016_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(E),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ),
    .Z(_0008_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1017_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q ),
    .A2(_0008_),
    .ZN(_0009_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1018_ (.A1(_0719_),
    .A2(_0858_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q ),
    .ZN(_0010_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1019_ (.I0(S2END[4]),
    .I1(W2END[4]),
    .I2(S4END[0]),
    .I3(WW4END[2]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ),
    .Z(_0011_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1020_ (.A1(_0719_),
    .A2(_0011_),
    .ZN(_0012_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1021_ (.I0(N2END[4]),
    .I1(E1END[2]),
    .I2(E2END[4]),
    .I3(E6END[0]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ),
    .Z(_0013_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1022_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q ),
    .A2(_0013_),
    .B(_0720_),
    .ZN(_0014_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1023_ (.A1(_0009_),
    .A2(_0010_),
    .B1(_0012_),
    .B2(_0014_),
    .ZN(\Inst_LUT4AB_switch_matrix.JS2BEG3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1024_ (.A1(_0009_),
    .A2(_0010_),
    .B1(_0012_),
    .B2(_0014_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q ),
    .ZN(_0015_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1025_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q ),
    .A2(W2MID[4]),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q ),
    .ZN(_0016_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1026_ (.I(_0016_),
    .ZN(_0017_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1027_ (.I0(N2MID[4]),
    .I1(E2MID[4]),
    .I2(W2MID[4]),
    .I3(\Inst_LUT4AB_switch_matrix.JS2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q ),
    .Z(_0018_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1028_ (.A1(_0015_),
    .A2(_0017_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q ),
    .C(_0857_),
    .ZN(_0019_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1029_ (.I0(N2MID[5]),
    .I1(E2MID[5]),
    .I2(S2MID[5]),
    .I3(W2MID[5]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit31.Q ),
    .Z(_0020_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1030_ (.A1(_0721_),
    .A2(_0020_),
    .B(_0725_),
    .ZN(_0021_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1031_ (.A1(_0019_),
    .A2(_0021_),
    .ZN(_0022_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1032_ (.A1(_0855_),
    .A2(_0022_),
    .ZN(_0023_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1033_ (.A1(_0850_),
    .A2(_0854_),
    .B1(_0019_),
    .B2(_0021_),
    .ZN(_0024_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1034_ (.I0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .I1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .S(_0834_),
    .Z(_0025_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1035_ (.I0(_0835_),
    .I1(_0025_),
    .S(_0811_),
    .Z(_0026_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1036_ (.I0(A),
    .I1(D),
    .I2(C),
    .I3(E),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ),
    .Z(_0027_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1037_ (.A1(_0728_),
    .A2(_0027_),
    .ZN(_0028_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1038_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ),
    .Z(_0029_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1039_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q ),
    .A2(_0029_),
    .B(_0729_),
    .ZN(_0030_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1040_ (.I0(N1END[0]),
    .I1(E2END[2]),
    .I2(N2END[2]),
    .I3(E6END[0]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ),
    .Z(_0031_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1041_ (.I0(S2END[2]),
    .I1(W2END[2]),
    .I2(S4END[2]),
    .I3(W6END[0]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ),
    .Z(_0032_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1042_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q ),
    .A2(_0032_),
    .ZN(_0033_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1043_ (.A1(_0728_),
    .A2(_0031_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q ),
    .ZN(_0034_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1044_ (.A1(_0028_),
    .A2(_0030_),
    .B1(_0033_),
    .B2(_0034_),
    .ZN(\Inst_LUT4AB_switch_matrix.JW2BEG1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1045_ (.I0(N4END[0]),
    .I1(E6END[0]),
    .I2(S4END[0]),
    .I3(\Inst_LUT4AB_switch_matrix.JW2BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit0.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit1.Q ),
    .Z(_0035_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1046_ (.I0(N2END[0]),
    .I1(S2END[0]),
    .I2(E2END[0]),
    .I3(WW4END[3]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit1.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit0.Q ),
    .Z(_0036_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1047_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(E),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ),
    .Z(_0037_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1048_ (.A1(_0726_),
    .A2(_0037_),
    .ZN(_0038_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1049_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_AB ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ),
    .Z(_0039_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1050_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q ),
    .A2(_0039_),
    .B(_0727_),
    .ZN(_0040_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1051_ (.I0(N1END[2]),
    .I1(E2END[4]),
    .I2(N2END[4]),
    .I3(E6END[0]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ),
    .Z(_0041_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1052_ (.I0(S2END[4]),
    .I1(W2END[4]),
    .I2(S4END[0]),
    .I3(WW4END[2]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ),
    .Z(_0042_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1053_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q ),
    .A2(_0042_),
    .ZN(_0043_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1054_ (.A1(_0726_),
    .A2(_0041_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q ),
    .ZN(_0044_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1055_ (.A1(_0038_),
    .A2(_0040_),
    .B1(_0043_),
    .B2(_0044_),
    .ZN(\Inst_LUT4AB_switch_matrix.JW2BEG3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1056_ (.I0(N2MID[0]),
    .I1(E2MID[0]),
    .I2(S2MID[0]),
    .I3(\Inst_LUT4AB_switch_matrix.JW2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit1.Q ),
    .Z(_0045_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1057_ (.I0(N2MID[1]),
    .I1(E2MID[1]),
    .I2(S2MID[1]),
    .I3(W2MID[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit1.Q ),
    .Z(_0046_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1058_ (.I(_0046_),
    .ZN(_0047_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1059_ (.I0(_0045_),
    .I1(_0046_),
    .I2(_0036_),
    .I3(_0035_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit8.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q ),
    .Z(_0048_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1060_ (.I0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .I1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .S(_0834_),
    .Z(_0049_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1061_ (.I0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .I1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .S(_0834_),
    .Z(_0050_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1062_ (.I0(_0049_),
    .I1(_0050_),
    .S(_0811_),
    .Z(_0051_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1063_ (.I0(_0026_),
    .I1(_0051_),
    .S(_0023_),
    .Z(_0052_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1064_ (.A1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .A2(_0834_),
    .Z(_0053_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1065_ (.I0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .I1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .S(_0834_),
    .Z(_0054_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1066_ (.A1(_0730_),
    .A2(_0834_),
    .B(_0811_),
    .ZN(_0055_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1067_ (.A1(_0811_),
    .A2(_0054_),
    .B1(_0055_),
    .B2(_0053_),
    .ZN(_0056_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1068_ (.A1(_0023_),
    .A2(_0056_),
    .ZN(_0057_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1069_ (.I0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .I1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .S(_0834_),
    .Z(_0058_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1070_ (.I0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .I1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .S(_0834_),
    .Z(_0059_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1071_ (.I0(_0059_),
    .I1(_0058_),
    .S(_0811_),
    .Z(_0060_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1072_ (.A1(_0023_),
    .A2(_0060_),
    .ZN(_0061_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1073_ (.A1(_0048_),
    .A2(_0061_),
    .ZN(_0062_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1074_ (.A1(_0048_),
    .A2(_0052_),
    .B1(_0057_),
    .B2(_0062_),
    .ZN(_0063_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1075_ (.A1(\Inst_LA_LUT4c_frame_config_dffesr.LUT_flop ),
    .A2(\Inst_LA_LUT4c_frame_config_dffesr.c_out_mux ),
    .ZN(_0064_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1076_ (.A1(\Inst_LA_LUT4c_frame_config_dffesr.c_out_mux ),
    .A2(_0063_),
    .B(_0064_),
    .ZN(A),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1077_ (.A1(_0736_),
    .A2(_0045_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q ),
    .ZN(_0065_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1078_ (.A1(_0736_),
    .A2(_0047_),
    .B(_0065_),
    .ZN(_0066_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1079_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit18.Q ),
    .A2(_0035_),
    .ZN(_0067_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1080_ (.A1(_0736_),
    .A2(_0036_),
    .ZN(_0068_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1081_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q ),
    .A2(_0067_),
    .A3(_0068_),
    .ZN(_0069_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1082_ (.A1(_0066_),
    .A2(_0069_),
    .ZN(_0070_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1083_ (.A1(_0066_),
    .A2(_0069_),
    .Z(_0071_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1084_ (.I0(_0018_),
    .I1(_0020_),
    .I2(_0851_),
    .I3(_0849_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit16.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit17.Q ),
    .Z(_0072_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1085_ (.I(_0072_),
    .ZN(_0073_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1086_ (.I0(_0795_),
    .I1(_0800_),
    .I2(_0810_),
    .I3(_0809_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit15.Q ),
    .Z(_0074_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1087_ (.I(_0074_),
    .ZN(_0075_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1088_ (.A1(_0073_),
    .A2(_0074_),
    .ZN(_0076_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1089_ (.A1(_0072_),
    .A2(_0075_),
    .ZN(_0077_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1090_ (.A1(_0072_),
    .A2(_0074_),
    .ZN(_0078_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1091_ (.A1(_0073_),
    .A2(_0075_),
    .ZN(_0079_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1092_ (.A1(_0072_),
    .A2(_0074_),
    .ZN(_0080_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1093_ (.A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .A2(_0077_),
    .B1(_0079_),
    .B2(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .ZN(_0081_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1094_ (.A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .A2(_0076_),
    .B1(_0080_),
    .B2(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .C(_0071_),
    .ZN(_0082_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1095_ (.I0(_0820_),
    .I1(_0821_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q ),
    .Z(_0083_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1096_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q ),
    .A2(_0832_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit13.Q ),
    .ZN(_0084_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1097_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q ),
    .A2(_0830_),
    .B(_0084_),
    .ZN(_0085_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1098_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit13.Q ),
    .A2(_0083_),
    .B(_0735_),
    .ZN(_0086_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1099_ (.A1(_0811_),
    .A2(_0024_),
    .ZN(_0087_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1100_ (.A1(_0811_),
    .A2(_0024_),
    .B(Ci),
    .ZN(_0088_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1101_ (.A1(_0735_),
    .A2(_0087_),
    .A3(_0088_),
    .B1(_0085_),
    .B2(_0086_),
    .ZN(_0089_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _1102_ (.A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .A2(_0076_),
    .B1(_0077_),
    .B2(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .C1(_0080_),
    .C2(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .ZN(_0090_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1103_ (.I(_0090_),
    .ZN(_0091_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1104_ (.A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .A2(_0079_),
    .B(_0091_),
    .C(_0070_),
    .ZN(_0092_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1105_ (.A1(_0081_),
    .A2(_0082_),
    .B(_0092_),
    .ZN(_0093_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1106_ (.A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .A2(_0076_),
    .B1(_0077_),
    .B2(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .ZN(_0094_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1107_ (.A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .A2(_0079_),
    .B1(_0080_),
    .B2(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .C(_0071_),
    .ZN(_0095_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _1108_ (.A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .A2(_0076_),
    .B1(_0077_),
    .B2(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .C1(_0079_),
    .C2(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .ZN(_0096_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1109_ (.I(_0096_),
    .ZN(_0097_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1110_ (.A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .A2(_0080_),
    .B(_0097_),
    .C(_0070_),
    .ZN(_0098_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1111_ (.A1(_0094_),
    .A2(_0095_),
    .B(_0098_),
    .ZN(_0099_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1112_ (.I0(_0093_),
    .I1(_0099_),
    .S(_0089_),
    .Z(_0100_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1113_ (.I0(_0100_),
    .I1(\Inst_LB_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(\Inst_LB_LUT4c_frame_config_dffesr.c_out_mux ),
    .Z(B),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1114_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ),
    .Z(_0101_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1115_ (.A1(_0742_),
    .A2(_0101_),
    .ZN(_0102_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1116_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ),
    .Z(_0103_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1117_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q ),
    .A2(_0103_),
    .B(_0743_),
    .ZN(_0104_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1118_ (.I0(S1END[1]),
    .I1(S2END[5]),
    .I2(S1END[3]),
    .I3(W1END[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ),
    .Z(_0105_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1119_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q ),
    .A2(_0105_),
    .ZN(_0106_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1120_ (.I0(N1END[1]),
    .I1(N2END[5]),
    .I2(E1END[1]),
    .I3(E2END[5]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ),
    .Z(_0107_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1121_ (.A1(_0742_),
    .A2(_0107_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q ),
    .ZN(_0108_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1122_ (.A1(_0102_),
    .A2(_0104_),
    .B1(_0106_),
    .B2(_0108_),
    .ZN(\Inst_LUT4AB_switch_matrix.E2BEG4 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1123_ (.I0(N2MID[2]),
    .I1(W2MID[2]),
    .I2(E2MID[2]),
    .I3(\Inst_LUT4AB_switch_matrix.E2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit5.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit4.Q ),
    .Z(_0109_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1124_ (.I0(N2MID[3]),
    .I1(E2MID[3]),
    .I2(S2MID[3]),
    .I3(W2MID[3]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit4.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit5.Q ),
    .Z(_0110_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1125_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_AD ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ),
    .Z(_0111_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1126_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q ),
    .A2(_0111_),
    .ZN(_0112_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1127_ (.I0(A),
    .I1(B),
    .I2(D),
    .I3(E),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ),
    .Z(_0113_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1128_ (.A1(_0744_),
    .A2(_0113_),
    .B(_0745_),
    .ZN(_0114_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1129_ (.I0(N1END[1]),
    .I1(N4END[3]),
    .I2(N2END[3]),
    .I3(E2END[3]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ),
    .Z(_0115_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1130_ (.I0(E6END[1]),
    .I1(S2END[3]),
    .I2(W2END[3]),
    .I3(W6END[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ),
    .Z(_0116_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1131_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q ),
    .A2(_0116_),
    .ZN(_0117_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1132_ (.A1(_0744_),
    .A2(_0115_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q ),
    .ZN(_0118_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1133_ (.A1(_0112_),
    .A2(_0114_),
    .B1(_0117_),
    .B2(_0118_),
    .ZN(\Inst_LUT4AB_switch_matrix.E2BEG2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1134_ (.I(\Inst_LUT4AB_switch_matrix.E2BEG2 ),
    .ZN(_0119_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1135_ (.I0(N4END[2]),
    .I1(E2END[2]),
    .I2(W2END[7]),
    .I3(\Inst_LUT4AB_switch_matrix.E2BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit4.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit5.Q ),
    .Z(_0120_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1136_ (.I0(N2END[2]),
    .I1(E2END[2]),
    .I2(S2END[2]),
    .I3(WW4END[2]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit4.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit5.Q ),
    .Z(_0121_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1137_ (.I0(_0109_),
    .I1(_0110_),
    .I2(_0121_),
    .I3(_0120_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit3.Q ),
    .Z(_0122_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1138_ (.I(_0122_),
    .ZN(_0123_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1139_ (.I0(A),
    .I1(B),
    .I2(D),
    .I3(E),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ),
    .Z(_0124_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1140_ (.A1(_0748_),
    .A2(_0124_),
    .ZN(_0125_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1141_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_AB ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ),
    .Z(_0126_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1142_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q ),
    .A2(_0126_),
    .B(_0749_),
    .ZN(_0127_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1143_ (.I0(NN4END[3]),
    .I1(E1END[1]),
    .I2(E2END[3]),
    .I3(E6END[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ),
    .Z(_0128_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1144_ (.A1(_0748_),
    .A2(_0128_),
    .ZN(_0129_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1145_ (.I0(S2END[3]),
    .I1(W2END[3]),
    .I2(S4END[3]),
    .I3(W6END[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ),
    .Z(_0130_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1146_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q ),
    .A2(_0130_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit5.Q ),
    .ZN(_0131_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1147_ (.A1(_0125_),
    .A2(_0127_),
    .B1(_0129_),
    .B2(_0131_),
    .ZN(\Inst_LUT4AB_switch_matrix.JS2BEG2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1148_ (.I0(NN4END[1]),
    .I1(EE4END[1]),
    .I2(S4END[1]),
    .I3(\Inst_LUT4AB_switch_matrix.JS2BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit7.Q ),
    .Z(_0132_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1149_ (.I0(N2END[4]),
    .I1(E2END[4]),
    .I2(SS4END[2]),
    .I3(W2END[4]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit7.Q ),
    .Z(_0133_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1150_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ),
    .Z(_0134_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1151_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ),
    .Z(_0135_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1152_ (.A1(_0746_),
    .A2(_0135_),
    .ZN(_0136_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1153_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q ),
    .A2(_0134_),
    .B(_0747_),
    .ZN(_0137_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1154_ (.I0(N1END[1]),
    .I1(N2END[5]),
    .I2(E1END[1]),
    .I3(E2END[5]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ),
    .Z(_0138_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1155_ (.I0(S1END[1]),
    .I1(S2END[5]),
    .I2(W1END[1]),
    .I3(W1END[3]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ),
    .Z(_0139_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1156_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q ),
    .A2(_0139_),
    .ZN(_0140_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1157_ (.A1(_0746_),
    .A2(_0138_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit13.Q ),
    .ZN(_0141_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1158_ (.A1(_0136_),
    .A2(_0137_),
    .B1(_0140_),
    .B2(_0141_),
    .ZN(\Inst_LUT4AB_switch_matrix.JS2BEG4 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1159_ (.I0(N2MID[4]),
    .I1(E2MID[4]),
    .I2(S2MID[4]),
    .I3(\Inst_LUT4AB_switch_matrix.JS2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q ),
    .Z(_0142_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1160_ (.I0(N2MID[5]),
    .I1(E2MID[5]),
    .I2(S2MID[5]),
    .I3(W2MID[5]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit7.Q ),
    .Z(_0143_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1161_ (.I0(_0142_),
    .I1(_0143_),
    .I2(_0133_),
    .I3(_0132_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit4.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit5.Q ),
    .Z(_0144_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1162_ (.A1(_0122_),
    .A2(_0144_),
    .ZN(_0145_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1163_ (.A1(_0122_),
    .A2(_0144_),
    .Z(_0146_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1164_ (.A1(_0122_),
    .A2(_0144_),
    .ZN(_0147_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1165_ (.I0(_0109_),
    .I1(_0110_),
    .I2(_0121_),
    .I3(_0120_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit24.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit25.Q ),
    .Z(_0148_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1166_ (.I(_0148_),
    .ZN(_0149_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1167_ (.I0(_0142_),
    .I1(_0143_),
    .I2(_0133_),
    .I3(_0132_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit27.Q ),
    .Z(_0150_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1168_ (.A1(_0148_),
    .A2(_0150_),
    .Z(_0151_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1169_ (.A1(_0148_),
    .A2(_0150_),
    .Z(_0152_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1170_ (.I(_0152_),
    .ZN(_0153_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1171_ (.A1(_0078_),
    .A2(_0087_),
    .A3(_0088_),
    .B(_0080_),
    .ZN(_0154_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1172_ (.A1(_0151_),
    .A2(_0154_),
    .B(_0152_),
    .ZN(_0155_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1173_ (.A1(_0122_),
    .A2(_0144_),
    .B1(_0151_),
    .B2(_0154_),
    .C(_0152_),
    .ZN(_0156_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1174_ (.I0(N4END[3]),
    .I1(W2END[3]),
    .I2(E2END[3]),
    .I3(\Inst_LUT4AB_switch_matrix.JN2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit10.Q ),
    .Z(_0157_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1175_ (.I0(N2END[7]),
    .I1(S2END[7]),
    .I2(EE4END[2]),
    .I3(W2END[7]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit10.Q ),
    .Z(_0158_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1176_ (.I0(E),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_AD ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ),
    .Z(_0159_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1177_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q ),
    .A2(_0159_),
    .ZN(_0160_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1178_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ),
    .Z(_0161_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1179_ (.A1(_0753_),
    .A2(_0161_),
    .B(_0754_),
    .ZN(_0162_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1180_ (.I0(N1END[2]),
    .I1(N2END[6]),
    .I2(E1END[2]),
    .I3(E2END[6]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ),
    .Z(_0163_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1181_ (.I0(S1END[2]),
    .I1(W1END[0]),
    .I2(S2END[6]),
    .I3(W1END[2]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ),
    .Z(_0164_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1182_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q ),
    .A2(_0164_),
    .ZN(_0165_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1183_ (.A1(_0753_),
    .A2(_0163_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q ),
    .ZN(_0166_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1184_ (.A1(_0160_),
    .A2(_0162_),
    .B1(_0165_),
    .B2(_0166_),
    .ZN(\Inst_LUT4AB_switch_matrix.JN2BEG5 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1185_ (.I0(N2MID[6]),
    .I1(W2MID[6]),
    .I2(E2MID[6]),
    .I3(\Inst_LUT4AB_switch_matrix.JN2BEG5 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q ),
    .Z(_0167_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1186_ (.A1(W2MID[7]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q ),
    .ZN(_0168_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1187_ (.A1(_0712_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q ),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit11.Q ),
    .C(_0168_),
    .ZN(_0169_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1188_ (.A1(E2MID[7]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q ),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit11.Q ),
    .ZN(_0170_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1189_ (.A1(_0711_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q ),
    .B(_0170_),
    .ZN(_0171_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1190_ (.A1(_0169_),
    .A2(_0171_),
    .ZN(_0172_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1191_ (.A1(_0169_),
    .A2(_0171_),
    .Z(_0173_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1192_ (.I0(_0167_),
    .I1(_0173_),
    .I2(_0158_),
    .I3(_0157_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q ),
    .Z(_0174_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1193_ (.A1(_0755_),
    .A2(_0174_),
    .ZN(_0175_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1194_ (.A1(_0755_),
    .A2(_0145_),
    .A3(_0156_),
    .B(_0175_),
    .ZN(_0176_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1195_ (.I0(NN4END[2]),
    .I1(S4END[2]),
    .I2(E2END[2]),
    .I3(\Inst_LUT4AB_switch_matrix.E2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit13.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q ),
    .Z(_0177_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1196_ (.I0(N2END[3]),
    .I1(S2END[3]),
    .I2(E2END[3]),
    .I3(WW4END[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit13.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q ),
    .Z(_0178_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1197_ (.I0(E),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_AB ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ),
    .Z(_0179_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1198_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ),
    .Z(_0180_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1199_ (.A1(_0758_),
    .A2(_0180_),
    .ZN(_0181_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1200_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q ),
    .A2(_0179_),
    .B(_0759_),
    .ZN(_0182_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1201_ (.I0(S1END[0]),
    .I1(S1END[2]),
    .I2(S2END[6]),
    .I3(W1END[2]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ),
    .Z(_0183_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1202_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q ),
    .A2(_0183_),
    .ZN(_0184_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1203_ (.I0(N1END[2]),
    .I1(N2END[6]),
    .I2(E1END[2]),
    .I3(E2END[6]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ),
    .Z(_0185_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1204_ (.A1(_0758_),
    .A2(_0185_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q ),
    .ZN(_0186_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1205_ (.A1(_0181_),
    .A2(_0182_),
    .B1(_0184_),
    .B2(_0186_),
    .ZN(\Inst_LUT4AB_switch_matrix.E2BEG5 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1206_ (.I0(N2MID[2]),
    .I1(S2MID[2]),
    .I2(E2MID[2]),
    .I3(\Inst_LUT4AB_switch_matrix.E2BEG5 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit13.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q ),
    .Z(_0187_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1207_ (.A1(W2MID[3]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit12.Q ),
    .ZN(_0188_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1208_ (.A1(_0716_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit12.Q ),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit13.Q ),
    .C(_0188_),
    .ZN(_0189_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1209_ (.I0(N2MID[3]),
    .I1(E2MID[3]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit12.Q ),
    .Z(_0190_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1210_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit13.Q ),
    .A2(_0190_),
    .B(_0189_),
    .ZN(_0191_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1211_ (.I(_0191_),
    .ZN(_0192_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1212_ (.I0(_0187_),
    .I1(_0192_),
    .I2(_0178_),
    .I3(_0177_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit12.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit13.Q ),
    .Z(_0193_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1213_ (.I0(N4END[1]),
    .I1(SS4END[1]),
    .I2(W2END[4]),
    .I3(\Inst_LUT4AB_switch_matrix.JS2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit15.Q ),
    .Z(_0194_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1214_ (.I0(N2END[5]),
    .I1(E2END[5]),
    .I2(SS4END[1]),
    .I3(W2END[5]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit15.Q ),
    .Z(_0195_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1215_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ),
    .Z(_0196_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1216_ (.A1(_0760_),
    .A2(_0196_),
    .ZN(_0197_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1217_ (.I0(E),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ),
    .Z(_0198_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1218_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q ),
    .A2(_0198_),
    .B(_0761_),
    .ZN(_0199_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1219_ (.I0(N1END[2]),
    .I1(N2END[6]),
    .I2(E1END[2]),
    .I3(E2END[6]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ),
    .Z(_0200_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1220_ (.I0(S1END[2]),
    .I1(W1END[0]),
    .I2(S2END[6]),
    .I3(W1END[2]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ),
    .Z(_0201_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1221_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q ),
    .A2(_0201_),
    .ZN(_0202_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1222_ (.A1(_0760_),
    .A2(_0200_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q ),
    .ZN(_0203_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1223_ (.A1(_0197_),
    .A2(_0199_),
    .B1(_0202_),
    .B2(_0203_),
    .ZN(\Inst_LUT4AB_switch_matrix.JS2BEG5 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1224_ (.I0(N2MID[4]),
    .I1(W2MID[4]),
    .I2(S2MID[4]),
    .I3(\Inst_LUT4AB_switch_matrix.JS2BEG5 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit15.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit14.Q ),
    .Z(_0204_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1225_ (.I0(N2MID[5]),
    .I1(E2MID[5]),
    .I2(S2MID[5]),
    .I3(W2MID[5]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit15.Q ),
    .Z(_0205_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1226_ (.I0(_0204_),
    .I1(_0205_),
    .I2(_0195_),
    .I3(_0194_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q ),
    .Z(_0206_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1227_ (.I(_0206_),
    .ZN(_0207_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1228_ (.A1(_0193_),
    .A2(_0206_),
    .ZN(_0208_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1229_ (.A1(_0193_),
    .A2(_0207_),
    .ZN(_0209_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1230_ (.A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .A2(_0193_),
    .A3(_0207_),
    .ZN(_0210_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1231_ (.A1(_0193_),
    .A2(_0206_),
    .ZN(_0211_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1232_ (.A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .A2(_0209_),
    .B1(_0211_),
    .B2(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .ZN(_0212_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1233_ (.A1(_0756_),
    .A2(_0208_),
    .B(_0210_),
    .C(_0212_),
    .ZN(_0213_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1234_ (.I0(EE4END[3]),
    .I1(WW4END[1]),
    .I2(S4END[0]),
    .I3(\Inst_LUT4AB_switch_matrix.JW2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit17.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit16.Q ),
    .Z(_0214_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1235_ (.I0(NN4END[2]),
    .I1(E2END[1]),
    .I2(S2END[1]),
    .I3(W2END[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit16.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit17.Q ),
    .Z(_0215_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1236_ (.I(_0215_),
    .ZN(_0216_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1237_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ),
    .Z(_0217_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1238_ (.I0(E),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ),
    .Z(_0218_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1239_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q ),
    .A2(_0218_),
    .ZN(_0219_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1240_ (.A1(_0762_),
    .A2(_0217_),
    .B(_0763_),
    .ZN(_0220_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1241_ (.I0(N1END[2]),
    .I1(N2END[6]),
    .I2(E1END[2]),
    .I3(E2END[6]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ),
    .Z(_0221_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1242_ (.I0(S1END[0]),
    .I1(S1END[2]),
    .I2(S2END[6]),
    .I3(W1END[2]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ),
    .Z(_0222_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1243_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q ),
    .A2(_0222_),
    .ZN(_0223_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1244_ (.A1(_0762_),
    .A2(_0221_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q ),
    .ZN(_0224_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1245_ (.A1(_0219_),
    .A2(_0220_),
    .B1(_0223_),
    .B2(_0224_),
    .ZN(\Inst_LUT4AB_switch_matrix.JW2BEG5 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1246_ (.I0(E2MID[0]),
    .I1(S2MID[0]),
    .I2(W2MID[0]),
    .I3(\Inst_LUT4AB_switch_matrix.JW2BEG5 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit16.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit17.Q ),
    .Z(_0225_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1247_ (.I0(N2MID[1]),
    .I1(E2MID[1]),
    .I2(S2MID[1]),
    .I3(W2MID[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit17.Q ),
    .Z(_0226_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1248_ (.I(_0226_),
    .ZN(_0227_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1249_ (.I0(_0225_),
    .I1(_0226_),
    .I2(_0215_),
    .I3(_0214_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q ),
    .Z(_0228_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1250_ (.A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .A2(_0193_),
    .ZN(_0229_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1251_ (.A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .A2(_0209_),
    .B1(_0211_),
    .B2(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .ZN(_0230_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1252_ (.A1(_0757_),
    .A2(_0208_),
    .B1(_0229_),
    .B2(_0206_),
    .C(_0230_),
    .ZN(_0231_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1253_ (.I0(_0231_),
    .I1(_0213_),
    .S(_0176_),
    .Z(_0232_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1254_ (.I0(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .I1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .I2(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .I3(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .S0(_0193_),
    .S1(_0206_),
    .Z(_0233_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1255_ (.A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .A2(_0193_),
    .A3(_0207_),
    .Z(_0234_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1256_ (.A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .A2(_0209_),
    .B1(_0211_),
    .B2(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .C(_0234_),
    .ZN(_0235_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1257_ (.A1(_0765_),
    .A2(_0208_),
    .B(_0235_),
    .ZN(_0236_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1258_ (.I0(_0236_),
    .I1(_0233_),
    .S(_0176_),
    .Z(_0237_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1259_ (.I0(_0232_),
    .I1(_0237_),
    .S(_0228_),
    .Z(_0238_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1260_ (.I0(_0238_),
    .I1(\Inst_LE_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(\Inst_LE_LUT4c_frame_config_dffesr.c_out_mux ),
    .Z(E),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1261_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ),
    .Z(_0239_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1262_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_AB ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ),
    .Z(_0240_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1263_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q ),
    .A2(_0240_),
    .ZN(_0241_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1264_ (.A1(_0737_),
    .A2(_0239_),
    .B(_0738_),
    .ZN(_0242_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1265_ (.I0(S1END[1]),
    .I1(S2END[5]),
    .I2(W1END[1]),
    .I3(W1END[3]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ),
    .Z(_0243_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1266_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q ),
    .A2(_0243_),
    .ZN(_0244_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1267_ (.I0(N1END[1]),
    .I1(N2END[5]),
    .I2(E1END[1]),
    .I3(E2END[5]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ),
    .Z(_0245_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1268_ (.A1(_0737_),
    .A2(_0245_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q ),
    .ZN(_0246_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1269_ (.A1(_0241_),
    .A2(_0242_),
    .B1(_0244_),
    .B2(_0246_),
    .ZN(\Inst_LUT4AB_switch_matrix.JN2BEG4 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1270_ (.I0(E2MID[6]),
    .I1(S2MID[6]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit2.Q ),
    .Z(_0247_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1271_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit2.Q ),
    .A2(\Inst_LUT4AB_switch_matrix.JN2BEG4 ),
    .ZN(_0248_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1272_ (.A1(_0708_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit2.Q ),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit3.Q ),
    .C(_0248_),
    .ZN(_0249_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1273_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit3.Q ),
    .A2(_0247_),
    .B(_0249_),
    .ZN(_0250_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1274_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q ),
    .A2(_0250_),
    .ZN(_0251_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1275_ (.I0(N2MID[7]),
    .I1(E2MID[7]),
    .I2(S2MID[7]),
    .I3(W2MID[7]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit3.Q ),
    .Z(_0252_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1276_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q ),
    .A2(_0252_),
    .B(_0251_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q ),
    .ZN(_0253_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1277_ (.I0(A),
    .I1(B),
    .I2(D),
    .I3(E),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ),
    .Z(_0254_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1278_ (.A1(_0740_),
    .A2(_0254_),
    .ZN(_0255_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1279_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ),
    .Z(_0256_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1280_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q ),
    .A2(_0256_),
    .B(_0741_),
    .ZN(_0257_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1281_ (.I0(N2END[3]),
    .I1(N4END[3]),
    .I2(E1END[1]),
    .I3(E2END[3]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ),
    .Z(_0258_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1282_ (.I0(E6END[1]),
    .I1(S2END[3]),
    .I2(W2END[3]),
    .I3(WW4END[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ),
    .Z(_0259_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1283_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q ),
    .A2(_0259_),
    .ZN(_0260_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1284_ (.A1(_0740_),
    .A2(_0258_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q ),
    .ZN(_0261_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1285_ (.A1(_0255_),
    .A2(_0257_),
    .B1(_0260_),
    .B2(_0261_),
    .ZN(\Inst_LUT4AB_switch_matrix.JN2BEG2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1286_ (.I0(E2END[3]),
    .I1(WW4END[2]),
    .I2(SS4END[3]),
    .I3(\Inst_LUT4AB_switch_matrix.JN2BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit3.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q ),
    .Z(_0262_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1287_ (.A1(W2END[6]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit2.Q ),
    .ZN(_0263_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1288_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit2.Q ),
    .A2(_0739_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit3.Q ),
    .C(_0263_),
    .ZN(_0264_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1289_ (.I0(NN4END[3]),
    .I1(E2END[6]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit2.Q ),
    .Z(_0265_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1290_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit3.Q ),
    .A2(_0265_),
    .B(_0264_),
    .ZN(_0266_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1291_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q ),
    .A2(_0266_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q ),
    .ZN(_0267_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1292_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q ),
    .A2(_0262_),
    .B(_0267_),
    .ZN(_0268_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1293_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.c_I0mux ),
    .A2(_0253_),
    .A3(_0268_),
    .ZN(_0269_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1294_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.c_I0mux ),
    .A2(_0154_),
    .Z(_0270_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1295_ (.A1(_0269_),
    .A2(_0270_),
    .ZN(_0271_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1296_ (.A1(_0149_),
    .A2(_0150_),
    .ZN(_0272_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1297_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .A2(_0151_),
    .B1(_0272_),
    .B2(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .ZN(_0273_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1298_ (.A1(_0149_),
    .A2(_0150_),
    .Z(_0274_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1299_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .A2(_0153_),
    .B1(_0274_),
    .B2(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .ZN(_0275_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1300_ (.A1(_0273_),
    .A2(_0275_),
    .ZN(_0276_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1301_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .A2(_0151_),
    .B1(_0274_),
    .B2(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .ZN(_0277_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1302_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .A2(_0153_),
    .B1(_0272_),
    .B2(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .ZN(_0278_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1303_ (.A1(_0277_),
    .A2(_0278_),
    .B(_0271_),
    .ZN(_0279_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1304_ (.I0(A),
    .I1(B),
    .I2(D),
    .I3(E),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ),
    .Z(_0280_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1305_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ),
    .Z(_0281_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1306_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q ),
    .A2(_0281_),
    .ZN(_0282_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1307_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q ),
    .A2(_0282_),
    .ZN(_0283_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1308_ (.A1(_0752_),
    .A2(_0280_),
    .B(_0283_),
    .ZN(_0284_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1309_ (.I0(N1END[1]),
    .I1(N2END[3]),
    .I2(EE4END[3]),
    .I3(E6END[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ),
    .Z(_0285_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1310_ (.I0(S4END[3]),
    .I1(W2END[3]),
    .I2(SS4END[3]),
    .I3(W6END[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ),
    .Z(_0286_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1311_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q ),
    .A2(_0286_),
    .Z(_0287_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1312_ (.A1(_0752_),
    .A2(_0285_),
    .B(_0287_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q ),
    .ZN(_0288_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1313_ (.A1(_0284_),
    .A2(_0288_),
    .ZN(\Inst_LUT4AB_switch_matrix.JW2BEG2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1314_ (.I0(N4END[0]),
    .I1(W6END[0]),
    .I2(SS4END[0]),
    .I3(\Inst_LUT4AB_switch_matrix.JW2BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit9.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q ),
    .Z(_0289_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1315_ (.I0(N2END[0]),
    .I1(S2END[0]),
    .I2(EE4END[1]),
    .I3(W2END[0]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit9.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q ),
    .Z(_0290_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1316_ (.I(_0290_),
    .ZN(_0291_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1317_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ),
    .Z(_0292_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1318_ (.A1(_0750_),
    .A2(_0292_),
    .ZN(_0293_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1319_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_AD ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ),
    .Z(_0294_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1320_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q ),
    .A2(_0294_),
    .B(_0751_),
    .ZN(_0295_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1321_ (.I0(N1END[1]),
    .I1(N2END[5]),
    .I2(E1END[1]),
    .I3(E2END[5]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ),
    .Z(_0296_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1322_ (.I0(S1END[1]),
    .I1(S2END[5]),
    .I2(S1END[3]),
    .I3(W1END[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ),
    .Z(_0297_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1323_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q ),
    .A2(_0297_),
    .ZN(_0298_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1324_ (.A1(_0750_),
    .A2(_0296_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q ),
    .ZN(_0299_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1325_ (.A1(_0293_),
    .A2(_0295_),
    .B1(_0298_),
    .B2(_0299_),
    .ZN(\Inst_LUT4AB_switch_matrix.JW2BEG4 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1326_ (.I0(N2MID[0]),
    .I1(S2MID[0]),
    .I2(W2MID[0]),
    .I3(\Inst_LUT4AB_switch_matrix.JW2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit9.Q ),
    .Z(_0300_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1327_ (.I0(N2MID[1]),
    .I1(E2MID[1]),
    .I2(S2MID[1]),
    .I3(W2MID[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit8.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit9.Q ),
    .Z(_0301_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1328_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q ),
    .A2(_0289_),
    .ZN(_0302_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1329_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q ),
    .A2(_0291_),
    .B(_0302_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q ),
    .ZN(_0303_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1330_ (.I0(_0300_),
    .I1(_0301_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q ),
    .Z(_0304_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1331_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q ),
    .A2(_0304_),
    .B(_0303_),
    .ZN(_0305_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1332_ (.I(_0305_),
    .ZN(_0306_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1333_ (.A1(_0271_),
    .A2(_0276_),
    .B(_0279_),
    .C(_0306_),
    .ZN(_0307_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1334_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .A2(_0151_),
    .B1(_0274_),
    .B2(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .ZN(_0308_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1335_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .A2(_0153_),
    .B1(_0272_),
    .B2(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .ZN(_0309_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1336_ (.A1(_0308_),
    .A2(_0309_),
    .ZN(_0310_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1337_ (.A1(_0271_),
    .A2(_0310_),
    .ZN(_0311_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1338_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .A2(_0153_),
    .B1(_0274_),
    .B2(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .ZN(_0312_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1339_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .A2(_0151_),
    .B1(_0272_),
    .B2(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .ZN(_0313_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1340_ (.A1(_0312_),
    .A2(_0313_),
    .ZN(_0314_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1341_ (.A1(_0269_),
    .A2(_0270_),
    .A3(_0314_),
    .B(_0305_),
    .ZN(_0315_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1342_ (.A1(_0311_),
    .A2(_0315_),
    .B(_0307_),
    .ZN(_0316_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1343_ (.I0(_0316_),
    .I1(\Inst_LC_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(\Inst_LC_LUT4c_frame_config_dffesr.c_out_mux ),
    .Z(C),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1344_ (.A1(_0145_),
    .A2(_0156_),
    .A3(_0208_),
    .B(_0211_),
    .ZN(_0317_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1345_ (.I0(_0167_),
    .I1(_0173_),
    .I2(_0158_),
    .I3(_0157_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit20.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q ),
    .Z(_0318_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1346_ (.I0(_0318_),
    .I1(_0317_),
    .S(\Inst_LF_LUT4c_frame_config_dffesr.c_I0mux ),
    .Z(_0319_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1347_ (.I0(_0204_),
    .I1(_0205_),
    .I2(_0195_),
    .I3(_0194_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit24.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q ),
    .Z(_0320_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1348_ (.I(_0320_),
    .ZN(_0321_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1349_ (.I0(_0187_),
    .I1(_0192_),
    .I2(_0178_),
    .I3(_0177_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit23.Q ),
    .Z(_0322_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1350_ (.A1(_0320_),
    .A2(_0322_),
    .Z(_0323_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1351_ (.A1(_0320_),
    .A2(_0322_),
    .ZN(_0324_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1352_ (.I(_0324_),
    .ZN(_0325_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1353_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .A2(_0323_),
    .B1(_0324_),
    .B2(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .ZN(_0326_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1354_ (.A1(_0321_),
    .A2(_0322_),
    .ZN(_0327_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1355_ (.A1(_0321_),
    .A2(_0322_),
    .ZN(_0328_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1356_ (.I(_0328_),
    .ZN(_0329_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1357_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .A2(_0327_),
    .B1(_0329_),
    .B2(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .ZN(_0330_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1358_ (.A1(_0326_),
    .A2(_0330_),
    .ZN(_0331_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1359_ (.A1(_0319_),
    .A2(_0331_),
    .Z(_0332_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1360_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q ),
    .A2(_0214_),
    .ZN(_0333_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1361_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q ),
    .A2(_0216_),
    .B(_0333_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q ),
    .ZN(_0334_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1362_ (.I0(_0225_),
    .I1(_0226_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q ),
    .Z(_0335_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1363_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q ),
    .A2(_0335_),
    .B(_0334_),
    .ZN(_0336_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1364_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .A2(_0323_),
    .B1(_0324_),
    .B2(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .ZN(_0337_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1365_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .A2(_0327_),
    .B1(_0329_),
    .B2(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .ZN(_0338_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1366_ (.A1(_0337_),
    .A2(_0338_),
    .B(_0319_),
    .ZN(_0339_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1367_ (.A1(_0332_),
    .A2(_0336_),
    .A3(_0339_),
    .Z(_0340_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1368_ (.A1(_0767_),
    .A2(_0319_),
    .ZN(_0341_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1369_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .A2(_0319_),
    .B(_0324_),
    .C(_0341_),
    .ZN(_0342_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1370_ (.I0(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .I1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .S(_0319_),
    .Z(_0343_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1371_ (.A1(_0766_),
    .A2(_0319_),
    .ZN(_0344_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1372_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .A2(_0319_),
    .B(_0327_),
    .C(_0344_),
    .ZN(_0345_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1373_ (.I0(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .I1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .S(_0319_),
    .Z(_0346_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1374_ (.A1(_0329_),
    .A2(_0343_),
    .B1(_0346_),
    .B2(_0323_),
    .ZN(_0347_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1375_ (.A1(_0336_),
    .A2(_0342_),
    .A3(_0345_),
    .A4(_0347_),
    .ZN(_0348_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1376_ (.A1(_0340_),
    .A2(_0348_),
    .ZN(_0349_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1377_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.LUT_flop ),
    .A2(\Inst_LF_LUT4c_frame_config_dffesr.c_out_mux ),
    .ZN(_0350_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1378_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.c_out_mux ),
    .A2(_0349_),
    .B(_0350_),
    .ZN(F),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1379_ (.A1(_0317_),
    .A2(_0323_),
    .B(_0325_),
    .ZN(_0351_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1380_ (.I0(E),
    .I1(H),
    .I2(F),
    .I3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ),
    .Z(_0352_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1381_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q ),
    .A2(_0352_),
    .ZN(_0353_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1382_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ),
    .Z(_0354_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1383_ (.A1(_0731_),
    .A2(_0354_),
    .B(_0732_),
    .ZN(_0355_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1384_ (.I0(N1END[3]),
    .I1(N2END[7]),
    .I2(E1END[3]),
    .I3(E2END[7]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ),
    .Z(_0356_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1385_ (.I0(S1END[3]),
    .I1(W1END[1]),
    .I2(S2END[7]),
    .I3(W1END[3]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ),
    .Z(_0357_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1386_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q ),
    .A2(_0357_),
    .ZN(_0358_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1387_ (.A1(_0731_),
    .A2(_0356_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q ),
    .ZN(_0359_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1388_ (.A1(_0353_),
    .A2(_0355_),
    .B1(_0358_),
    .B2(_0359_),
    .ZN(\Inst_LUT4AB_switch_matrix.JN2BEG6 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1389_ (.I0(N2MID[6]),
    .I1(E2MID[6]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q ),
    .Z(_0360_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1390_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q ),
    .A2(\Inst_LUT4AB_switch_matrix.JN2BEG6 ),
    .ZN(_0361_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1391_ (.A1(_0707_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q ),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit19.Q ),
    .C(_0361_),
    .ZN(_0362_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1392_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit19.Q ),
    .A2(_0360_),
    .B(_0362_),
    .ZN(_0363_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1393_ (.I0(N2MID[7]),
    .I1(E2MID[7]),
    .I2(S2MID[7]),
    .I3(W2MID[7]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit19.Q ),
    .Z(_0364_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1394_ (.I0(N4END[3]),
    .I1(EE4END[0]),
    .I2(S4END[3]),
    .I3(\Inst_LUT4AB_switch_matrix.JN2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit19.Q ),
    .Z(_0365_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1395_ (.I0(N2END[7]),
    .I1(E2END[7]),
    .I2(S2END[7]),
    .I3(WW4END[0]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit19.Q ),
    .Z(_0366_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1396_ (.I(_0366_),
    .ZN(_0367_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1397_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q ),
    .A2(_0364_),
    .ZN(_0368_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1398_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q ),
    .A2(_0363_),
    .B(_0368_),
    .ZN(_0369_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1399_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q ),
    .A2(_0365_),
    .ZN(_0370_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1400_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q ),
    .A2(_0367_),
    .B(_0370_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit31.Q ),
    .ZN(_0371_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1401_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit31.Q ),
    .A2(_0369_),
    .B(_0371_),
    .C(_0768_),
    .ZN(_0372_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1402_ (.A1(_0768_),
    .A2(_0351_),
    .B(_0372_),
    .ZN(_0373_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1403_ (.I0(N4END[2]),
    .I1(W2END[2]),
    .I2(SS4END[2]),
    .I3(\Inst_LUT4AB_switch_matrix.E2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit21.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit20.Q ),
    .Z(_0374_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1404_ (.I0(N2END[3]),
    .I1(SS4END[0]),
    .I2(E2END[3]),
    .I3(W2END[3]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit21.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit20.Q ),
    .Z(_0375_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1405_ (.I0(E),
    .I1(H),
    .I2(F),
    .I3(\Inst_LUT4AB_switch_matrix.M_AD ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ),
    .Z(_0376_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1406_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ),
    .Z(_0377_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1407_ (.A1(_0769_),
    .A2(_0377_),
    .ZN(_0378_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1408_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q ),
    .A2(_0376_),
    .B(_0770_),
    .ZN(_0379_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1409_ (.I0(S1END[1]),
    .I1(S1END[3]),
    .I2(S2END[7]),
    .I3(W1END[3]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ),
    .Z(_0380_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1410_ (.I0(N1END[3]),
    .I1(N2END[7]),
    .I2(E1END[3]),
    .I3(E2END[7]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ),
    .Z(_0381_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1411_ (.A1(_0769_),
    .A2(_0381_),
    .ZN(_0382_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1412_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q ),
    .A2(_0380_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q ),
    .ZN(_0383_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1413_ (.A1(_0378_),
    .A2(_0379_),
    .B1(_0382_),
    .B2(_0383_),
    .ZN(\Inst_LUT4AB_switch_matrix.E2BEG6 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1414_ (.I0(N2MID[2]),
    .I1(W2MID[2]),
    .I2(S2MID[2]),
    .I3(\Inst_LUT4AB_switch_matrix.E2BEG6 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit21.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit20.Q ),
    .Z(_0384_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1415_ (.I0(N2MID[3]),
    .I1(E2MID[3]),
    .I2(S2MID[3]),
    .I3(W2MID[3]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit20.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit21.Q ),
    .Z(_0385_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1416_ (.I0(_0384_),
    .I1(_0385_),
    .I2(_0375_),
    .I3(_0374_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit0.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit1.Q ),
    .Z(_0386_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1417_ (.I(_0386_),
    .ZN(_0387_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1418_ (.I0(E6END[1]),
    .I1(S4END[1]),
    .I2(WW4END[3]),
    .I3(\Inst_LUT4AB_switch_matrix.JS2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit23.Q ),
    .Z(_0388_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1419_ (.I0(NN4END[1]),
    .I1(S2END[5]),
    .I2(E2END[5]),
    .I3(W2END[5]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit22.Q ),
    .Z(_0389_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1420_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ),
    .Z(_0390_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1421_ (.A1(_0771_),
    .A2(_0390_),
    .ZN(_0391_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1422_ (.I0(E),
    .I1(H),
    .I2(F),
    .I3(\Inst_LUT4AB_switch_matrix.M_AB ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ),
    .Z(_0392_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1423_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q ),
    .A2(_0392_),
    .B(_0772_),
    .ZN(_0393_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1424_ (.I0(N1END[3]),
    .I1(N2END[7]),
    .I2(E1END[3]),
    .I3(E2END[7]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ),
    .Z(_0394_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1425_ (.I0(S1END[3]),
    .I1(W1END[1]),
    .I2(S2END[7]),
    .I3(W1END[3]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ),
    .Z(_0395_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1426_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q ),
    .A2(_0395_),
    .ZN(_0396_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1427_ (.A1(_0771_),
    .A2(_0394_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q ),
    .ZN(_0397_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1428_ (.A1(_0391_),
    .A2(_0393_),
    .B1(_0396_),
    .B2(_0397_),
    .ZN(\Inst_LUT4AB_switch_matrix.JS2BEG6 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1429_ (.I0(E2MID[4]),
    .I1(W2MID[4]),
    .I2(S2MID[4]),
    .I3(\Inst_LUT4AB_switch_matrix.JS2BEG6 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q ),
    .Z(_0398_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1430_ (.I0(N2MID[5]),
    .I1(E2MID[5]),
    .I2(S2MID[5]),
    .I3(W2MID[5]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit23.Q ),
    .Z(_0399_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1431_ (.I0(_0398_),
    .I1(_0399_),
    .I2(_0389_),
    .I3(_0388_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit3.Q ),
    .Z(_0400_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1432_ (.A1(_0386_),
    .A2(_0400_),
    .ZN(_0401_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1433_ (.A1(_0387_),
    .A2(_0400_),
    .ZN(_0402_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1434_ (.A1(_0386_),
    .A2(_0400_),
    .ZN(_0403_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1435_ (.I0(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .I1(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .I2(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .I3(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .S0(_0386_),
    .S1(_0400_),
    .Z(_0404_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1436_ (.I0(NN4END[0]),
    .I1(W2END[0]),
    .I2(E6END[0]),
    .I3(\Inst_LUT4AB_switch_matrix.JW2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit25.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit24.Q ),
    .Z(_0405_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1437_ (.I0(N2END[1]),
    .I1(EE4END[3]),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit24.Q ),
    .Z(_0406_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1438_ (.A1(W2END[1]),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit24.Q ),
    .ZN(_0407_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1439_ (.A1(_0764_),
    .A2(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit24.Q ),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit25.Q ),
    .C(_0407_),
    .ZN(_0408_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1440_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit25.Q ),
    .A2(_0406_),
    .B(_0408_),
    .ZN(_0409_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1441_ (.I(_0409_),
    .ZN(_0410_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1442_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ),
    .Z(_0411_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1443_ (.A1(_0773_),
    .A2(_0411_),
    .Z(_0412_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1444_ (.I0(E),
    .I1(H),
    .I2(F),
    .I3(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ),
    .Z(_0413_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1445_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q ),
    .A2(_0413_),
    .B(_0412_),
    .ZN(_0414_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1446_ (.I0(S1END[1]),
    .I1(S1END[3]),
    .I2(S2END[7]),
    .I3(W1END[3]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ),
    .Z(_0415_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1447_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q ),
    .A2(_0415_),
    .ZN(_0416_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1448_ (.I0(N1END[3]),
    .I1(N2END[7]),
    .I2(E1END[3]),
    .I3(E2END[7]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ),
    .Z(_0417_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1449_ (.A1(_0773_),
    .A2(_0417_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q ),
    .ZN(_0418_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1450_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q ),
    .A2(_0414_),
    .B1(_0416_),
    .B2(_0418_),
    .ZN(\Inst_LUT4AB_switch_matrix.JW2BEG6 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1451_ (.I0(N2MID[0]),
    .I1(E2MID[0]),
    .I2(W2MID[0]),
    .I3(\Inst_LUT4AB_switch_matrix.JW2BEG6 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit25.Q ),
    .Z(_0419_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1452_ (.I0(N2MID[1]),
    .I1(E2MID[1]),
    .I2(S2MID[1]),
    .I3(W2MID[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit25.Q ),
    .Z(_0420_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1453_ (.I0(_0419_),
    .I1(_0420_),
    .I2(_0410_),
    .I3(_0405_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit4.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit5.Q ),
    .Z(_0421_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1454_ (.A1(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .A2(_0387_),
    .A3(_0400_),
    .ZN(_0422_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1455_ (.A1(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .A2(_0402_),
    .B1(_0403_),
    .B2(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .ZN(_0423_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1456_ (.A1(_0774_),
    .A2(_0401_),
    .B(_0422_),
    .C(_0423_),
    .ZN(_0424_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1457_ (.I0(_0424_),
    .I1(_0404_),
    .S(_0373_),
    .Z(_0425_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1458_ (.I0(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .I1(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .I2(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .I3(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .S0(_0386_),
    .S1(_0400_),
    .Z(_0426_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1459_ (.I0(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .I1(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .I2(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .I3(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .S0(_0386_),
    .S1(_0400_),
    .Z(_0427_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1460_ (.I0(_0427_),
    .I1(_0426_),
    .S(_0373_),
    .Z(_0428_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1461_ (.I0(_0428_),
    .I1(_0425_),
    .S(_0421_),
    .Z(_0429_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1462_ (.I0(_0429_),
    .I1(\Inst_LG_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(\Inst_LG_LUT4c_frame_config_dffesr.c_out_mux ),
    .Z(G),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1463_ (.A1(_0317_),
    .A2(_0323_),
    .B1(_0386_),
    .B2(_0400_),
    .C(_0325_),
    .ZN(_0430_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1464_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q ),
    .A2(_0364_),
    .ZN(_0431_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1465_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q ),
    .A2(_0363_),
    .B(_0431_),
    .ZN(_0432_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1466_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q ),
    .A2(_0365_),
    .ZN(_0433_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1467_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q ),
    .A2(_0367_),
    .B(_0433_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q ),
    .ZN(_0434_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1468_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q ),
    .A2(_0432_),
    .B(_0434_),
    .C(_0775_),
    .ZN(_0435_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1469_ (.A1(_0775_),
    .A2(_0401_),
    .A3(_0430_),
    .B(_0435_),
    .ZN(_0436_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1470_ (.I0(_0398_),
    .I1(_0399_),
    .I2(_0389_),
    .I3(_0388_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit12.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit13.Q ),
    .Z(_0437_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1471_ (.I(_0437_),
    .ZN(_0438_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1472_ (.I0(_0384_),
    .I1(_0385_),
    .I2(_0375_),
    .I3(_0374_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit10.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit11.Q ),
    .Z(_0439_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1473_ (.I(_0439_),
    .ZN(_0440_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1474_ (.A1(_0437_),
    .A2(_0440_),
    .ZN(_0441_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1475_ (.A1(_0438_),
    .A2(_0439_),
    .ZN(_0442_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1476_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .A2(_0441_),
    .B1(_0442_),
    .B2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .ZN(_0443_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1477_ (.A1(_0438_),
    .A2(_0440_),
    .ZN(_0444_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1478_ (.A1(_0437_),
    .A2(_0439_),
    .ZN(_0445_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1479_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .A2(_0444_),
    .B1(_0445_),
    .B2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .ZN(_0446_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1480_ (.A1(_0443_),
    .A2(_0446_),
    .ZN(_0447_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1481_ (.I0(_0419_),
    .I1(_0420_),
    .I2(_0410_),
    .I3(_0405_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit15.Q ),
    .Z(_0448_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1482_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .A2(_0441_),
    .B1(_0444_),
    .B2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .ZN(_0449_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1483_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .A2(_0442_),
    .B1(_0445_),
    .B2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .ZN(_0450_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1484_ (.A1(_0449_),
    .A2(_0450_),
    .ZN(_0451_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1485_ (.I0(_0451_),
    .I1(_0447_),
    .S(_0436_),
    .Z(_0452_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1486_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .A2(_0441_),
    .B1(_0445_),
    .B2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .ZN(_0453_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1487_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .A2(_0442_),
    .B1(_0444_),
    .B2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .ZN(_0454_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1488_ (.A1(_0453_),
    .A2(_0454_),
    .ZN(_0455_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1489_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .A2(_0441_),
    .B1(_0444_),
    .B2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .ZN(_0456_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1490_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .A2(_0442_),
    .B1(_0445_),
    .B2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .ZN(_0457_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1491_ (.A1(_0456_),
    .A2(_0457_),
    .ZN(_0458_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1492_ (.I0(_0458_),
    .I1(_0455_),
    .S(_0436_),
    .Z(_0459_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1493_ (.I0(_0459_),
    .I1(_0452_),
    .S(_0448_),
    .Z(_0460_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1494_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.c_out_mux ),
    .A2(_0460_),
    .ZN(_0461_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1495_ (.A1(_0776_),
    .A2(\Inst_LH_LUT4c_frame_config_dffesr.c_out_mux ),
    .B(_0461_),
    .ZN(H),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1496_ (.I0(\Inst_LUT4AB_switch_matrix.JN2BEG6 ),
    .I1(\Inst_LUT4AB_switch_matrix.E2BEG6 ),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit22.Q ),
    .Z(_0462_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1497_ (.I0(\Inst_LUT4AB_switch_matrix.JS2BEG6 ),
    .I1(\Inst_LUT4AB_switch_matrix.JW2BEG6 ),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit22.Q ),
    .Z(_0463_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1498_ (.I0(_0462_),
    .I1(_0463_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit23.Q ),
    .Z(_0464_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1499_ (.I0(\Inst_LUT4AB_switch_matrix.JN2BEG4 ),
    .I1(\Inst_LUT4AB_switch_matrix.JS2BEG4 ),
    .I2(\Inst_LUT4AB_switch_matrix.E2BEG4 ),
    .I3(\Inst_LUT4AB_switch_matrix.JW2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit18.Q ),
    .Z(_0465_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1500_ (.I0(_0464_),
    .I1(_0465_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q ),
    .Z(_0466_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1501_ (.I0(E),
    .I1(F),
    .S(_0466_),
    .Z(\Inst_LUT4AB_switch_matrix.M_EF ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1502_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q ),
    .A2(_0252_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q ),
    .ZN(_0467_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1503_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q ),
    .A2(_0250_),
    .B(_0467_),
    .ZN(_0468_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1504_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q ),
    .A2(_0262_),
    .ZN(_0469_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1505_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q ),
    .A2(_0266_),
    .B(_0469_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q ),
    .ZN(_0470_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1506_ (.A1(_0468_),
    .A2(_0470_),
    .ZN(_0471_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1507_ (.I0(_0471_),
    .I1(_0155_),
    .S(\Inst_LD_LUT4c_frame_config_dffesr.c_I0mux ),
    .Z(_0472_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1508_ (.A1(_0123_),
    .A2(_0144_),
    .ZN(_0473_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1509_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .A2(_0146_),
    .B1(_0473_),
    .B2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .ZN(_0474_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1510_ (.A1(_0123_),
    .A2(_0144_),
    .Z(_0475_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1511_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .A2(_0147_),
    .B1(_0475_),
    .B2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .ZN(_0476_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1512_ (.A1(_0474_),
    .A2(_0476_),
    .ZN(_0477_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1513_ (.A1(_0472_),
    .A2(_0477_),
    .ZN(_0478_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1514_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .A2(_0146_),
    .B1(_0475_),
    .B2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .ZN(_0479_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1515_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .A2(_0147_),
    .B1(_0473_),
    .B2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .ZN(_0480_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1516_ (.A1(_0479_),
    .A2(_0480_),
    .B(_0472_),
    .ZN(_0481_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1517_ (.I(_0481_),
    .ZN(_0482_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1518_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit6.Q ),
    .A2(_0289_),
    .ZN(_0483_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1519_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit6.Q ),
    .A2(_0291_),
    .B(_0483_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit7.Q ),
    .ZN(_0484_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1520_ (.I0(_0300_),
    .I1(_0301_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit6.Q ),
    .Z(_0485_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1521_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit7.Q ),
    .A2(_0485_),
    .B(_0484_),
    .ZN(_0486_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1522_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .A2(_0146_),
    .B1(_0147_),
    .B2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .ZN(_0487_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1523_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .A2(_0473_),
    .B1(_0475_),
    .B2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .ZN(_0488_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1524_ (.A1(_0487_),
    .A2(_0488_),
    .B(_0472_),
    .ZN(_0489_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1525_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .A2(_0146_),
    .B1(_0147_),
    .B2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .ZN(_0490_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1526_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .A2(_0473_),
    .B1(_0475_),
    .B2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .ZN(_0491_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1527_ (.A1(_0490_),
    .A2(_0491_),
    .ZN(_0492_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1528_ (.A1(_0472_),
    .A2(_0492_),
    .Z(_0493_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1529_ (.A1(_0486_),
    .A2(_0489_),
    .A3(_0493_),
    .ZN(_0494_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1530_ (.A1(_0478_),
    .A2(_0482_),
    .A3(_0486_),
    .B(_0494_),
    .ZN(_0495_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1531_ (.I0(_0495_),
    .I1(\Inst_LD_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(\Inst_LD_LUT4c_frame_config_dffesr.c_out_mux ),
    .Z(D),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1532_ (.I0(\Inst_LUT4AB_switch_matrix.JN2BEG5 ),
    .I1(\Inst_LUT4AB_switch_matrix.E2BEG5 ),
    .I2(\Inst_LUT4AB_switch_matrix.JS2BEG5 ),
    .I3(\Inst_LUT4AB_switch_matrix.JW2BEG5 ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit21.Q ),
    .Z(_0496_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1533_ (.I0(_0465_),
    .I1(_0496_),
    .S(_0783_),
    .Z(_0497_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1534_ (.I0(C),
    .I1(D),
    .S(_0497_),
    .Z(_0498_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1535_ (.I0(\Inst_LUT4AB_switch_matrix.M_AB ),
    .I1(_0498_),
    .S(_0496_),
    .Z(_0499_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1536_ (.I0(_0498_),
    .I1(_0499_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.M_AD ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1537_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ),
    .Z(_0500_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1538_ (.I0(E),
    .I1(G),
    .I2(F),
    .I3(\Inst_LUT4AB_switch_matrix.M_AD ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ),
    .Z(_0501_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1539_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q ),
    .A2(_0501_),
    .ZN(_0502_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1540_ (.A1(_0781_),
    .A2(_0500_),
    .B(_0782_),
    .ZN(_0503_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1541_ (.I0(N1END[0]),
    .I1(N2END[0]),
    .I2(E1END[0]),
    .I3(E2END[0]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ),
    .Z(_0504_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1542_ (.I0(S1END[0]),
    .I1(W1END[0]),
    .I2(S2END[0]),
    .I3(W1END[2]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ),
    .Z(_0505_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1543_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q ),
    .A2(_0505_),
    .ZN(_0506_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1544_ (.A1(_0781_),
    .A2(_0504_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q ),
    .ZN(_0507_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1545_ (.A1(_0502_),
    .A2(_0503_),
    .B1(_0506_),
    .B2(_0507_),
    .ZN(\Inst_LUT4AB_switch_matrix.JS2BEG7 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1546_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ),
    .Z(_0508_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1547_ (.I(_0508_),
    .ZN(_0509_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1548_ (.I0(E),
    .I1(G),
    .I2(F),
    .I3(\Inst_LUT4AB_switch_matrix.M_AB ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ),
    .Z(_0510_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1549_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q ),
    .A2(_0510_),
    .ZN(_0511_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1550_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q ),
    .A2(_0509_),
    .B(_0511_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q ),
    .ZN(_0512_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1551_ (.I0(N1END[0]),
    .I1(NN4END[0]),
    .I2(E1END[0]),
    .I3(E2END[0]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ),
    .Z(_0513_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1552_ (.I0(S1END[0]),
    .I1(S1END[2]),
    .I2(S2END[0]),
    .I3(W1END[0]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ),
    .Z(_0514_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1553_ (.I0(_0513_),
    .I1(_0514_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q ),
    .Z(_0515_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1554_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q ),
    .A2(_0515_),
    .B(_0512_),
    .ZN(_0516_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1555_ (.I(_0516_),
    .ZN(\Inst_LUT4AB_switch_matrix.JW2BEG7 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1556_ (.I0(E),
    .I1(G),
    .I2(F),
    .I3(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ),
    .Z(_0517_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1557_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ),
    .Z(_0518_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1558_ (.A1(_0777_),
    .A2(_0518_),
    .ZN(_0519_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1559_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q ),
    .A2(_0517_),
    .B(_0778_),
    .ZN(_0520_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1560_ (.I0(N1END[0]),
    .I1(N2END[0]),
    .I2(E1END[0]),
    .I3(EE4END[0]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ),
    .Z(_0521_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1561_ (.A1(_0777_),
    .A2(_0521_),
    .ZN(_0522_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1562_ (.I0(S1END[0]),
    .I1(W1END[0]),
    .I2(S2END[0]),
    .I3(W1END[2]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ),
    .Z(_0523_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1563_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q ),
    .A2(_0523_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q ),
    .ZN(_0524_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1564_ (.A1(_0519_),
    .A2(_0520_),
    .B1(_0522_),
    .B2(_0524_),
    .ZN(\Inst_LUT4AB_switch_matrix.JN2BEG7 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1565_ (.I0(A),
    .I1(B),
    .I2(C),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ),
    .Z(_0525_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1566_ (.I0(E),
    .I1(G),
    .I2(F),
    .I3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ),
    .Z(_0526_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1567_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q ),
    .A2(_0526_),
    .ZN(_0527_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1568_ (.A1(_0779_),
    .A2(_0525_),
    .B(_0780_),
    .ZN(_0528_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1569_ (.I0(S1END[0]),
    .I1(S1END[2]),
    .I2(SS4END[0]),
    .I3(WW4END[0]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ),
    .Z(_0529_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1570_ (.I0(N1END[0]),
    .I1(N2END[0]),
    .I2(E1END[0]),
    .I3(E2END[0]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ),
    .Z(_0530_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1571_ (.A1(_0779_),
    .A2(_0530_),
    .ZN(_0531_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1572_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q ),
    .A2(_0529_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q ),
    .ZN(_0532_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1573_ (.A1(_0527_),
    .A2(_0528_),
    .B1(_0531_),
    .B2(_0532_),
    .ZN(\Inst_LUT4AB_switch_matrix.E2BEG7 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1574_ (.I(\Inst_LUT4AB_switch_matrix.E2BEG7 ),
    .ZN(_0533_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1575_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q ),
    .A2(_0533_),
    .ZN(_0534_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1576_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q ),
    .A2(\Inst_LUT4AB_switch_matrix.JN2BEG7 ),
    .B(_0534_),
    .ZN(_0535_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1577_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q ),
    .A2(_0516_),
    .ZN(_0536_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1578_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q ),
    .A2(\Inst_LUT4AB_switch_matrix.JS2BEG7 ),
    .B(_0536_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q ),
    .ZN(_0537_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1579_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q ),
    .A2(_0535_),
    .B(_0537_),
    .ZN(_0538_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1580_ (.I0(_0538_),
    .I1(_0496_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q ),
    .Z(_0539_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1581_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ),
    .A2(_0466_),
    .Z(_0540_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1582_ (.A1(_0783_),
    .A2(_0539_),
    .B(_0540_),
    .ZN(_0541_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1583_ (.I0(H),
    .I1(G),
    .S(_0541_),
    .Z(_0542_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1584_ (.I0(\Inst_LUT4AB_switch_matrix.M_EF ),
    .I1(_0542_),
    .S(_0539_),
    .Z(_0543_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1585_ (.I0(_0499_),
    .I1(_0543_),
    .S(_0538_),
    .Z(_0544_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1586_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q ),
    .A2(_0544_),
    .ZN(_0545_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1587_ (.A1(_0783_),
    .A2(_0543_),
    .ZN(_0546_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1588_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ),
    .A2(_0542_),
    .ZN(_0547_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1589_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q ),
    .A2(_0546_),
    .A3(_0547_),
    .B(_0545_),
    .ZN(\Inst_LUT4AB_switch_matrix.M_AH ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1590_ (.I0(A),
    .I1(B),
    .S(_0465_),
    .Z(\Inst_LUT4AB_switch_matrix.M_AB ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1591_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_AD ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ),
    .Z(_0548_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1592_ (.A1(_0784_),
    .A2(_0548_),
    .ZN(_0549_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1593_ (.I0(B),
    .I1(D),
    .I2(C),
    .I3(E),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ),
    .Z(_0550_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1594_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q ),
    .A2(_0550_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q ),
    .ZN(_0551_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1595_ (.I0(S2END[1]),
    .I1(W2END[1]),
    .I2(S4END[1]),
    .I3(W6END[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ),
    .Z(_0552_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1596_ (.A1(_0784_),
    .A2(_0552_),
    .ZN(_0553_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1597_ (.I0(N1END[3]),
    .I1(E2END[1]),
    .I2(N2END[1]),
    .I3(E6END[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ),
    .Z(_0554_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1598_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q ),
    .A2(_0554_),
    .ZN(_0555_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1599_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q ),
    .A2(_0553_),
    .A3(_0555_),
    .B1(_0549_),
    .B2(_0551_),
    .ZN(\Inst_LUT4AB_switch_matrix.JW2BEG0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1600_ (.I0(B),
    .I1(D),
    .I2(C),
    .I3(E),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ),
    .Z(_0556_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1601_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ),
    .Z(_0557_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1602_ (.I(_0557_),
    .ZN(_0558_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1603_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q ),
    .A2(_0558_),
    .ZN(_0559_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1604_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q ),
    .A2(_0556_),
    .B(_0559_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q ),
    .ZN(_0560_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1605_ (.I0(NN4END[1]),
    .I1(E2END[1]),
    .I2(E1END[3]),
    .I3(E6END[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ),
    .Z(_0561_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1606_ (.I0(S2END[1]),
    .I1(W2END[1]),
    .I2(S4END[1]),
    .I3(W6END[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ),
    .Z(_0562_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1607_ (.I(_0562_),
    .ZN(_0563_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1608_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q ),
    .A2(_0563_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q ),
    .ZN(_0564_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1609_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q ),
    .A2(_0561_),
    .B(_0564_),
    .ZN(_0565_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1610_ (.A1(_0560_),
    .A2(_0565_),
    .ZN(\Inst_LUT4AB_switch_matrix.JS2BEG0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1611_ (.I0(B),
    .I1(D),
    .I2(C),
    .I3(E),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ),
    .Z(_0566_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1612_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q ),
    .A2(_0566_),
    .ZN(_0567_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1613_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ),
    .Z(_0568_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1614_ (.A1(_0785_),
    .A2(_0568_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q ),
    .ZN(_0569_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1615_ (.I0(N1END[3]),
    .I1(N2END[1]),
    .I2(N4END[1]),
    .I3(EE4END[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ),
    .Z(_0570_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1616_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q ),
    .A2(_0570_),
    .ZN(_0571_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1617_ (.I0(E6END[1]),
    .I1(W2END[1]),
    .I2(S2END[1]),
    .I3(W6END[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ),
    .Z(_0572_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1618_ (.A1(_0785_),
    .A2(_0572_),
    .ZN(_0573_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1619_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q ),
    .A2(_0571_),
    .A3(_0573_),
    .B1(_0567_),
    .B2(_0569_),
    .ZN(\Inst_LUT4AB_switch_matrix.E2BEG0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1620_ (.I0(B),
    .I1(D),
    .I2(C),
    .I3(E),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ),
    .Z(_0574_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1621_ (.I0(F),
    .I1(G),
    .I2(H),
    .I3(\Inst_LUT4AB_switch_matrix.M_AB ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ),
    .Z(_0575_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1622_ (.I(_0575_),
    .ZN(_0576_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1623_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q ),
    .A2(_0576_),
    .ZN(_0577_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1624_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q ),
    .A2(_0574_),
    .B(_0577_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q ),
    .ZN(_0578_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1625_ (.I0(E6END[1]),
    .I1(SS4END[1]),
    .I2(W2END[1]),
    .I3(W6END[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ),
    .Z(_0579_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1626_ (.I(_0579_),
    .ZN(_0580_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1627_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q ),
    .A2(_0580_),
    .ZN(_0581_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1628_ (.I0(N2END[1]),
    .I1(E1END[3]),
    .I2(N4END[1]),
    .I3(E2END[1]),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ),
    .Z(_0582_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1629_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q ),
    .A2(_0582_),
    .B(_0581_),
    .ZN(_0583_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1630_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q ),
    .A2(_0583_),
    .B(_0578_),
    .ZN(\Inst_LUT4AB_switch_matrix.JN2BEG0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1631_ (.I0(E1END[2]),
    .I1(W1END[2]),
    .I2(A),
    .I3(B),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ),
    .Z(_0584_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1632_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q ),
    .A2(_0584_),
    .ZN(_0585_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1633_ (.I0(C),
    .I1(D),
    .I2(E),
    .I3(F),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ),
    .Z(_0586_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1634_ (.A1(_0786_),
    .A2(_0586_),
    .ZN(_0587_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1635_ (.I0(_0018_),
    .I1(_0142_),
    .I2(_0204_),
    .I3(_0398_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ),
    .Z(_0588_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1636_ (.A1(_0786_),
    .A2(_0588_),
    .ZN(_0589_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1637_ (.I0(G),
    .I1(H),
    .I2(\Inst_LUT4AB_switch_matrix.M_AD ),
    .I3(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ),
    .Z(_0590_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1638_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q ),
    .A2(_0590_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q ),
    .ZN(_0591_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1639_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q ),
    .A2(_0585_),
    .A3(_0587_),
    .B1(_0589_),
    .B2(_0591_),
    .ZN(\Inst_LUT4AB_switch_matrix.W6BEG1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1640_ (.I0(E1END[3]),
    .I1(W1END[3]),
    .I2(A),
    .I3(B),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ),
    .Z(_0592_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1641_ (.I0(C),
    .I1(D),
    .I2(E),
    .I3(F),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ),
    .Z(_0593_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1642_ (.I0(_0800_),
    .I1(_0110_),
    .I2(_0192_),
    .I3(_0385_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ),
    .Z(_0594_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1643_ (.I0(G),
    .I1(H),
    .I2(\Inst_LUT4AB_switch_matrix.M_AB ),
    .I3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ),
    .Z(_0595_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1644_ (.I0(_0592_),
    .I1(_0593_),
    .I2(_0595_),
    .I3(_0594_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit29.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.W6BEG0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1645_ (.I0(E),
    .I1(_0204_),
    .I2(_0398_),
    .I3(_0851_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit24.Q ),
    .Z(_0596_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1646_ (.I0(N1END[1]),
    .I1(S1END[1]),
    .I2(W1END[1]),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit24.Q ),
    .Z(_0597_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1647_ (.I0(_0597_),
    .I1(_0596_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit25.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.WW4BEG3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1648_ (.I0(C),
    .I1(_0192_),
    .I2(_0385_),
    .I3(_0133_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q ),
    .Z(_0598_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1649_ (.I0(N1END[0]),
    .I1(W1END[0]),
    .I2(S1END[0]),
    .I3(B),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q ),
    .Z(_0599_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1650_ (.I0(_0599_),
    .I1(_0598_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit22.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.WW4BEG2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1651_ (.I0(H),
    .I1(_0018_),
    .I2(_0142_),
    .I3(_0195_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q ),
    .Z(_0600_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1652_ (.I0(N1END[3]),
    .I1(S1END[3]),
    .I2(W1END[3]),
    .I3(A),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q ),
    .Z(_0601_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1653_ (.I0(_0601_),
    .I1(_0600_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit19.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.WW4BEG1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1654_ (.I0(G),
    .I1(_0800_),
    .I2(_0110_),
    .I3(_0389_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q ),
    .Z(_0602_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1655_ (.I0(N1END[2]),
    .I1(S1END[2]),
    .I2(W1END[2]),
    .I3(F),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q ),
    .Z(_0603_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1656_ (.I0(_0603_),
    .I1(_0602_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit16.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.WW4BEG0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1657_ (.I0(E),
    .I1(_0204_),
    .I2(_0398_),
    .I3(_0036_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q ),
    .Z(_0604_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1658_ (.I0(N1END[1]),
    .I1(E1END[1]),
    .I2(W1END[1]),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q ),
    .Z(_0605_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1659_ (.I0(_0605_),
    .I1(_0604_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit5.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.SS4BEG3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1660_ (.I0(C),
    .I1(_0192_),
    .I2(_0385_),
    .I3(_0290_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q ),
    .Z(_0606_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1661_ (.I0(N1END[0]),
    .I1(W1END[0]),
    .I2(E1END[0]),
    .I3(B),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q ),
    .Z(_0607_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1662_ (.I0(_0607_),
    .I1(_0606_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit2.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.SS4BEG2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1663_ (.I0(H),
    .I1(_0018_),
    .I2(_0142_),
    .I3(_0215_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q ),
    .Z(_0608_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1664_ (.I0(N1END[3]),
    .I1(E1END[3]),
    .I2(W1END[3]),
    .I3(A),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q ),
    .Z(_0609_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1665_ (.I0(_0609_),
    .I1(_0608_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.SS4BEG1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1666_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ),
    .A2(_0409_),
    .ZN(_0610_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1667_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ),
    .A2(_0110_),
    .B(_0610_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q ),
    .ZN(_0611_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1668_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ),
    .A2(_0799_),
    .ZN(_0612_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1669_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ),
    .A2(G),
    .B(_0612_),
    .ZN(_0613_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1670_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q ),
    .A2(_0613_),
    .B(_0611_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q ),
    .ZN(_0614_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1671_ (.I0(N1END[2]),
    .I1(W1END[2]),
    .I2(E1END[2]),
    .I3(F),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ),
    .Z(_0615_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1672_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q ),
    .A2(_0615_),
    .B(_0614_),
    .ZN(_0616_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1673_ (.I(_0616_),
    .ZN(\Inst_LUT4AB_switch_matrix.SS4BEG0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1674_ (.I0(E1END[2]),
    .I1(W1END[2]),
    .I2(A),
    .I3(B),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ),
    .Z(_0617_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1675_ (.I0(C),
    .I1(D),
    .I2(E),
    .I3(F),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ),
    .Z(_0618_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1676_ (.I0(_0617_),
    .I1(_0618_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q ),
    .Z(_0619_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1677_ (.I0(G),
    .I1(H),
    .I2(\Inst_LUT4AB_switch_matrix.M_AD ),
    .I3(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ),
    .Z(_0620_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1678_ (.I0(_0018_),
    .I1(_0142_),
    .I2(_0204_),
    .I3(_0398_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ),
    .Z(_0621_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1679_ (.I0(_0620_),
    .I1(_0621_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q ),
    .Z(_0622_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1680_ (.I0(_0619_),
    .I1(_0622_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit9.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.E6BEG1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1681_ (.I0(E1END[3]),
    .I1(W1END[3]),
    .I2(A),
    .I3(B),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ),
    .Z(_0623_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1682_ (.I0(C),
    .I1(D),
    .I2(E),
    .I3(F),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ),
    .Z(_0624_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1683_ (.I0(_0800_),
    .I1(_0110_),
    .I2(_0192_),
    .I3(_0385_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ),
    .Z(_0625_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1684_ (.I0(G),
    .I1(H),
    .I2(\Inst_LUT4AB_switch_matrix.M_AB ),
    .I3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ),
    .Z(_0626_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1685_ (.I0(_0623_),
    .I1(_0624_),
    .I2(_0626_),
    .I3(_0625_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit5.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.E6BEG0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1686_ (.I0(E),
    .I1(_0204_),
    .I2(_0398_),
    .I3(_0831_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q ),
    .Z(_0627_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1687_ (.I0(N1END[1]),
    .I1(E1END[1]),
    .I2(S1END[1]),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q ),
    .Z(_0628_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1688_ (.I0(_0628_),
    .I1(_0627_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit1.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.EE4BEG3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1689_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q ),
    .A2(_0266_),
    .ZN(_0629_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1690_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q ),
    .A2(_0385_),
    .B(_0629_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q ),
    .ZN(_0630_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1691_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q ),
    .A2(_0191_),
    .ZN(_0631_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1692_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q ),
    .A2(C),
    .B(_0631_),
    .ZN(_0632_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1693_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q ),
    .A2(_0632_),
    .B(_0630_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q ),
    .ZN(_0633_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1694_ (.I0(N1END[0]),
    .I1(S1END[0]),
    .I2(E1END[0]),
    .I3(B),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q ),
    .Z(_0634_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1695_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q ),
    .A2(_0634_),
    .B(_0633_),
    .ZN(_0635_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1696_ (.I(_0635_),
    .ZN(\Inst_LUT4AB_switch_matrix.EE4BEG2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1697_ (.I0(H),
    .I1(_0018_),
    .I2(_0142_),
    .I3(_0158_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q ),
    .Z(_0636_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1698_ (.I0(N1END[3]),
    .I1(E1END[3]),
    .I2(S1END[3]),
    .I3(A),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q ),
    .Z(_0637_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1699_ (.I0(_0637_),
    .I1(_0636_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit27.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.EE4BEG1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1700_ (.I0(G),
    .I1(_0800_),
    .I2(_0110_),
    .I3(_0366_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q ),
    .Z(_0638_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1701_ (.I0(N1END[2]),
    .I1(S1END[2]),
    .I2(E1END[2]),
    .I3(F),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q ),
    .Z(_0639_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1702_ (.I0(_0639_),
    .I1(_0638_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit24.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.EE4BEG0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1703_ (.I0(E),
    .I1(_0204_),
    .I2(_0398_),
    .I3(_0810_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit12.Q ),
    .Z(_0640_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1704_ (.I0(N1END[1]),
    .I1(E1END[1]),
    .I2(W1END[1]),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit12.Q ),
    .Z(_0641_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1705_ (.I0(_0641_),
    .I1(_0640_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit13.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.NN4BEG3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1706_ (.I0(C),
    .I1(_0192_),
    .I2(_0385_),
    .I3(_0121_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q ),
    .Z(_0642_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1707_ (.I0(N1END[0]),
    .I1(W1END[0]),
    .I2(E1END[0]),
    .I3(B),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q ),
    .Z(_0643_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1708_ (.I0(_0643_),
    .I1(_0642_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit10.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.NN4BEG2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1709_ (.I0(H),
    .I1(_0018_),
    .I2(_0142_),
    .I3(_0178_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q ),
    .Z(_0644_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1710_ (.I0(N1END[3]),
    .I1(E1END[3]),
    .I2(W1END[3]),
    .I3(A),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q ),
    .Z(_0645_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1711_ (.I0(_0645_),
    .I1(_0644_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit7.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.NN4BEG1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1712_ (.I0(G),
    .I1(_0800_),
    .I2(_0110_),
    .I3(_0375_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q ),
    .Z(_0646_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1713_ (.I0(N1END[2]),
    .I1(W1END[2]),
    .I2(E1END[2]),
    .I3(F),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q ),
    .Z(_0647_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1714_ (.I0(_0647_),
    .I1(_0646_),
    .S(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit4.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.NN4BEG0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1715_ (.I0(A),
    .I1(_0020_),
    .I2(\Inst_LUT4AB_switch_matrix.JS2BEG2 ),
    .I3(_0830_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit12.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit13.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.W1BEG3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1716_ (.I0(H),
    .I1(\Inst_LUT4AB_switch_matrix.JS2BEG1 ),
    .I2(_0385_),
    .I3(_0405_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit10.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.W1BEG2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1717_ (.I0(G),
    .I1(_0173_),
    .I2(\Inst_LUT4AB_switch_matrix.JS2BEG0 ),
    .I3(_0194_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit8.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit9.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.W1BEG1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1718_ (.I0(F),
    .I1(\Inst_LUT4AB_switch_matrix.JS2BEG3 ),
    .I2(_0301_),
    .I3(_0120_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit7.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit6.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.W1BEG0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1719_ (.I0(S2END[1]),
    .I1(S4END[0]),
    .I2(W6END[0]),
    .I3(D),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit24.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit25.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.S4BEG3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1720_ (.I0(S2END[0]),
    .I1(W6END[1]),
    .I2(S4END[3]),
    .I3(C),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit22.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.S4BEG2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1721_ (.I0(E6END[0]),
    .I1(S4END[2]),
    .I2(S2END[3]),
    .I3(B),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit21.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit20.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.S4BEG1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1722_ (.I0(E6END[1]),
    .I1(S4END[1]),
    .I2(S2END[2]),
    .I3(A),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit18.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.S4BEG0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1723_ (.I0(H),
    .I1(_0020_),
    .I2(\Inst_LUT4AB_switch_matrix.E2BEG2 ),
    .I3(_0830_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit16.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit17.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.S1BEG3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1724_ (.I0(G),
    .I1(\Inst_LUT4AB_switch_matrix.E2BEG1 ),
    .I2(_0385_),
    .I3(_0405_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit15.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit14.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.S1BEG2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1725_ (.I0(F),
    .I1(_0173_),
    .I2(\Inst_LUT4AB_switch_matrix.E2BEG0 ),
    .I3(_0194_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit12.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit13.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.S1BEG1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1726_ (.I0(E),
    .I1(\Inst_LUT4AB_switch_matrix.E2BEG3 ),
    .I2(_0301_),
    .I3(_0120_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit11.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit10.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.S1BEG0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1727_ (.I0(G),
    .I1(_0020_),
    .I2(\Inst_LUT4AB_switch_matrix.JN2BEG2 ),
    .I3(_0830_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit20.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit21.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.E1BEG3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1728_ (.I0(F),
    .I1(\Inst_LUT4AB_switch_matrix.JN2BEG1 ),
    .I2(_0385_),
    .I3(_0405_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit18.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.E1BEG2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1729_ (.I0(E),
    .I1(_0173_),
    .I2(\Inst_LUT4AB_switch_matrix.JN2BEG0 ),
    .I3(_0194_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit16.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit17.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.E1BEG1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1730_ (.I0(D),
    .I1(\Inst_LUT4AB_switch_matrix.JN2BEG3 ),
    .I2(_0301_),
    .I3(_0120_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit15.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit14.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.E1BEG0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1731_ (.I0(N2END[1]),
    .I1(W6END[0]),
    .I2(N4END[0]),
    .I3(H),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit1.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit0.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.N4BEG3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1732_ (.I0(N2END[0]),
    .I1(N4END[3]),
    .I2(W6END[1]),
    .I3(G),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit30.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit31.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.N4BEG2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1733_ (.I0(N2END[3]),
    .I1(N4END[2]),
    .I2(E6END[0]),
    .I3(F),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit28.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit29.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.N4BEG1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1734_ (.I0(N2END[2]),
    .I1(N4END[1]),
    .I2(E6END[1]),
    .I3(E),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit26.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit27.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.N4BEG0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1735_ (.I0(F),
    .I1(_0020_),
    .I2(\Inst_LUT4AB_switch_matrix.JW2BEG2 ),
    .I3(_0830_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit24.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit25.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.N1BEG3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1736_ (.I0(E),
    .I1(\Inst_LUT4AB_switch_matrix.JW2BEG1 ),
    .I2(_0385_),
    .I3(_0405_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit23.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit22.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.N1BEG2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1737_ (.I0(D),
    .I1(_0173_),
    .I2(\Inst_LUT4AB_switch_matrix.JW2BEG0 ),
    .I3(_0194_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit20.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit21.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.N1BEG1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1738_ (.I0(C),
    .I1(\Inst_LUT4AB_switch_matrix.JW2BEG3 ),
    .I2(_0301_),
    .I3(_0120_),
    .S0(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit19.Q ),
    .S1(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit18.Q ),
    .Z(\Inst_LUT4AB_switch_matrix.N1BEG0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1739_ (.A1(_0401_),
    .A2(_0430_),
    .B(_0445_),
    .ZN(_0648_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1740_ (.A1(_0444_),
    .A2(_0648_),
    .Z(net1),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1741_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ),
    .A2(_0419_),
    .ZN(_0649_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1742_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ),
    .A2(_0047_),
    .B(_0649_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q ),
    .ZN(_0650_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1743_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ),
    .A2(_0301_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q ),
    .ZN(_0651_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1744_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ),
    .A2(_0227_),
    .B(_0651_),
    .ZN(_0652_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1745_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ),
    .A2(\Inst_LUT4AB_switch_matrix.JN2BEG2 ),
    .ZN(_0653_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1746_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ),
    .A2(_0119_),
    .B(_0653_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q ),
    .ZN(_0654_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1747_ (.A1(_0284_),
    .A2(_0288_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ),
    .ZN(_0655_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1748_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ),
    .A2(\Inst_LUT4AB_switch_matrix.JS2BEG2 ),
    .B(_0655_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q ),
    .ZN(_0656_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1749_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q ),
    .A2(_0656_),
    .ZN(_0657_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1750_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q ),
    .A2(_0650_),
    .A3(_0652_),
    .B1(_0654_),
    .B2(_0657_),
    .ZN(_0658_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1751_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit17.Q ),
    .A2(_0658_),
    .ZN(_0659_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1752_ (.A1(_0733_),
    .A2(_0363_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q ),
    .ZN(_0660_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1753_ (.A1(_0733_),
    .A2(_0821_),
    .B(_0660_),
    .ZN(_0661_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1754_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ),
    .A2(_0252_),
    .B(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q ),
    .ZN(_0662_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1755_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ),
    .A2(_0172_),
    .B(_0662_),
    .ZN(_0663_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1756_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q ),
    .A2(_0663_),
    .ZN(_0664_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1757_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ),
    .A2(\Inst_LUT4AB_switch_matrix.JS2BEG1 ),
    .Z(_0665_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1758_ (.A1(_0733_),
    .A2(\Inst_LUT4AB_switch_matrix.JW2BEG1 ),
    .B(_0665_),
    .C(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q ),
    .ZN(_0666_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1759_ (.A1(_0733_),
    .A2(\Inst_LUT4AB_switch_matrix.E2BEG1 ),
    .ZN(_0667_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1760_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q ),
    .A2(_0667_),
    .ZN(_0668_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1761_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ),
    .A2(\Inst_LUT4AB_switch_matrix.JN2BEG1 ),
    .B(_0668_),
    .ZN(_0669_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1762_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q ),
    .A2(_0666_),
    .A3(_0669_),
    .Z(_0670_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1763_ (.A1(_0661_),
    .A2(_0664_),
    .B(_0670_),
    .ZN(_0671_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1764_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit16.Q ),
    .A2(_0671_),
    .ZN(_0672_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1765_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit16.Q ),
    .A2(_0671_),
    .B(_0460_),
    .ZN(_0673_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1766_ (.A1(\Inst_LH_LUT4c_frame_config_dffesr.c_reset_value ),
    .A2(_0672_),
    .B(_0659_),
    .ZN(_0674_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1767_ (.A1(_0776_),
    .A2(_0659_),
    .B1(_0673_),
    .B2(_0674_),
    .ZN(_0000_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1768_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit10.Q ),
    .A2(_0671_),
    .ZN(_0675_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1769_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit11.Q ),
    .A2(_0658_),
    .ZN(_0676_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1770_ (.A1(_0063_),
    .A2(_0675_),
    .ZN(_0677_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1771_ (.A1(\Inst_LA_LUT4c_frame_config_dffesr.c_reset_value ),
    .A2(_0675_),
    .B(_0676_),
    .C(_0677_),
    .ZN(_0678_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1772_ (.A1(_0734_),
    .A2(_0676_),
    .B(_0678_),
    .ZN(_0001_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1773_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit21.Q ),
    .A2(_0658_),
    .Z(_0679_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1774_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit20.Q ),
    .A2(_0671_),
    .ZN(_0680_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1775_ (.I0(\Inst_LB_LUT4c_frame_config_dffesr.c_reset_value ),
    .I1(_0100_),
    .S(_0680_),
    .Z(_0681_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1776_ (.I0(_0681_),
    .I1(\Inst_LB_LUT4c_frame_config_dffesr.LUT_flop ),
    .S(_0679_),
    .Z(_0002_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1777_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit31.Q ),
    .A2(_0658_),
    .Z(_0682_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1778_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.LUT_flop ),
    .A2(_0682_),
    .ZN(_0683_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1779_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit30.Q ),
    .A2(_0671_),
    .ZN(_0684_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1780_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit30.Q ),
    .A2(_0671_),
    .B(_0316_),
    .ZN(_0685_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1781_ (.A1(\Inst_LC_LUT4c_frame_config_dffesr.c_reset_value ),
    .A2(_0684_),
    .ZN(_0686_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1782_ (.A1(_0682_),
    .A2(_0685_),
    .A3(_0686_),
    .B(_0683_),
    .ZN(_0003_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1783_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit9.Q ),
    .A2(_0658_),
    .Z(_0687_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1784_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.LUT_flop ),
    .A2(_0687_),
    .ZN(_0688_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1785_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit8.Q ),
    .A2(_0671_),
    .ZN(_0689_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1786_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit8.Q ),
    .A2(_0671_),
    .B(_0495_),
    .ZN(_0690_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1787_ (.A1(\Inst_LD_LUT4c_frame_config_dffesr.c_reset_value ),
    .A2(_0689_),
    .ZN(_0691_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1788_ (.A1(_0687_),
    .A2(_0690_),
    .A3(_0691_),
    .B(_0688_),
    .ZN(_0004_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1789_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit19.Q ),
    .A2(_0658_),
    .Z(_0692_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1790_ (.A1(\Inst_LE_LUT4c_frame_config_dffesr.LUT_flop ),
    .A2(_0692_),
    .ZN(_0693_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1791_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit18.Q ),
    .A2(_0671_),
    .ZN(_0694_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1792_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit18.Q ),
    .A2(_0671_),
    .B(_0238_),
    .ZN(_0695_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1793_ (.A1(\Inst_LE_LUT4c_frame_config_dffesr.c_reset_value ),
    .A2(_0694_),
    .ZN(_0696_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1794_ (.A1(_0692_),
    .A2(_0695_),
    .A3(_0696_),
    .B(_0693_),
    .ZN(_0005_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1795_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit29.Q ),
    .A2(_0658_),
    .Z(_0697_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1796_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.LUT_flop ),
    .A2(_0697_),
    .ZN(_0698_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1797_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit28.Q ),
    .A2(_0671_),
    .ZN(_0699_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1798_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit28.Q ),
    .A2(_0671_),
    .B(_0348_),
    .C(_0340_),
    .ZN(_0700_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1799_ (.A1(\Inst_LF_LUT4c_frame_config_dffesr.c_reset_value ),
    .A2(_0699_),
    .ZN(_0701_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1800_ (.A1(_0697_),
    .A2(_0700_),
    .A3(_0701_),
    .B(_0698_),
    .ZN(_0006_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1801_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit7.Q ),
    .A2(_0658_),
    .Z(_0702_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1802_ (.A1(\Inst_LG_LUT4c_frame_config_dffesr.LUT_flop ),
    .A2(_0702_),
    .ZN(_0703_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1803_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit6.Q ),
    .A2(_0671_),
    .ZN(_0704_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1804_ (.A1(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit6.Q ),
    .A2(_0671_),
    .B(_0429_),
    .ZN(_0705_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1805_ (.A1(\Inst_LG_LUT4c_frame_config_dffesr.c_reset_value ),
    .A2(_0704_),
    .ZN(_0706_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1806_ (.A1(_0702_),
    .A2(_0705_),
    .A3(_0706_),
    .B(_0703_),
    .ZN(_0007_),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1807_ (.D(FrameData[24]),
    .E(FrameStrobe[19]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1808_ (.D(FrameData[25]),
    .E(FrameStrobe[19]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1809_ (.D(FrameData[26]),
    .E(FrameStrobe[19]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1810_ (.D(FrameData[27]),
    .E(FrameStrobe[19]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1811_ (.D(FrameData[28]),
    .E(FrameStrobe[19]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1812_ (.D(FrameData[29]),
    .E(FrameStrobe[19]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1813_ (.D(FrameData[30]),
    .E(FrameStrobe[19]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1814_ (.D(FrameData[31]),
    .E(FrameStrobe[19]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1815_ (.D(FrameData[0]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1816_ (.D(FrameData[1]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1817_ (.D(FrameData[2]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1818_ (.D(FrameData[3]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1819_ (.D(FrameData[4]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1820_ (.D(FrameData[5]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1821_ (.D(FrameData[6]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1822_ (.D(FrameData[7]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1823_ (.D(FrameData[8]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.c_out_mux ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1824_ (.D(FrameData[9]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.c_I0mux ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1825_ (.D(FrameData[10]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.c_reset_value ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1826_ (.D(FrameData[11]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1827_ (.D(FrameData[12]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1828_ (.D(FrameData[13]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1829_ (.D(FrameData[14]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1830_ (.D(FrameData[15]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1831_ (.D(FrameData[16]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1832_ (.D(FrameData[17]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1833_ (.D(FrameData[18]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1834_ (.D(FrameData[19]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1835_ (.D(FrameData[20]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1836_ (.D(FrameData[21]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1837_ (.D(FrameData[22]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1838_ (.D(FrameData[23]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1839_ (.D(FrameData[24]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1840_ (.D(FrameData[25]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1841_ (.D(FrameData[26]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1842_ (.D(FrameData[27]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.c_out_mux ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1843_ (.D(FrameData[28]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.c_I0mux ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1844_ (.D(FrameData[29]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.c_reset_value ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1845_ (.D(FrameData[30]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1846_ (.D(FrameData[31]),
    .E(FrameStrobe[18]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1847_ (.D(FrameData[0]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1848_ (.D(FrameData[1]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1849_ (.D(FrameData[2]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1850_ (.D(FrameData[3]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1851_ (.D(FrameData[4]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1852_ (.D(FrameData[5]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1853_ (.D(FrameData[6]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1854_ (.D(FrameData[7]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1855_ (.D(FrameData[8]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1856_ (.D(FrameData[9]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1857_ (.D(FrameData[10]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1858_ (.D(FrameData[11]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1859_ (.D(FrameData[12]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1860_ (.D(FrameData[13]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1861_ (.D(FrameData[14]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.c_out_mux ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1862_ (.D(FrameData[15]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.c_I0mux ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1863_ (.D(FrameData[16]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.c_reset_value ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1864_ (.D(FrameData[17]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1865_ (.D(FrameData[18]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1866_ (.D(FrameData[19]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1867_ (.D(FrameData[20]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1868_ (.D(FrameData[21]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1869_ (.D(FrameData[22]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1870_ (.D(FrameData[23]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1871_ (.D(FrameData[24]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1872_ (.D(FrameData[25]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1873_ (.D(FrameData[26]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1874_ (.D(FrameData[27]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1875_ (.D(FrameData[28]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1876_ (.D(FrameData[29]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1877_ (.D(FrameData[30]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1878_ (.D(FrameData[31]),
    .E(FrameStrobe[17]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1879_ (.D(FrameData[0]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1880_ (.D(FrameData[1]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.c_out_mux ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1881_ (.D(FrameData[2]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.c_I0mux ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1882_ (.D(FrameData[3]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.c_reset_value ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1883_ (.D(FrameData[4]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1884_ (.D(FrameData[5]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1885_ (.D(FrameData[6]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1886_ (.D(FrameData[7]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1887_ (.D(FrameData[8]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1888_ (.D(FrameData[9]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1889_ (.D(FrameData[10]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1890_ (.D(FrameData[11]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1891_ (.D(FrameData[12]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1892_ (.D(FrameData[13]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1893_ (.D(FrameData[14]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1894_ (.D(FrameData[15]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1895_ (.D(FrameData[16]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1896_ (.D(FrameData[17]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1897_ (.D(FrameData[18]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1898_ (.D(FrameData[19]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1899_ (.D(FrameData[20]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.c_out_mux ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1900_ (.D(FrameData[21]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.c_I0mux ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1901_ (.D(FrameData[22]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.c_reset_value ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1902_ (.D(FrameData[23]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1903_ (.D(FrameData[24]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1904_ (.D(FrameData[25]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1905_ (.D(FrameData[26]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1906_ (.D(FrameData[27]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1907_ (.D(FrameData[28]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1908_ (.D(FrameData[29]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1909_ (.D(FrameData[30]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1910_ (.D(FrameData[31]),
    .E(FrameStrobe[16]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1911_ (.D(FrameData[0]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1912_ (.D(FrameData[1]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1913_ (.D(FrameData[2]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1914_ (.D(FrameData[3]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1915_ (.D(FrameData[4]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1916_ (.D(FrameData[5]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1917_ (.D(FrameData[6]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1918_ (.D(FrameData[7]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.c_out_mux ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1919_ (.D(FrameData[8]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.c_I0mux ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1920_ (.D(FrameData[9]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.c_reset_value ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1921_ (.D(FrameData[10]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1922_ (.D(FrameData[11]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1923_ (.D(FrameData[12]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1924_ (.D(FrameData[13]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1925_ (.D(FrameData[14]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1926_ (.D(FrameData[15]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1927_ (.D(FrameData[16]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1928_ (.D(FrameData[17]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1929_ (.D(FrameData[18]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1930_ (.D(FrameData[19]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1931_ (.D(FrameData[20]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1932_ (.D(FrameData[21]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1933_ (.D(FrameData[22]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1934_ (.D(FrameData[23]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1935_ (.D(FrameData[24]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1936_ (.D(FrameData[25]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1937_ (.D(FrameData[26]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.c_out_mux ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1938_ (.D(FrameData[27]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.c_I0mux ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1939_ (.D(FrameData[28]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.c_reset_value ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1940_ (.D(FrameData[29]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1941_ (.D(FrameData[30]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1942_ (.D(FrameData[31]),
    .E(FrameStrobe[15]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1943_ (.D(FrameData[0]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1944_ (.D(FrameData[1]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1945_ (.D(FrameData[2]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1946_ (.D(FrameData[3]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1947_ (.D(FrameData[4]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1948_ (.D(FrameData[5]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1949_ (.D(FrameData[6]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1950_ (.D(FrameData[7]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1951_ (.D(FrameData[8]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1952_ (.D(FrameData[9]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1953_ (.D(FrameData[10]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1954_ (.D(FrameData[11]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1955_ (.D(FrameData[12]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1956_ (.D(FrameData[13]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.c_out_mux ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1957_ (.D(FrameData[14]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.c_I0mux ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1958_ (.D(FrameData[15]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.c_reset_value ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1959_ (.D(FrameData[16]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1960_ (.D(FrameData[17]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1961_ (.D(FrameData[18]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit18.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1962_ (.D(FrameData[19]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit19.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1963_ (.D(FrameData[20]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit20.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1964_ (.D(FrameData[21]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit21.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1965_ (.D(FrameData[22]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit22.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1966_ (.D(FrameData[23]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit23.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1967_ (.D(FrameData[24]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit24.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1968_ (.D(FrameData[25]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit25.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1969_ (.D(FrameData[26]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit26.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1970_ (.D(FrameData[27]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit27.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1971_ (.D(FrameData[28]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit28.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1972_ (.D(FrameData[29]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit29.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1973_ (.D(FrameData[30]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit30.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1974_ (.D(FrameData[31]),
    .E(FrameStrobe[14]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame14_bit31.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1975_ (.D(FrameData[0]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit0.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1976_ (.D(FrameData[1]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit1.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1977_ (.D(FrameData[2]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1978_ (.D(FrameData[3]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1979_ (.D(FrameData[4]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit4.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1980_ (.D(FrameData[5]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1981_ (.D(FrameData[6]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1982_ (.D(FrameData[7]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit7.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1983_ (.D(FrameData[8]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1984_ (.D(FrameData[9]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1985_ (.D(FrameData[10]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit10.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1986_ (.D(FrameData[11]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1987_ (.D(FrameData[12]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit12.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1988_ (.D(FrameData[13]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit13.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1989_ (.D(FrameData[14]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit14.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1990_ (.D(FrameData[15]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit15.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1991_ (.D(FrameData[16]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit16.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1992_ (.D(FrameData[17]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit17.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1993_ (.D(FrameData[18]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit18.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1994_ (.D(FrameData[19]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit19.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1995_ (.D(FrameData[20]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit20.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1996_ (.D(FrameData[21]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit21.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1997_ (.D(FrameData[22]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1998_ (.D(FrameData[23]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _1999_ (.D(FrameData[24]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit24.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2000_ (.D(FrameData[25]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2001_ (.D(FrameData[26]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2002_ (.D(FrameData[27]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit27.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2003_ (.D(FrameData[28]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2004_ (.D(FrameData[29]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2005_ (.D(FrameData[30]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2006_ (.D(FrameData[31]),
    .E(FrameStrobe[13]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2007_ (.D(FrameData[0]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2008_ (.D(FrameData[1]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit1.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2009_ (.D(FrameData[2]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2010_ (.D(FrameData[3]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2011_ (.D(FrameData[4]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2012_ (.D(FrameData[5]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit5.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2013_ (.D(FrameData[6]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2014_ (.D(FrameData[7]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2015_ (.D(FrameData[8]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2016_ (.D(FrameData[9]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit9.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2017_ (.D(FrameData[10]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit10.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2018_ (.D(FrameData[11]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit11.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2019_ (.D(FrameData[12]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit12.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2020_ (.D(FrameData[13]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit13.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2021_ (.D(FrameData[14]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit14.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2022_ (.D(FrameData[15]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit15.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2023_ (.D(FrameData[16]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit16.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2024_ (.D(FrameData[17]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit17.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2025_ (.D(FrameData[18]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit18.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2026_ (.D(FrameData[19]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit19.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2027_ (.D(FrameData[20]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit20.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2028_ (.D(FrameData[21]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit21.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2029_ (.D(FrameData[22]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit22.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2030_ (.D(FrameData[23]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit23.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2031_ (.D(FrameData[24]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit24.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2032_ (.D(FrameData[25]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit25.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2033_ (.D(FrameData[26]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2034_ (.D(FrameData[27]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2035_ (.D(FrameData[28]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2036_ (.D(FrameData[29]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2037_ (.D(FrameData[30]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2038_ (.D(FrameData[31]),
    .E(FrameStrobe[12]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2039_ (.D(FrameData[0]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2040_ (.D(FrameData[1]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2041_ (.D(FrameData[2]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit2.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2042_ (.D(FrameData[3]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2043_ (.D(FrameData[4]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2044_ (.D(FrameData[5]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit5.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2045_ (.D(FrameData[6]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit6.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2046_ (.D(FrameData[7]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit7.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2047_ (.D(FrameData[8]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit8.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2048_ (.D(FrameData[9]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit9.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2049_ (.D(FrameData[10]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit10.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2050_ (.D(FrameData[11]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit11.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2051_ (.D(FrameData[12]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit12.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2052_ (.D(FrameData[13]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit13.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2053_ (.D(FrameData[14]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2054_ (.D(FrameData[15]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2055_ (.D(FrameData[16]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit16.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2056_ (.D(FrameData[17]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2057_ (.D(FrameData[18]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2058_ (.D(FrameData[19]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit19.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2059_ (.D(FrameData[20]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2060_ (.D(FrameData[21]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2061_ (.D(FrameData[22]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit22.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2062_ (.D(FrameData[23]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2063_ (.D(FrameData[24]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit24.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2064_ (.D(FrameData[25]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit25.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2065_ (.D(FrameData[26]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2066_ (.D(FrameData[27]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2067_ (.D(FrameData[28]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2068_ (.D(FrameData[29]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit29.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2069_ (.D(FrameData[30]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2070_ (.D(FrameData[31]),
    .E(FrameStrobe[11]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2071_ (.D(FrameData[0]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2072_ (.D(FrameData[1]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2073_ (.D(FrameData[2]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit2.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2074_ (.D(FrameData[3]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit3.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2075_ (.D(FrameData[4]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit4.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2076_ (.D(FrameData[5]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit5.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2077_ (.D(FrameData[6]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2078_ (.D(FrameData[7]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit7.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2079_ (.D(FrameData[8]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit8.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2080_ (.D(FrameData[9]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2081_ (.D(FrameData[10]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit10.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2082_ (.D(FrameData[11]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit11.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2083_ (.D(FrameData[12]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2084_ (.D(FrameData[13]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit13.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2085_ (.D(FrameData[14]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit14.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2086_ (.D(FrameData[15]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit15.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2087_ (.D(FrameData[16]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit16.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2088_ (.D(FrameData[17]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit17.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2089_ (.D(FrameData[18]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit18.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2090_ (.D(FrameData[19]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2091_ (.D(FrameData[20]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit20.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2092_ (.D(FrameData[21]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit21.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2093_ (.D(FrameData[22]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2094_ (.D(FrameData[23]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2095_ (.D(FrameData[24]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit24.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2096_ (.D(FrameData[25]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit25.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2097_ (.D(FrameData[26]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit26.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2098_ (.D(FrameData[27]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit27.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2099_ (.D(FrameData[28]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2100_ (.D(FrameData[29]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2101_ (.D(FrameData[30]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit30.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2102_ (.D(FrameData[31]),
    .E(FrameStrobe[10]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame10_bit31.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2103_ (.D(FrameData[0]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2104_ (.D(FrameData[1]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2105_ (.D(FrameData[2]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit2.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2106_ (.D(FrameData[3]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit3.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2107_ (.D(FrameData[4]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit4.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2108_ (.D(FrameData[5]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit5.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2109_ (.D(FrameData[6]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit6.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2110_ (.D(FrameData[7]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit7.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2111_ (.D(FrameData[8]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit8.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2112_ (.D(FrameData[9]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit9.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2113_ (.D(FrameData[10]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit10.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2114_ (.D(FrameData[11]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2115_ (.D(FrameData[12]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit12.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2116_ (.D(FrameData[13]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit13.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2117_ (.D(FrameData[14]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit14.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2118_ (.D(FrameData[15]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2119_ (.D(FrameData[16]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2120_ (.D(FrameData[17]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2121_ (.D(FrameData[18]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit18.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2122_ (.D(FrameData[19]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit19.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2123_ (.D(FrameData[20]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit20.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2124_ (.D(FrameData[21]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2125_ (.D(FrameData[22]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit22.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2126_ (.D(FrameData[23]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit23.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2127_ (.D(FrameData[24]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit24.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2128_ (.D(FrameData[25]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2129_ (.D(FrameData[26]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2130_ (.D(FrameData[27]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2131_ (.D(FrameData[28]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit28.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2132_ (.D(FrameData[29]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit29.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2133_ (.D(FrameData[30]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2134_ (.D(FrameData[31]),
    .E(FrameStrobe[9]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame9_bit31.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2135_ (.D(FrameData[0]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit0.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2136_ (.D(FrameData[1]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit1.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2137_ (.D(FrameData[2]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit2.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2138_ (.D(FrameData[3]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit3.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2139_ (.D(FrameData[4]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit4.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2140_ (.D(FrameData[5]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit5.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2141_ (.D(FrameData[6]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit6.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2142_ (.D(FrameData[7]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit7.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2143_ (.D(FrameData[8]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2144_ (.D(FrameData[9]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2145_ (.D(FrameData[10]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit10.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2146_ (.D(FrameData[11]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit11.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2147_ (.D(FrameData[12]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit12.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2148_ (.D(FrameData[13]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit13.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2149_ (.D(FrameData[14]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit14.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2150_ (.D(FrameData[15]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit15.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2151_ (.D(FrameData[16]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit16.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2152_ (.D(FrameData[17]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit17.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2153_ (.D(FrameData[18]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit18.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2154_ (.D(FrameData[19]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit19.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2155_ (.D(FrameData[20]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2156_ (.D(FrameData[21]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit21.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2157_ (.D(FrameData[22]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit22.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2158_ (.D(FrameData[23]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit23.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2159_ (.D(FrameData[24]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2160_ (.D(FrameData[25]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2161_ (.D(FrameData[26]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit26.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2162_ (.D(FrameData[27]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit27.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2163_ (.D(FrameData[28]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit28.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2164_ (.D(FrameData[29]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit29.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2165_ (.D(FrameData[30]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2166_ (.D(FrameData[31]),
    .E(FrameStrobe[8]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2167_ (.D(FrameData[0]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2168_ (.D(FrameData[1]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit1.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2169_ (.D(FrameData[2]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit2.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2170_ (.D(FrameData[3]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit3.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2171_ (.D(FrameData[4]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit4.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2172_ (.D(FrameData[5]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit5.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2173_ (.D(FrameData[6]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2174_ (.D(FrameData[7]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2175_ (.D(FrameData[8]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2176_ (.D(FrameData[9]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit9.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2177_ (.D(FrameData[10]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2178_ (.D(FrameData[11]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit11.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2179_ (.D(FrameData[12]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2180_ (.D(FrameData[13]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit13.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2181_ (.D(FrameData[14]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit14.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2182_ (.D(FrameData[15]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit15.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2183_ (.D(FrameData[16]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit16.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2184_ (.D(FrameData[17]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit17.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2185_ (.D(FrameData[18]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2186_ (.D(FrameData[19]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit19.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2187_ (.D(FrameData[20]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit20.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2188_ (.D(FrameData[21]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit21.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2189_ (.D(FrameData[22]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2190_ (.D(FrameData[23]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit23.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2191_ (.D(FrameData[24]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2192_ (.D(FrameData[25]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit25.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2193_ (.D(FrameData[26]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit26.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2194_ (.D(FrameData[27]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit27.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2195_ (.D(FrameData[28]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit28.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2196_ (.D(FrameData[29]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit29.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2197_ (.D(FrameData[30]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit30.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2198_ (.D(FrameData[31]),
    .E(FrameStrobe[7]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame7_bit31.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2199_ (.D(FrameData[0]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2200_ (.D(FrameData[1]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit1.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2201_ (.D(FrameData[2]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit2.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2202_ (.D(FrameData[3]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit3.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2203_ (.D(FrameData[4]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit4.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2204_ (.D(FrameData[5]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit5.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2205_ (.D(FrameData[6]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit6.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2206_ (.D(FrameData[7]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit7.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2207_ (.D(FrameData[8]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit8.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2208_ (.D(FrameData[9]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit9.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2209_ (.D(FrameData[10]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2210_ (.D(FrameData[11]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit11.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2211_ (.D(FrameData[12]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit12.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2212_ (.D(FrameData[13]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit13.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2213_ (.D(FrameData[14]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit14.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2214_ (.D(FrameData[15]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit15.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2215_ (.D(FrameData[16]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2216_ (.D(FrameData[17]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit17.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2217_ (.D(FrameData[18]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2218_ (.D(FrameData[19]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit19.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2219_ (.D(FrameData[20]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit20.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2220_ (.D(FrameData[21]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit21.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2221_ (.D(FrameData[22]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2222_ (.D(FrameData[23]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit23.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2223_ (.D(FrameData[24]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2224_ (.D(FrameData[25]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit25.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2225_ (.D(FrameData[26]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit26.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2226_ (.D(FrameData[27]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit27.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2227_ (.D(FrameData[28]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit28.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2228_ (.D(FrameData[29]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit29.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2229_ (.D(FrameData[30]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit30.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2230_ (.D(FrameData[31]),
    .E(FrameStrobe[6]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame6_bit31.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2231_ (.D(FrameData[0]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit0.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2232_ (.D(FrameData[1]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit1.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2233_ (.D(FrameData[2]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit2.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2234_ (.D(FrameData[3]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit3.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2235_ (.D(FrameData[4]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit4.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2236_ (.D(FrameData[5]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit5.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2237_ (.D(FrameData[6]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit6.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2238_ (.D(FrameData[7]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit7.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2239_ (.D(FrameData[8]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2240_ (.D(FrameData[9]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit9.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2241_ (.D(FrameData[10]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit10.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2242_ (.D(FrameData[11]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit11.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2243_ (.D(FrameData[12]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2244_ (.D(FrameData[13]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit13.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2245_ (.D(FrameData[14]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2246_ (.D(FrameData[15]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit15.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2247_ (.D(FrameData[16]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit16.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2248_ (.D(FrameData[17]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit17.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2249_ (.D(FrameData[18]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit18.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2250_ (.D(FrameData[19]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit19.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2251_ (.D(FrameData[20]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit20.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2252_ (.D(FrameData[21]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit21.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2253_ (.D(FrameData[22]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit22.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2254_ (.D(FrameData[23]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit23.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2255_ (.D(FrameData[24]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit24.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2256_ (.D(FrameData[25]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit25.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2257_ (.D(FrameData[26]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2258_ (.D(FrameData[27]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2259_ (.D(FrameData[28]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2260_ (.D(FrameData[29]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2261_ (.D(FrameData[30]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2262_ (.D(FrameData[31]),
    .E(FrameStrobe[5]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2263_ (.D(FrameData[0]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2264_ (.D(FrameData[1]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2265_ (.D(FrameData[2]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2266_ (.D(FrameData[3]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2267_ (.D(FrameData[4]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2268_ (.D(FrameData[5]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2269_ (.D(FrameData[6]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2270_ (.D(FrameData[7]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2271_ (.D(FrameData[8]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2272_ (.D(FrameData[9]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2273_ (.D(FrameData[10]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2274_ (.D(FrameData[11]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2275_ (.D(FrameData[12]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2276_ (.D(FrameData[13]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2277_ (.D(FrameData[14]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2278_ (.D(FrameData[15]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2279_ (.D(FrameData[16]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2280_ (.D(FrameData[17]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2281_ (.D(FrameData[18]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2282_ (.D(FrameData[19]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2283_ (.D(FrameData[20]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2284_ (.D(FrameData[21]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2285_ (.D(FrameData[22]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2286_ (.D(FrameData[23]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2287_ (.D(FrameData[24]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2288_ (.D(FrameData[25]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2289_ (.D(FrameData[26]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2290_ (.D(FrameData[27]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2291_ (.D(FrameData[28]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2292_ (.D(FrameData[29]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2293_ (.D(FrameData[30]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2294_ (.D(FrameData[31]),
    .E(FrameStrobe[4]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2295_ (.D(FrameData[0]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2296_ (.D(FrameData[1]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2297_ (.D(FrameData[2]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2298_ (.D(FrameData[3]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2299_ (.D(FrameData[4]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2300_ (.D(FrameData[5]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2301_ (.D(FrameData[6]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2302_ (.D(FrameData[7]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2303_ (.D(FrameData[8]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2304_ (.D(FrameData[9]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit9.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2305_ (.D(FrameData[10]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2306_ (.D(FrameData[11]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2307_ (.D(FrameData[12]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2308_ (.D(FrameData[13]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2309_ (.D(FrameData[14]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2310_ (.D(FrameData[15]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2311_ (.D(FrameData[16]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2312_ (.D(FrameData[17]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2313_ (.D(FrameData[18]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2314_ (.D(FrameData[19]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2315_ (.D(FrameData[20]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2316_ (.D(FrameData[21]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2317_ (.D(FrameData[22]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2318_ (.D(FrameData[23]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2319_ (.D(FrameData[24]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2320_ (.D(FrameData[25]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2321_ (.D(FrameData[26]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2322_ (.D(FrameData[27]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2323_ (.D(FrameData[28]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2324_ (.D(FrameData[29]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2325_ (.D(FrameData[30]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2326_ (.D(FrameData[31]),
    .E(FrameStrobe[3]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2327_ (.D(FrameData[0]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2328_ (.D(FrameData[1]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2329_ (.D(FrameData[2]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2330_ (.D(FrameData[3]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2331_ (.D(FrameData[4]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2332_ (.D(FrameData[5]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit5.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2333_ (.D(FrameData[6]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2334_ (.D(FrameData[7]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2335_ (.D(FrameData[8]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2336_ (.D(FrameData[9]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2337_ (.D(FrameData[10]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2338_ (.D(FrameData[11]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2339_ (.D(FrameData[12]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2340_ (.D(FrameData[13]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit13.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2341_ (.D(FrameData[14]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2342_ (.D(FrameData[15]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2343_ (.D(FrameData[16]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2344_ (.D(FrameData[17]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2345_ (.D(FrameData[18]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2346_ (.D(FrameData[19]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2347_ (.D(FrameData[20]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2348_ (.D(FrameData[21]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2349_ (.D(FrameData[22]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2350_ (.D(FrameData[23]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2351_ (.D(FrameData[24]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2352_ (.D(FrameData[25]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2353_ (.D(FrameData[26]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2354_ (.D(FrameData[27]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2355_ (.D(FrameData[28]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2356_ (.D(FrameData[29]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2357_ (.D(FrameData[30]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2358_ (.D(FrameData[31]),
    .E(FrameStrobe[2]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2359_ (.D(FrameData[0]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2360_ (.D(FrameData[1]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2361_ (.D(FrameData[2]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2362_ (.D(FrameData[3]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2363_ (.D(FrameData[4]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2364_ (.D(FrameData[5]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2365_ (.D(FrameData[6]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2366_ (.D(FrameData[7]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2367_ (.D(FrameData[8]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2368_ (.D(FrameData[9]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2369_ (.D(FrameData[10]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2370_ (.D(FrameData[11]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2371_ (.D(FrameData[12]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2372_ (.D(FrameData[13]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2373_ (.D(FrameData[14]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2374_ (.D(FrameData[15]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2375_ (.D(FrameData[16]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2376_ (.D(FrameData[17]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2377_ (.D(FrameData[18]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2378_ (.D(FrameData[19]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2379_ (.D(FrameData[20]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2380_ (.D(FrameData[21]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2381_ (.D(FrameData[22]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2382_ (.D(FrameData[23]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2383_ (.D(FrameData[24]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2384_ (.D(FrameData[25]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2385_ (.D(FrameData[26]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit26.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2386_ (.D(FrameData[27]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit27.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2387_ (.D(FrameData[28]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit28.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2388_ (.D(FrameData[29]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit29.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2389_ (.D(FrameData[30]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2390_ (.D(FrameData[31]),
    .E(FrameStrobe[1]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame1_bit31.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2391_ (.D(FrameData[0]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit0.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2392_ (.D(FrameData[1]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit1.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2393_ (.D(FrameData[2]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2394_ (.D(FrameData[3]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit3.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2395_ (.D(FrameData[4]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit4.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2396_ (.D(FrameData[5]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit5.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2397_ (.D(FrameData[6]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit6.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2398_ (.D(FrameData[7]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit7.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2399_ (.D(FrameData[8]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2400_ (.D(FrameData[9]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit9.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2401_ (.D(FrameData[10]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit10.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2402_ (.D(FrameData[11]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit11.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2403_ (.D(FrameData[12]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2404_ (.D(FrameData[13]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit13.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2405_ (.D(FrameData[14]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit14.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2406_ (.D(FrameData[15]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit15.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2407_ (.D(FrameData[16]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit16.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2408_ (.D(FrameData[17]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit17.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2409_ (.D(FrameData[18]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit18.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2410_ (.D(FrameData[19]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit19.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2411_ (.D(FrameData[20]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit20.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2412_ (.D(FrameData[21]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit21.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2413_ (.D(FrameData[22]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2414_ (.D(FrameData[23]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit23.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2415_ (.D(FrameData[24]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit24.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2416_ (.D(FrameData[25]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit25.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2417_ (.D(FrameData[26]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2418_ (.D(FrameData[27]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2419_ (.D(FrameData[28]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2420_ (.D(FrameData[29]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2421_ (.D(FrameData[30]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__latq_1 _2422_ (.D(FrameData[31]),
    .E(FrameStrobe[0]),
    .Q(\Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2423_ (.D(_0000_),
    .CLK(clknet_1_1__leaf_UserCLK_regs),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.LUT_flop ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2424_ (.D(_0001_),
    .CLK(clknet_1_0__leaf_UserCLK_regs),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.LUT_flop ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2425_ (.D(_0002_),
    .CLK(clknet_1_0__leaf_UserCLK_regs),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.LUT_flop ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2426_ (.D(_0003_),
    .CLK(clknet_1_0__leaf_UserCLK_regs),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.LUT_flop ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2427_ (.D(_0004_),
    .CLK(clknet_1_0__leaf_UserCLK_regs),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.LUT_flop ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2428_ (.D(_0005_),
    .CLK(clknet_1_1__leaf_UserCLK_regs),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.LUT_flop ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2429_ (.D(_0006_),
    .CLK(clknet_1_1__leaf_UserCLK_regs),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.LUT_flop ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2430_ (.D(_0007_),
    .CLK(clknet_1_1__leaf_UserCLK_regs),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.LUT_flop ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2431_ (.I(\Inst_LUT4AB_switch_matrix.E1BEG0 ),
    .Z(net2),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2432_ (.I(\Inst_LUT4AB_switch_matrix.E1BEG1 ),
    .Z(net3),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2433_ (.I(\Inst_LUT4AB_switch_matrix.E1BEG2 ),
    .Z(net4),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2434_ (.I(\Inst_LUT4AB_switch_matrix.E1BEG3 ),
    .Z(net5),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2435_ (.I(\Inst_LUT4AB_switch_matrix.E2BEG0 ),
    .Z(net6),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2436_ (.I(\Inst_LUT4AB_switch_matrix.E2BEG1 ),
    .Z(net7),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2437_ (.I(\Inst_LUT4AB_switch_matrix.E2BEG2 ),
    .Z(net8),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2438_ (.I(\Inst_LUT4AB_switch_matrix.E2BEG3 ),
    .Z(net9),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2439_ (.I(\Inst_LUT4AB_switch_matrix.E2BEG4 ),
    .Z(net10),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2440_ (.I(\Inst_LUT4AB_switch_matrix.E2BEG5 ),
    .Z(net11),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2441_ (.I(\Inst_LUT4AB_switch_matrix.E2BEG6 ),
    .Z(net12),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2442_ (.I(\Inst_LUT4AB_switch_matrix.E2BEG7 ),
    .Z(net13),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2443_ (.I(E2MID[0]),
    .Z(net14),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2444_ (.I(E2MID[1]),
    .Z(net15),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2445_ (.I(E2MID[2]),
    .Z(net16),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2446_ (.I(E2MID[3]),
    .Z(net17),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2447_ (.I(E2MID[4]),
    .Z(net18),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2448_ (.I(E2MID[5]),
    .Z(net19),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2449_ (.I(E2MID[6]),
    .Z(net20),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2450_ (.I(E2MID[7]),
    .Z(net21),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2451_ (.I(E6END[2]),
    .Z(net22),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2452_ (.I(E6END[3]),
    .Z(net25),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2453_ (.I(E6END[4]),
    .Z(net26),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2454_ (.I(E6END[5]),
    .Z(net27),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2455_ (.I(E6END[6]),
    .Z(net28),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2456_ (.I(E6END[7]),
    .Z(net29),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2457_ (.I(E6END[8]),
    .Z(net30),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2458_ (.I(E6END[9]),
    .Z(net31),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2459_ (.I(E6END[10]),
    .Z(net32),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2460_ (.I(E6END[11]),
    .Z(net33),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2461_ (.I(\Inst_LUT4AB_switch_matrix.E6BEG0 ),
    .Z(net23),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2462_ (.I(\Inst_LUT4AB_switch_matrix.E6BEG1 ),
    .Z(net24),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2463_ (.I(EE4END[4]),
    .Z(net34),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2464_ (.I(EE4END[5]),
    .Z(net41),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2465_ (.I(EE4END[6]),
    .Z(net42),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2466_ (.I(EE4END[7]),
    .Z(net43),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2467_ (.I(EE4END[8]),
    .Z(net44),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2468_ (.I(EE4END[9]),
    .Z(net45),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2469_ (.I(EE4END[10]),
    .Z(net46),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2470_ (.I(EE4END[11]),
    .Z(net47),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2471_ (.I(EE4END[12]),
    .Z(net48),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2472_ (.I(EE4END[13]),
    .Z(net49),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2473_ (.I(EE4END[14]),
    .Z(net35),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2474_ (.I(EE4END[15]),
    .Z(net36),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2475_ (.I(\Inst_LUT4AB_switch_matrix.EE4BEG0 ),
    .Z(net37),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2476_ (.I(\Inst_LUT4AB_switch_matrix.EE4BEG1 ),
    .Z(net38),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2477_ (.I(\Inst_LUT4AB_switch_matrix.EE4BEG2 ),
    .Z(net39),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2478_ (.I(\Inst_LUT4AB_switch_matrix.EE4BEG3 ),
    .Z(net40),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2479_ (.I(FrameData[0]),
    .Z(net50),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2480_ (.I(FrameData[1]),
    .Z(net61),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2481_ (.I(FrameData[2]),
    .Z(net72),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2482_ (.I(FrameData[3]),
    .Z(net75),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2483_ (.I(FrameData[4]),
    .Z(net76),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2484_ (.I(FrameData[5]),
    .Z(net77),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2485_ (.I(FrameData[6]),
    .Z(net78),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2486_ (.I(FrameData[7]),
    .Z(net79),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2487_ (.I(FrameData[8]),
    .Z(net80),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2488_ (.I(FrameData[9]),
    .Z(net81),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2489_ (.I(FrameData[10]),
    .Z(net51),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2490_ (.I(FrameData[11]),
    .Z(net52),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2491_ (.I(FrameData[12]),
    .Z(net53),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2492_ (.I(FrameData[13]),
    .Z(net54),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2493_ (.I(FrameData[14]),
    .Z(net55),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2494_ (.I(FrameData[15]),
    .Z(net56),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2495_ (.I(FrameData[16]),
    .Z(net57),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2496_ (.I(FrameData[17]),
    .Z(net58),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2497_ (.I(FrameData[18]),
    .Z(net59),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2498_ (.I(FrameData[19]),
    .Z(net60),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2499_ (.I(FrameData[20]),
    .Z(net62),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2500_ (.I(FrameData[21]),
    .Z(net63),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2501_ (.I(FrameData[22]),
    .Z(net64),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2502_ (.I(FrameData[23]),
    .Z(net65),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2503_ (.I(FrameData[24]),
    .Z(net66),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2504_ (.I(FrameData[25]),
    .Z(net67),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2505_ (.I(FrameData[26]),
    .Z(net68),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2506_ (.I(FrameData[27]),
    .Z(net69),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2507_ (.I(FrameData[28]),
    .Z(net70),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2508_ (.I(FrameData[29]),
    .Z(net71),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2509_ (.I(FrameData[30]),
    .Z(net73),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2510_ (.I(FrameData[31]),
    .Z(net74),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2511_ (.I(FrameStrobe[0]),
    .Z(net82),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2512_ (.I(FrameStrobe[1]),
    .Z(net93),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2513_ (.I(FrameStrobe[2]),
    .Z(net94),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2514_ (.I(FrameStrobe[3]),
    .Z(net95),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2515_ (.I(FrameStrobe[4]),
    .Z(net96),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2516_ (.I(FrameStrobe[5]),
    .Z(net97),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2517_ (.I(FrameStrobe[6]),
    .Z(net98),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2518_ (.I(FrameStrobe[7]),
    .Z(net99),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2519_ (.I(FrameStrobe[8]),
    .Z(net100),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2520_ (.I(FrameStrobe[9]),
    .Z(net101),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2521_ (.I(FrameStrobe[10]),
    .Z(net83),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2522_ (.I(FrameStrobe[11]),
    .Z(net84),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2523_ (.I(FrameStrobe[12]),
    .Z(net85),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2524_ (.I(FrameStrobe[13]),
    .Z(net86),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2525_ (.I(FrameStrobe[14]),
    .Z(net87),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2526_ (.I(FrameStrobe[15]),
    .Z(net88),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2527_ (.I(FrameStrobe[16]),
    .Z(net89),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2528_ (.I(FrameStrobe[17]),
    .Z(net90),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2529_ (.I(FrameStrobe[18]),
    .Z(net91),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2530_ (.I(FrameStrobe[19]),
    .Z(net92),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2531_ (.I(\Inst_LUT4AB_switch_matrix.N1BEG0 ),
    .Z(net102),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2532_ (.I(\Inst_LUT4AB_switch_matrix.N1BEG1 ),
    .Z(net103),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2533_ (.I(\Inst_LUT4AB_switch_matrix.N1BEG2 ),
    .Z(net104),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2534_ (.I(\Inst_LUT4AB_switch_matrix.N1BEG3 ),
    .Z(net105),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2535_ (.I(\Inst_LUT4AB_switch_matrix.JN2BEG0 ),
    .Z(net106),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2536_ (.I(\Inst_LUT4AB_switch_matrix.JN2BEG1 ),
    .Z(net107),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2537_ (.I(\Inst_LUT4AB_switch_matrix.JN2BEG2 ),
    .Z(net108),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2538_ (.I(\Inst_LUT4AB_switch_matrix.JN2BEG3 ),
    .Z(net109),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2539_ (.I(\Inst_LUT4AB_switch_matrix.JN2BEG4 ),
    .Z(net110),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2540_ (.I(\Inst_LUT4AB_switch_matrix.JN2BEG5 ),
    .Z(net111),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2541_ (.I(\Inst_LUT4AB_switch_matrix.JN2BEG6 ),
    .Z(net112),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2542_ (.I(\Inst_LUT4AB_switch_matrix.JN2BEG7 ),
    .Z(net113),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2543_ (.I(N2MID[0]),
    .Z(net114),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2544_ (.I(N2MID[1]),
    .Z(net115),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2545_ (.I(N2MID[2]),
    .Z(net116),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2546_ (.I(N2MID[3]),
    .Z(net117),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2547_ (.I(N2MID[4]),
    .Z(net118),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2548_ (.I(N2MID[5]),
    .Z(net119),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2549_ (.I(N2MID[6]),
    .Z(net120),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2550_ (.I(N2MID[7]),
    .Z(net121),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2551_ (.I(N4END[4]),
    .Z(net122),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2552_ (.I(N4END[5]),
    .Z(net129),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2553_ (.I(N4END[6]),
    .Z(net130),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2554_ (.I(N4END[7]),
    .Z(net131),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2555_ (.I(N4END[8]),
    .Z(net132),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2556_ (.I(N4END[9]),
    .Z(net133),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2557_ (.I(N4END[10]),
    .Z(net134),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2558_ (.I(N4END[11]),
    .Z(net135),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2559_ (.I(N4END[12]),
    .Z(net136),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2560_ (.I(N4END[13]),
    .Z(net137),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2561_ (.I(N4END[14]),
    .Z(net123),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2562_ (.I(N4END[15]),
    .Z(net124),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2563_ (.I(\Inst_LUT4AB_switch_matrix.N4BEG0 ),
    .Z(net125),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2564_ (.I(\Inst_LUT4AB_switch_matrix.N4BEG1 ),
    .Z(net126),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2565_ (.I(\Inst_LUT4AB_switch_matrix.N4BEG2 ),
    .Z(net127),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2566_ (.I(\Inst_LUT4AB_switch_matrix.N4BEG3 ),
    .Z(net128),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2567_ (.I(NN4END[4]),
    .Z(net138),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2568_ (.I(NN4END[5]),
    .Z(net145),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2569_ (.I(NN4END[6]),
    .Z(net146),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2570_ (.I(NN4END[7]),
    .Z(net147),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2571_ (.I(NN4END[8]),
    .Z(net148),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2572_ (.I(NN4END[9]),
    .Z(net149),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2573_ (.I(NN4END[10]),
    .Z(net150),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2574_ (.I(NN4END[11]),
    .Z(net151),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2575_ (.I(NN4END[12]),
    .Z(net152),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2576_ (.I(NN4END[13]),
    .Z(net153),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2577_ (.I(NN4END[14]),
    .Z(net139),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2578_ (.I(NN4END[15]),
    .Z(net140),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2579_ (.I(\Inst_LUT4AB_switch_matrix.NN4BEG0 ),
    .Z(net141),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2580_ (.I(\Inst_LUT4AB_switch_matrix.NN4BEG1 ),
    .Z(net142),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2581_ (.I(\Inst_LUT4AB_switch_matrix.NN4BEG2 ),
    .Z(net143),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2582_ (.I(\Inst_LUT4AB_switch_matrix.NN4BEG3 ),
    .Z(net144),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2583_ (.I(\Inst_LUT4AB_switch_matrix.S1BEG0 ),
    .Z(net154),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2584_ (.I(\Inst_LUT4AB_switch_matrix.S1BEG1 ),
    .Z(net155),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2585_ (.I(\Inst_LUT4AB_switch_matrix.S1BEG2 ),
    .Z(net156),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2586_ (.I(\Inst_LUT4AB_switch_matrix.S1BEG3 ),
    .Z(net157),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2587_ (.I(\Inst_LUT4AB_switch_matrix.JS2BEG0 ),
    .Z(net158),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2588_ (.I(\Inst_LUT4AB_switch_matrix.JS2BEG1 ),
    .Z(net159),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2589_ (.I(\Inst_LUT4AB_switch_matrix.JS2BEG2 ),
    .Z(net160),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2590_ (.I(\Inst_LUT4AB_switch_matrix.JS2BEG3 ),
    .Z(net161),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2591_ (.I(\Inst_LUT4AB_switch_matrix.JS2BEG4 ),
    .Z(net162),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2592_ (.I(\Inst_LUT4AB_switch_matrix.JS2BEG5 ),
    .Z(net163),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2593_ (.I(\Inst_LUT4AB_switch_matrix.JS2BEG6 ),
    .Z(net164),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2594_ (.I(\Inst_LUT4AB_switch_matrix.JS2BEG7 ),
    .Z(net165),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2595_ (.I(S2MID[0]),
    .Z(net166),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2596_ (.I(S2MID[1]),
    .Z(net167),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2597_ (.I(S2MID[2]),
    .Z(net168),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2598_ (.I(S2MID[3]),
    .Z(net169),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2599_ (.I(S2MID[4]),
    .Z(net170),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2600_ (.I(S2MID[5]),
    .Z(net171),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2601_ (.I(S2MID[6]),
    .Z(net172),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2602_ (.I(S2MID[7]),
    .Z(net173),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2603_ (.I(S4END[4]),
    .Z(net174),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2604_ (.I(S4END[5]),
    .Z(net181),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2605_ (.I(S4END[6]),
    .Z(net182),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2606_ (.I(S4END[7]),
    .Z(net183),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2607_ (.I(S4END[8]),
    .Z(net184),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2608_ (.I(S4END[9]),
    .Z(net185),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2609_ (.I(S4END[10]),
    .Z(net186),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2610_ (.I(S4END[11]),
    .Z(net187),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2611_ (.I(S4END[12]),
    .Z(net188),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2612_ (.I(S4END[13]),
    .Z(net189),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2613_ (.I(S4END[14]),
    .Z(net175),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2614_ (.I(S4END[15]),
    .Z(net176),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2615_ (.I(\Inst_LUT4AB_switch_matrix.S4BEG0 ),
    .Z(net177),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2616_ (.I(\Inst_LUT4AB_switch_matrix.S4BEG1 ),
    .Z(net178),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2617_ (.I(\Inst_LUT4AB_switch_matrix.S4BEG2 ),
    .Z(net179),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2618_ (.I(\Inst_LUT4AB_switch_matrix.S4BEG3 ),
    .Z(net180),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2619_ (.I(SS4END[4]),
    .Z(net190),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2620_ (.I(SS4END[5]),
    .Z(net197),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2621_ (.I(SS4END[6]),
    .Z(net198),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2622_ (.I(SS4END[7]),
    .Z(net199),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2623_ (.I(SS4END[8]),
    .Z(net200),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2624_ (.I(SS4END[9]),
    .Z(net201),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2625_ (.I(SS4END[10]),
    .Z(net202),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2626_ (.I(SS4END[11]),
    .Z(net203),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2627_ (.I(SS4END[12]),
    .Z(net204),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2628_ (.I(SS4END[13]),
    .Z(net205),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2629_ (.I(SS4END[14]),
    .Z(net191),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2630_ (.I(SS4END[15]),
    .Z(net192),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2631_ (.I(\Inst_LUT4AB_switch_matrix.SS4BEG0 ),
    .Z(net193),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2632_ (.I(\Inst_LUT4AB_switch_matrix.SS4BEG1 ),
    .Z(net194),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2633_ (.I(\Inst_LUT4AB_switch_matrix.SS4BEG2 ),
    .Z(net195),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2634_ (.I(\Inst_LUT4AB_switch_matrix.SS4BEG3 ),
    .Z(net196),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2635_ (.I(clknet_1_0__leaf_UserCLK),
    .Z(net206),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2636_ (.I(\Inst_LUT4AB_switch_matrix.W1BEG0 ),
    .Z(net207),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2637_ (.I(\Inst_LUT4AB_switch_matrix.W1BEG1 ),
    .Z(net208),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2638_ (.I(\Inst_LUT4AB_switch_matrix.W1BEG2 ),
    .Z(net209),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2639_ (.I(\Inst_LUT4AB_switch_matrix.W1BEG3 ),
    .Z(net210),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2640_ (.I(\Inst_LUT4AB_switch_matrix.JW2BEG0 ),
    .Z(net211),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2641_ (.I(\Inst_LUT4AB_switch_matrix.JW2BEG1 ),
    .Z(net212),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2642_ (.I(\Inst_LUT4AB_switch_matrix.JW2BEG2 ),
    .Z(net213),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2643_ (.I(\Inst_LUT4AB_switch_matrix.JW2BEG3 ),
    .Z(net214),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2644_ (.I(\Inst_LUT4AB_switch_matrix.JW2BEG4 ),
    .Z(net215),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2645_ (.I(\Inst_LUT4AB_switch_matrix.JW2BEG5 ),
    .Z(net216),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2646_ (.I(\Inst_LUT4AB_switch_matrix.JW2BEG6 ),
    .Z(net217),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2647_ (.I(\Inst_LUT4AB_switch_matrix.JW2BEG7 ),
    .Z(net218),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2648_ (.I(W2MID[0]),
    .Z(net219),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2649_ (.I(W2MID[1]),
    .Z(net220),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2650_ (.I(W2MID[2]),
    .Z(net221),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2651_ (.I(W2MID[3]),
    .Z(net222),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2652_ (.I(W2MID[4]),
    .Z(net223),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2653_ (.I(W2MID[5]),
    .Z(net224),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2654_ (.I(W2MID[6]),
    .Z(net225),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2655_ (.I(W2MID[7]),
    .Z(net226),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2656_ (.I(W6END[2]),
    .Z(net227),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2657_ (.I(W6END[3]),
    .Z(net230),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2658_ (.I(W6END[4]),
    .Z(net231),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2659_ (.I(W6END[5]),
    .Z(net232),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2660_ (.I(W6END[6]),
    .Z(net233),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2661_ (.I(W6END[7]),
    .Z(net234),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2662_ (.I(W6END[8]),
    .Z(net235),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2663_ (.I(W6END[9]),
    .Z(net236),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2664_ (.I(W6END[10]),
    .Z(net237),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2665_ (.I(W6END[11]),
    .Z(net238),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2666_ (.I(\Inst_LUT4AB_switch_matrix.W6BEG0 ),
    .Z(net228),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2667_ (.I(\Inst_LUT4AB_switch_matrix.W6BEG1 ),
    .Z(net229),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2668_ (.I(WW4END[4]),
    .Z(net239),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2669_ (.I(WW4END[5]),
    .Z(net246),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2670_ (.I(WW4END[6]),
    .Z(net247),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2671_ (.I(WW4END[7]),
    .Z(net248),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2672_ (.I(WW4END[8]),
    .Z(net249),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2673_ (.I(WW4END[9]),
    .Z(net250),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2674_ (.I(WW4END[10]),
    .Z(net251),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2675_ (.I(WW4END[11]),
    .Z(net252),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2676_ (.I(WW4END[12]),
    .Z(net253),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2677_ (.I(WW4END[13]),
    .Z(net254),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2678_ (.I(WW4END[14]),
    .Z(net240),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2679_ (.I(WW4END[15]),
    .Z(net241),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2680_ (.I(\Inst_LUT4AB_switch_matrix.WW4BEG0 ),
    .Z(net242),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2681_ (.I(\Inst_LUT4AB_switch_matrix.WW4BEG1 ),
    .Z(net243),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2682_ (.I(\Inst_LUT4AB_switch_matrix.WW4BEG2 ),
    .Z(net244),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2683_ (.I(\Inst_LUT4AB_switch_matrix.WW4BEG3 ),
    .Z(net245),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Right_62 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Right_63 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Right_64 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Right_65 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Right_66 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Right_67 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Right_68 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Right_69 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Right_70 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_71 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_72 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_73 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_74 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_75 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_76 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_77 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_78 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_79 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_80 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_81 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_82 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_83 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_84 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_85 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_86 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_87 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_88 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_89 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_90 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_91 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_92 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_93 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_94 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_95 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_96 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_97 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_98 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_99 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_100 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_101 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_102 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_103 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_104 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_105 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_106 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_107 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_108 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_109 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_110 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_111 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_112 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_113 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_114 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_115 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_116 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_117 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_118 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_119 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_120 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_121 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_122 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_123 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_124 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_125 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_126 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_127 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_128 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_129 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_130 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_131 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_132 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Left_133 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Left_134 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Left_135 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Left_136 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Left_137 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Left_138 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Left_139 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Left_140 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Left_141 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_142 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_143 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_144 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_145 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_146 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_147 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_148 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_149 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_150 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_151 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_152 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_153 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_154 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_155 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_156 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_157 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_158 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_159 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_160 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_161 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_162 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_163 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_164 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_165 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_166 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_167 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_168 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_169 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_170 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_171 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_172 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_173 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_174 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_175 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_176 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_177 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_178 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_179 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_180 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_181 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_182 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_183 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_184 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_185 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_186 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_187 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_188 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_189 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_190 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_191 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_192 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_193 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_194 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_195 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_196 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_197 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_198 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_199 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_200 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_201 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_202 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_203 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_204 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_205 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_206 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_207 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_208 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_209 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_210 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_211 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_212 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_213 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_214 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_215 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_216 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_217 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_218 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_219 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_220 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_221 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_222 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_223 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_224 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_225 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_226 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_227 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_228 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_229 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_230 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_231 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_232 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_233 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_234 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_235 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_236 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_237 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_238 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_239 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_240 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_241 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_242 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_243 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_244 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_245 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_246 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_247 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_248 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_249 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_250 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_251 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_252 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_253 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_254 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_255 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_256 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_257 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_258 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_259 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_260 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_261 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_262 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_263 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_264 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_265 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_266 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_267 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_268 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_269 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_270 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_271 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_272 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_273 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_274 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_275 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_276 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_277 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_278 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_279 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_280 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_281 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_282 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_283 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_284 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_285 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_286 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_287 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_288 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_289 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_290 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_291 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_292 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_293 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_294 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_295 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_296 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_297 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_298 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_299 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_300 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_301 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_302 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_303 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_304 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_305 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_306 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_307 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_308 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_309 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_310 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_311 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_312 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_313 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_314 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_315 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_316 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_317 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_318 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_319 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_320 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_321 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_322 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_323 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_324 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_325 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_326 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_327 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_328 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_329 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_330 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_331 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_332 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_333 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_334 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_335 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_336 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_337 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_338 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_339 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_340 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_341 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_342 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_343 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_344 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_345 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_346 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_347 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_348 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_349 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_350 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_351 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_352 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_353 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_354 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_355 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_356 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_357 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_358 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_359 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_360 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_361 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_362 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_363 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_364 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_365 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_366 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_367 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_368 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_369 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_370 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_371 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_372 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_373 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_374 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_375 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_376 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_377 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_378 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_379 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_380 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_381 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_382 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_383 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_384 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_385 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_386 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_387 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_388 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_389 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_390 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_391 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_392 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_393 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_394 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_395 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_396 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_397 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_398 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_399 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_400 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_401 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_402 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_403 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_404 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_405 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_406 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_407 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_408 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_409 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_410 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_411 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_412 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_413 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_414 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_415 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_416 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_417 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_418 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_419 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_420 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_421 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_422 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_423 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_424 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_425 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_426 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_427 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_428 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_429 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_430 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_431 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_432 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_433 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_434 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_435 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_436 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_437 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_438 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_439 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_440 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_441 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_442 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_443 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_444 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_445 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_446 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_447 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_448 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_449 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_450 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_451 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_452 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_453 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_454 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_455 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_456 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_457 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_458 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_459 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_460 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_461 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_462 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_463 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_464 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_465 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_466 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_467 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_468 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_469 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_470 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_471 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_472 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_473 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_474 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_475 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_476 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_477 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_478 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_479 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_480 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_481 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_482 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_483 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_484 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_485 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_486 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_487 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_488 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_489 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_490 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_491 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_492 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_493 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_494 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_495 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_496 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_497 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_498 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_499 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_500 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_501 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_502 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_503 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_504 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_505 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_506 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_507 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_508 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_509 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_510 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_511 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_512 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_513 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_514 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_515 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_516 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_517 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_518 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_519 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_520 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_521 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_522 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_523 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_524 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_525 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_526 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_527 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_528 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_529 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_530 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_531 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_532 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_533 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_534 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_535 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_536 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_537 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_538 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_539 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_540 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_541 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_542 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_543 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_544 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_545 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_546 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_547 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_548 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_549 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_550 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_551 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_552 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_553 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_554 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_555 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_556 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_557 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_558 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_559 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_560 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_561 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_562 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_563 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_564 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_565 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_566 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_567 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_568 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_569 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_570 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_571 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_572 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_573 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_574 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_575 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_576 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_577 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_578 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_579 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_580 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_581 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_582 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_583 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_584 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_585 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_586 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_587 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_588 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_589 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_590 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_591 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_592 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_593 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_594 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_595 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_596 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_597 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_598 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_599 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_600 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_601 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_602 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_603 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_604 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_605 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_606 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_607 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_608 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_609 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_610 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_611 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_612 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_613 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_614 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_615 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_616 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_617 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_618 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_619 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_620 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_621 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_622 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_623 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_624 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_625 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_626 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_627 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_628 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_629 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_630 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_631 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_632 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_633 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_634 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_635 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_636 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_637 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_638 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_639 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_640 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_641 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_642 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_643 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_644 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_645 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_646 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_647 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_648 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_649 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_650 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_651 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_652 (.VDD(VDD),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output1 (.I(net1),
    .Z(Co),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output2 (.I(net2),
    .Z(E1BEG[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output3 (.I(net3),
    .Z(E1BEG[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output4 (.I(net4),
    .Z(E1BEG[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output5 (.I(net5),
    .Z(E1BEG[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output6 (.I(net6),
    .Z(E2BEG[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output7 (.I(net7),
    .Z(E2BEG[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output8 (.I(net8),
    .Z(E2BEG[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output9 (.I(net9),
    .Z(E2BEG[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output10 (.I(net10),
    .Z(E2BEG[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output11 (.I(net11),
    .Z(E2BEG[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output12 (.I(net12),
    .Z(E2BEG[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output13 (.I(net13),
    .Z(E2BEG[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output14 (.I(net14),
    .Z(E2BEGb[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output15 (.I(net15),
    .Z(E2BEGb[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output16 (.I(net16),
    .Z(E2BEGb[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output17 (.I(net17),
    .Z(E2BEGb[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output18 (.I(net18),
    .Z(E2BEGb[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output19 (.I(net19),
    .Z(E2BEGb[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output20 (.I(net20),
    .Z(E2BEGb[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output21 (.I(net21),
    .Z(E2BEGb[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output22 (.I(net22),
    .Z(E6BEG[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output23 (.I(net23),
    .Z(E6BEG[10]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output24 (.I(net24),
    .Z(E6BEG[11]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output25 (.I(net25),
    .Z(E6BEG[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output26 (.I(net26),
    .Z(E6BEG[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output27 (.I(net27),
    .Z(E6BEG[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output28 (.I(net28),
    .Z(E6BEG[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output29 (.I(net29),
    .Z(E6BEG[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output30 (.I(net30),
    .Z(E6BEG[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output31 (.I(net31),
    .Z(E6BEG[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output32 (.I(net32),
    .Z(E6BEG[8]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output33 (.I(net33),
    .Z(E6BEG[9]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output34 (.I(net34),
    .Z(EE4BEG[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output35 (.I(net35),
    .Z(EE4BEG[10]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output36 (.I(net36),
    .Z(EE4BEG[11]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output37 (.I(net37),
    .Z(EE4BEG[12]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output38 (.I(net38),
    .Z(EE4BEG[13]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output39 (.I(net39),
    .Z(EE4BEG[14]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output40 (.I(net40),
    .Z(EE4BEG[15]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output41 (.I(net41),
    .Z(EE4BEG[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output42 (.I(net42),
    .Z(EE4BEG[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output43 (.I(net43),
    .Z(EE4BEG[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output44 (.I(net44),
    .Z(EE4BEG[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output45 (.I(net45),
    .Z(EE4BEG[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output46 (.I(net46),
    .Z(EE4BEG[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output47 (.I(net47),
    .Z(EE4BEG[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output48 (.I(net48),
    .Z(EE4BEG[8]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output49 (.I(net49),
    .Z(EE4BEG[9]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output50 (.I(net50),
    .Z(FrameData_O[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output51 (.I(net51),
    .Z(FrameData_O[10]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output52 (.I(net52),
    .Z(FrameData_O[11]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output53 (.I(net53),
    .Z(FrameData_O[12]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output54 (.I(net54),
    .Z(FrameData_O[13]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output55 (.I(net55),
    .Z(FrameData_O[14]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output56 (.I(net56),
    .Z(FrameData_O[15]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output57 (.I(net57),
    .Z(FrameData_O[16]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output58 (.I(net58),
    .Z(FrameData_O[17]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output59 (.I(net59),
    .Z(FrameData_O[18]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output60 (.I(net60),
    .Z(FrameData_O[19]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output61 (.I(net61),
    .Z(FrameData_O[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output62 (.I(net62),
    .Z(FrameData_O[20]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output63 (.I(net63),
    .Z(FrameData_O[21]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output64 (.I(net64),
    .Z(FrameData_O[22]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output65 (.I(net65),
    .Z(FrameData_O[23]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output66 (.I(net66),
    .Z(FrameData_O[24]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output67 (.I(net67),
    .Z(FrameData_O[25]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output68 (.I(net68),
    .Z(FrameData_O[26]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output69 (.I(net69),
    .Z(FrameData_O[27]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output70 (.I(net70),
    .Z(FrameData_O[28]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output71 (.I(net71),
    .Z(FrameData_O[29]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output72 (.I(net72),
    .Z(FrameData_O[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output73 (.I(net73),
    .Z(FrameData_O[30]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output74 (.I(net74),
    .Z(FrameData_O[31]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output75 (.I(net75),
    .Z(FrameData_O[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output76 (.I(net76),
    .Z(FrameData_O[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output77 (.I(net77),
    .Z(FrameData_O[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output78 (.I(net78),
    .Z(FrameData_O[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output79 (.I(net79),
    .Z(FrameData_O[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output80 (.I(net80),
    .Z(FrameData_O[8]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output81 (.I(net81),
    .Z(FrameData_O[9]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output82 (.I(net82),
    .Z(FrameStrobe_O[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output83 (.I(net83),
    .Z(FrameStrobe_O[10]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output84 (.I(net84),
    .Z(FrameStrobe_O[11]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output85 (.I(net85),
    .Z(FrameStrobe_O[12]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output86 (.I(net86),
    .Z(FrameStrobe_O[13]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output87 (.I(net87),
    .Z(FrameStrobe_O[14]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output88 (.I(net88),
    .Z(FrameStrobe_O[15]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output89 (.I(net89),
    .Z(FrameStrobe_O[16]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output90 (.I(net90),
    .Z(FrameStrobe_O[17]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output91 (.I(net91),
    .Z(FrameStrobe_O[18]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output92 (.I(net92),
    .Z(FrameStrobe_O[19]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output93 (.I(net93),
    .Z(FrameStrobe_O[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output94 (.I(net94),
    .Z(FrameStrobe_O[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output95 (.I(net95),
    .Z(FrameStrobe_O[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output96 (.I(net96),
    .Z(FrameStrobe_O[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output97 (.I(net97),
    .Z(FrameStrobe_O[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output98 (.I(net98),
    .Z(FrameStrobe_O[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output99 (.I(net99),
    .Z(FrameStrobe_O[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output100 (.I(net100),
    .Z(FrameStrobe_O[8]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output101 (.I(net101),
    .Z(FrameStrobe_O[9]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output102 (.I(net102),
    .Z(N1BEG[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output103 (.I(net103),
    .Z(N1BEG[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output104 (.I(net104),
    .Z(N1BEG[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output105 (.I(net105),
    .Z(N1BEG[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output106 (.I(net106),
    .Z(N2BEG[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output107 (.I(net107),
    .Z(N2BEG[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output108 (.I(net108),
    .Z(N2BEG[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output109 (.I(net109),
    .Z(N2BEG[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output110 (.I(net110),
    .Z(N2BEG[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output111 (.I(net111),
    .Z(N2BEG[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output112 (.I(net112),
    .Z(N2BEG[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output113 (.I(net113),
    .Z(N2BEG[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output114 (.I(net114),
    .Z(N2BEGb[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output115 (.I(net115),
    .Z(N2BEGb[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output116 (.I(net116),
    .Z(N2BEGb[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output117 (.I(net117),
    .Z(N2BEGb[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output118 (.I(net118),
    .Z(N2BEGb[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output119 (.I(net119),
    .Z(N2BEGb[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output120 (.I(net120),
    .Z(N2BEGb[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output121 (.I(net121),
    .Z(N2BEGb[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output122 (.I(net122),
    .Z(N4BEG[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output123 (.I(net123),
    .Z(N4BEG[10]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output124 (.I(net124),
    .Z(N4BEG[11]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output125 (.I(net125),
    .Z(N4BEG[12]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output126 (.I(net126),
    .Z(N4BEG[13]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output127 (.I(net127),
    .Z(N4BEG[14]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output128 (.I(net128),
    .Z(N4BEG[15]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output129 (.I(net129),
    .Z(N4BEG[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output130 (.I(net130),
    .Z(N4BEG[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output131 (.I(net131),
    .Z(N4BEG[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output132 (.I(net132),
    .Z(N4BEG[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output133 (.I(net133),
    .Z(N4BEG[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output134 (.I(net134),
    .Z(N4BEG[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output135 (.I(net135),
    .Z(N4BEG[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output136 (.I(net136),
    .Z(N4BEG[8]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output137 (.I(net137),
    .Z(N4BEG[9]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output138 (.I(net138),
    .Z(NN4BEG[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output139 (.I(net139),
    .Z(NN4BEG[10]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output140 (.I(net140),
    .Z(NN4BEG[11]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output141 (.I(net141),
    .Z(NN4BEG[12]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output142 (.I(net142),
    .Z(NN4BEG[13]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output143 (.I(net143),
    .Z(NN4BEG[14]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output144 (.I(net144),
    .Z(NN4BEG[15]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output145 (.I(net145),
    .Z(NN4BEG[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output146 (.I(net146),
    .Z(NN4BEG[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output147 (.I(net147),
    .Z(NN4BEG[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output148 (.I(net148),
    .Z(NN4BEG[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output149 (.I(net149),
    .Z(NN4BEG[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output150 (.I(net150),
    .Z(NN4BEG[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output151 (.I(net151),
    .Z(NN4BEG[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output152 (.I(net152),
    .Z(NN4BEG[8]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output153 (.I(net153),
    .Z(NN4BEG[9]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output154 (.I(net154),
    .Z(S1BEG[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output155 (.I(net155),
    .Z(S1BEG[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output156 (.I(net156),
    .Z(S1BEG[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output157 (.I(net157),
    .Z(S1BEG[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output158 (.I(net158),
    .Z(S2BEG[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output159 (.I(net159),
    .Z(S2BEG[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output160 (.I(net160),
    .Z(S2BEG[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output161 (.I(net161),
    .Z(S2BEG[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output162 (.I(net162),
    .Z(S2BEG[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output163 (.I(net163),
    .Z(S2BEG[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output164 (.I(net164),
    .Z(S2BEG[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output165 (.I(net165),
    .Z(S2BEG[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output166 (.I(net166),
    .Z(S2BEGb[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output167 (.I(net167),
    .Z(S2BEGb[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output168 (.I(net168),
    .Z(S2BEGb[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output169 (.I(net169),
    .Z(S2BEGb[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output170 (.I(net170),
    .Z(S2BEGb[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output171 (.I(net171),
    .Z(S2BEGb[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output172 (.I(net172),
    .Z(S2BEGb[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output173 (.I(net173),
    .Z(S2BEGb[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output174 (.I(net174),
    .Z(S4BEG[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output175 (.I(net175),
    .Z(S4BEG[10]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output176 (.I(net176),
    .Z(S4BEG[11]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output177 (.I(net177),
    .Z(S4BEG[12]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output178 (.I(net178),
    .Z(S4BEG[13]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output179 (.I(net179),
    .Z(S4BEG[14]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output180 (.I(net180),
    .Z(S4BEG[15]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output181 (.I(net181),
    .Z(S4BEG[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output182 (.I(net182),
    .Z(S4BEG[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output183 (.I(net183),
    .Z(S4BEG[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output184 (.I(net184),
    .Z(S4BEG[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output185 (.I(net185),
    .Z(S4BEG[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output186 (.I(net186),
    .Z(S4BEG[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output187 (.I(net187),
    .Z(S4BEG[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output188 (.I(net188),
    .Z(S4BEG[8]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output189 (.I(net189),
    .Z(S4BEG[9]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output190 (.I(net190),
    .Z(SS4BEG[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output191 (.I(net191),
    .Z(SS4BEG[10]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output192 (.I(net192),
    .Z(SS4BEG[11]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output193 (.I(net193),
    .Z(SS4BEG[12]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output194 (.I(net194),
    .Z(SS4BEG[13]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output195 (.I(net195),
    .Z(SS4BEG[14]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output196 (.I(net196),
    .Z(SS4BEG[15]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output197 (.I(net197),
    .Z(SS4BEG[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output198 (.I(net198),
    .Z(SS4BEG[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output199 (.I(net199),
    .Z(SS4BEG[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output200 (.I(net200),
    .Z(SS4BEG[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output201 (.I(net201),
    .Z(SS4BEG[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output202 (.I(net202),
    .Z(SS4BEG[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output203 (.I(net203),
    .Z(SS4BEG[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output204 (.I(net204),
    .Z(SS4BEG[8]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output205 (.I(net205),
    .Z(SS4BEG[9]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output206 (.I(net206),
    .Z(UserCLKo),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output207 (.I(net207),
    .Z(W1BEG[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output208 (.I(net208),
    .Z(W1BEG[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output209 (.I(net209),
    .Z(W1BEG[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output210 (.I(net210),
    .Z(W1BEG[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output211 (.I(net211),
    .Z(W2BEG[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output212 (.I(net212),
    .Z(W2BEG[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output213 (.I(net213),
    .Z(W2BEG[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output214 (.I(net214),
    .Z(W2BEG[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output215 (.I(net215),
    .Z(W2BEG[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output216 (.I(net216),
    .Z(W2BEG[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output217 (.I(net217),
    .Z(W2BEG[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output218 (.I(net218),
    .Z(W2BEG[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output219 (.I(net219),
    .Z(W2BEGb[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output220 (.I(net220),
    .Z(W2BEGb[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output221 (.I(net221),
    .Z(W2BEGb[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output222 (.I(net222),
    .Z(W2BEGb[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output223 (.I(net223),
    .Z(W2BEGb[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output224 (.I(net224),
    .Z(W2BEGb[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output225 (.I(net225),
    .Z(W2BEGb[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output226 (.I(net226),
    .Z(W2BEGb[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output227 (.I(net227),
    .Z(W6BEG[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output228 (.I(net228),
    .Z(W6BEG[10]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output229 (.I(net229),
    .Z(W6BEG[11]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output230 (.I(net230),
    .Z(W6BEG[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output231 (.I(net231),
    .Z(W6BEG[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output232 (.I(net232),
    .Z(W6BEG[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output233 (.I(net233),
    .Z(W6BEG[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output234 (.I(net234),
    .Z(W6BEG[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output235 (.I(net235),
    .Z(W6BEG[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output236 (.I(net236),
    .Z(W6BEG[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output237 (.I(net237),
    .Z(W6BEG[8]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output238 (.I(net238),
    .Z(W6BEG[9]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output239 (.I(net239),
    .Z(WW4BEG[0]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output240 (.I(net240),
    .Z(WW4BEG[10]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output241 (.I(net241),
    .Z(WW4BEG[11]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output242 (.I(net242),
    .Z(WW4BEG[12]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output243 (.I(net243),
    .Z(WW4BEG[13]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output244 (.I(net244),
    .Z(WW4BEG[14]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output245 (.I(net245),
    .Z(WW4BEG[15]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output246 (.I(net246),
    .Z(WW4BEG[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output247 (.I(net247),
    .Z(WW4BEG[2]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output248 (.I(net248),
    .Z(WW4BEG[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output249 (.I(net249),
    .Z(WW4BEG[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output250 (.I(net250),
    .Z(WW4BEG[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output251 (.I(net251),
    .Z(WW4BEG[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output252 (.I(net252),
    .Z(WW4BEG[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output253 (.I(net253),
    .Z(WW4BEG[8]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 output254 (.I(net254),
    .Z(WW4BEG[9]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_regs_0_UserCLK (.I(UserCLK),
    .Z(UserCLK_regs),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_UserCLK (.I(UserCLK),
    .Z(clknet_0_UserCLK),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_0__f_UserCLK (.I(clknet_0_UserCLK),
    .Z(clknet_1_0__leaf_UserCLK),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_UserCLK_regs (.I(UserCLK_regs),
    .Z(clknet_0_UserCLK_regs),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_0__f_UserCLK_regs (.I(clknet_0_UserCLK_regs),
    .Z(clknet_1_0__leaf_UserCLK_regs),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_1__f_UserCLK_regs (.I(clknet_0_UserCLK_regs),
    .Z(clknet_1_1__leaf_UserCLK_regs),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_1 (.I(E6END[3]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_2 (.I(E6END[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_3 (.I(E6END[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_4 (.I(EE4END[13]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_5 (.I(EE4END[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_6 (.I(EE4END[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_7 (.I(EE4END[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_8 (.I(EE4END[8]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_9 (.I(EE4END[9]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_10 (.I(\Inst_LUT4AB_switch_matrix.JW2BEG2 ),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_11 (.I(N4END[10]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_12 (.I(N4END[11]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_13 (.I(N4END[12]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_14 (.I(N4END[13]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_15 (.I(N4END[14]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_16 (.I(N4END[15]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_17 (.I(N4END[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_18 (.I(N4END[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_19 (.I(N4END[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_20 (.I(N4END[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_21 (.I(N4END[8]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_22 (.I(N4END[9]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_23 (.I(NN4END[10]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_24 (.I(NN4END[11]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_25 (.I(NN4END[12]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_26 (.I(NN4END[13]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_27 (.I(NN4END[14]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_28 (.I(NN4END[15]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_29 (.I(NN4END[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_30 (.I(NN4END[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_31 (.I(NN4END[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_32 (.I(NN4END[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_33 (.I(NN4END[8]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_34 (.I(NN4END[9]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_35 (.I(SS4END[10]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_36 (.I(SS4END[11]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_37 (.I(SS4END[12]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_38 (.I(SS4END[13]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_39 (.I(SS4END[14]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_40 (.I(SS4END[15]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_41 (.I(SS4END[4]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_42 (.I(SS4END[5]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_43 (.I(SS4END[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_44 (.I(SS4END[7]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_45 (.I(SS4END[8]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_46 (.I(SS4END[9]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_47 (.I(net230),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_48 (.I(net237),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_49 (.I(net234),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_50 (.I(net248),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_51 (.I(B),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_52 (.I(EE4END[15]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_53 (.I(N4END[13]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_54 (.I(SS4END[12]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_55 (.I(W2MID[6]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_56 (.I(net233),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_57 (.I(net236),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_58 (.I(W6END[1]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_59 (.I(net251),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_60 (.I(N4END[13]),
    .VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_264 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_271 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_360 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_370 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_378 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_384 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_396 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_402 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_410 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_438 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_450 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_466 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_474 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_478 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_494 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_498 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_277 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_279 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_288 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_322 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_349 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_364 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_374 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_418 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_446 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_478 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_486 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_498 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_249 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_288 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_310 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_314 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_329 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_362 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_372 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_441 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_449 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_453 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_457 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_473 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_278 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_294 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_348 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_376 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_383 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_389 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_401 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_411 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_419 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_428 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_460 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_476 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_498 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_166 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_223 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_279 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_312 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_314 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_323 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_383 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_393 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_401 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_427 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_443 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_451 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_457 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_465 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_475 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_492 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_176 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_332 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_334 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_372 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_374 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_395 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_407 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_415 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_419 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_422 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_454 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_462 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_466 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_474 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_492 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_133 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_233 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_279 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_283 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_314 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_349 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_387 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_427 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_444 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_452 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_454 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_457 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_461 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_494 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_498 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_86 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_238 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_246 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_282 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_284 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_327 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_329 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_352 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_373 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_377 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_398 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_419 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_422 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_430 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_432 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_488 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_498 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_211 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_219 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_240 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_287 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_317 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_321 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_374 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_402 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_406 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_447 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_477 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_498 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_30 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_128 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_253 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_257 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_259 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_282 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_290 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_343 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_347 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_349 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_372 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_374 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_488 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_498 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_238 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_257 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_265 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_269 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_290 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_294 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_300 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_308 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_312 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_314 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_317 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_325 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_327 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_366 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_374 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_378 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_425 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_427 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_448 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_472 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_156 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_205 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_264 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_282 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_290 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_292 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_313 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_352 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_419 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_442 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_444 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_485 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_489 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_492 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_51 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_213 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_221 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_252 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_254 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_313 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_317 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_341 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_362 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_364 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_387 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_395 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_496 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_498 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_74 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_165 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_228 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_277 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_279 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_282 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_299 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_329 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_352 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_356 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_361 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_401 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_405 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_408 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_485 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_489 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_492 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_71 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_251 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_272 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_280 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_284 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_286 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_293 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_317 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_339 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_341 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_374 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_382 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_384 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_407 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_411 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_413 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_496 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_498 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_302 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_310 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_356 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_378 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_386 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_419 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_436 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_438 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_467 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_488 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_492 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_198 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_233 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_313 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_317 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_338 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_342 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_344 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_355 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_363 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_387 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_403 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_440 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_469 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_473 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_498 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_126 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_232 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_282 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_304 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_308 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_329 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_380 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_396 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_400 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_417 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_419 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_487 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_489 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_492 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_171 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_226 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_242 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_267 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_271 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_273 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_314 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_317 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_371 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_379 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_383 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_407 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_409 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_428 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_430 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_497 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_220 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_274 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_278 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_282 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_290 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_294 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_347 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_349 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_392 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_394 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_434 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_498 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_116 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_120 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_255 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_308 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_312 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_314 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_337 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_345 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_369 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_387 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_497 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_121 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_206 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_237 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_245 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_267 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_275 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_279 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_282 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_374 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_408 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_422 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_424 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_469 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_498 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_14 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_185 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_218 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_304 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_312 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_314 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_362 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_384 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_452 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_454 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_496 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_498 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_76 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_131 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_178 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_182 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_277 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_279 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_297 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_299 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_332 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_348 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_437 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_498 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_53 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_113 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_134 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_255 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_259 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_312 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_314 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_369 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_391 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_432 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_434 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_457 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_498 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_45 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_49 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_254 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_256 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_277 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_279 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_342 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_349 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_362 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_370 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_374 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_437 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_487 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_489 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_498 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_100 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_125 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_242 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_255 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_259 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_313 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_317 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_321 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_328 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_381 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_387 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_395 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_399 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_421 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_453 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_469 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_490 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_492 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_168 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_232 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_266 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_274 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_278 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_282 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_342 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_352 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_406 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_468 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_489 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_498 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_99 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_141 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_239 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_243 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_251 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_305 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_313 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_317 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_325 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_329 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_362 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_364 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_453 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_489 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_192 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_200 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_322 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_346 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_422 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_449 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_473 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_477 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_488 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_498 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_46 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_48 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_222 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_224 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_251 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_259 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_263 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_284 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_314 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_337 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_341 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_360 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_382 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_384 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_387 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_395 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_399 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_457 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_461 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_498 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_80 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_117 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_270 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_274 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_282 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_366 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_399 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_477 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_479 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_498 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_195 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_238 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_242 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_267 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_322 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_364 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_387 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_391 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_437 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_158 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_191 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_269 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_277 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_279 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_282 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_332 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_413 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_489 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_492 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_27 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_83 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_184 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_249 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_302 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_304 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_325 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_346 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_373 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_387 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_399 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_403 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_475 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_497 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_16 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_226 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_228 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_249 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_253 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_282 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_284 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_392 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_469 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_488 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_498 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_41 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_103 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_237 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_263 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_271 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_312 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_314 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_325 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_395 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_431 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_433 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_454 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_457 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_459 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_480 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_497 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_68 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_92 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_96 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_119 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_196 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_220 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_224 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_226 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_259 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_333 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_349 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_352 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_367 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_369 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_385 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_387 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_408 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_454 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_456 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_485 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_498 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_193 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_226 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_242 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_255 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_302 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_304 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_317 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_384 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_395 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_403 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_468 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_489 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_497 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_62 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_64 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_79 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_147 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_220 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_224 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_258 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_282 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_336 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_344 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_348 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_352 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_405 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_413 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_498 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_155 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_227 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_243 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_303 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_327 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_361 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_363 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_384 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_395 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_397 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_430 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_490 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_492 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_111 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_137 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_144 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_202 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_218 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_271 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_279 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_282 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_290 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_292 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_333 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_349 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_372 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_376 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_378 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_419 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_442 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_498 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_115 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_263 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_296 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_304 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_325 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_383 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_387 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_420 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_465 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_486 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_106 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_118 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_276 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_282 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_290 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_292 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_325 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_327 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_348 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_372 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_466 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_468 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_489 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_498 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_25 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_230 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_238 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_242 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_298 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_314 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_369 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_407 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_409 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_445 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_447 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_489 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_187 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_189 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_266 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_274 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_278 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_342 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_352 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_356 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_422 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_466 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_498 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_23 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_33 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_102 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_167 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_228 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_255 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_257 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_310 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_314 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_337 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_345 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_367 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_379 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_383 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_424 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_132 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_150 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_154 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_282 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_290 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_292 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_345 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_349 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_352 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_488 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_498 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_22 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_32 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_77 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_181 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_183 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_204 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_268 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_276 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_300 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_308 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_312 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_314 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_317 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_321 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_382 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_384 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_387 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_393 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_431 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_452 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_454 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_457 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_484 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_67 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_105 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_255 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_276 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_282 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_348 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_362 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_418 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_488 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_498 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_164 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_172 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_251 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_309 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_342 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_407 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_409 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_439 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_465 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_220 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_222 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_243 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_282 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_326 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_348 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_360 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_401 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_403 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_468 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_492 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_89 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_162 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_251 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_313 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_317 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_384 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_433 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_468 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_497 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_151 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_153 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_227 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_278 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_302 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_304 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_377 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_489 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_498 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_6 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_57 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_61 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_82 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_84 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_161 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_169 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_308 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_337 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_498 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_148 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_201 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_248 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_302 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_304 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_362 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_418 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_437 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_439 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_492 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_73 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_75 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_314 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_336 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_407 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_454 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_463 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_496 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_498 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_4 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_63 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_199 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_207 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_209 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_216 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_269 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_322 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_382 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_384 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_422 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_451 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_453 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_468 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_489 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_492 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_122 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_124 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_157 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_232 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_240 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_244 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_251 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_283 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_403 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_497 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_8 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_10 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_268 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_317 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_338 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_422 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_492 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_173 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_233 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_263 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_285 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_287 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_314 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_317 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_418 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_450 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_454 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_139 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_255 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_279 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_282 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_322 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_343 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_442 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_464 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_466 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_487 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_489 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_498 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_233 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_241 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_255 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_357 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_359 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_383 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_431 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_433 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_454 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_52 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_54 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_78 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_194 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_276 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_307 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_348 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_398 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_400 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_417 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_419 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_483 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_492 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_98 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_109 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_146 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_170 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_243 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_337 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_339 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_387 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_410 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_412 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_442 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_463 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_465 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_483 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_496 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_498 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_24 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_26 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_35 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_208 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_279 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_302 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_367 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_397 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_399 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_432 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_469 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_471 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_492 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_13 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_43 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_149 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_177 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_213 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_243 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_267 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_312 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_314 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_395 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_437 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_463 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_479 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_69 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_97 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_159 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_175 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_179 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_232 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_253 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_269 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_282 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_284 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_305 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_316 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_422 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_442 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_461 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_487 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_489 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_492 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_37 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_39 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_60 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_87 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_91 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_107 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_130 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_136 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_174 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_247 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_263 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_267 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_269 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_312 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_314 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_325 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_327 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_383 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_457 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_485 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_72 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_114 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_123 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_127 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_236 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_238 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_257 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_261 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_349 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_352 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_402 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_404 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_417 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_419 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_498 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_70 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_104 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_138 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_142 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_163 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_180 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_186 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_190 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_203 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_212 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_214 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_233 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_237 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_264 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_274 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_278 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_303 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_305 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_326 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_348 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_376 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_440 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_474 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_478 (.VDD(VDD),
    .VNW(VDD),
    .VPW(VSS),
    .VSS(VSS));
endmodule
